library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 2**16) of integer;

  constant input_wght : mem := (
    -- bias
    -2634, -108, 222, 3427, 194, -1576, 1538, -444, 159, 365, 

    -- weights
    -- filter=0 channel=0
    0, 0, -1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 3, 1, 1, 1, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 1, 3, 0, 0, 0, 1, 1, 0, -1, 0, -1, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 2, 2, 0, 0, 0, 0, -1, -1, 0, -2, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 2, 2, 1, 1, 2, 1, 0, 0, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 3, 1, 0, 1, 2, 0, 1, 0, 0, -1, 0, -1, -1, -1, 0, -2, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 3, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 1, 1, 2, 1, 1, 0, 0, 0, 0, -1, -2, -2, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 2, 1, 0, 1, 3, 1, 2, 0, -1, 0, -1, 0, 0, -1, -2, -1, -1, 0, -1, 0, -1, -1, 0, 1, 1, 0, 2, 2, 2, 1, 1, 0, 0, 1, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 2, 0, 1, 2, 2, 1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 2, 0, 0, 0, 1, 2, 3, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 2, 2, 2, 2, 2, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 2, 0, 2, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, -1, 0, -1, 1, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, 2, 2, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 2, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, -2, -2, -1, -3, -4, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 1, 1, 0, 0, 0, -2, -2, -2, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, 1, 1, 1, 0, 0, 0, -2, -2, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, -1, 1, 1, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, -1, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 2, 2, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 2, 0, 1, 2, 3, 2, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, 1, 2, 1, 3, 3, 2, 0, 2, 0, 0, -1, 0, 0, -1, 0, -1, 0, 1, 1, 1, 2, 3, 0, 1, 0, 1, 2, 1, 0, 1, 2, 0, 0, 1, 0, 0, 0, -1, 0, -2, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, 0, 2, 1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -2, 0, 0, 0, 0, 1, 0, 0, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, -1, -3, -4, -3, -3, -3, -4, -2, -3, -3, -1, -3, -3, -3, -4, -3, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, -4, -4, -4, -3, -4, -3, -2, -2, -2, 0, -2, 0, -2, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, -4, -3, -2, -3, -4, -4, -2, -1, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, -3, -4, -3, -3, -2, -4, -3, -1, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, -4, -3, -3, -2, -2, -3, -3, -2, -2, -1, -2, 0, -2, -2, -2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -5, -4, -1, -1, -1, -3, -2, -3, -1, -2, -2, -1, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, -3, -3, -3, -2, -3, -2, -3, -1, -1, -3, -2, -3, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -2, -2, -2, -2, -2, -3, -2, -2, -3, -1, -3, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, -2, -3, -2, -3, -2, -3, -2, -3, -1, -1, -1, -2, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -3, -2, -3, -1, -4, -2, -3, -1, 0, -1, -1, -2, -1, -1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, -3, -2, -2, -2, -1, -2, -1, -3, -2, -2, -1, 0, 0, -2, -2, 0, -1, 1, 1, 0, 0, -1, -1, 1, 2, 0, -2, -2, -1, -2, -3, -1, -1, -1, -2, -2, 0, -1, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 1, 2, -3, -4, -4, -1, -1, -2, -2, -1, -2, -1, 0, -1, 0, -1, -1, -1, 0, 2, 3, 1, 0, -1, 0, 0, 0, 3, -2, -3, -2, -4, -2, -2, -1, -2, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, -1, 0, 2, -4, -4, -2, -3, -2, -3, -3, -1, 0, -1, -1, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 2, -4, -2, -3, -2, -3, -4, -3, -1, -3, -1, 0, 0, 0, -2, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 2, -3, -4, -1, -2, -3, -3, -2, -2, -2, -1, 0, -1, -2, -1, -2, -1, -1, 1, 0, 0, 1, 0, 0, 1, 0, 2, -4, -4, -2, -2, -3, -3, -3, -2, 0, -2, 0, 0, -1, -2, -2, -2, 0, 0, 0, 0, 1, 0, 1, 0, 0, 2, -5, -4, -3, -2, -3, -3, -1, 0, -1, 0, -2, -1, 0, -1, -2, -2, 0, -1, 0, 2, 1, 0, 1, 0, 0, 2, -4, -3, -3, -2, -1, -3, -2, -2, -3, -1, -1, -2, -2, -2, -2, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 2, -4, -3, -2, -3, -2, -2, -2, -2, -1, -2, -1, -3, -3, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 3, -3, -2, -4, -3, -2, -3, -1, -1, -2, -2, -2, -2, -2, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 2, 1, -4, -3, -2, -3, -4, -4, -2, -1, -2, -3, 0, -2, -1, 0, -1, 0, 0, -1, -1, 1, 0, 0, 1, 2, 1, 2, -5, -3, -4, -5, -4, -4, -3, -2, -1, -2, -1, -1, -2, -1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 2, 3, -3, -4, -4, -5, -4, -3, -2, -3, -1, -2, -1, -2, -2, -1, -1, 0, -1, -1, 0, 1, 0, 1, 2, 2, 2, 1, -4, -3, -5, -4, -5, -5, -4, -2, -3, -3, -3, -3, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 2, 3, 3, 2, 0, -1, 0, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, -1, 0, -1, 0, -1, -2, 0, 0, -1, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, -2, -2, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -2, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -2, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, -1, -1, 0, -1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, -2, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -2, -2, -2, -1, -2, 0, -1, 0, 1, 0, 1, 1, 0, 2, 1, 2, 1, 1, 1, 1, 0, 0, -1, -2, -1, -1, -3, -1, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, -2, -2, -3, -1, -3, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, -1, -2, -2, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 2, 0, 1, 1, 0, 0, -1, -1, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 1, 2, 1, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 1, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 1, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, -2, 0, 0, -1, -2, -2, 0, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -2, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, -1, -1, 0, -1, -1, 0, -2, -2, -3, -3, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, -2, -1, -2, -2, -2, -2, -2, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -3, -3, -3, -1, -1, -1, -1, -2, 0, -1, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -3, -2, -3, -3, -1, -2, -2, -2, 0, 0, 0, -1, -1, -1, 0, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 2, 2, 3, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 2, 2, 1, 1, 0, 2, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 1, 1, 1, 2, 2, 2, 0, 1, 1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 0, 1, 1, 2, 1, 1, 2, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, -2, 0, -1, -1, 0, 0, 0, 0, 1, 3, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 3, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -2, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 1, 2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -2, -1, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, -1, -2, 0, 0, -1, 0, 1, 1, 1, 1, 2, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -2, -1, 0, 0, -2, -3, -2, 0, 1, 1, 0, 1, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, -2, -1, -1, 0, 0, 1, 0, 1, 0, 1, 1, 2, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 2, 2, 2, 2, 2, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 1, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 1, 2, 1, 3, 2, 3, 4, -1, -1, -1, 0, 0, 0, -1, 0, 1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 3, 2, 1, 3, 3, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 1, 0, 1, 2, 1, 2, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 2, 2, 1, 3, 2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 2, 1, 1, 2, 3, 3, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 3, 1, 1, 2, 3, 1, -2, -3, -2, -4, -4, -3, -3, -1, -1, 0, -1, -1, -2, -2, 0, 0, 2, 2, 3, 2, 3, 2, 2, 1, 3, 2, -4, -2, -3, -1, -3, -3, -1, -2, 0, 0, 0, 0, 0, -1, 0, 0, 2, 4, 3, 2, 1, 1, 0, 2, 2, 1, -3, -1, -2, 0, -1, -1, -1, -1, 0, -1, 0, 1, 0, 0, 0, 1, 2, 5, 3, 2, 1, 1, 0, 0, 1, 3, -4, -2, -1, 0, 0, 0, -2, -1, -1, 0, 0, 0, 1, 0, -1, 1, 3, 4, 5, 4, 3, 3, 0, 0, 0, 0, -4, -2, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 1, 0, -1, 0, 2, 3, 3, 2, 3, 3, 0, 1, 1, 1, -2, -3, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 2, 4, 3, 2, 1, 3, 1, 0, 0, -4, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, 0, 2, 4, 3, 3, 1, 2, 1, 1, 0, -2, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -3, -2, 0, 1, 3, 3, 0, 2, 0, 0, 0, 0, -3, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, -3, -1, -1, 0, 0, 1, 1, 2, 0, 0, 0, 0, 1, -2, 0, 0, 0, 0, 0, -1, -1, -1, -3, 0, 0, 0, -1, -2, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, -1, 0, -2, -2, -3, 0, -2, -1, -2, -3, -2, -2, 0, 0, 1, 1, 0, 0, 0, 0, 2, -2, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, 0, -2, -3, -3, -2, -3, 0, 1, 1, 2, 0, -1, 0, 1, 4, -1, 0, -1, -1, -1, 0, -1, -2, -1, -1, -2, 0, -2, -1, -2, -3, -1, 0, 0, 2, 0, 0, -1, 0, 0, 3, -1, 0, 0, 0, 0, 0, 0, -2, -1, 0, -2, 0, -3, -3, -2, -4, -3, -1, 0, 0, 0, 1, 0, -1, 0, 3, 0, -1, -1, 0, 0, -1, 0, -2, -2, -1, -1, 0, -1, -2, -2, -2, -3, 0, 0, 0, 0, 0, -2, -1, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -2, -3, -2, -2, -1, 0, 0, 0, 0, -1, 0, 0, 3, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -3, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, -1, -2, -1, -1, -1, -1, 1, 1, 0, 0, 0, -1, -1, 0, 1, -1, -1, 0, -1, 0, 0, 0, 1, 1, 1, -1, -2, -2, 0, 0, 0, 0, 1, 1, 1, 1, -1, -1, -1, 0, 0, -2, -1, -1, -1, 0, -1, 1, 2, 2, 0, -2, -2, -2, -3, -1, 0, 0, 1, 1, 2, 2, 0, 0, 0, 0, 1, -1, -3, -1, 0, -1, 0, 0, 0, 1, 0, -2, -1, -3, -2, 0, 0, 2, 2, 1, 0, 0, 2, 1, 0, 2, 1, -1, -1, -1, 0, -1, -2, -1, -1, 0, 0, 0, -1, -3, -2, -1, 0, 1, 1, 2, 1, 0, 0, 0, 1, 2, 1, -1, 0, -2, -1, -1, -1, -1, 0, 0, -2, -1, -1, -1, -1, -1, 0, 0, 1, 2, 1, 3, 1, 0, 1, 1, 1, -1, -2, 0, -2, -1, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 2, 2, 2, 2, 2, 2, 1, -2, -1, 0, 0, -3, -3, -1, -1, -1, 0, -1, 0, 0, 1, 0, 2, 3, 1, 1, 4, 4, 1, 1, 2, 1, 2, -4, -1, -2, -1, -3, -3, -3, -1, 0, 0, 0, 0, 0, 0, 0, 3, 3, 3, 0, 3, 4, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 2, 2, 1, 4, 5, 6, 6, 7, 6, 4, 3, 2, 0, 0, -2, 0, 1, 0, 0, 0, -2, -1, -4, -1, -1, -1, 0, 0, 2, 3, 3, 4, 6, 4, 5, 5, 4, 1, 0, 0, -1, 0, 1, 1, 0, 0, -2, -2, -4, -2, -3, -1, -2, 0, 0, 2, 2, 3, 4, 5, 4, 2, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -2, 0, -2, -2, -1, 1, 0, 1, 2, 2, 4, 2, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 2, 1, 2, 0, -1, 0, -1, 0, -1, 0, 1, 0, 3, 2, 0, 1, 3, 2, 0, 1, 0, 0, 2, 1, 1, 2, 2, 3, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 2, 1, 3, 2, 2, 2, 0, 0, 0, 0, 1, 1, 1, 4, 3, 2, 0, 0, 0, 0, 1, 0, 0, 0, 2, 0, 0, 3, 2, 3, 1, 1, 1, 0, 1, 1, 0, 1, 3, 4, 3, 3, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 2, 1, 1, 2, 1, 0, 0, 0, 2, 2, 2, 1, 3, 3, 4, 4, 0, 1, 2, 1, 1, 2, 2, 4, 3, 2, 2, 1, 2, 2, 0, 0, 0, 0, 1, 2, 2, 3, 2, 4, 3, 5, 2, 3, 1, 2, 2, 3, 3, 5, 3, 3, 4, 1, 3, 0, 0, 0, 0, 0, 1, 0, 2, 2, 4, 4, 4, 5, 1, 2, 3, 3, 3, 3, 5, 5, 3, 3, 3, 2, 2, 1, 0, 0, 0, 0, 0, 1, 2, 4, 4, 4, 5, 6, 1, 1, 3, 2, 2, 2, 2, 4, 2, 1, 0, 0, 0, 0, 0, -1, -1, -1, -2, 0, 1, 2, 4, 3, 5, 7, 0, 1, 1, 1, 0, 1, 3, 2, 0, 1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 3, 4, 4, 6, 0, 0, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 3, 2, 3, 3, 5, 4, 0, 0, 0, 1, 1, 1, 3, 2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 2, 2, 2, 2, 2, 2, 3, 0, 0, 0, 1, 0, 2, 1, 2, 1, -1, -1, 0, 2, 2, 0, 2, 0, 1, 2, 2, 4, 3, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 2, 2, 0, 0, 1, 2, 2, 2, 1, 2, 2, 3, 2, 0, 0, 0, -2, 0, -1, 1, 1, 0, 0, 0, 1, 2, 0, 2, 0, 0, 0, 1, 0, 2, 1, 1, 1, 2, 2, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 3, 3, 2, 2, 0, 1, 0, 0, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 2, 2, 3, 2, 2, 2, 2, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 3, 2, 3, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, -2, -2, -3, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 3, 1, 1, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, 0, -2, 0, 0, 0, 1, 0, 1, 3, 4, 3, 4, 3, 1, 0, 0, -2, -1, -1, -1, -1, -1, -1, -2, 0, 0, -1, 0, -1, 0, 1, 0, 2, 2, 4, 3, 2, 3, 1, 1, -1, -1, -4, -2, -1, 0, -2, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, -2, -2, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 1, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 1, 2, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 1, 0, 1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 2, 3, 1, 0, 0, 0, 0, 0, 2, 3, 4, 4, 5, 5, 6, 7, 7, 5, 4, 3, 0, -2, -2, -2, 0, 0, 0, 0, -1, -2, -2, -1, -1, 0, 0, 1, 1, 3, 4, 3, 5, 6, 5, 5, 5, 3, 0, 0, -1, -2, -1, 1, 0, 0, 0, -1, -1, -4, -4, -4, -1, 0, 0, 1, 1, 3, 3, 5, 5, 4, 2, 3, 0, -1, -1, 0, 0, 1, 1, 0, 0, -1, -2, -2, -3, -2, -2, -1, -1, 0, 0, 1, 1, 4, 3, 3, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, 1, 3, 1, 1, 1, 1, 1, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 2, 2, 1, 0, -1, -1, 0, 0, 0, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 2, 3, 2, 4, -1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 2, 3, 3, 3, 4, -1, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 2, 2, 0, 0, 0, -1, 1, 0, 0, 3, 3, 3, 4, 0, 0, 2, 1, 0, 0, 1, 0, 0, 0, 1, 0, 2, 1, 0, 0, -1, 0, 0, 0, 1, 2, 1, 2, 4, 7, 0, 0, 1, 3, 2, 1, 1, 1, 1, 2, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 2, 1, 2, 3, 5, 7, 0, 1, 2, 2, 2, 2, 2, 3, 3, 1, 2, 2, 0, 0, -1, -2, 0, -1, -1, 0, 1, 2, 2, 5, 6, 6, 0, 1, 3, 2, 3, 4, 3, 4, 4, 3, 2, 0, 0, 0, -2, -2, -1, -3, 0, 0, 2, 3, 3, 5, 7, 7, 0, 2, 2, 2, 2, 4, 3, 4, 3, 2, 0, 0, 0, -1, -1, -1, -2, -1, -3, -1, 0, 2, 4, 6, 6, 8, 0, 1, 0, 2, 2, 3, 2, 3, 1, 0, -1, -1, -1, -1, 0, -3, -2, -3, -1, -2, 1, 3, 4, 4, 5, 6, -1, 1, 1, 2, 1, 3, 3, 1, 0, 0, 0, 0, -1, 0, -1, -1, -3, -2, 0, 0, 0, 3, 4, 4, 5, 6, 1, 0, 0, 0, 0, 3, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 4, 0, 1, 0, 0, 1, 0, 2, 1, 0, -1, -1, 0, 2, 2, 1, 2, 0, 1, 0, 1, 1, 0, 1, 0, 3, 2, 0, 0, 0, 1, 1, 1, 2, 2, 2, 1, 1, 0, 2, 3, 2, 1, 1, 1, 2, 1, 1, 2, 1, 1, 2, 1, 1, 0, 0, -1, 0, 0, 0, 3, 2, 1, 2, 2, 2, 3, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 2, 2, -1, -1, -1, 0, -1, 0, 1, 1, 2, 2, 0, 2, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 0, 0, -1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 1, 2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 1, 0, 3, 2, 2, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 1, 1, 1, 2, 2, 2, 2, 0, 1, -1, 0, 0, 1, 0, 0, 0, 0, -1, -2, -2, -1, -2, -1, 0, 0, 0, 1, 1, 2, 1, 2, 2, 3, 1, 1, -2, -3, -2, -1, 0, 0, 0, 0, -2, -1, 0, -2, -1, -1, 1, 1, 2, 2, 1, 2, 3, 3, 4, 2, 0, 0, -2, -4, -4, -1, -2, -1, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -2, -1, -2, -3, -1, -2, -2, -1, -1, -2, -1, 0, -2, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -2, -2, -3, -2, -1, -2, -2, -1, -2, -3, -2, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -3, -1, 0, -2, -3, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, -2, -1, -2, -1, -1, -2, -2, -1, 0, -2, -1, -1, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, -1, -2, -2, -2, -1, -2, -2, -3, -3, -3, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -2, -1, -1, -1, -2, -1, -1, -3, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -2, -1, -2, -2, -2, -2, -1, -1, 0, -2, -1, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, 0, -1, -3, -1, -2, -2, -2, -1, -1, -2, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, -2, -2, -2, 0, -3, -1, -1, -1, 0, -1, -2, -2, -1, -1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -2, -2, 0, -1, -1, -1, -2, -2, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, 0, -1, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -2, -2, -1, 0, -1, 0, 0, -1, -1, 1, 0, 1, 1, 0, 0, 0, 2, 0, 0, 1, 0, 0, -1, -1, -2, -1, 0, 0, 0, -3, -3, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -2, 0, 0, -1, -1, -1, -2, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 2, 0, 1, 1, 0, 0, -1, -1, -1, 0, 0, -2, 0, -2, -3, -1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 1, 0, -1, -1, -1, -1, -1, -3, -3, -1, -1, -1, -3, -2, -1, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -2, -1, -3, -4, -3, -2, -1, -2, -2, -2, -2, -2, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -2, -3, -2, -2, -3, -1, -1, -1, -3, -2, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, -3, -3, -2, -3, -3, -2, -3, -2, -3, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -3, -3, -3, -3, -4, -4, -2, -2, -3, -2, -3, -1, -2, 0, 0, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -3, -4, -4, -2, -2, -2, -3, -1, -2, 0, -2, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, -3, -3, -3, -2, -2, -3, -2, -4, -3, -1, -2, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -2, -3, -2, -2, -3, -4, -2, -1, -2, -3, -4, -2, -2, -3, -1, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -3, -2, -1, -3, -3, -2, -2, -3, -3, -2, -1, -2, -2, -1, -1, -2, -2, -2, -1, -1, 0, 0, 0, -2, -2, -2, -2, -3, -2, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -2, -1, -1, -1, 0, -1, -1, 0, 0, 0, 2, 2, 1, 1, 1, 0, 0, 0, -2, -2, 0, -1, 0, -1, 0, -1, -2, -1, -1, -1, -3, -1, 0, 0, 1, 1, 2, 2, 1, 0, 0, 1, -1, -1, 0, -2, -1, 0, -1, 0, 1, 1, 0, 0, 0, -2, -1, -1, -1, 0, -1, 0, 1, 2, 2, 1, 1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, 0, -2, -1, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 1, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 0, 3, 0, 0, 0, 1, 0, 2, 2, 1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 2, 0, 0, 1, 1, 0, 1, 2, 1, 1, 2, 2, 1, 2, 0, 0, 0, 0, -1, 0, 0, 1, 2, 1, 1, 0, 2, 0, 0, 2, 0, 0, 2, 2, 2, 1, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, 2, 0, 1, 0, 1, 2, 0, 1, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 1, 2, 1, 0, 0, 0, 1, 0, 2, 3, 1, 2, 1, 1, 1, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 2, 3, 2, 3, 2, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 1, 0, 0, 2, 0, 0, 2, 1, 0, 3, 3, 2, 1, 0, 1, 1, 2, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 1, 3, 2, 3, 2, 1, 0, 1, 3, 3, 0, 1, 0, 0, 1, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 2, 1, 3, 2, 1, 1, 1, 2, 2, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, 2, 2, 1, 0, 0, 0, 1, 1, 2, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 2, 1, 1, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 1, 1, -1, 0, -1, 0, 0, 2, 0, 3, 3, 3, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 1, 1, 1, 2, 3, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, -3, -2, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 1, 1, 0, -2, -1, 0, 0, 0, 0, 0, 0, -3, -2, -1, -2, 0, 0, 1, 1, 1, 1, 3, 2, 2, 2, 1, 0, 0, 0, -2, 0, 0, -1, 0, 0, 0, -2, -3, -1, -2, -1, -2, 0, 0, 1, 0, 2, 2, 3, 3, 2, 1, 1, 0, -2, -3, -3, 0, -2, 0, -1, -2, 0, -2, 0, -2, 0, 0, 0, 0, 0, 0, 2, 1, 2, 2, 1, 0, 0, 0, -1, -3, 0, -1, 0, 0, 0, 0, -2, -1, 0, -1, -1, -1, -1, 0, 0, 2, 1, 2, 2, 3, 2, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, -2, 0, -2, -1, 0, 0, 0, 1, 1, 2, 3, 2, 1, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, -1, 1, 0, 3, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -2, -2, 0, 0, -1, 0, 0, 1, 1, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -2, 0, 0, 0, -1, 0, -1, 0, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, -1, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 1, 2, 0, 0, 1, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 2, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 0, 0, 0, 1, 0, 1, 0, 1, 1, 2, 2, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 1, 2, 2, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 0, 1, 0, 1, 1, 0, 1, 1, 2, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 2, 2, 0, 1, 1, 0, 0, 0, 2, 0, 2, 1, 0, 1, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 1, 1, 1, 2, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 1, 2, 2, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 2, 2, 1, 1, 0, 1, 1, 0, 1, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 1, 2, 1, 1, 0, 1, 0, 2, 1, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 2, 2, 0, 0, 0, -1, 0, 0, 1, 2, 2, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 3, 3, 2, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 0, 2, 3, 3, 1, 3, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -2, -1, -2, 0, 1, 0, 1, 1, 1, 3, 1, 3, 2, 1, 1, 1, -1, 1, 0, 0, 0, -1, -1, 0, -2, -1, -1, -1, -1, 1, 0, 1, 1, 2, 3, 2, 4, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -2, 0, -1, 0, 0, 1, 2, 1, 2, 2, 2, 1, 1, 1, 0, 0, -2, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 2, 2, 1, 2, 4, 2, 1, 2, 1, 0, 0, -2, 2, 2, 2, 1, 1, 0, -1, -3, -2, -1, -1, 0, 1, 2, 3, 4, 4, 5, 4, 3, 3, 1, 0, -1, -2, -4, 1, 0, 1, 0, 0, -1, -2, -4, -4, -3, -2, -1, -1, 1, 2, 3, 5, 3, 4, 5, 2, 0, 0, -1, 0, 0, 3, 1, 0, 0, 0, -1, -1, -3, -2, -3, 0, -2, -1, 0, 2, 2, 2, 3, 2, 2, 2, 1, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, -1, -1, -1, -1, 0, -2, 0, -1, 1, 2, 2, 3, 2, 1, 1, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 2, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, -1, -1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 2, 0, 1, 0, 0, 1, 0, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, 3, 2, 1, 0, 0, 0, 0, 2, 1, 1, 1, 1, 2, 1, 1, 1, 1, 0, 0, 0, 1, 0, 1, 2, 2, 3, 1, 2, 1, 1, 0, 1, 0, 2, 2, 3, 1, 3, 0, 2, 1, 1, 2, 2, 2, 2, 2, 1, 0, 2, 0, 1, 0, 1, 1, 0, 1, 1, 1, 1, 2, 2, 3, 4, 1, 0, 0, 1, 1, 3, 3, 2, 3, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 4, 3, 4, 2, 0, 2, 1, 2, 4, 5, 4, 4, 3, 3, 2, 1, 0, -1, -1, -1, 0, 0, 0, 0, 2, 2, 3, 4, 4, 2, 1, 2, 1, 4, 4, 6, 6, 4, 3, 3, 1, 0, -1, 0, -1, -2, -2, -2, -1, 1, 1, 4, 6, 5, 6, 3, 2, 1, 1, 2, 3, 6, 4, 3, 3, 1, 0, -1, 0, 0, -2, -2, -2, -2, 0, 0, 2, 4, 5, 6, 4, 2, 2, 1, 3, 2, 4, 2, 4, 3, 2, 1, 0, 0, 0, -1, -3, -1, -2, -3, 0, 0, 2, 4, 4, 6, 5, 2, 0, 2, 1, 3, 3, 2, 2, 1, 0, -1, 0, 0, 0, -1, -2, -1, -1, -1, 0, 0, 1, 2, 3, 4, 4, 1, 0, 0, 0, 2, 1, 2, 1, 0, 0, 0, 0, 1, 1, 0, -2, 0, 0, 0, 1, 0, 3, 2, 4, 4, 5, 0, 0, 1, 0, 2, 1, 2, 0, 1, -1, 1, 0, 1, 1, 1, 1, 1, 0, 1, 2, 2, 1, 3, 1, 4, 3, 0, 0, 0, -1, 1, 1, 2, 1, 0, 0, 1, 1, 1, 3, 3, 2, 0, 1, 3, 3, 3, 0, 0, 2, 4, 2, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 2, 3, 3, 1, 1, 1, 3, 2, 2, 0, 2, 1, 1, 3, 0, 0, -1, 0, -1, 1, 1, 0, 1, 1, 0, 1, 1, 2, 2, 2, 0, 0, 2, 3, 3, 0, 1, 1, 2, 2, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 2, 0, 1, 1, 3, 3, 3, 1, 1, 2, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, -2, -2, 0, 1, 2, 2, 1, 1, 3, 3, 3, 4, 2, 1, 1, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, -2, -2, -2, 0, 1, 0, 2, 2, 4, 5, 3, 3, 5, 3, 1, 0, 0, -1, 2, 0, 1, 0, 0, -1, 0, -1, -2, -3, -2, -1, 1, 1, 2, 0, 4, 6, 4, 3, 3, 1, 1, 0, 0, -2, 2, 0, 0, 0, 0, 0, 0, -1, -3, -1, -2, 0, -1, 1, 1, 1, 3, 6, 5, 5, 4, 2, 0, -1, -2, -4, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 4, 5, 4, 2, 0, 0, -1, -1, -5, -6, 0, -1, -1, 0, -1, -1, -2, -1, -1, 0, 0, 0, 1, 1, 2, 5, 3, 4, 4, 4, 3, 1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, -2, -1, -2, 0, 0, 0, 1, 2, 1, 3, 3, 4, 4, 3, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, -2, -1, -1, 0, 0, 1, 1, 1, 3, 3, 3, 2, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 3, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 2, 1, 2, 1, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 0, -1, 0, 0, 0, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 1, 1, 1, 2, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 1, 2, 1, 2, 2, 2, 0, 0, 0, 1, 1, 0, 2, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 1, 1, 3, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 2, 0, 1, 1, 3, 0, 0, 1, 2, 2, 2, 2, 0, 1, 0, 0, 0, 0, 0, -1, -2, -2, -1, 0, 0, 2, 0, 0, 0, 1, 4, 1, 1, 3, 3, 2, 3, 1, 1, 2, 0, 0, 0, -1, -2, -3, -2, -3, 0, 0, 0, 0, 0, 1, 1, 4, 5, 1, 2, 1, 1, 2, 1, 2, 1, 0, 1, 1, 0, 0, -3, -2, -3, -3, -3, -2, 0, 0, 1, 1, 2, 4, 6, 1, 2, 2, 0, 1, 1, 1, 0, 0, 0, -1, -1, -1, -3, -3, -3, -4, -4, -2, 0, 0, 2, 1, 2, 5, 5, 1, 0, 1, 2, 0, 1, 1, 0, 1, 0, 0, -1, -2, -4, -2, -2, -4, -2, -1, -2, -1, 0, 1, 3, 3, 3, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -3, -2, -2, -3, -3, -1, -1, 0, 1, 0, 1, 4, 5, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, -1, 0, -1, -2, -2, -3, -3, -1, -2, -1, 1, 1, 1, 2, 3, 3, -1, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, -1, 0, -1, -1, -1, -1, -1, 0, 0, 1, 1, 0, 0, 2, 3, 0, 0, 1, 0, 0, 1, 2, 2, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 2, 0, 1, 0, 0, 3, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 2, 2, -1, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, -1, -2, -1, -1, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -1, 0, -1, -1, -1, -1, 0, -2, 0, 0, 0, 1, 1, 1, 0, 1, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -1, -2, -2, -1, 0, 0, 1, 2, 1, 2, 3, 1, 1, 1, 0, 2, -1, 0, 0, 0, -1, 0, -2, -1, -1, 0, -1, -1, 0, 0, 1, 1, 2, 2, 3, 3, 3, 3, 2, 1, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 2, 0, 2, 3, 3, 3, 4, 3, 2, 1, 1, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 3, 2, 4, 4, 4, 5, 3, 3, 3, 1, -1, -1, 0, 4, 3, 1, 1, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 2, 3, 2, 2, 1, 3, 1, 0, 1, 0, -1, -1, 3, 2, 2, 1, 0, -1, 0, -2, -3, -2, -1, -2, -1, 0, 0, 2, 1, 2, 4, 3, 2, 1, 0, 0, 0, 0, 4, 3, 2, 1, 0, -1, -1, -1, -3, -3, -3, -2, -1, 0, 0, 1, 2, 3, 1, 3, 1, 2, 0, 1, 0, 1, 3, 3, 1, 1, 1, 0, 0, 0, -1, 0, -1, -2, -2, 0, 0, 1, 1, 1, 2, 2, 3, 1, 1, 1, 0, 0, 3, 3, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, -2, -1, -1, 1, 0, 0, 2, 2, 1, 0, 1, 0, 1, 1, 2, 1, 2, 1, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 2, 0, 1, 1, 0, 0, 1, 2, 1, 1, 2, 1, 0, 1, 1, 1, 0, 1, 1, 0, -1, 0, 0, 0, 1, 1, 2, 2, 1, 2, 1, 1, 1, 1, 1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 4, 1, 0, 0, 0, 0, 1, 0, 2, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 3, 4, 4, 0, 0, 0, 0, 1, 2, 3, 3, 1, 2, 2, 2, 0, -1, -1, -2, 0, 0, 0, -1, 1, 1, 3, 2, 4, 4, 0, 0, 0, 0, 1, 2, 4, 3, 4, 4, 2, 0, 0, -2, -3, -2, -1, 0, 0, 0, 1, 1, 3, 3, 4, 6, 2, 0, 1, 1, 2, 3, 3, 5, 4, 4, 3, 1, -2, -2, -2, -2, -3, 0, 0, 0, 0, 1, 4, 5, 4, 5, 1, 1, 2, 2, 1, 4, 4, 5, 4, 4, 2, 0, 0, -1, -3, -4, -3, -2, -1, 0, 0, 0, 2, 5, 5, 5, 1, 0, 2, 0, 2, 3, 4, 4, 4, 2, 0, 0, -2, -4, -3, -3, -4, -4, -1, 0, 1, 2, 2, 5, 5, 5, 2, 2, 1, 2, 1, 1, 3, 2, 2, 0, 0, -1, -3, -3, -4, -3, -3, -2, -1, 0, 0, 0, 2, 4, 5, 5, 3, 0, 0, 1, 2, 2, 2, 2, 0, 0, 0, 0, -1, -3, -3, -3, -1, 0, 0, 0, 1, 2, 2, 4, 3, 4, 1, 1, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 2, 2, 3, 3, 3, 1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 3, 3, 2, 2, 2, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 1, 1, 1, 2, 2, 2, 2, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 1, 2, 0, 2, 2, 2, 0, 0, 0, 1, 1, 0, 2, 0, 0, -1, -1, 0, 0, 1, 0, 1, 2, 1, 1, 2, 1, 2, 0, 1, 1, 2, 1, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 2, 3, 2, 1, 2, 1, 1, 2, 2, 1, 1, 1, 1, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 2, 0, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, -2, 0, 0, -1, 0, 1, 3, 3, 2, 2, 1, 1, 1, 1, 0, 3, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -2, -1, 0, -1, -1, 0, 3, 3, 2, 2, 1, 2, 1, 0, -1, 1, 0, 0, 1, 0, 1, 1, 0, -1, -1, -1, -2, -2, -1, -1, 0, 1, 1, 2, 2, 1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 2, 1, 2, 4, 3, 4, 4, 3, 2, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, -1, 0, -1, 0, 0, 2, 2, 1, 1, 2, 3, 1, 2, 0, -1, -1, 0, -2, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 1, 1, 1, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 2, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 2, 1, 0, 2, 1, 2, 2, 1, 1, 2, 1, 1, 0, 1, 1, 0, -1, -1, -2, 0, 0, 0, 0, 2, 0, 1, 1, 1, 0, 1, 2, 2, 3, 3, 1, 2, 1, 1, 0, 0, 1, 0, 0, -2, -1, -2, -1, 0, 0, 1, 1, 1, 0, 2, 1, 1, 1, 1, 2, 0, 1, 2, 1, 0, 0, 0, 0, 0, -2, -2, -3, -1, -2, 0, 0, 0, 0, 1, 0, 2, 1, 2, 2, 1, 2, 1, 1, 2, 0, 0, 0, 0, -1, -1, -2, -2, -2, -2, 0, -1, 0, 1, 2, 0, 1, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, -1, -1, -2, -1, -2, -1, -3, -1, -1, 0, 0, 0, 1, 2, 3, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 2, 0, 2, 0, 1, 2, 0, 2, 0, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 1, 0, 1, 1, 1, 1, 2, 1, 2, 2, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 2, 2, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 2, 0, 1, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 1, 1, 0, 0, 1, -1, 1, 0, 1, 0, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 2, 1, 2, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 2, 3, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, -2, 0, -2, -1, -1, 1, 0, 0, 0, 2, 2, 3, 3, 3, 2, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, -2, 0, 0, 0, 0, 1, 1, 2, 3, 3, 3, 2, 3, 1, 1, -1, -3, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 3, 3, 2, 3, 4, 3, 3, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 2, 1, 3, 3, 4, 4, 2, 3, 3, 2, 0, -1, -2, -2, -1, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, 1, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, -1, 0, 0, 1, -1, 1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, -1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, -1, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 1, 1, 1, 0, 0, 1, 1, 1, 1, 2, 2, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 0, 1, 0, 2, 1, 2, 2, 2, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 1, 0, 1, 1, 0, 2, 2, 2, 1, 2, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 2, 0, 0, 2, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 2, 2, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 1, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 1, 1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, -1, -1, -1, 0, -1, 0, 0, 1, 0, 1, 1, 2, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 1, 2, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 0, 2, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 2, 2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 2, 1, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 2, 0, 1, 3, 2, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 2, 1, 1, 3, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 2, 0, 1, 1, 1, 0, 0, 2, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 2, 0, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 1, 2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, -2, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -1, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -2, 0, -2, 0, -1, -1, 0, -1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -2, 0, -2, 0, -1, 0, 0, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -2, 0, -1, -1, -1, -1, 1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -2, -2, -1, -2, 0, -1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, -1, 0, 1, 1, 0, 1, -1, 0, -1, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, -2, -1, 0, -2, -1, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -2, -2, -2, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 2, 1, 1, 2, 1, 1, 2, 0, 0, -5, -7, -5, -6, -3, -3, 0, -1, -1, 0, -1, 0, -2, -3, -1, -1, 1, 2, 0, 0, 1, 2, 2, 1, 1, -1, -3, -4, -3, -3, -1, -1, 0, -1, 0, -1, 0, 0, -3, -3, -2, -2, -1, 0, 0, 0, -1, 0, 3, 0, 0, 0, -1, -2, -2, -1, 0, 0, 1, -1, -1, 0, 0, 0, -2, -3, -2, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, -1, -3, -2, -2, -1, -3, -3, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -3, -2, -2, -1, -2, -2, -3, -2, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, -3, -2, -1, 0, 0, -1, -1, 0, 0, 3, 2, 0, 0, -1, -1, 0, 1, 0, -3, -2, -1, 0, -2, -1, 0, 0, -2, -2, -2, -2, 0, 0, 0, 0, 1, 3, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, -1, 0, -2, -1, -3, -3, -4, -3, -1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -4, -2, -3, -2, 0, -1, 0, 0, 0, 0, -1, -3, 0, 1, 3, 3, 0, -1, -1, -1, -1, 0, -1, 0, -1, -3, -3, -2, -2, 0, 0, 0, 0, 0, 0, 1, -1, -1, 1, 1, 0, 0, 0, -1, -1, -3, -1, 0, -1, -2, -1, -4, -2, -2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, -2, -3, -3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 2, 1, 2, 0, 0, -1, -1, 0, -3, -3, -4, -6, -3, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 1, 1, 2, 1, 0, 0, -1, 0, -1, -1, -3, -2, -4, -3, -4, -1, 0, 0, -2, -1, -1, -1, -2, 0, 0, 1, 0, 2, 0, 0, -2, -2, -1, -2, -3, -3, -2, -3, -2, -4, -1, -1, -2, -2, -2, 0, -1, -2, -1, -1, 1, 0, 0, -1, 0, -1, -2, -2, -3, -2, -4, -3, -4, -3, -2, -2, -1, -3, -2, 0, -1, 0, 0, -1, 0, -1, 0, -2, -2, 0, 0, -1, -3, -3, -2, -3, -4, -2, -2, -3, -3, -1, -2, -3, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -2, -4, -2, -3, -3, -2, -1, -1, -3, -1, -1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, -3, -3, -3, -4, -4, -2, -4, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 1, 3, 2, 2, 1, 1, -1, -2, -2, -2, -4, -3, -3, -4, -3, -4, -2, 0, -3, 0, 0, 0, 0, 0, 1, 2, 2, 4, 3, 4, 2, 0, 0, -2, -1, -3, -3, -4, -5, -3, -3, -3, -3, -2, -1, 0, 0, 0, 2, 0, 1, 4, 5, 5, 3, 1, 0, 0, 0, -2, -1, -4, -6, -3, -5, -4, -4, -4, -3, -2, -3, -1, 0, 0, 1, 1, 1, 3, 3, 3, 3, 2, 1, 0, -1, -2, -1, -4, -5, -5, -6, -7, -6, -6, -4, 0, -1, -2, 0, 1, 2, 2, 1, 2, 4, 3, 3, 3, 0, -1, -2, 0, -3, -3, -4, -6, -5, -7, -7, -5, -3, -1, -2, -1, 1, 1, 0, 1, 0, 2, 2, 1, 3, 1, 0, -2, -2, -1, -3, -5, -6, -5, -6, -6, -4, -2, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, -2, -2, -2, -5, -4, -5, -4, -5, -4, -3, -1, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, -1, 0, -1, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 1, -1, -2, -2, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, -1, 1, 0, 2, 4, 4, 2, 3, 3, 2, 0, -1, -1, -3, -2, 0, 0, 0, -2, -1, -3, -1, -1, -2, -2, -1, 0, -1, 1, 1, 2, 2, 3, 3, 0, 0, 0, -1, -2, -2, -1, 0, 0, -1, -1, -2, -1, 0, -1, -3, -3, -3, -1, 0, 0, 0, 2, 1, 2, 2, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -2, -3, -2, -2, -2, 0, 0, 0, 1, 1, 2, 3, 0, 1, 0, -1, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, -2, 0, 0, 2, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 1, 2, 1, 0, 0, 0, 2, 0, -1, 0, -1, 0, 0, 0, 0, 1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 2, 0, 1, 1, 0, 2, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 2, 1, 1, 0, 1, 2, 0, 0, 2, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 1, 3, 2, 1, 2, 1, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 2, 2, 2, 3, 3, 3, 3, 2, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 3, 2, 2, 2, 2, 1, 1, 0, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 2, 1, 2, 2, 2, 2, 3, 2, 3, 2, 0, 1, 0, -2, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 3, 3, 3, 3, 1, 2, 2, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 0, 2, 1, 1, 2, 3, 2, 1, 0, 2, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 2, 1, 3, 3, 2, 2, 1, 0, 1, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 2, 4, 3, 0, 1, 1, 0, 2, 2, 0, 2, 0, 1, 1, 2, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 3, 1, 1, 2, 1, 0, 0, 2, 1, 3, 2, 2, 2, 2, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, 0, 1, 2, 3, 2, 2, 1, 2, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 3, 2, 2, 2, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 2, 4, 4, 4, 2, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -3, -2, 0, 0, 0, 1, 2, 3, 4, 3, 4, 3, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -2, -2, -2, -2, -2, 0, 0, 0, 0, 3, 3, 4, 4, 3, 4, 1, 1, 0, -1, 0, -1, 0, -1, -2, -2, 0, -2, -2, -2, -1, 0, 1, 1, 0, 1, 2, 3, 3, 4, 4, 2, 0, 0, -1, -2, -2, -1, -1, 0, 0, -2, -3, -2, -2, -2, -1, -1, 0, 0, 2, 3, 4, 3, 4, 4, 2, 2, 0, 0, -3, -1, 0, -1, 0, 0, -1, -1, -1, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -2, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -4, -3, -2, -2, -4, -3, -3, -2, -1, -2, -1, 0, 0, 1, 2, 1, 3, 3, 5, 6, 3, 4, 3, 1, 3, 3, -3, -3, -3, -1, -1, -2, 0, -1, -2, -2, 0, -1, 0, 1, 0, 1, 3, 4, 6, 5, 3, 3, 2, 1, 2, 1, -3, 0, 0, 0, -1, 0, 0, -1, -1, -3, -1, 0, 0, -1, 0, 1, 1, 4, 5, 4, 4, 3, 1, 1, 0, 1, -3, -1, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, 0, 0, -2, -1, 1, 1, 3, 3, 3, 2, 1, 2, 2, 2, -4, -2, 0, 0, 0, 2, 0, 0, 0, -2, 0, 0, -1, -1, -1, 0, 0, 0, 2, 1, 4, 2, 2, 3, 1, 3, -3, -1, 0, 0, 1, 1, 1, 0, 1, 0, -1, 0, 0, -1, -1, -2, -1, 0, 2, 2, 3, 2, 3, 4, 2, 0, -1, 0, 1, 0, 0, 2, 2, 0, -1, 0, -1, 0, 0, -2, -2, -4, -3, 0, 0, 1, 2, 1, 2, 3, 2, 0, 0, 1, 1, 0, 3, 2, 2, 0, -1, 0, -1, -3, -3, -3, -4, -2, -3, 0, 1, 1, 1, 2, 1, 1, 1, 0, 0, 1, 1, 3, 2, 1, 1, 0, 0, -3, -2, -3, -3, -3, -3, -4, -3, -2, 0, 2, 2, 1, 1, 1, 0, 2, 0, 3, 2, 3, 1, 2, 1, 0, -1, -2, -2, -2, -4, -2, -5, -4, -3, -2, 0, 0, 0, 2, 1, 1, 2, 3, 2, 1, 3, 1, 1, 1, 1, -1, -2, 0, -1, -2, -3, -5, -4, -5, -3, -1, 0, 0, 1, 1, 2, 0, 2, 3, 1, 2, 2, 0, 1, 1, 1, -1, 0, 0, -3, -4, -5, -5, -5, -6, -5, -4, 0, 0, 0, 2, 0, 0, 1, 2, 1, 2, 1, 1, 0, 1, 0, -1, 0, -1, -1, -3, -4, -5, -5, -5, -6, -4, -2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -3, -3, -4, -5, -6, -6, -4, -2, -1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -3, -3, -3, -5, -5, -3, -2, 0, -1, 0, 0, 1, 1, 1, 0, -1, 1, 0, 0, 0, 0, 1, 1, 2, 1, -1, -1, -2, -4, -4, -3, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 1, 0, 0, -3, -2, -2, -3, -4, -2, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, -2, -4, -3, -2, -2, 0, 1, 2, 2, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 2, 2, 0, -3, -3, -3, -3, -1, -1, 2, 0, 2, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -2, -1, -4, -3, -2, -1, 0, 2, 1, 2, 3, 1, 0, 1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -2, -2, -2, -2, -3, 0, 0, 2, 3, 3, 2, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, -2, -1, -1, -1, -1, 2, 3, 2, 2, 3, 3, 2, 1, 0, 2, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -2, 0, -1, 0, 0, 1, 1, 2, 5, 4, 3, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -2, -1, -1, 0, -1, -1, 0, 1, 2, 3, 3, 4, 4, 4, 3, 4, 2, 0, 0, -2, -1, -1, -2, -1, 0, -2, -1, -1, 0, 0, 0, 0, 2, 2, 2, 4, 5, 5, 5, 5, 4, 2, 0, 0, 0, -4, -4, -3, -2, 0, 0, 0, 0, -1, 0, 0, 1, 2, 3, 3, 3, 5, 5, 5, 4, 5, 3, 3, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, -1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 1, 1, 0, 1, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -8, -7, -7, -8, -7, -7, -6, -6, -6, -7, -7, -7, -8, -9, -6, -3, -1, -2, -1, -1, -1, -1, 0, 1, 0, -1, -7, -7, -8, -7, -6, -8, -6, -6, -5, -5, -4, -4, -7, -7, -4, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, -6, -5, -6, -5, -6, -5, -6, -5, -5, -3, -3, -3, -5, -6, -2, -2, 0, -2, -1, -1, 0, -1, -1, -1, -2, -2, -6, -6, -5, -5, -6, -6, -5, -5, -3, -4, -4, -3, -3, -4, -2, -2, -1, 0, 0, -2, 0, 0, 0, 0, -2, -1, -6, -6, -3, -3, -4, -6, -6, -4, -3, -2, -2, -3, -3, -3, -2, -2, 0, 0, 0, -1, 0, 1, 0, 0, -2, 0, -7, -6, -3, -5, -4, -7, -6, -5, -2, -2, -3, -2, -3, -3, -1, 0, 0, 1, 0, 0, 0, 1, 1, 0, -1, -1, -4, -4, -5, -4, -6, -6, -5, -3, -3, -1, -3, -2, 0, -1, 0, 0, 2, 2, 1, 0, 1, 0, 0, 0, -1, 0, -6, -5, -5, -4, -5, -4, -3, -2, -2, -2, -1, -2, 0, 0, 0, 2, 2, 1, 2, 2, 0, -1, 0, 0, 0, -1, -6, -5, -5, -4, -4, -4, -3, -1, -1, 0, 0, 1, 1, 0, 2, 1, 2, 3, 1, 1, 1, 0, 0, 0, 0, -1, -4, -4, -4, -4, -3, -4, -3, 0, 0, 0, 2, 1, 1, 1, 3, 2, 2, 4, 2, 1, 0, -1, -1, 0, 0, 0, -6, -4, -4, -5, -4, -4, -1, 0, 1, 1, 2, 2, 2, 3, 4, 2, 2, 6, 4, 2, 0, 0, 0, 0, 0, 0, -5, -5, -3, -4, -4, -4, -1, 1, 1, 1, 2, 4, 4, 5, 3, 3, 4, 5, 4, 3, 1, 0, -2, 0, 0, 0, -5, -4, -5, -3, -4, -1, -1, 0, 1, 2, 3, 4, 4, 5, 4, 3, 4, 6, 5, 3, 0, 0, -2, 0, 0, 0, -4, -6, -5, -5, -3, -2, 0, 1, 1, 2, 3, 5, 5, 6, 3, 4, 6, 5, 5, 3, 1, 0, 0, 0, 0, 1, -4, -4, -5, -2, -2, -2, -1, 0, 2, 3, 4, 5, 6, 4, 5, 4, 5, 6, 4, 2, 3, 0, 0, 0, 0, 0, -4, -3, -3, -3, -3, -2, -1, -1, 0, 1, 2, 4, 6, 4, 4, 5, 6, 6, 4, 2, 2, 0, -1, -1, 0, -1, -6, -3, -3, -2, -3, -3, -3, 0, 0, 1, 2, 3, 4, 4, 4, 3, 3, 3, 2, 1, 1, 0, -1, -2, 0, 0, -5, -5, -3, -3, -2, -1, -3, 0, 0, 0, 2, 4, 2, 4, 4, 4, 2, 3, 1, 1, 0, 0, 0, 0, -1, 0, -5, -4, -2, -2, -2, -2, -2, -1, 0, 0, 0, 0, 1, 2, 1, 2, 2, 3, 1, 1, 1, 0, -1, -1, 0, 0, -5, -3, -2, -4, -2, -3, -1, 0, 0, 0, -1, -1, -1, 1, 0, 2, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -4, -5, -5, -3, -4, -4, -4, -1, -1, -1, -1, -1, -1, 0, 0, 3, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -5, -5, -3, -5, -5, -4, -4, -2, -3, -2, -3, -2, -2, -1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 1, 0, -1, -5, -4, -4, -5, -5, -5, -4, -5, -4, -2, -2, -2, -2, -3, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, -4, -6, -5, -6, -6, -6, -4, -5, -4, -3, -3, -3, -3, -1, -2, -1, -2, -2, -1, 0, 0, -1, 0, 0, 0, -1, -5, -4, -6, -6, -7, -5, -6, -6, -5, -5, -3, -3, -5, -2, -2, -2, -2, -1, -2, 0, 0, -1, 0, 1, 0, 0, -6, -6, -7, -8, -7, -6, -7, -7, -6, -8, -7, -7, -5, -5, -2, -2, -2, -1, -2, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, -1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, -2, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 2, 1, 0, -1, 0, -1, -1, 0, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 1, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, -1, 0, -1, -1, 1, 0, 0, 0, 0, -1, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, -2, -1, -3, -2, -3, -4, -2, -4, -2, -3, -2, -4, -3, -4, -2, -2, -1, 0, 1, 0, 0, -2, 0, -2, -3, -1, -2, -2, -2, -3, -2, -4, -4, -2, -2, -3, -2, -2, -2, -3, -2, -1, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -1, -2, -1, -3, -2, -3, -3, -4, -3, -2, -2, -2, -4, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, -2, -1, -3, -1, -2, -3, -3, -1, -1, -1, -3, -2, -4, -3, -1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -3, -2, -1, 0, -2, -2, -2, -1, 0, 0, -1, -3, -2, -2, -2, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -2, -1, -1, -1, -1, -1, -2, -2, 0, 0, -1, -1, -1, -3, -3, -3, -2, 0, 1, 1, 0, 0, 0, 1, -1, 0, -1, -1, -1, -2, -2, -1, -2, -1, -2, 0, -1, -1, 0, 0, -1, 0, -1, 0, 1, 0, 0, 1, 0, 0, 1, 0, -2, -1, -2, -2, -1, -2, -2, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -2, -1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 1, 1, 2, 1, 2, 0, 1, 0, 2, 1, 1, 1, 0, 1, 1, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 1, 2, 3, 2, 2, 0, 2, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 1, 0, 3, 3, 2, 2, 1, 3, 1, 1, 0, 0, 1, 3, 2, 1, -1, -1, 0, 0, 1, -2, -1, 0, 0, 0, 0, 3, 2, 4, 2, 2, 2, 1, 2, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, 1, 2, 0, 3, 1, 3, 3, 2, 2, 1, 0, 0, 0, 2, 1, 1, 0, -1, -1, 0, 1, 0, -1, -1, -1, 0, 1, 1, 2, 3, 3, 3, 4, 4, 1, 1, 1, 1, 2, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, -2, -1, 0, -1, 0, 2, 2, 2, 3, 3, 2, 3, 2, 0, 1, 1, 2, 3, 3, 0, 0, 0, 0, 0, 1, -2, 0, 0, 0, 0, 1, 1, 2, 2, 2, 1, 1, 2, 2, 1, 1, 2, 1, 2, 1, 2, 0, 0, 0, 0, 0, -2, -2, -1, 0, 0, 0, 2, 1, 1, 1, 1, 1, 0, 1, 0, 3, 3, 2, 3, 2, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 2, 1, 3, 1, 1, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 3, 2, 1, 1, 2, 0, 0, -1, -1, 0, -1, -2, -2, -2, -2, 0, -1, 0, 0, 0, -1, 0, -1, -2, 0, 1, 1, 2, 2, 2, 3, 1, 0, 0, -1, 0, -1, 0, -2, -1, -1, -2, 0, -1, -1, -1, -1, -2, -2, -3, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, 0, -1, -1, -2, -1, -2, -2, -3, -1, -1, -2, -2, 0, -3, -3, -3, -1, 0, 0, 0, 0, 2, 2, 0, 1, 0, 0, -1, 0, -3, -2, -2, -2, -2, -3, -1, -2, -3, -3, -4, -2, -2, -1, 0, 0, -1, 0, 1, 2, 2, 0, 0, 0, 0, -2, -1, -2, -2, -2, -2, -3, -4, -4, -3, -5, -3, -2, -3, -2, -2, -1, 0, 1, 0, 1, 0, 0, -1, 0, 0, -1, -1, -1, -2, -3, -4, -3, -4, -4, -5, -5, -4, -5, -4, -3, -2, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -3, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, -1, 0, -1, 0, 0, 0, -1, 1, 1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, -4, -2, -2, -2, -2, 0, 0, 0, 1, 1, 1, 4, 4, 4, 3, 4, 6, 5, 7, 6, 3, 0, -1, -2, -1, 0, -3, -2, 0, -2, -1, 0, -1, 0, 0, 0, 1, 1, 2, 4, 2, 3, 3, 6, 5, 4, 1, 1, -2, 0, -1, 0, -2, 0, -1, 0, 0, 0, -1, 0, -1, -2, 0, 1, 0, 1, 0, 1, 3, 4, 4, 3, 1, 1, 0, -2, 0, -2, -3, -2, -1, 0, 1, 1, 0, 0, -1, -2, -1, 0, 0, 1, 0, 0, 1, 3, 3, 3, 1, 1, 0, -1, 0, -1, -3, -2, 0, 0, 0, 0, 1, 2, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -1, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, -3, -3, -3, 0, 0, 0, 1, 1, 2, 1, 0, -2, -1, 0, 0, 1, 0, 1, 2, 1, 1, 0, 0, 0, 1, 0, -2, -3, -3, -3, 0, 0, 0, 1, 2, 0, -1, 0, -2, -1, 0, 2, 1, 3, 2, 2, 0, 0, -1, 0, 0, 0, 0, -2, -3, -2, 0, -1, -1, 1, 0, 1, 0, 0, 0, 0, 2, 2, 3, 2, 3, 0, -1, -1, -1, 0, 1, -1, -1, -2, -3, -2, -1, 0, 0, 0, 1, 0, -1, 0, 0, 1, 4, 3, 2, 3, 2, 0, -2, -3, -2, 0, 0, -2, -2, -3, -4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 4, 4, 2, 1, 1, 0, -1, -2, 0, 0, -2, -3, -4, -5, -3, -2, 0, 0, 0, 0, -1, 0, 0, 1, 2, 1, 2, 2, 3, 1, 1, 0, -1, -3, -1, 0, -1, -3, -3, -3, -4, -3, 0, 0, 0, 1, 0, -1, 0, 1, 0, 2, 1, 2, 1, 0, 1, 0, -1, -1, -1, -2, -2, -3, -3, -5, -5, -4, -1, -1, 1, 0, 0, 0, 0, 0, 0, 2, 3, 3, 1, 0, 0, 0, -1, 0, 0, -1, -2, -5, -4, -3, -3, -5, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 1, 0, -1, 0, 0, 0, -1, -3, -3, -5, -3, -4, -2, 0, 1, 0, -1, -1, 0, 1, 0, 1, 2, 0, 0, 2, 1, 2, 0, 0, 0, 0, 0, -1, -3, -3, -4, -3, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 1, 0, 1, 0, 0, 0, -3, -3, -2, -2, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 2, 1, 0, 1, 1, 2, 2, 0, 0, -2, -2, -3, -3, -2, -3, -1, 0, 0, 0, 0, -2, -3, -3, -2, -1, -1, 0, 0, 0, 1, 2, 3, 2, 2, -1, 0, -1, -1, -1, -1, -1, 0, 1, 1, 0, 0, -2, -2, -3, -2, -1, 0, -1, 0, 0, 0, 0, 1, 2, 0, 0, 0, -2, -2, -2, -1, -1, 0, -1, 1, 1, 0, 0, -2, -2, -2, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, -1, -1, -2, -2, 0, 0, 0, 0, 2, 0, 0, -1, -2, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, 1, 0, 1, 2, 1, 0, -1, -2, -2, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 2, 0, 0, 0, -1, 0, 1, 0, 1, 1, 1, 2, 1, 0, -1, -1, -1, 0, 0, -1, 0, -1, -2, -1, 0, 1, 1, 0, 2, 0, 0, 0, 3, 1, 3, 2, 4, 2, 1, -1, -2, -2, -3, -1, 0, 0, -1, -1, -2, -2, -1, 1, 1, 1, 2, 3, 4, 3, 5, 4, 5, 3, 5, 3, 1, 0, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 3, 2, 5, 6, 6, 6, 5, 5, 4, 4, 0, -1, -2, -3, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, -1, -2, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, 1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, -1, 0, 1, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -2, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 1, 0, -1, -2, -1, 0, 1, 1, 0, 2, 1, 1, 2, 2, 2, 0, -1, -2, -3, -3, -3, -2, -1, -1, -2, -1, 0, 0, -2, -1, -1, 0, -1, 0, 0, 1, 1, 1, 2, 3, 1, 1, -1, -2, -2, -2, 0, -1, 0, 0, -2, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, -1, 0, -1, -1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, -2, -1, 0, 0, -1, -2, 0, -1, 0, 0, 1, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, -2, -1, -1, -1, -1, 0, 0, 0, -2, 0, 0, -1, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, -1, -1, -1, 0, -1, 1, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, -1, -2, 0, 0, 1, 0, 1, -1, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -2, 0, 0, 0, 0, -1, 0, -2, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, -1, -1, -2, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, -3, -2, -2, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, -2, -2, -1, 0, -2, -1, -1, -1, -2, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -2, -1, -2, -1, -2, -2, -1, -1, -1, -2, 0, 0, -1, -1, 0, 1, 0, 0, 0, -2, -1, -1, 0, -1, 0, 0, -2, -1, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -3, -1, -2, -2, -1, -1, -2, -2, -1, 0, 0, -1, 0, 0, 0, 1, 0, -1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -3, -1, -2, 0, 0, -1, 0, -1, -1, -1, 0, 0, 1, 0, 1, 0, 1, 2, 1, 0, 0, 0, -1, -3, -1, -1, -3, -2, -2, -2, 0, -3, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, -1, -1, -1, -2, -1, -2, -2, -2, -2, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, -1, -2, 0, -2, -3, -4, -3, -3, -2, -3, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, -1, 0, 0, -2, -2, -2, -3, -2, -3, -4, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, -2, -3, -3, -2, -1, -2, -2, -1, 0, 0, 0, -1, 0, 0, 0, -2, -1, 0, 0, -1, 0, 0, 0, -2, -1, -2, -3, -2, -3, -1, -2, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 1, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, -2, -3, -3, -3, -1, -2, -2, -1, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, -2, -3, -2, -3, -2, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, -2, -2, -2, -3, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 1, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 2, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 2, 1, 2, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 2, 0, 0, 0, 2, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 2, 0, 1, 1, 1, 1, 0, 0, 2, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -1, -2, -2, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -2, 0, -2, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, -1, -1, -1, -2, -2, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, -1, -1, -1, -2, -1, 0, -1, -2, -1, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -1, -1, -2, -3, 0, 0, 0, 0, -2, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, 0, -1, -1, -1, -1, -2, -1, -1, -2, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, -2, -1, -1, -1, -2, 0, -2, -2, -2, -2, -2, -2, 0, 0, 0, 0, -2, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -3, -4, -5, -4, -3, -4, -3, -3, -4, -4, -3, -1, -2, 0, -2, -2, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -4, -4, -3, -4, -4, -2, -4, -2, -3, -2, -3, -2, -2, -2, -2, -2, -1, -1, 0, 1, 1, 1, 1, -1, 0, -1, -2, -4, -3, -2, -3, -3, -2, -1, -2, 0, 0, -1, -1, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, -3, -2, -1, -1, 0, -1, -2, -1, -1, 0, -1, -1, -2, 0, -1, -2, -1, -1, 1, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -2, -1, -2, -2, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, 0, -2, -2, 0, 0, 0, 0, -2, -1, -2, -1, -1, 0, -1, 0, 0, 1, 1, 2, 0, 1, 1, -1, 0, 0, 0, -1, 0, -2, -1, 0, 0, 0, -1, -2, 0, 0, -1, 0, 0, 1, 1, 2, 3, 1, 0, 2, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -3, -1, -1, -1, -2, 0, 0, 0, 1, 2, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 2, 0, -1, -1, -2, 0, -1, -2, 0, 0, 1, 0, 0, 0, 2, 0, 0, 1, 1, 2, 1, 1, 0, 1, 0, 2, 0, 0, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 2, 1, 1, 0, 0, -1, 0, 0, 0, -1, -2, -2, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 3, 2, 2, 3, 2, 1, 1, 0, 0, 0, 1, 0, -1, -1, -2, -1, -1, -1, 0, 1, 0, 1, 1, 1, 2, 2, 2, 4, 3, 3, 1, 3, 2, 0, 0, 0, 0, 0, 0, -2, -2, -2, -1, -1, -1, 0, 0, 0, 0, 1, 2, 2, 1, 2, 3, 3, 2, 1, 1, 1, 0, 1, 0, 0, 0, -2, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 2, 2, 2, 3, 3, 0, 1, 1, 0, 1, 1, 0, 0, -1, -1, -1, -1, -1, -2, 0, -2, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 2, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, -3, -2, 0, -2, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, 0, 0, -1, -1, -1, -1, 0, -1, -2, -1, -2, -2, -1, -2, -1, 0, 0, 0, 1, 0, 1, 1, 0, -1, -1, 0, 0, -2, -1, 0, 0, 0, -1, 0, -2, -3, -2, -1, -3, -1, -1, 0, 0, 0, 0, 0, 2, 0, 0, -1, 0, -2, 0, -2, -1, 0, -1, 0, -1, -2, -3, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, -2, -2, -2, -2, -2, -2, 0, -1, -3, -2, -1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -2, -2, -1, -3, -2, 0, -2, -1, -2, -3, -1, -1, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, -2, 0, -3, -2, -3, -2, -1, -1, -1, -1, -2, -1, -1, -1, -2, -3, -2, -1, -2, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, -2, -3, -2, -3, -3, -3, 0, -2, -2, -1, -2, -2, -2, -2, -1, -2, -1, -1, -1, 0, -1, -2, -2, -2, -2, -1, -4, -2, -2, -3, -2, -1, -2, -2, -1, -1, -3, -3, -3, -2, -3, -3, -1, -2, -2, -2, -1, -3, -2, -3, -2, -3, -4, -2, -3, -3, -1, -1, 0, -2, -2, -3, -2, -2, -2, -2, -3, -2, -2, -2, -2, -2, -3, -3, -2, -1, -2, -3, -2, -2, -2, -3, -3, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, -2, 0, 0, -1, 0, 1, 1, 2, 4, 4, 3, 3, 1, 0, -1, 0, -2, -1, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, -2, -1, 0, 0, 0, 1, 3, 2, 3, 3, 2, 1, -1, 0, -2, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, -1, -2, -2, 0, -1, 0, 0, 1, 2, 3, 1, 1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, -1, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, -1, -1, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 2, 2, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 1, 1, 2, 1, 2, 2, 1, 2, 1, 0, 1, 1, 0, 0, -1, 1, 1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 1, 0, 2, 1, 1, 1, 2, 0, 2, 0, 0, -1, 0, 0, 0, 2, 0, 1, 1, 0, 1, 0, 2, 0, 1, 2, 2, 2, 1, 1, 3, 2, 0, 2, 1, 0, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, 1, 2, 1, 0, 0, 1, 1, 0, 2, 2, 3, 1, 1, 0, 2, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 3, 0, 2, 0, 2, 1, 1, 2, 2, 1, 1, 0, 0, 0, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 1, 1, 2, 3, 2, 2, 2, 0, 0, 1, 0, 0, -1, -2, -1, -2, -1, 0, 1, 0, 1, 3, 2, 0, 2, 2, 0, 2, 2, 3, 2, 2, 2, 1, 2, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 2, 2, 0, 1, 1, 2, 2, 3, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 1, 2, 0, 1, 1, 2, 2, 2, 3, 1, 2, 1, 2, 1, 2, 1, 2, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 2, 3, 2, 2, 1, 0, 0, 1, 0, 1, 2, 1, 0, 1, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 1, 0, 1, 0, 1, 1, 1, 0, 2, 1, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 2, 3, 2, 2, 2, 2, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 3, 2, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, -2, -1, 0, 0, 0, 1, 2, 2, 4, 4, 2, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, -2, -1, 0, 1, 0, 2, 3, 2, 4, 4, 4, 2, 1, 0, 0, -2, 0, -1, 0, -1, -1, -2, -1, -1, -1, -1, -1, -2, 0, 0, 0, 1, 2, 3, 4, 5, 3, 3, 0, 0, -1, -3, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -2, 0, 0, 0, 1, 3, 3, 4, 5, 5, 3, 2, 1, 0, -3, -2, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 5, 5, 3, 3, 1, 1, 0, 0, -2, -4, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 1, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 1, 0, 1, 1, 1, -1, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, -2, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, -1, 1, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -2, -1, 0, 0, -2, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, 0, -1, -1, 0, 0, 0, 0, 0, -3, -1, -1, -1, 0, -2, 0, -1, 0, 0, 0, 1, 0, 0, 1, 2, 1, 2, 3, 5, 4, 1, 1, 1, 0, 1, -3, -2, -2, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 2, 2, 2, 1, 1, 0, -1, 0, -1, -2, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 2, 1, 1, 0, 0, 1, 1, 0, -2, -3, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, 0, 1, 0, 1, 0, 2, 0, 1, 0, -2, -2, 0, 0, 1, 0, 2, 0, 1, 1, 0, 0, 1, 0, 0, -1, 0, -1, 0, 1, 0, 0, 1, 2, 1, 0, -2, -1, -1, 1, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, -1, 1, 1, 1, 0, 1, 1, 1, 0, -1, -1, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 2, 2, 0, 1, 0, 0, 0, 0, 0, -1, -1, -2, -2, 0, 1, 0, -1, 0, 1, 1, 0, 0, 1, 2, 1, 2, 2, 1, 2, 1, -1, 0, -1, 0, -1, 0, -2, -3, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 2, 1, 0, 1, 2, 0, 0, -1, 0, 0, 0, -3, -4, -2, -1, -1, 0, 1, 0, 1, 0, 0, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -4, -2, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, -1, -2, -3, -2, -2, -2, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -4, -1, -3, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -2, -2, -2, -1, -2, -1, -1, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -2, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 2, 2, 0, -1, 0, -1, -1, -2, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 1, 0, 1, 0, 1, 2, 2, 2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, -1, -1, 0, 0, 2, 1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 1, -1, -1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 2, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 2, 3, 2, 1, 3, 1, 2, 0, 0, -1, -2, -1, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 1, 1, 2, 3, 2, 3, 3, 2, 0, -1, 0, -1, -2, 0, 0, 1, 0, -1, 0, 0, 0, 1, 1, 2, 2, 1, 1, 3, 4, 4, 2, 2, 1, 3, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, -1, -1, 0, 0, 0, 1, 0, 1, 2, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, -2, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, -1, 0, 0, 0, -1, -1, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, -6, -5, -4, -5, -5, -5, -5, -4, -4, -5, -4, -6, -6, -4, -5, -2, -2, 0, 0, 3, 3, 2, 2, 4, 5, 5, -6, -6, -5, -3, -3, -3, -3, -3, -2, -2, -2, -3, -4, -4, -3, -3, -2, 0, 0, 1, 3, 2, 3, 3, 5, 4, -6, -6, -5, -4, -4, -3, -2, -3, -3, -3, -3, -3, -2, -1, -1, -2, 0, -1, 0, 1, 2, 1, 3, 3, 4, 5, -6, -5, -3, -2, -2, -2, -3, -1, -1, -2, -2, -3, -3, -3, -3, -2, 0, 0, 1, 2, 1, 0, 1, 3, 3, 2, -6, -3, -3, -2, -4, -3, -3, -3, -1, -1, -2, -4, -2, -3, -4, -3, -1, 0, 2, 2, 3, 2, 2, 2, 4, 3, -4, -5, -2, -2, -2, -2, -3, -3, -1, -2, -3, -3, -3, -3, -5, -3, 0, 0, 2, 2, 2, 1, 2, 3, 3, 4, -4, -3, -2, -4, -4, -3, -2, -2, -2, -3, -4, -4, -2, -4, -4, -2, -1, 1, 0, 2, 1, 2, 3, 2, 5, 4, -4, -2, -2, -3, -4, -4, -2, -2, -3, -2, -3, -1, -2, -1, -4, -2, -3, -1, 1, 0, 0, 2, 2, 3, 4, 3, -2, -2, -2, -2, -2, -2, -2, -3, -2, -3, -3, -1, -3, -2, -2, -2, -1, 0, 1, 1, 0, 2, 2, 3, 3, 3, -4, -4, -3, -3, -3, -2, -1, -2, -1, -1, -2, -3, -1, -1, -1, -2, -1, 0, 0, 2, 1, 1, 1, 3, 3, 4, -3, -3, -3, -3, -2, -3, -2, -1, -2, -1, -2, -1, -1, -1, -2, -1, 0, 0, 1, 0, 1, 0, 2, 3, 3, 4, -3, -4, -2, -1, -2, -2, 0, 0, 0, -2, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 2, 2, 3, 4, -2, -4, -2, -2, -3, -3, -1, -2, -2, 0, 0, -1, 0, 0, -1, -1, 0, 0, 3, 2, 1, 0, 0, 4, 3, 3, -2, -4, -3, -1, -3, -1, 0, -1, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, 1, 3, 2, 1, 1, 3, 3, 4, -2, -3, -2, -1, -1, -2, 0, -1, -1, 0, -1, 0, 0, -2, -2, 0, -1, 1, 2, 2, 3, 1, 1, 1, 4, 3, -2, -3, -2, -2, -2, -3, -2, -1, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 1, 1, 3, 2, 0, 3, 3, 4, -3, -3, -3, -2, -1, -3, -2, -1, -2, 0, 0, -2, -2, -4, -3, -3, 0, 0, 2, 3, 2, 3, 3, 3, 2, 3, -5, -3, -2, -1, -1, -2, -1, -1, -2, -1, -1, -1, -4, -3, -2, -3, -2, 0, 1, 3, 3, 2, 2, 2, 3, 5, -4, -3, -3, -1, -1, -1, -2, -2, 0, 0, -2, -1, -2, -3, -5, -3, -2, 0, 1, 4, 3, 3, 3, 4, 4, 5, -4, -3, -2, -2, -1, -2, -1, -2, -1, -1, -2, -4, -3, -2, -3, -4, -3, -1, 0, 2, 1, 4, 3, 3, 4, 5, -4, -3, -4, -3, -2, -2, -1, -2, -1, -2, -4, -3, -3, -2, -1, -2, -2, -1, 0, 1, 2, 2, 4, 4, 5, 4, -5, -3, -4, -3, -2, -2, -2, -2, -2, -2, -2, -4, -3, -2, -3, -3, -3, 0, 1, 1, 2, 3, 4, 5, 5, 5, -5, -3, -4, -3, -2, -2, -1, -3, -1, -3, -2, -2, -4, -3, -2, -1, -3, -1, 0, 2, 2, 3, 6, 5, 5, 5, -4, -5, -4, -4, -5, -4, -4, -3, -2, -3, -3, -3, -2, -3, -3, -4, -3, 0, 0, 2, 2, 5, 6, 5, 6, 6, -4, -6, -4, -4, -5, -5, -4, -4, -4, -2, -3, -3, -2, -3, -2, -1, -2, 0, 0, 2, 4, 3, 5, 5, 6, 7, -6, -5, -5, -6, -7, -6, -5, -5, -3, -5, -4, -4, -4, -2, -1, -1, 0, 0, 0, 2, 5, 5, 4, 7, 7, 6, -2, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, -1, 1, 0, 1, 1, 1, 2, 1, 2, 1, 1, 3, -2, -2, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 1, 1, 3, 2, 3, 0, 0, 2, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 2, 3, 2, 2, 1, 2, 1, 1, 1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, 1, 2, 2, 2, 2, 1, 0, 2, 2, 0, -1, -1, 1, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 2, 0, 1, 0, 1, 2, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, -2, -1, -1, -2, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, -1, -1, 0, 0, -1, 0, 0, -2, -1, -2, -1, -1, -2, -2, -2, -2, 0, 1, 0, 1, 0, 2, 1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, -3, -1, -2, -2, -3, -2, -3, -2, -1, 0, 1, 0, 1, 0, 0, 2, 2, 0, 0, 1, 1, 0, 0, -1, -2, -2, -2, -1, -3, -2, -2, -2, -4, -3, -1, -1, -1, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, -1, 0, 0, 0, -2, -3, -3, -1, -2, -3, -3, -3, -3, -1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, 0, -2, -1, -1, -3, -2, -3, -5, -4, -1, 0, -1, -1, 0, 0, 0, 1, 2, 1, 1, 0, 0, -1, 0, 0, -1, -2, -1, -3, -2, -2, -3, -5, -3, -2, -3, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -3, -3, -4, -5, -4, -3, -2, -2, 0, -1, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, -3, -2, -3, -5, -5, -2, -2, -2, -1, 0, 0, 0, 0, 2, 2, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -2, -3, -2, -4, -4, -3, -1, -1, 0, -1, -1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, -3, -3, -3, -3, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, -3, -4, -4, -3, -2, 0, 0, 0, 1, 1, 0, 0, 0, 2, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -2, -3, -3, -3, -3, -1, 0, 0, 1, 1, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -2, -3, -2, -4, -3, -2, -1, 0, 0, 1, 1, 1, 1, 1, 0, 1, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, -2, -2, -3, -3, -3, -1, 0, 0, 0, 0, 2, 2, 2, 0, 3, 1, -1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, -3, 0, 0, 0, 0, 1, 0, 1, 0, 2, 2, 4, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -2, -1, -1, 0, 0, 1, 1, 2, 1, 2, 2, 2, 4, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 1, 2, 1, 3, 3, 2, 3, 1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 2, 3, 3, 1, 3, 2, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 3, 1, 3, 3, 3, 4, 2, 4, -2, -1, -2, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 1, 2, 3, 2, 2, 3, 3, 3, 3, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, -1, 0, 0, -2, -1, -1, 0, -1, -1, -1, 0, 1, 2, 1, 2, 2, 2, 1, 1, 1, 1, 0, 0, -1, -1, 0, -1, 0, -1, -1, -2, -1, -1, -2, -1, -1, 1, 1, 1, 3, 2, 3, 2, 3, 3, 3, 1, 2, 0, 1, 0, 0, 0, -2, -2, -1, -1, -2, -1, -1, -1, -1, -1, 1, 1, 1, 2, 2, 3, 3, 2, 1, 2, 3, 3, 1, 1, 0, 0, 0, -2, -3, -2, -1, -2, -1, -2, -2, -2, 0, 0, 0, 1, 1, 2, 3, 4, 4, 4, 5, 3, 2, 0, 0, -1, -2, -1, -2, -4, -1, -1, -1, 0, -1, 0, 0, 2, 1, 0, 1, 3, 3, 2, 2, 4, 4, 5, 3, 2, 0, 0, 0, -2, -4, -3, -3, -2, -2, 0, -1, -2, 0, 0, 0, 0, 0, 1, 4, 1, 3, 4, 5, 4, 4, 2, 0, -1, -1, -2, -4, -4, -4, -2, -3, -1, -2, 0, 0, 0, -1, 0, 0, 3, 3, 2, 2, 3, 6, 5, 3, 1, 0, -1, 0, -1, -2, -3, -4, -3, -4, -3, -2, 0, 0, 0, 0, 0, 0, 3, 3, 2, 3, 3, 5, 5, 2, 3, 2, 0, -1, -1, -3, -3, -2, -3, -2, -3, -2, -1, 0, 0, -1, 0, 2, 1, 3, 1, 4, 4, 5, 5, 2, 2, 2, 0, 0, 0, -1, -2, -4, -4, -4, -3, -2, 0, 0, 0, -1, 0, 1, 2, 1, 3, 4, 5, 7, 6, 2, 2, 1, 0, 0, 0, -1, -3, -3, -4, -3, -2, -3, -1, 0, -1, 0, 0, 0, 1, 2, 1, 5, 4, 7, 5, 4, 1, 0, 0, 1, -1, -1, -2, -3, -5, -2, -3, 0, 0, -1, -2, -2, 0, 1, 2, 1, 2, 4, 4, 5, 7, 3, 2, 2, 0, 0, -1, -1, -3, -5, -5, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 3, 3, 4, 4, 5, 4, 2, 0, 0, 0, -2, -2, -3, -5, -5, -2, -2, 0, 0, 0, 0, -1, -1, 0, 2, 2, 1, 2, 4, 5, 5, 2, 2, 2, -1, 0, -1, -1, -1, -3, -4, -2, -2, 0, -2, 0, 0, -1, 0, 1, 1, 3, 2, 3, 5, 4, 2, 3, 2, 2, -1, 0, -1, 0, 0, -3, -3, -3, -2, -1, -1, 0, -1, -1, 0, 2, 3, 3, 1, 3, 3, 5, 2, 2, 2, 1, 0, -1, 0, 0, -1, -1, -2, -3, -1, -1, 0, -1, 0, -2, -2, 1, 2, 2, 3, 4, 4, 5, 1, 1, 2, 0, -2, -2, 0, -1, 0, -2, -2, -4, -2, -1, 0, 0, 0, -3, -1, 0, 0, 0, 0, 4, 4, 3, 2, 3, 2, -1, -1, -2, 0, -1, 0, 0, -1, -4, -2, -2, 0, -1, 0, -1, -3, -1, 0, 1, 1, 2, 3, 2, 2, 3, 2, 0, 0, -3, -1, -1, -1, 0, 0, -2, -2, -1, -1, -1, 0, -1, -2, -1, 0, 1, 1, 2, 2, 1, 2, 1, 0, 0, 0, -3, -2, -2, -2, -1, 0, -2, -1, 0, 0, -1, 0, -2, -1, 0, 0, 0, 2, 2, 2, 2, 1, 1, 0, 0, -1, 0, -2, -4, -2, -1, -1, -3, -2, 0, -1, 0, 0, -2, 0, -1, -2, -1, 0, 0, 2, 2, 0, 2, 0, 0, 0, -1, -2, -2, -2, -1, 0, -2, -2, 0, 0, -1, 0, -2, -2, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -2, -1, -2, -2, 0, -3, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, -3, -3, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -2, -2, 0, -2, 0, -1, -1, -1, -1, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -2, -3, -3, -3, -2, -1, -1, -1, -1, 0, 0, -1, -1, 0, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -3, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, -2, -2, -2, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, -2, -1, 0, 0, 1, 0, 1, 2, 0, 2, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, -1, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, -1, 0, -2, -1, -2, -2, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 1, 0, 1, 0, -1, 0, 2, 1, 0, 0, 0, 0, 0, -2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -2, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 2, 0, 0, 1, 1, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 2, 1, 2, 2, 1, 0, 0, 1, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -2, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, -1, -2, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -2, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, -2, -1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 1, -1, 0, -1, -1, -3, -2, -1, -1, 0, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, 0, 0, -1, -2, -2, -2, -1, -1, -1, -1, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, -2, -1, -2, -1, -3, -3, -2, -2, -1, -2, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 2, 1, 0, 0, -1, 0, -1, -2, -2, -1, -2, -3, -2, -4, -4, -3, -3, -1, -1, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -2, -1, -2, -3, -3, -3, -4, -3, -2, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -2, -3, -2, -4, -3, -3, -2, -3, -1, -1, -1, 0, -2, -1, 0, -2, -1, 0, 0, -1, 0, 0, 0, -2, -2, -1, -1, -4, -2, -3, -4, -3, -1, -2, -1, -2, -1, -1, -1, 0, -1, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -2, 0, -2, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, 0, -2, -2, 0, 0, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, -2, -2, 0, -2, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, -1, -1, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, -1, -2, -1, 0, 0, 0, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, -2, -2, -1, -2, -1, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -2, -1, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -2, -1, -2, -2, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -2, -2, -2, -2, -1, -2, 0, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -2, -2, -2, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, -2, -1, -2, -2, -1, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -2, 0, 0, -1, 0, -1, 0, 1, -2, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, -1, 0, -1, 1, 2, 1, 2, 3, 5, 6, 5, 7, 7, 6, 5, 2, 0, -1, -2, -1, 0, 0, 0, -1, 0, -2, 0, -1, 0, -1, 0, 1, 3, 1, 2, 4, 5, 6, 7, 4, 2, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -2, 0, 1, 1, 2, 3, 4, 5, 5, 4, 1, 0, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 3, 3, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 2, 0, 0, 0, 0, -2, 0, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 1, 0, 0, 0, 2, 2, 1, 1, 0, 0, -2, -2, -1, 0, 2, 2, 2, 3, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, -1, -1, 1, 1, 1, 1, 1, 0, 1, 1, 0, 2, 1, 2, 0, -1, 0, 0, -1, 0, 0, 2, 1, 1, 0, 3, 0, 1, 0, 1, 0, 3, 1, 1, 1, 0, 2, 1, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 2, 2, 0, 3, 1, 1, 1, 0, 0, 2, 2, 0, -1, -1, 0, 0, 0, 0, 2, 2, 1, 2, 2, 4, 1, 0, 1, 1, 3, 1, 2, 1, 1, 0, 0, 1, 0, -1, -2, -1, -1, 0, 0, 1, 1, 2, 1, 2, 3, 5, 1, 2, 2, 3, 3, 2, 2, 2, 0, 0, 1, 2, 0, -1, -2, -1, -1, -1, 0, 0, 1, 0, 0, 2, 5, 5, 1, 1, 2, 1, 2, 1, 2, 1, 0, 1, 2, 0, -1, -2, -2, -1, -3, -2, 0, 0, 0, 1, 1, 3, 5, 7, 1, 1, 1, 2, 1, 1, 2, 0, 0, 1, 0, 0, 0, -3, -3, -4, -3, -3, -1, 0, 2, 1, 2, 3, 4, 5, 1, 0, 0, 2, 2, 2, 2, 2, 0, 0, 1, 0, -1, -1, -1, -2, -3, -2, 0, 0, 0, 1, 2, 1, 3, 4, 0, 1, 0, 0, 1, 3, 3, 2, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 4, 5, 0, 0, 0, 0, 0, 3, 1, 1, 1, 0, 2, 1, 2, 0, 0, -1, -1, -1, 1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 1, 3, 3, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 3, 1, 1, 2, 0, 0, 2, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, -1, 0, 1, 3, 1, 2, 1, 1, 0, 0, 1, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, -1, -1, 0, 1, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 3, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 4, 4, 2, 3, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 4, 5, 3, 2, 3, 1, 0, 0, -2, -2, 0, -1, -1, -2, -1, 0, -1, -2, 0, 0, 1, 0, 1, 3, 2, 3, 5, 5, 5, 5, 2, 1, 0, -2, -2, -2, -1, -1, 0, 0, 0, -1, -1, 0, 1, 0, 0, 2, 3, 2, 5, 6, 6, 4, 5, 3, 2, 0, -1, -3, -3, -4, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, -1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, -1, -1, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, 1, 2, 2, 1, 3, 3, 2, 2, 2, 1, -1, -1, 0, 1, -1, 0, -2, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 2, 3, 1, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 1, -1, -1, 0, 0, 1, 0, 0, 1, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, -2, -2, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, -2, -2, -1, -1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, -1, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 1, -1, -1, 0, 0, 0, 0, 2, 1, 0, 1, 0, -1, 0, 1, 2, 1, 2, 1, 1, -1, 0, 0, 1, 0, 1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 2, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 1, 1, 2, 1, 0, 2, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, -1, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, -2, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, -2, 0, -1, -1, 0, -1, -1, 0, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, -1, -2, -1, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 2, 0, 0, -1, 0, 0, -2, 0, -1, 0, -1, 0, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, -1, 1, 1, 1, 0, 1, 1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, -1, 0, 1, 1, 0, 1, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, -2, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 3, 2, 0, 0, -1, -1, -2, -1, -1, -7, -5, -5, -4, -5, -6, -4, -3, -3, -5, -4, -4, -4, -4, -5, -3, -3, -1, 0, 0, 1, 3, 3, 5, 4, 6, -6, -6, -6, -3, -5, -2, -2, -3, -2, -3, -3, -3, -1, -3, -3, -2, -3, -1, 0, 0, 2, 2, 3, 4, 4, 5, -5, -6, -4, -3, -3, -3, -2, -3, -3, -1, -1, -2, -2, 0, -3, -2, -3, 0, -1, 0, 1, 1, 1, 3, 4, 4, -5, -5, -4, -3, -4, -2, -1, -2, -2, -1, -3, -3, -3, -1, -1, -4, -2, -1, 0, 0, 1, 1, 0, 2, 1, 4, -4, -4, -5, -3, -4, -4, -3, -2, -1, -2, -3, -4, -2, -2, -1, -2, -1, -1, -1, -1, 0, 1, 1, 1, 1, 2, -4, -3, -5, -3, -3, -3, -2, -3, -2, -2, -3, -3, -2, -2, -2, -3, -3, -1, 0, 0, 0, 0, 0, 0, 1, 2, -5, -5, -4, -3, -2, -2, -3, -2, -3, -2, -4, -4, -3, -2, -4, -1, -2, -1, -2, -1, 0, 0, 1, 0, 2, 2, -3, -4, -2, -4, -2, -2, -2, -3, -2, -2, -2, -2, -2, -3, -2, -3, -3, -3, -2, -1, 0, 0, 1, 1, 1, 2, -3, -2, -3, -4, -3, -3, -1, -3, -3, -2, -2, -1, -1, -2, -2, -3, -3, -3, -2, -1, 0, 0, 0, 0, 2, 3, -3, -2, -3, -2, -2, -2, -3, -3, -1, -1, -2, -3, -3, -1, -2, -1, -1, -1, -2, -1, -1, 0, 1, 1, 1, 1, -4, -2, -3, -3, -2, -1, -1, -2, -2, -2, -2, -1, -2, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 3, 2, -3, -2, -3, -2, -3, -3, -2, -1, 0, -2, -2, -1, -1, -2, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 3, 3, -3, -3, -2, -4, -4, -2, -2, -2, -1, 0, -1, -1, -2, -1, 0, 0, 1, 1, 0, -1, -1, -1, -1, 2, 2, 2, -3, -3, -2, -3, -3, -3, -1, -2, -1, -1, -1, -2, 0, -2, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 3, -3, -3, -1, -1, -1, -3, -2, -1, -2, -2, 0, -1, -1, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 2, 3, -4, -3, -1, -2, -1, -3, -3, -2, -1, -1, -1, 0, -2, -2, -3, -2, -2, -1, 0, 1, 0, 1, 0, 0, 1, 2, -3, -2, -2, -3, -2, -2, -1, -2, -2, -1, -2, -2, -2, -4, -3, -5, -4, -3, -1, 1, 0, 1, 1, 0, 1, 4, -2, -4, -4, -2, -3, -3, -3, -2, -2, -2, -1, -3, -4, -4, -5, -6, -5, -4, 0, 1, 0, 1, 0, 2, 3, 4, -5, -3, -4, -3, -1, -1, -1, -2, -2, -2, -2, -1, -3, -4, -6, -5, -6, -3, -2, 0, 0, 1, 1, 2, 2, 5, -5, -2, -4, -4, -2, -2, -3, -2, -2, -3, -2, -3, -5, -4, -6, -6, -5, -4, -2, -2, -1, 0, 1, 1, 4, 4, -5, -3, -4, -3, -3, -3, -3, -3, -2, -2, -4, -4, -4, -5, -4, -6, -7, -4, -3, -2, 0, 0, 1, 3, 3, 5, -4, -3, -5, -2, -5, -4, -3, -4, -1, -3, -4, -4, -3, -3, -4, -5, -6, -5, -4, -2, 0, 0, 2, 3, 3, 6, -4, -4, -5, -3, -3, -3, -4, -4, -2, -3, -4, -4, -3, -5, -5, -5, -6, -3, -3, -3, 0, 0, 2, 2, 3, 5, -5, -6, -5, -5, -6, -5, -4, -2, -3, -4, -3, -4, -5, -5, -6, -4, -5, -3, -3, -2, 0, 1, 2, 4, 4, 4, -6, -5, -6, -6, -6, -6, -5, -5, -2, -2, -5, -3, -4, -3, -4, -5, -5, -2, -2, 0, 0, 1, 4, 3, 5, 6, -5, -5, -6, -7, -6, -6, -4, -4, -4, -5, -5, -6, -4, -4, -4, -3, -3, -1, -1, 0, 2, 2, 4, 6, 6, 5, -1, 0, 0, -1, -2, 0, 0, 0, 0, -1, -1, 0, -2, -1, 0, 0, 0, 1, 2, 1, 1, 2, 2, 0, 0, 1, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 3, 2, 1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 3, 1, 1, 0, 1, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 2, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, -2, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, -2, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -2, -1, -1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 2, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 2, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 2, 2, 1, 0, 0, 2, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 2, 1, 1, 0, 2, 1, 2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 1, 1, 2, 2, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 2, -1, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, -2, -1, 0, 1, 0, 0, 1, 0, 2, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, -2, -1, 0, 0, 0, 1, 0, 0, 1, 2, 2, 2, 0, 1, 1, 1, -1, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, 1, 0, 0, 0, 0, 1, 1, 2, 1, 0, -1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 2, 1, 1, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 2, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 2, 2, 0, 2, 0, 0, 1, 0, 0, 2, -1, 0, -1, 0, 1, 1, 0, 2, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 2, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, 2, 1, 2, 1, 0, 1, 0, 2, 1, 0, 0, 1, 0, 2, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 1, 2, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 2, 0, 2, -1, 0, 0, 0, 0, 2, 0, 1, 1, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 2, 0, 1, 1, 2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 2, 1, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 2, 2, 2, 1, 1, -1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 1, 1, 1, 0, 0, 1, 0, 1, 2, 2, 0, 1, 0, 1, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, -1, 0, -1, -1, -1, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 1, 0, 1, -1, -2, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 2, 1, 1, 1, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 2, 1, 1, -1, -1, -2, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 0, 2, 2, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, -2, -1, -2, -2, -2, -2, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 2, 0, 0, 0, 0, -2, -3, -2, -3, -1, 0, -2, 0, 0, -1, 0, 1, 1, 0, 0, 0, 1, 2, 1, 2, 2, 1, 1, 0, 1, 0, -2, -2, -2, -2, -2, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 2, 2, 0, 0, 0, 0, 0, -1, -2, 0, -2, -1, -2, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 2, 0, 1, 0, 1, 0, 0, 0, 1, 1, -1, -1, -1, -1, 0, -1, 0, 0, 1, 0, 2, 3, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 2, 2, 3, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, -2, 0, -1, 0, 0, 0, 0, 1, 2, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 2, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 0, -1, 1, 0, 0, 1, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 1, 1, 2, 1, 1, 0, 0, 1, 1, 1, 1, 0, 1, 0, 1, 1, 3, 0, 1, 0, 0, 0, 2, 1, 2, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 1, 2, 2, 2, 0, 2, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 1, 2, 3, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, -1, -1, 0, 1, 0, 1, 1, 2, 3, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, -1, -1, -2, 0, 0, 0, 0, 1, 2, 1, 1, 3, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 3, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 3, 1, 0, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 1, 1, 1, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 2, 0, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, 1, 2, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, 1, 1, 1, 1, 2, 2, 1, 1, 1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 2, 1, 0, 1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 2, 1, 2, 2, 2, 2, 2, 3, 2, 1, 0, -1, 0, -2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 0, 1, 2, 2, 1, 2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 2, 3, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -2, -2, -1, -1, 0, 0, 0, 0, 1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, -2, -1, -1, -2, -1, -2, -2, 0, 0, -1, 0, -1, 1, 0, 1, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -2, -2, 0, -1, -1, -2, -2, -1, -2, 0, -1, -1, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, -2, 0, 0, 0, -1, -1, 0, -2, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 2, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 1, 1, 1, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 1, 0, 2, 1, 1, 0, 0, 0, 1, 1, 0, 0, -1, 1, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, -1, 0, -1, 1, 1, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 1, 1, 2, 0, 0, 2, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 1, 2, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 2, 0, 0, 0, 1, 2, 2, 2, 1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 2, 1, 1, 3, 3, 2, 2, 0, 0, 0, 0, -1, 0, -1, -1, -1, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 3, 2, 0, 0, -2, -2, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, -2, -1, 0, 0, 1, 1, 2, 3, 2, 2, 0, 0, 0, -1, -1, 0, 0, 0, 0, -2, -1, -1, -2, -2, -1, -1, 0, 0, -1, 0, 0, 2, 1, 2, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, -1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, -2, 0, 0, 2, 2, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, -1, 0, 1, 2, 1, 1, 1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, -2, 0, 0, -1, 0, 1, 0, 0, 0, 0, 2, 0, 1, 1, 1, 0, 0, 0, 1, 2, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 2, 0, 1, 2, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 2, 2, 1, 0, 0, 1, 0, 0, 2, 1, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 2, 1, 1, 1, 2, 1, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 2, 2, 3, 2, 3, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 1, 0, 1, 1, 1, 2, 3, 1, 4, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 1, 1, 2, 3, 2, 1, 3, 4, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 2, 0, 0, 0, 1, 1, 1, 0, 2, 1, 1, 3, 2, 3, 1, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, -1, 1, 0, 0, 1, 1, 0, 1, 2, 2, 1, 3, 2, 3, 3, 1, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 2, 3, 2, 2, 3, 2, 2, 1, 1, 0, 0, 2, 0, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 3, 2, 1, 1, 1, 1, 1, 1, 2, 2, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 1, 1, 1, 3, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 2, 2, 3, 3, 3, 2, 3, 2, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 3, 3, 2, 3, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 2, 3, 4, 3, 1, 1, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, -2, 0, -1, 0, -2, -1, -2, 0, 0, 1, 1, 2, 4, 2, 3, 2, 2, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, -2, -2, 0, 0, 0, 1, 2, 2, 3, 3, 2, 2, 1, 2, 1, 0, -1, 0, 0, -1, 0, -1, -2, -1, -1, -2, -2, 0, -1, -1, 0, 1, 1, 2, 1, 3, 4, 3, 1, 0, 0, 0, -1, 0, 0, -1, 0, -2, -2, -1, -1, -1, -1, -1, -1, -1, 0, 1, 0, 3, 3, 2, 2, 1, 1, 0, -1, -2, -2, 3, 3, 3, 1, 2, 1, -1, -2, -2, -3, -3, -3, -1, 0, 0, 2, 1, 2, 1, 1, 1, 2, 0, -1, -3, -4, 4, 2, 2, 0, 0, -1, -2, -2, -3, -4, -3, -3, -2, -1, -1, 1, 0, 0, 2, 2, 2, 3, 1, 0, -1, -3, 3, 1, 1, 0, 0, -1, -2, -3, -4, -2, -4, -2, -3, -3, -1, 1, 1, 1, 1, 3, 3, 2, 2, 0, 1, 0, 3, 2, 1, 1, -1, 0, -2, -3, -2, -2, 0, -2, -1, -1, 0, 0, 0, 1, 2, 1, 1, 1, 1, 1, 0, 0, 3, 2, 0, 1, 0, -2, 0, -2, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 2, 1, 2, 1, 0, 0, 0, 0, 3, 1, 0, 2, 0, 0, -1, 0, 0, 2, 2, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 2, 1, 2, 2, 0, 0, 0, -1, -1, 0, 0, 2, 4, 2, 1, 1, 1, 2, 0, 1, 1, 0, 0, 0, 0, 0, 2, 0, 2, 0, 1, 0, 0, 0, 0, 0, 1, 1, 4, 2, 2, 0, 1, 0, 1, 1, 0, 0, 0, 1, 2, 3, 3, 3, 0, 0, 0, -1, 0, 0, 1, 1, 3, 2, 2, 1, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 2, 3, 3, 1, 0, -1, 0, 0, 0, 2, 1, 3, 3, 2, 2, 2, 0, 0, 0, -1, 0, 0, 0, -1, 1, 1, 2, 3, 3, 2, 0, 0, -1, 0, 1, 3, 2, 4, 4, 3, 1, 0, 0, -2, -2, 0, -1, -1, -1, 0, 1, 1, 4, 3, 2, 2, 0, 0, 0, 1, 2, 3, 5, 5, 6, 3, 2, 0, -1, -1, -1, -1, -2, -3, -2, -1, 0, 2, 2, 4, 3, 1, 2, 2, 2, 1, 2, 3, 4, 4, 4, 4, 2, 2, -1, -1, -3, -3, -3, -4, -3, -2, 0, 2, 4, 3, 3, 2, 2, 2, 2, 3, 2, 3, 5, 4, 3, 4, 2, 0, 0, -1, -1, -1, -2, -4, -2, -1, 0, 0, 3, 4, 4, 2, 0, 1, 0, 0, 1, 2, 3, 1, 1, 2, 0, 0, 0, -1, -2, -1, -2, -3, -1, -1, 0, 0, 2, 3, 3, 2, 2, 1, 1, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, 0, -1, -1, -2, -1, -1, 0, 0, 2, 3, 2, 2, 3, 2, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 3, 2, 4, 2, 2, 0, -1, 0, 0, 2, 2, 1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 2, 2, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 2, 1, 1, 0, 0, 1, 0, 2, 1, 0, 1, 1, 3, 2, 2, 0, 0, 0, 1, 1, 1, 0, -1, -1, 1, 0, 3, 3, 2, 1, 1, 1, 2, 2, 0, 2, 2, 0, 2, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 3, 3, 3, 2, 0, 0, 1, 0, 2, 1, 0, 1, 1, 0, 1, 2, 1, 0, 0, 0, 2, 0, 0, -1, 0, 1, 3, 3, 1, 1, 0, 0, 2, 2, 1, 2, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, 2, 1, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 2, 3, 1, 2, 1, 0, 1, 1, 1, 1, 2, 0, 1, 2, 2, 2, 0, -1, -2, -1, -2, 0, 0, -1, 0, 0, 2, 2, 2, 1, 0, 0, 0, 0, -1, 4, 3, 0, 2, 1, 1, 2, 0, -1, -2, -2, -2, -1, -2, -2, -1, 0, 1, 2, 2, 2, 1, 0, 0, -2, 0, 2, 3, 3, 2, 4, 3, 3, 2, 0, -1, 0, -3, -1, -3, -2, 0, 0, 2, 1, 3, 0, 0, 0, -3, -3, -3, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, -1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, -1, -1, -1, 0, 1, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, -1, -2, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -2, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -2, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, -1, 0, -1, -2, -3, -2, -4, -3, -4, -3, -3, -2, 0, -1, 0, -2, -2, -2, -5, -5, -5, -5, -6, -6, 1, 0, -1, -3, -1, -3, -3, -3, -3, -3, -3, -3, -4, -2, -2, -2, -1, -1, -3, -3, -2, -2, -3, -4, -3, -4, 3, 0, 0, -1, -1, -2, -3, -1, -3, -5, -5, -4, -4, -3, -3, -2, -3, -2, -1, -1, -1, -2, -2, -2, -4, -3, 3, 0, 0, -2, -1, -2, -1, -2, -2, -2, -4, -3, -3, -2, -4, -4, -3, -2, -3, -2, -1, -1, -2, -2, -4, -4, 2, 1, 0, 0, -2, -1, -2, -2, -2, -2, -3, -2, -3, -2, -3, -2, -4, -3, -1, -2, 0, 0, -2, -1, -2, -4, 2, 2, 0, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, -2, -2, -2, -3, -2, -2, -1, 0, 0, -2, -2, -3, -2, 1, 1, 0, 0, 0, -1, 1, 0, 1, 1, 1, 1, 1, 0, 0, -1, -1, -1, -2, 0, -1, 0, -1, -2, -1, -2, 2, 0, 0, 0, 1, 0, 0, 2, 0, 2, 2, 3, 2, 2, 1, 1, 0, 0, -2, 0, 0, 0, 0, -2, -1, -1, 1, 1, 2, 0, 1, 3, 2, 3, 3, 2, 2, 4, 3, 2, 0, 0, 0, 0, -1, -2, 0, 1, 1, 0, 0, -2, 1, 0, 0, 1, 2, 4, 4, 3, 4, 4, 4, 3, 1, 1, 0, 2, 2, 0, 0, 0, -1, 1, 0, 0, 0, -2, 1, 0, 1, 0, 3, 3, 3, 4, 3, 4, 4, 4, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 2, 0, 0, -2, 0, 1, 0, 2, 3, 4, 4, 6, 6, 3, 4, 3, 2, 0, 0, 2, 2, 0, 0, -2, 0, 0, 0, 1, -1, -2, 2, 1, 1, 1, 3, 5, 7, 5, 6, 6, 6, 4, 3, 1, 0, 2, 2, 0, -1, 0, 0, 1, 0, 0, -2, -3, 2, 0, 1, 2, 3, 5, 5, 4, 6, 5, 3, 3, 1, 1, 1, 3, 1, 1, 0, 0, 1, 1, 0, 0, 0, -4, 1, 1, 0, 2, 3, 3, 3, 3, 4, 6, 4, 3, 2, 2, 1, 3, 2, 2, 1, 1, 0, 0, 0, -1, -3, -5, 2, 2, 0, 0, 2, 3, 4, 3, 4, 3, 2, 2, 2, 2, 0, 1, 2, 2, 1, 0, 1, 0, 0, -2, -2, -4, 2, 0, 0, 0, 0, 1, 2, 4, 3, 3, 2, 2, 1, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, -3, -5, 0, 0, 0, 0, 0, 0, 1, 3, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -4, 1, 1, 1, 0, 0, 1, 1, 1, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -2, -1, -2, 0, -2, -4, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, -1, -1, -1, -2, -1, -3, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 0, -1, 0, -1, -2, -2, -1, 0, -1, -2, -2, -4, -4, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, 1, 0, 0, -2, -2, -2, 0, -1, -2, -2, -1, -2, -3, -4, 1, 0, 0, -1, 1, 0, 0, -1, -2, -1, -1, 0, 0, 0, -1, -3, -1, -2, -2, -1, 0, 0, -1, -2, -2, -3, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -2, -3, -4, -3, 0, 0, -1, -1, 0, -1, -3, -4, -4, 1, 0, 0, 0, 0, 0, 0, -2, -3, -2, -4, -2, -5, -4, -4, -2, -1, -1, -1, 0, -1, 0, 0, -2, -4, -4, 0, 0, 0, 0, 0, -1, -1, -3, -3, -4, -4, -6, -6, -5, -4, -3, -1, 0, 0, 0, -1, 0, -3, -3, -4, -5, -2, -2, 0, 0, -1, -1, 0, 0, -1, 1, 0, 2, 1, 3, 3, 4, 3, 4, 4, 4, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 2, 2, 3, 3, 4, 4, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -2, 0, -1, 1, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 1, 2, 0, 0, 0, 1, -2, -1, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, -2, 0, -1, 0, 0, 1, 2, 1, 1, 0, -1, -1, -1, 0, 0, 2, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 1, 1, 2, 0, 1, 1, -1, 0, 0, 0, 0, 1, 2, 0, 0, 0, -1, 0, 1, 1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, 2, 0, 1, 0, -1, 0, -1, 0, 2, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 2, 2, 0, 0, 0, 3, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 1, 1, 2, 0, 0, 2, 2, 1, 2, 1, 2, 1, 0, 0, 0, -1, 0, -2, -2, -1, 0, 0, 0, 0, 2, 2, 0, 2, 3, 0, 1, 2, 1, 2, 2, 0, 1, 0, 0, 0, 0, -1, -1, -2, -2, -1, -2, -1, 0, 1, 0, 0, 2, 3, 4, -1, 0, 1, 1, 2, 2, 0, 2, 0, 0, 0, -1, 0, 0, -2, -1, -3, -3, -2, 0, 0, 1, 1, 2, 2, 2, 0, 0, 1, 0, 1, 0, 1, 1, 0, -2, 0, -1, 0, -1, -2, -2, -3, -2, -2, 0, 0, 0, 1, 2, 3, 3, 0, 0, 0, 1, 1, 0, 1, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, -3, -2, 0, 0, 2, 0, 1, 1, 2, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -2, 0, 1, 0, 0, 0, 0, 2, 0, -1, 0, 1, 0, 0, 2, 0, 0, 0, -1, 1, 0, -1, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, -1, -1, 0, -1, -1, -1, -1, 0, 0, 1, 0, -1, 1, -1, 0, 1, 0, 0, 0, 0, 1, 0, 2, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, 1, 1, 0, 0, -1, 1, -2, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 2, 2, 2, 2, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 2, 0, 2, 2, 2, 2, 3, 2, 2, 0, 1, -1, 0, -1, -3, -2, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 2, 3, 4, 2, 1, 0, 2, 1, 0, -1, -1, -5, -4, -5, -5, -4, -4, -4, -3, -3, -4, -4, -3, -3, -5, -3, -1, 0, 0, 2, 1, 1, 1, 3, 2, 3, 3, -4, -3, -4, -2, -3, -3, -3, -2, -3, -2, -3, -3, -2, -3, -1, -1, 0, 0, 1, 2, 3, 2, 2, 0, 1, 3, -5, -4, -4, -3, -2, -4, -4, -3, -3, -2, -3, -3, -2, -2, -2, 0, 1, 0, 1, 2, 1, 2, 0, 1, 0, 2, -4, -4, -2, -3, -2, -2, -2, -2, -2, -1, -2, -2, -2, -1, 0, 0, 1, 1, 2, 1, 2, 0, 2, 2, 2, 2, -4, -4, -2, -2, -1, -2, -1, -2, -1, -2, -2, -1, -3, -1, -2, -2, 0, 1, 1, 2, 3, 2, 1, 0, 2, 0, -5, -2, -1, -3, -1, -2, -1, -1, -1, -1, -2, -3, -1, -3, -1, -2, -1, 2, 1, 1, 2, 1, 1, 1, 1, 1, -3, -3, -3, -1, -3, -1, -3, -1, 0, -1, -1, -3, -3, -1, -1, -1, 0, 0, 1, 0, 1, 2, 1, 1, 0, 1, -4, -2, -3, -2, -1, -2, -3, -2, -2, -3, -2, -1, -3, -1, -3, -1, 0, 0, 2, 0, 0, 1, 0, 1, 1, 0, -3, -3, -1, -3, -2, -2, -2, -3, -2, -2, -1, -1, -2, -2, -1, -1, 0, 1, 0, 0, 2, 1, 1, 0, 1, 0, -2, -1, -1, -1, -3, -3, -1, -3, -2, -1, 0, 0, -1, -2, -2, -1, 0, 0, 2, 2, 0, 1, 0, 1, 2, 1, -3, -1, -1, -2, -3, -1, -2, -2, -2, -2, 0, 0, 0, 0, 0, -2, -1, 1, 0, 0, 2, 0, 1, 0, 2, 1, -2, -2, -1, -3, -2, -3, -1, -1, -1, -1, -1, -1, -1, -1, -2, -2, 0, 1, 2, 3, 1, 0, 0, 0, 2, 1, -2, -1, -3, -3, -1, -1, -2, -1, 0, -2, 0, -1, 0, -2, 0, -1, -1, 0, 1, 1, 0, 1, 0, 1, 1, 2, -4, -2, -2, -1, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, -3, -1, -3, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, -4, -2, -2, -2, -2, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -2, -2, -3, -2, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 2, 1, 0, 0, 0, 0, 0, 1, -2, -2, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, -3, -3, -3, -1, -2, -2, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 1, 2, 3, 0, 0, 0, 1, 0, -2, -3, -2, -2, -1, -2, -1, -1, 0, -1, -1, -2, -1, -1, 0, 0, 1, 1, 0, 1, 2, 0, 0, 1, 1, 2, -3, -3, -2, -1, 0, -2, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 2, 2, 0, 0, 0, 1, 2, -2, -2, -2, -2, -2, -2, -3, -1, -2, -2, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 2, 2, 2, 1, 2, 2, -2, -3, -2, -2, -3, -3, -1, -2, -2, -1, -1, 0, -2, 0, 0, 0, 2, 0, 0, 2, 1, 2, 1, 1, 3, 0, -4, -4, -3, -3, -4, -3, -3, -1, -1, -3, 0, -1, 0, 0, -1, 0, 0, 0, 1, 2, 1, 2, 2, 2, 2, 1, -4, -3, -2, -4, -2, -3, -2, -2, -2, -2, -3, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 3, 3, 2, 2, -3, -3, -3, -4, -4, -4, -4, -4, -3, -3, -2, -3, -2, 0, 0, -1, 0, 1, 2, 2, 2, 2, 2, 2, 3, 3, 4, 3, 2, 1, 1, 1, -1, -3, -2, -3, -3, 0, -1, 1, 3, 4, 4, 6, 6, 7, 5, 5, 3, 3, 1, 0, 2, 3, 2, 2, 0, 0, -1, -3, -4, -3, -4, -2, -1, 0, 0, 2, 5, 6, 7, 6, 7, 5, 5, 3, 1, 1, 3, 1, 0, 1, 0, -1, -2, -2, -2, -3, -3, -2, -3, 0, 0, 2, 3, 4, 5, 4, 6, 5, 5, 3, 2, 1, 4, 1, 1, 1, 1, 0, 0, -1, -2, -2, -2, -2, -3, -1, 0, 1, 3, 3, 4, 5, 5, 3, 4, 2, 3, 1, 4, 2, 2, 2, 1, 0, 0, -1, 0, 0, 0, -2, 0, 0, -1, 1, 3, 3, 3, 3, 4, 2, 1, 2, 3, 4, 3, 2, 2, 2, 1, 0, 0, 0, 1, 0, 2, 1, 0, 0, -1, 1, 1, 3, 2, 2, 3, 1, 1, 3, 2, 3, 2, 0, 0, 2, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 1, 0, 2, 1, 1, 1, 1, 1, 1, 2, 4, 4, 2, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 3, 2, 2, 2, 2, 3, 3, 6, 4, 0, 0, 0, 0, 1, 2, 2, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 3, 4, 5, 5, 5, 0, 0, 1, 1, 1, 3, 3, 4, 2, 2, 3, 0, 0, 0, -2, 0, -2, 0, 1, 0, 3, 3, 5, 5, 7, 6, 0, 1, 0, 0, 2, 4, 4, 6, 6, 2, 2, 1, 0, -3, -3, -3, -3, -1, 0, 0, 1, 3, 5, 5, 7, 6, 0, 1, 1, 2, 3, 5, 6, 5, 6, 4, 1, 0, -1, -3, -4, -4, -2, -2, -1, 0, 1, 3, 6, 6, 6, 8, 0, 2, 2, 2, 3, 4, 6, 4, 4, 2, 0, 0, 0, -3, -3, -4, -4, -4, -1, 0, 2, 4, 6, 7, 7, 8, 2, 1, 3, 3, 3, 4, 4, 4, 3, 3, 1, -2, -2, -2, -5, -5, -4, -4, 0, -1, 0, 4, 5, 7, 6, 6, 1, 0, 0, 1, 2, 2, 2, 2, 2, 1, 0, -2, -3, -3, -3, -2, -3, -1, 0, 0, 1, 2, 5, 6, 6, 7, 1, 0, 1, 1, 2, 2, 1, 2, 0, 0, 0, -1, 0, -1, -3, -2, 0, 0, 1, 0, 1, 3, 5, 5, 6, 5, 0, -1, 0, 0, 2, 1, 2, 0, 0, -1, -2, -2, 0, 0, 0, -1, 0, 0, 2, 3, 4, 4, 5, 5, 5, 5, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 2, 3, 4, 3, 4, 6, 5, 5, 0, 0, -1, -1, 1, 0, 1, 1, 0, -1, -2, 0, 1, 1, 1, 0, 0, 2, 2, 2, 3, 3, 4, 6, 5, 5, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 2, 0, 1, 1, 1, 3, 3, 3, 3, 5, 5, 5, 5, 0, -1, -1, 0, 0, 0, 1, 1, -1, 0, 0, 0, 1, 0, 1, 0, 1, 2, 4, 5, 5, 4, 3, 3, 5, 5, 0, 0, -1, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, 1, 0, 2, 1, 2, 4, 4, 4, 5, 4, 5, 5, 5, 0, 0, 0, 0, 1, 2, 1, -1, -1, -2, -1, 0, 0, 1, 2, 1, 2, 3, 6, 6, 5, 5, 4, 3, 5, 2, 0, 0, 0, 1, 1, 1, 1, 0, -2, -2, -3, 0, 0, 0, 0, 2, 4, 3, 5, 7, 6, 5, 4, 4, 2, 2, 1, 0, 0, 1, 2, 2, 1, 0, -2, -2, -2, -1, 0, -1, 0, 1, 3, 5, 7, 7, 6, 5, 2, 3, 1, 2, 1, 0, 2, 1, 1, 3, 3, 0, 1, -1, -2, -2, 0, 0, 1, 0, 3, 6, 4, 6, 4, 4, 2, 2, 1, 0,
    -- filter=0 channel=1
    0, 0, -1, -2, -1, 1, 0, 0, 0, 1, 3, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 2, 2, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 2, 3, 1, 0, 0, 1, 0, 1, 0, 2, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 3, 1, 2, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 3, 2, 3, 0, 0, 1, 0, 0, 0, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 3, 2, 2, 1, 1, 1, 1, 2, 0, 1, 0, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 3, 3, 2, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 2, 1, 0, 0, 0, 2, 1, 3, 2, 2, 3, 1, 2, 1, 0, 0, 0, 1, 0, 1, 1, 0, 2, 1, -1, 0, 0, 0, 0, 0, 0, 2, 1, 3, 4, 3, 4, 2, 2, 2, 0, 1, 0, 0, 1, 2, 0, 2, 0, 0, 1, 1, 0, -1, 0, 0, 0, 1, 2, 1, 2, 3, 3, 3, 3, 2, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, -1, 0, 0, 0, 0, 1, 2, 1, 1, 3, 4, 2, 4, 3, 1, 1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 4, 2, 2, 4, 4, 1, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, -1, 1, 1, 0, 2, 1, 2, 1, 4, 2, 4, 4, 1, 2, 1, 0, 0, 0, 0, 0, 0, 2, 2, 0, -1, -1, 1, 0, 2, 1, 2, 1, 1, 3, 2, 4, 5, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 1, 1, 2, 2, 2, 1, 3, 3, 3, 2, 3, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, -2, 0, 0, 0, 0, 1, 1, 3, 3, 2, 2, 4, 4, 3, 1, 0, 1, 0, 0, 1, 0, 1, 0, 3, 0, 1, 0, 0, 1, 0, 0, 2, 1, 2, 2, 2, 2, 2, 3, 3, 2, 1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, -1, 0, 1, 1, 0, 0, 1, 2, 2, 3, 3, 2, 1, 3, 2, 0, 0, -1, 0, 1, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 1, 1, 3, 1, 2, 3, 1, 3, 1, 1, 1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, -1, 1, 1, 0, 0, 0, 3, 2, 1, 2, 3, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 0, 0, 0, 0, 1, 0, 2, 2, 1, 1, 2, 2, 1, 2, 0, 1, 0, 1, 0, 0, 0, 1, 0, 2, 0, 0, 0, -1, 0, 0, 1, 0, 1, 2, 1, 3, 2, 2, 2, 1, 1, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 1, 1, 1, 1, 1, 1, 1, 2, 2, 3, 3, 2, 2, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 2, 2, 2, 1, 3, 1, 1, 2, 2, 0, 0, 2, 0, 2, 1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 1, 0, 3, 2, 1, 3, 2, 1, 1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 1, 2, 3, 2, 1, 0, 2, 0, 0, 2, 2, 2, 1, 2, 1, 1, 0, 0, -2, -2, -3, -1, 0, 0, 0, 0, 0, -2, -2, -2, -2, -2, -1, -2, 0, 0, 1, 0, 0, 0, 1, 1, 2, 2, -3, -1, -2, 0, 0, 1, 0, 0, 0, -2, -2, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 1, 0, -2, -1, -2, 0, 0, 0, 0, -1, -1, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 2, 0, 0, -1, 0, -2, -1, 0, 0, 0, 1, 0, 0, 1, 2, 2, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, -2, -2, -2, 0, 0, 0, 1, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 0, 0, -1, 0, -2, 0, -1, 0, 0, 1, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 2, 0, 3, 1, 0, 2, 1, 2, 0, -1, 0, -1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 1, 1, 3, 1, 1, 3, 2, 0, 1, 0, 1, 1, 0, 0, 0, 0, -2, -2, -2, 0, -1, 0, 0, 0, 0, 0, 2, 2, 2, 1, 2, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 2, 3, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -2, -1, -1, 0, 0, 1, 0, 0, 0, 0, 2, 2, 2, 3, 3, 1, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, -2, -1, 0, 1, 0, 1, -1, 0, 0, 0, 1, 1, 1, 1, 3, 1, 3, 2, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 2, 1, 1, -1, 0, -1, 1, 1, 1, 1, 1, 3, 3, 0, 0, 1, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 2, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 2, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -2, -1, -2, -1, 0, -1, 0, 1, 0, 0, 0, 2, 1, 1, 2, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 2, -2, -1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 2, 2, 1, 2, 0, 2, 1, 3, 1, 4, 3, 2, 3, 0, 0, -1, -2, -3, -3, -2, 0, -1, 0, 1, 1, 0, 2, 2, 0, 1, 0, 0, 0, 1, 3, 3, 4, 2, 1, 0, -2, -3, -3, -3, -3, -1, 0, -1, -1, 0, 0, 0, 1, 2, 1, 0, 0, 0, 3, 2, 3, 2, 3, 1, 0, 0, -2, -2, -2, -2, -3, 0, 0, -2, -2, -1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 3, 3, 2, 2, 2, 0, -1, -3, -2, -3, -2, -2, -2, 0, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -2, -2, -1, -2, -3, -3, -3, -1, 0, -1, -2, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, -1, -2, -1, -1, -3, -2, -1, -2, -1, 0, -1, -1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 2, 0, 1, 1, 1, 0, -1, -2, -1, -1, -2, -1, -2, -2, -1, -2, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 2, 0, 1, 1, 0, 0, -1, 0, -1, -2, -1, -2, -3, -1, -3, -4, -2, 1, 1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 2, 2, 0, 0, 0, 0, -1, -2, -2, -2, -2, -2, -3, -4, -2, 0, 2, 2, 0, -1, -1, -1, 0, 0, 0, 1, 1, 3, 1, 0, -2, 0, 0, -1, -1, -2, -4, -4, -4, -3, -2, 0, 1, 1, 0, -2, -2, -2, -1, 0, 1, 0, 0, 3, 2, 0, -1, -2, 0, 0, 0, -2, -2, -2, -2, -4, -2, 0, 3, 2, 0, -2, -2, -3, -1, 0, 0, 1, 2, 1, 1, -2, -1, -1, -1, 0, 0, -1, -2, -3, -4, -3, -2, -2, 4, 1, 0, -2, -2, -2, -1, 0, 0, 2, 2, 2, 0, -2, -3, 0, 0, 0, 0, -1, -2, -4, -3, -3, -3, -2, 3, 1, 0, -3, -3, -3, -2, 0, -1, 0, 2, 3, 0, -2, -3, -1, 0, -1, -1, -1, -3, -4, -3, -3, -2, 0, 1, 0, -1, -2, -4, -2, -1, -2, -1, 0, 0, 1, 0, 0, -2, -1, -2, -1, -1, 0, -4, -2, -3, -1, -1, 0, 1, 0, -1, -1, -2, -1, -3, -3, -1, -2, 1, 1, 0, 0, -2, 0, -1, -1, 0, 0, -3, -3, -1, -1, -2, 0, 2, 1, 0, 0, -1, 0, -2, -2, -1, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, -1, -2, -2, -2, -1, -1, 0, 1, 2, 1, 0, 0, 0, -1, -2, -1, 0, 1, 2, 0, 0, -1, -1, -1, -2, -1, -2, -2, -2, -3, -1, 0, 0, 2, 2, 1, 0, 0, 1, 1, -1, -1, 0, 3, 2, 0, 0, -1, 0, 0, -2, -2, -1, -2, -1, -3, -3, -2, -1, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, -1, -2, -1, -2, -3, -2, -3, -2, -1, -2, -1, -2, -1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 0, -1, 0, -1, -2, -2, -2, -1, -3, -1, -1, 0, -1, 0, 2, 0, 0, 0, 0, 2, 2, 0, 0, 1, 0, 0, 0, -2, -3, -3, -3, -3, -3, -1, -3, -3, -1, 0, -1, -1, 1, 0, 2, 0, 1, 2, 3, 3, 0, 1, 1, 0, -1, -1, -3, -1, -2, -1, -1, -1, -4, -2, -1, -1, 0, 0, 1, 1, 0, 1, 1, 3, 3, 2, 2, 0, 1, 1, 0, -2, -1, -1, -1, -1, -2, -3, -2, -2, -1, 0, 0, 0, 2, 0, 1, 1, 2, 4, 3, 3, 3, 2, 2, 2, 0, -2, -2, -1, 0, -2, -3, -3, -1, 0, 0, 1, 0, 0, 2, 1, 1, 1, 1, 3, 4, 1, 3, 3, 2, 2, 1, -1, -1, -2, -1, 0, -2, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, -1, -1, -2, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, -1, -1, 0, 0, 0, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, -2, 0, -1, -1, 0, -2, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, -2, 0, -2, 0, -1, 0, 1, 0, 0, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, -1, -1, -2, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, -2, -2, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -3, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -2, -2, -1, -2, 0, -1, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, -2, 0, -1, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, -1, -3, -2, -1, -2, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -3, -3, -2, -2, -2, -2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -2, -3, -1, -1, 0, 0, 0, 0, 1, 0, -1, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -3, -1, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, -3, -1, -3, -1, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 2, 0, 1, 1, 1, 1, 1, 2, 3, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 2, 1, 1, 2, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, 0, -2, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -2, -2, -2, -2, 0, 0, 0, -1, 0, -1, -1, -2, 0, -3, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, -2, -2, -2, -3, -1, 0, -2, -1, -1, -1, 0, -2, -2, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -2, -1, -4, -2, -2, -1, 0, -1, -1, -1, -2, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -3, -2, -3, -1, -1, -1, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, -1, -1, -1, -2, -1, -3, -2, -2, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, -2, -2, -3, -3, -3, -2, -2, -2, -3, -3, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, -1, -2, -1, -2, -3, -3, -2, -2, -3, -2, -3, 0, -2, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, -2, -1, -2, -3, -3, -2, -2, -2, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -3, -3, -2, -1, -1, -1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -2, 0, 0, -1, 0, -1, -1, -1, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, 0, -2, -2, -1, -2, -2, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -2, -1, -2, -1, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -2, -2, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -2, -1, -1, -2, -3, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, -1, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, -3, -1, 0, -2, -1, -1, -1, -1, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -3, -2, 0, -2, -3, -1, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, -2, -1, -1, -3, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -3, -2, -2, -3, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 1, 0, 0, 0, 0, 0, 0, -2, -1, -2, -2, -2, -1, -1, -2, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -2, 0, -1, -2, -2, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, -2, -1, 0, -1, 0, 0, 0, 2, 2, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -2, 2, 1, 2, 0, 2, 2, 1, 1, 0, 1, 0, 1, 0, -1, -1, -2, -1, -1, -1, 0, 0, -2, -1, -2, -2, -1, 1, 2, 1, 1, 2, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, -2, -1, 0, -1, -1, 0, 0, -2, -2, -1, 2, 2, 1, 2, 2, 0, 0, 0, 2, 3, 2, 2, 1, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -2, -1, 3, 1, 0, 2, 2, 1, 0, 0, 1, 2, 3, 2, 1, 1, 2, 2, 0, 0, 1, 2, 1, 1, 0, 0, -1, -2, 1, 1, 2, 0, 0, 1, 0, 0, 0, 3, 2, 3, 2, 1, 1, 1, 1, 2, 1, 0, 2, 0, 0, 0, 0, -1, 3, 1, 0, 0, 1, 0, 1, 0, 0, 2, 3, 1, 3, 3, 2, 2, 1, 1, 2, 2, 1, 0, 1, 0, 0, 0, 3, 1, 0, 1, 1, 0, 0, 0, 1, 0, 1, 2, 3, 1, 2, 3, 2, 2, 0, 2, 0, 0, 0, -1, -2, -1, 1, 1, 0, 1, 0, 0, -1, 0, 1, 2, 1, 2, 3, 1, 4, 4, 2, 1, 1, 1, 0, 0, 0, 0, -1, -1, 2, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 3, 3, 2, 2, 2, 3, 1, 1, 1, 2, 0, 0, 0, -1, -2, 1, 1, 1, -1, 0, -1, 0, -1, -1, 1, 1, 2, 2, 3, 3, 1, 2, 1, 2, 2, 2, 0, 0, 0, -2, -1, 1, 1, 1, 0, -1, -1, -3, -1, -1, 1, 1, 2, 2, 3, 2, 2, 2, 3, 1, 2, 0, 0, 0, -2, -1, -3, 2, 0, 0, 0, 0, -3, -2, -1, 0, 0, 2, 3, 4, 4, 2, 2, 2, 2, 1, 1, 1, 0, 0, -1, -2, -2, 1, 0, 0, 0, -1, -2, -2, -3, 0, 0, 2, 3, 4, 3, 3, 2, 0, 3, 3, 1, 0, 0, 0, -2, -2, -3, 1, 0, 1, -1, -1, -2, -1, -1, 0, 0, 3, 2, 4, 3, 2, 2, 0, 2, 3, 1, 0, -1, -3, -3, -3, -1, 0, 0, 0, 0, 0, -2, -2, -1, -1, 0, 1, 3, 4, 4, 2, 1, 2, 1, 1, 2, 0, 0, -2, -1, -1, -1, 1, 0, 0, 0, -1, -2, -1, -3, 0, 1, 2, 3, 3, 4, 3, 3, 1, 2, 2, 2, 0, -1, -2, -2, -1, -2, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 3, 2, 4, 4, 2, 3, 2, 3, 2, 2, 2, 0, 0, -2, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 4, 3, 6, 3, 3, 3, 4, 4, 4, 2, 0, 0, -1, 0, -2, -1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 2, 3, 5, 6, 4, 3, 3, 3, 5, 3, 2, 1, 0, 0, -1, -1, -2, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 3, 4, 7, 5, 5, 2, 3, 4, 2, 2, 1, 0, -1, 0, -2, -1, 0, 2, 1, 1, 0, -1, 0, 0, 0, 0, 3, 4, 4, 4, 5, 3, 3, 1, 1, 2, 0, -1, 0, 0, -1, -1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 3, 2, 3, 3, 3, 3, 1, 1, 2, 0, 0, -1, -2, -2, -3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 2, 2, 0, 2, 0, 2, 0, 0, 0, -2, 0, -2, -2, 0, 0, 0, 0, -1, 0, 2, 1, 2, 2, 1, 0, 2, 1, 1, 1, 0, 0, 1, -1, -2, -1, -2, -1, -3, -2, 1, 0, 0, 0, 0, 1, 0, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -2, -2, -2, -1, 0, 1, 1, 0, 1, 0, 1, 2, 1, 1, 0, 0, 0, -1, 0, -2, 0, 0, -1, -1, -2, 0, -1, 0, 0, -2, 2, 3, 4, 3, 4, 4, 5, 6, 5, 3, 5, 2, 2, 0, -2, -1, -1, -1, -2, -2, 0, 1, 1, 3, 7, 8, 3, 4, 4, 2, 2, 3, 4, 6, 5, 5, 4, 4, 2, -1, -4, -4, -2, -3, -3, -2, 0, 0, -2, 1, 3, 5, 2, 2, 2, 3, 0, 0, 2, 4, 6, 4, 5, 6, 2, -1, -5, -6, -4, -4, -3, -2, -1, 1, -1, 0, 2, 6, 1, 2, 0, 0, 0, 0, 1, 2, 5, 5, 5, 6, 4, 0, -1, -5, -4, -4, -4, -2, 0, 1, 1, 1, 1, 5, 0, 0, 1, 0, -1, -1, -1, 2, 4, 6, 6, 7, 3, 1, 0, -1, -4, -2, -2, -1, 0, 1, 2, 1, 2, 4, 1, 0, 0, -1, 0, -2, -2, 0, 3, 4, 4, 5, 5, 2, 0, -1, -3, -3, -1, -1, 0, 1, 1, 1, 0, 3, 2, 1, 0, 1, -2, -3, -3, -1, 1, 4, 4, 6, 4, 2, 0, -1, 0, -2, -1, -2, -1, 0, 1, 0, 0, 3, 4, 2, 2, 0, -1, -3, -3, -2, 0, 3, 4, 4, 6, 2, 2, 0, 1, 0, 0, -1, -3, -2, 0, 0, -1, 0, 3, 2, 2, 0, -1, -3, -2, -3, 0, 1, 4, 3, 4, 4, 3, 3, 0, 0, 0, -1, -3, -2, -2, -1, 0, 0, 4, 2, 1, 1, -1, -4, -2, -2, 0, 1, 3, 3, 3, 4, 4, 2, 1, 0, 0, -2, -2, -3, -3, -1, -1, 0, 3, 1, 2, 0, -3, -5, -6, -4, 0, 0, 4, 4, 4, 4, 1, 2, 0, 1, 0, -1, -3, -2, -3, -1, 0, -1, 0, 0, 2, -1, -3, -7, -7, -5, -2, 1, 3, 4, 4, 4, 2, 1, 0, 0, -1, -2, -3, -2, -4, -3, 0, 0, 0, 0, 0, 0, -5, -7, -8, -5, -2, 0, 2, 5, 4, 3, 1, -1, -1, -2, -1, -2, -2, -3, -3, -3, 0, 0, 3, 2, 0, -1, -3, -6, -5, -4, -2, 0, 2, 5, 5, 4, 2, 0, 0, -2, -3, -1, -4, -4, -5, -3, -1, -1, 1, 0, 0, -2, -3, -5, -5, -7, -4, -1, 2, 4, 6, 3, 2, 1, 0, -1, -1, -2, -4, -6, -6, -3, -1, 0, 2, 0, 0, -2, -4, -3, -5, -4, -3, -1, 2, 5, 4, 4, 4, 2, 0, 0, 0, -2, -3, -5, -5, -2, -2, 0, 4, 2, 0, -3, -2, -3, -4, -5, -4, 0, 3, 6, 5, 2, 3, 2, 0, 0, 0, -2, -2, -3, -3, -2, 0, 1, 2, 2, -1, -1, -2, -4, -2, -3, -1, 0, 2, 6, 3, 3, 4, 2, 0, 0, -2, -2, -3, -3, -3, 0, 0, 3, 3, 2, 0, 0, -2, -1, -2, -1, -1, 0, 4, 5, 3, 4, 1, 0, 1, 0, -2, -2, -2, -1, -1, 1, 2, 5, 5, 3, 2, 0, -2, -2, -1, -1, 0, 1, 4, 7, 5, 4, 2, 0, -1, -1, -2, -1, -1, -1, 0, 1, 4, 4, 3, 3, 1, 1, -1, -1, 0, 0, 0, 1, 3, 6, 5, 3, 1, 0, 0, -1, -2, -3, -1, -1, -1, 0, 4, 4, 3, 2, 0, 1, -1, 0, 0, 0, 1, 2, 4, 4, 3, 3, -2, -1, -4, -2, -4, -3, -2, -1, -2, 0, 4, 6, 0, 0, 0, 0, -2, 0, 0, 1, 2, 2, 4, 3, 2, 1, -1, -3, -3, -4, -3, -2, -1, -2, -3, 0, 3, 5, 1, -1, -1, 0, -2, -1, 2, 1, 2, 3, 4, 5, 2, 0, -4, -4, -5, -4, -3, -2, -3, -2, -1, 0, 2, 6, 0, -1, 0, 0, -1, 0, 3, 2, 2, 4, 3, 5, 1, -1, -4, -5, -4, -5, -2, -2, -2, -3, -1, 0, 3, 5, 1, 1, 0, 0, 0, 2, 3, 2, 2, 2, 4, 4, 2, 0, -2, -5, -4, -3, -1, 0, -1, -1, -2, 0, 2, 7, -7, -4, 0, 4, 5, 6, 5, 4, 2, 1, 0, -4, -5, -6, -6, -4, -1, 0, -1, 0, 0, 0, 2, 1, 4, 6, -5, -2, 0, 3, 4, 2, 3, 2, 2, 1, 0, -1, -2, -1, -2, -1, -2, 0, 1, 0, -1, 0, 0, 0, 1, 3, -3, -3, -1, 1, 1, 3, 2, 2, 3, 1, 1, 0, 0, -1, -1, -1, -2, 1, 1, 0, 0, 0, -1, 0, 0, 3, -2, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 1, 2, 2, 1, 1, 1, 1, 2, 0, 1, 1, 0, 1, 2, 1, 0, 0, 1, 0, 1, 0, -1, -1, 1, 1, 3, 3, 2, 2, 1, 3, 2, 1, 2, 1, 0, 0, 0, 0, 0, 2, 1, 3, 2, 1, 0, 0, -2, -2, 0, 0, 2, 2, 3, 2, 3, 4, 1, 2, 0, 1, 0, -1, 0, 0, 0, 2, 4, 4, 1, 1, 0, 0, -3, -3, 0, 0, 0, 0, 0, 1, 3, 2, 0, 0, 1, 1, -1, -2, -1, -1, 0, 0, 3, 4, 2, 2, 0, -2, -2, -2, 0, 2, 1, 0, 2, 2, 3, 1, 0, 0, 1, 1, 0, -1, -1, -1, 0, 1, 4, 3, 1, 1, 0, 0, -1, 0, 0, 2, 0, 0, 0, 3, 3, 2, 3, 3, 0, 0, 0, -2, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 2, 3, 0, 1, 1, 3, 4, 3, 3, 1, 0, 0, 0, -1, -3, -2, 0, -1, 0, -1, 0, 0, 0, 1, 1, 3, 5, 3, 2, 2, 3, 3, 4, 3, 1, 2, 1, 0, -2, -2, -2, -2, -1, -2, -3, 0, 0, 2, 1, 3, 1, 4, 5, 4, 5, 4, 2, 2, 3, 2, 0, 0, 0, 0, -1, -3, -3, -1, 0, -3, 0, -1, 0, 2, 3, 1, 1, 3, 4, 6, 5, 2, 2, 3, 1, 1, 0, 0, 0, -2, -2, -1, -2, -1, 0, -1, 0, 0, 0, 2, 2, 1, 2, 2, 5, 3, 4, 2, 1, 2, 1, 1, 1, 1, 0, -2, -1, -2, -1, -1, 0, -1, 1, 1, 1, 0, 0, 0, 0, 0, 3, 3, 2, 3, 2, 2, 3, 4, 3, 1, 0, 0, 0, -1, -1, -3, -1, -2, 1, 1, 2, 2, 0, 0, 0, 0, 2, 2, 2, 1, 2, 1, 3, 3, 2, 2, 0, 0, 0, 0, -3, -2, 0, -2, 0, 2, 3, 1, 0, 0, -1, 0, 0, 1, 0, 2, 0, 2, 2, 4, 2, 2, 2, 0, 0, 0, -2, -1, 0, 0, 0, 1, 1, 1, 0, -2, 0, 0, 0, 0, 1, 2, 1, 0, 3, 4, 4, 3, 1, 2, 0, 0, 0, 0, 2, -1, 0, 2, 2, 0, -1, -3, -4, -1, 0, -1, 0, 1, 1, 2, 3, 4, 4, 3, 2, 1, 0, -2, -1, 0, 3, 0, 0, 2, 1, 1, -2, -5, -4, -3, -3, -2, 0, 1, 1, 1, 3, 4, 5, 3, 2, 0, 0, 0, 0, 1, 2, 0, 0, 2, 0, 0, -3, -4, -4, -5, -2, 0, 0, 1, 3, 3, 4, 4, 4, 1, 0, 0, 0, -1, 0, 2, 3, 0, 1, 1, 0, 0, 0, -2, -2, -2, 0, 0, 1, 1, 4, 3, 4, 2, 1, 0, 0, -1, -1, 0, 1, 2, 5, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 2, 3, 3, 1, 0, 0, 0, 0, -1, 0, 0, 1, 6, 0, 0, 0, 0, 0, -1, 1, 0, 2, 0, 1, 1, 0, 1, 1, 0, 0, 0, -1, -2, -2, 0, -3, -2, 0, 4, -2, 0, 0, 0, 0, 0, 1, 2, 3, 1, 1, 0, 0, -1, 0, -1, -1, -2, -3, -2, -1, -3, -2, -2, 0, 4, -2, -1, 0, 0, 0, 1, 1, 3, 2, 1, 0, -2, -3, -2, -3, -4, -2, -2, -1, -1, 0, 0, -1, -1, 0, 3, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 2, 0, 1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 1, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, -1, 1, 1, 1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, -1, 0, 1, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -2, -2, -1, -2, 0, -1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, -1, 0, -1, -2, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -7, -4, -1, 3, 5, 7, 6, 5, 3, 1, -1, -4, -5, -4, -4, -3, -2, 0, 0, -1, -1, 1, 3, 5, 8, 10, -5, -3, -1, 1, 3, 3, 3, 3, 0, 1, 0, -3, -2, -3, -3, -3, -2, 0, 0, 0, -2, -1, 0, 1, 2, 6, -4, -3, 0, 2, 2, 1, 2, 1, 2, 1, 1, 0, -1, 0, -2, -3, -1, -1, 0, -1, -2, -1, -2, 0, 1, 5, -3, -2, 0, 0, 1, 0, -1, 0, 1, 1, 2, 1, 2, 2, 0, -1, -2, 0, -1, 0, -1, 0, -2, 0, 1, 4, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, 1, 3, 3, 2, 1, 1, 1, 1, 0, -1, -2, -1, -1, 0, 2, 4, 2, 1, 1, 1, -1, -2, -4, -2, -1, 0, 0, 2, 2, 4, 2, 2, 1, 1, 0, -1, -2, -2, -2, -1, 0, 4, 4, 3, 3, 0, 0, -4, -3, -3, -2, 0, 0, 3, 2, 4, 2, 1, 0, 0, -1, -1, -2, -2, -3, 0, -1, 3, 5, 4, 4, 1, 0, -2, -4, -4, -2, 0, 0, 1, 3, 2, 2, 1, 0, 0, -2, -1, -1, -4, -4, -1, -2, 2, 5, 3, 1, 1, 0, -3, -3, -3, 0, 0, 1, 1, 1, 1, 1, 3, 1, 0, 0, 0, -1, -4, -5, -3, -1, 1, 3, 3, 0, 0, 0, -2, -2, -1, 0, 1, 2, 2, 2, 3, 3, 2, 4, 2, 1, 1, -1, -2, -3, -3, -1, 1, -1, 1, 1, -1, 0, 0, 0, 1, 2, 3, 3, 4, 2, 3, 3, 4, 3, 1, 1, 0, -1, -1, -2, -2, -2, 0, -2, -1, -1, 0, 0, 0, 0, 1, 1, 3, 5, 5, 5, 3, 2, 1, 1, 0, 0, 0, -3, -3, -4, -2, -3, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 3, 5, 4, 5, 4, 3, 0, -1, -2, -1, -1, -1, -2, -4, -3, -2, -2, -1, 0, 0, 0, 1, 0, 0, 0, 1, 3, 3, 5, 3, 2, 3, 2, 0, 0, -2, -2, -2, -1, -2, -4, -2, 0, -2, 0, 1, 0, 1, 0, -1, 0, 0, 3, 3, 3, 2, 2, 1, 2, 2, 2, 0, -1, -2, -2, -2, -3, -3, 0, -1, 1, 1, 1, 0, 0, -1, -1, 0, 2, 4, 2, 2, 1, 2, 2, 1, 2, 1, 0, -2, -2, -3, -2, -1, 0, 0, 1, 2, 1, 0, 0, -2, -1, 0, 0, 2, 2, 2, 2, 0, 2, 1, 1, 1, 1, 0, -1, -3, -3, -1, 1, 0, 1, 1, 2, 0, -2, -2, -2, 0, 0, 1, 0, 2, 0, 0, 1, 2, 2, 1, 0, 0, -2, -3, -2, -1, 3, 0, 2, 1, 1, 0, -3, -4, -3, -2, -1, -1, 1, 0, 0, 1, 1, 1, 2, 0, 0, 0, -1, -2, -1, 1, 5, 2, 2, 3, 2, -2, -3, -5, -7, -4, -2, -1, -1, -1, 1, 0, 2, 1, 1, 1, 1, 0, -1, -2, -1, 2, 7, 0, 2, 1, 1, -1, -4, -6, -5, -4, -1, 0, 0, 1, 2, 2, 2, 2, 2, 0, -1, -1, -2, -1, 0, 3, 7, 1, 0, 1, 0, 0, -3, -3, -4, -1, 0, 0, 1, 3, 1, 2, 3, 2, 0, -1, 0, -1, -2, -1, 1, 5, 10, 0, 0, 0, 0, -1, -2, -1, 0, 0, 2, 1, 3, 2, 1, 0, 1, -1, 0, -1, -3, -3, -2, -1, 0, 5, 10, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 1, 2, 2, 0, 0, 0, -3, -3, -2, -1, -2, -1, 1, 4, 10, -1, 0, 1, -1, -1, 0, 1, 1, 2, 0, 0, 0, 1, 0, 0, -1, -1, -3, -4, -3, -3, -1, -2, 0, 3, 9, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, -1, -1, -1, -1, -3, -2, -2, 0, -1, -1, -1, 1, 5, 11, 2, 3, 1, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 1, 3, 2, 4, 2, 3, 1, 2, 2, 1, 1, 1, 1, 1, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 1, 1, 2, 3, 4, 2, 1, 0, 2, 2, 2, 2, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 0, 2, 2, 0, 2, 2, 2, 4, 3, 2, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 1, 1, 2, 2, 3, 1, 1, 3, 3, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 2, 1, 1, 2, 2, 0, 2, 2, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 2, 3, 3, 3, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 1, 3, 4, 2, 3, 2, 2, 3, 3, 2, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 2, 2, 2, 1, 1, 1, 3, 3, 4, 2, 3, 2, 3, 2, 0, 0, 1, 0, 0, 0, -1, 0, -1, -2, -2, 0, 1, 1, 1, 3, 2, 1, 2, 2, 1, 3, 3, 3, 3, 3, 1, 2, 1, 0, 0, 0, 0, -1, -2, -1, 0, 0, 1, 1, 0, 3, 2, 1, 2, 2, 1, 3, 4, 3, 3, 3, 1, 1, 1, 0, -1, 0, 0, -1, -1, 0, -1, 0, 1, 1, 0, 1, 1, 0, 2, 2, 1, 2, 2, 4, 3, 4, 3, 1, 0, -1, -1, 0, 0, 0, -2, -1, -1, 0, -1, 0, 2, 2, 1, 2, 2, 2, 1, 2, 2, 4, 4, 3, 3, 0, 0, 0, 0, -2, -2, 0, -2, -2, 0, 0, 0, 1, 3, 1, 2, 0, 2, 1, 1, 1, 1, 2, 3, 3, 1, 0, 0, -1, 0, 0, -2, -1, -3, -2, 0, 0, 0, 2, 1, 1, 0, 0, 1, 0, 2, 2, 2, 1, 2, 3, 0, 0, 0, 0, 0, 0, -2, -2, -2, -1, -1, 0, 1, 1, 2, 2, 0, 1, 0, 1, 3, 1, 3, 2, 2, 2, 1, 1, 0, -1, -1, -1, -2, -2, -2, -2, -1, -1, 0, 1, 1, 1, 0, 1, 0, 2, 1, 2, 3, 4, 4, 3, 1, 0, 0, 0, 0, -1, -1, -2, 0, -2, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 2, 2, 3, 3, 2, 3, 2, 1, 0, 0, 1, 0, -1, -2, -1, -2, 0, 0, 2, 3, 1, 2, 0, 0, 0, 0, 1, 1, 1, 2, 2, 3, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 2, 4, 3, 2, 1, 1, 1, 0, 1, 3, 1, 3, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, -1, 0, 3, 2, 2, 2, 0, 0, 0, 0, 0, 2, 4, 3, 2, 0, 2, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 3, 2, 3, 2, 0, 1, 0, 0, 1, 3, 3, 3, 3, 0, 1, 1, 0, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 2, 2, 2, 1, 0, 0, 0, 0, 2, 2, 2, 2, 0, 2, 2, 2, 1, 0, 0, 0, 0, -2, -2, -1, 0, 0, 0, 2, 0, 0, 0, -1, -1, 1, 1, 3, 3, 0, 0, 2, 0, 2, 0, 0, 0, 0, -1, 0, -2, 0, -1, 0, 0, 1, 0, -1, -2, -2, 0, 2, 1, 1, 0, 2, -1, 1, 2, 2, 1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, -1, -1, -2, -2, 0, 1, 0, 0, 2, 0, 0, 1, 0, 3, 2, 2, 1, 1, 2, 0, 0, 0, -1, -1, -1, -2, 0, -1, -3, -2, -1, 0, 0, -1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -1, -3, -3, -2, -4, -3, 0, -1, -1, -2, 0, 0, 1, 3, -2, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, -2, -2, -2, -2, 0, -1, 0, 0, 0, 1, 2, -1, 0, 0, -1, -1, -1, 0, -2, 0, 0, 0, 1, 0, 1, -1, -2, -2, -1, 0, 0, 0, 0, 1, 0, 1, 2, 1, 0, 0, -1, 0, -2, -2, -1, -2, 1, 2, 3, 3, 2, 1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 2, 1, 2, 2, 1, 1, 0, -1, -3, -3, -1, 0, 1, 1, 3, 2, 2, 1, 0, 0, 0, -1, 0, 0, -1, 0, 2, 1, 1, 2, 1, 0, -1, -2, -3, -4, -2, 0, 0, 2, 1, 2, 1, 0, 0, -1, -1, -1, -1, -2, 0, -1, 0, 1, 1, 1, 2, 0, 0, -3, -3, -3, -4, -1, 0, 2, 1, 2, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, -2, -2, -3, -2, 0, 1, 0, 2, 2, 3, 3, 2, 1, 1, 0, 0, -2, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, -2, -3, 0, 0, 2, 1, 2, 2, 2, 2, 1, 2, 0, 0, 1, -2, -2, -3, -1, 0, 0, 0, 1, 0, 0, 0, -2, -1, 0, 0, 0, 2, 3, 2, 2, 1, 0, 0, 0, 0, 0, -2, -3, -2, -2, -1, 0, -1, 0, 0, 0, 0, -1, -2, -1, 0, 1, 4, 4, 4, 2, 1, 0, -1, -1, -2, 0, -2, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, 3, 4, 3, 3, 2, 1, 0, -1, -1, -1, -3, -2, -3, -3, -3, -2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 3, 3, 4, 2, 1, 1, 0, 0, 0, -1, 0, -1, -3, -3, -2, -1, 0, 1, 1, 2, 0, 1, 0, 0, 0, 1, 2, 3, 2, 1, 3, 1, 1, 0, 0, -1, -1, -1, -2, -4, -3, -1, 0, 0, 2, 0, 2, 1, 0, 0, 0, 0, 3, 3, 2, 3, 2, 1, 1, 0, 1, 0, 0, -2, -2, -2, -2, 0, 0, 2, 2, 0, 2, 0, 0, 0, -1, 1, 1, 1, 3, 2, 3, 1, 1, 0, 1, 0, -2, -1, -3, -2, -2, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 3, 1, 1, 1, 1, 1, 0, 0, -1, -1, -3, -3, 0, 1, 0, 1, 1, 1, 1, -1, -1, 0, -1, -1, 0, 1, 2, 1, 0, 2, 0, 0, 0, 0, -2, -1, 0, 0, 0, 2, 0, 1, 2, 0, 0, -1, -1, -1, -2, -1, 0, 0, 1, 0, 2, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 3, 0, 0, 1, 0, 0, -1, -2, -1, 0, 0, 1, 0, 1, 1, 0, 1, 0, -1, -1, -1, -3, -3, -2, 0, 0, 3, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 1, 1, 2, 1, 0, 1, 0, 0, -1, -1, -2, -3, -2, 0, 1, 4, 0, 1, 0, -1, -1, 0, 0, 1, 0, 2, 2, 1, 1, 0, 0, -1, -2, -3, -3, -2, -1, -2, -2, -1, 0, 3, 0, 0, 0, 0, -2, 0, 0, 0, 1, 2, 2, 2, 0, 0, 0, -2, -3, -4, -3, -3, -2, -2, -1, -2, 0, 4, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 1, 0, 0, 0, 0, -2, -1, -3, -4, -4, -3, -2, -1, -1, 0, 3, -1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, -1, -1, -2, -2, -2, -2, -1, 0, 0, 0, 1, 4, -2, -1, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, -2, -2, -1, 0, -1, 0, 0, 1, 0, 2, 3, 4, 4, 6, -2, -1, -1, 0, 0, 2, 3, 3, 2, 1, 1, 0, 0, -1, -1, -2, -1, 0, 0, 2, 0, 1, 2, 1, 3, 4, -1, 0, 0, 1, 2, 1, 1, 3, 2, 1, 0, 1, 0, 0, -2, -1, -3, -2, 0, 1, 1, 0, 0, 1, 1, 4, -2, 0, 0, 1, 1, 0, 1, 1, 2, 1, 2, 2, 1, 1, 1, 0, -1, -2, 0, 0, 0, 0, 1, 1, 2, 3, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 3, 3, 1, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 4, 3, 3, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 0, 1, 0, 0, 0, 0, -2, 0, 2, 3, 4, 2, 3, 3, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, 0, 0, 0, -2, -1, -1, 0, 2, 1, 4, 3, 4, 3, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 2, 1, 1, 0, 0, -2, -2, 0, 1, 1, 2, 4, 2, 3, 2, 2, 2, 1, 0, 0, -1, 0, -1, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 2, 2, 3, 4, 3, 4, 1, 1, 2, 0, 0, -1, 0, -2, -1, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 2, 3, 2, 2, 0, 0, -1, -1, -1, -1, -1, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 3, 3, 4, 4, 2, 4, 1, 0, 0, 0, 0, -2, -4, -2, -1, 0, -2, 0, -1, 0, 0, 1, 0, 0, 0, 2, 3, 3, 4, 4, 3, 4, 1, 0, -1, 0, 0, -2, -3, -2, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 2, 2, 4, 5, 4, 3, 3, 1, 0, -1, -1, -1, -2, -2, -2, -2, -1, -2, -1, 0, 0, 0, 0, -1, -1, 2, 3, 4, 4, 4, 3, 3, 2, 0, 0, -1, 0, -2, -1, -2, -3, -3, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 3, 5, 4, 3, 3, 3, 0, 0, 0, 0, -1, -3, -3, -4, -3, -1, -2, 0, 0, 0, 1, 0, -1, -1, 0, 1, 3, 4, 4, 2, 2, 3, 2, 0, 0, 0, -2, -2, -2, -4, -4, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 2, 2, 3, 3, 4, 1, 3, 0, 0, 0, 0, -1, -2, -3, -3, -3, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 3, 3, 2, 2, 3, 1, 0, 0, 1, 0, -2, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, -2, -3, -1, 0, 1, 3, 1, 3, 2, 3, 2, 0, 1, 0, -1, -3, -2, -1, 0, 2, 0, 1, 1, 2, 1, -1, -1, -2, 0, 1, 1, 2, 1, 2, 3, 3, 1, 0, 1, 0, -1, -2, -2, 0, 0, 3, 0, 1, 0, 0, 0, 0, -2, -2, -2, 0, 1, 2, 1, 1, 2, 1, 2, 0, -1, 0, -1, -3, -1, 0, 0, 1, -1, 0, 0, -1, 0, 0, 0, -2, -2, 0, 2, 2, 1, 3, 3, 2, 1, 0, -1, -1, -1, -2, -1, 0, 2, 2, -1, 0, -1, 0, -1, -1, -1, 0, -1, 0, 1, 1, 2, 0, 2, 0, 0, -1, -1, -1, -3, -2, 0, 0, 0, 3, -1, -1, 0, -2, -2, -1, -1, 0, 0, 1, 0, 1, 0, 1, -1, 0, -2, -3, -2, -2, -3, -2, 0, -1, 0, 3, -2, 0, -2, -2, -2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -2, -2, -2, -2, -1, -2, -2, 0, 0, 0, 3, -3, -2, -1, -1, -1, -1, -1, -1, 0, 0, 0, -2, -3, -3, -4, -2, -3, -3, -1, -2, 0, 0, 0, 0, 2, 5, -7, -5, -1, 0, 1, 0, -1, -1, -2, -5, -8, -9, -9, -7, -6, -7, -4, -4, -2, 0, -2, -2, -4, -1, -1, 1, -6, -4, -2, -1, 1, 0, 0, 0, -1, -4, -5, -5, -4, -5, -4, -4, -1, -2, 0, 0, -1, 0, -2, -1, -1, 0, -3, -2, 0, 0, 1, 0, 0, -2, -2, -1, -1, -1, 0, 0, 0, -1, 0, 1, 1, 0, -1, 0, -1, -1, 0, 1, -3, 0, 0, 1, 2, 1, 0, -1, 0, 0, 1, 3, 0, 0, 2, 2, 1, 1, 0, 1, 1, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 2, 4, 3, 3, 3, 5, 3, 2, 0, 0, 0, 0, -1, 0, 1, 2, 1, 0, 2, 1, 0, -1, -2, 0, 0, 2, 2, 3, 3, 3, 4, 4, 2, 1, 2, 0, 1, 0, 0, -1, 0, 0, 2, 2, 0, 0, -1, -1, -2, 0, 1, 3, 4, 4, 3, 3, 4, 2, 2, 1, 1, 2, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 2, 3, 3, 4, 4, 4, 4, 3, 3, 3, 0, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 2, 4, 5, 3, 6, 5, 4, 5, 4, 2, 0, 0, 0, 0, -2, -2, 0, -1, 0, -1, 0, 0, 1, 0, 2, 3, 4, 4, 5, 5, 5, 4, 3, 3, 2, 1, 0, 0, -3, -1, -3, -1, -2, -3, -1, 0, 0, 0, 2, 3, 1, 4, 6, 6, 6, 6, 6, 5, 3, 1, -1, 0, -2, -2, -3, -2, -3, -3, -1, -3, -3, -1, 1, 1, 2, 4, 4, 5, 6, 7, 6, 6, 7, 4, 1, 1, -1, -1, -2, -3, -2, -3, -2, -2, -2, -3, -2, 0, 1, 3, 3, 3, 3, 6, 5, 8, 6, 8, 6, 6, 1, 1, 0, -1, -1, -3, -2, -3, -1, -1, -1, -3, 0, 1, 3, 4, 2, 4, 4, 5, 6, 6, 6, 7, 4, 4, 3, 1, 0, 1, 0, 0, 0, -1, -2, -1, -1, -3, 0, 2, 3, 4, 2, 4, 5, 6, 6, 5, 5, 5, 4, 6, 5, 2, 2, 1, 0, 0, 0, -2, -1, -2, -1, -1, 0, 2, 4, 4, 1, 2, 4, 6, 5, 5, 5, 5, 5, 4, 5, 3, 1, 2, 1, 0, -1, -2, -3, -2, 0, -3, -1, 0, 3, 2, 1, 1, 3, 3, 3, 4, 4, 5, 5, 3, 5, 2, 4, 2, 0, 0, -1, -2, -3, -1, 0, -3, 0, 2, 1, 1, 0, 1, 1, 1, 2, 3, 5, 3, 2, 2, 3, 4, 4, 3, 1, 1, 0, -1, -1, 0, 1, -3, 0, 2, 2, 0, 0, 0, 0, 0, 3, 2, 2, 3, 2, 3, 4, 4, 4, 4, 2, 0, -1, -1, 0, -1, 2, -2, 0, 0, 0, 0, -1, -3, -1, 0, 2, 3, 2, 4, 3, 5, 5, 4, 4, 3, 0, 1, 0, -1, 0, 0, 2, -1, -1, 0, 0, 0, -1, -2, 0, 1, 2, 1, 4, 5, 4, 4, 5, 4, 1, 2, 0, -1, 0, 0, 0, 0, 4, -2, 0, -2, -1, 0, -1, -1, 0, 1, 2, 2, 2, 4, 4, 4, 2, 1, 1, 1, 0, 0, 0, -1, -1, 0, 3, -1, -1, -1, -1, -2, -1, 0, 0, 1, 1, 1, 1, 0, 2, 2, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, 3, -2, -2, -2, -2, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -4, -2, 0, 2, -2, -3, -3, -2, -2, -2, 0, 0, 0, -1, -2, -3, -4, -3, -1, 0, 0, -1, -2, -2, -3, -2, -4, -1, 0, 4, -3, -3, -4, -3, -3, -3, 0, 0, -1, -4, -5, -8, -9, -8, -6, -4, -3, -1, -2, -1, 0, 0, 0, 0, 2, 5, -1, 0, 2, 3, 5, 4, 4, 3, 2, 0, -2, -2, -2, -3, -3, -4, -2, -1, -1, -1, -1, -1, 1, 1, 4, 9, -1, 0, 0, 1, 2, 1, 0, 0, 2, 1, 0, 0, 0, -1, -2, -3, -4, -1, -2, -1, -3, 0, 0, 0, 2, 5, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 3, 1, 2, 0, -1, -1, -1, -3, -2, -2, -1, -1, 0, 1, 1, 4, 0, 0, 0, 0, 0, -1, -2, 0, 1, 3, 4, 3, 2, 1, 1, 0, -1, -1, -1, -3, -2, -2, 0, 0, 1, 4, 3, 0, 1, 0, -2, -3, -4, -1, 0, 3, 3, 4, 3, 3, 1, 0, 0, -1, -2, -2, -3, -1, -1, 0, 2, 3, 4, 3, 1, 0, -3, -4, -3, -2, 0, 2, 2, 3, 3, 2, 3, 0, -1, -1, -3, -2, -4, -4, -1, -1, 0, 1, 3, 2, 1, 0, -2, -4, -3, -2, -1, 1, 2, 4, 4, 2, 3, 0, 0, -1, -3, -4, -4, -5, -2, -1, 0, 2, 4, 2, 0, 0, -2, -3, -4, -2, 0, 0, 3, 3, 3, 2, 2, 1, 0, 0, -2, -4, -3, -5, -4, -3, 0, 2, 2, 0, 0, 0, -1, -2, -3, -2, 0, 1, 2, 2, 3, 1, 3, 2, 1, 1, 0, 0, -3, -2, -4, -4, 0, 0, 0, 0, 0, -1, -2, -2, -2, -2, 0, 1, 4, 3, 4, 3, 3, 2, 2, 0, 0, -1, -2, -3, -4, -3, -1, 0, 0, -2, -2, -3, -2, -4, -2, -2, 0, 1, 5, 5, 5, 3, 1, 1, 1, 0, 0, 0, -3, -3, -3, -4, -1, 0, -2, -2, -3, -2, -2, -3, -4, -1, 0, 1, 4, 6, 5, 3, 3, 1, 0, 0, 0, -2, -4, -3, -3, -2, -1, 0, -2, -1, -2, -2, -4, -3, -2, -2, 0, 3, 4, 4, 3, 3, 1, 1, 0, -2, -1, -2, -4, -4, -4, -2, -2, 0, 0, 0, 0, -1, -3, -4, -3, -2, 0, 2, 3, 4, 4, 3, 2, 2, 0, -1, -2, -3, -2, -3, -5, -3, -2, -1, -1, 0, -1, -1, -3, -3, -3, -1, -1, 2, 4, 4, 2, 3, 3, 2, 2, 0, 0, -2, -3, -3, -5, -3, -1, 0, 1, 0, 0, -1, -3, -4, -4, -3, 0, 0, 2, 3, 2, 1, 2, 3, 2, 0, 1, 0, -3, -4, -4, -3, -2, 1, 0, 1, -1, 0, -3, -2, -2, -2, 0, 1, 3, 3, 3, 0, 0, 2, 0, 1, 0, 0, -3, -3, -4, -2, 0, 2, 0, 0, 1, -2, -2, -4, -3, -3, 0, 0, 1, 2, 2, 1, 1, 1, 2, 2, 0, -1, -3, -3, -4, -1, 0, 2, 0, 2, 1, -1, -3, -4, -4, -4, -2, 0, 2, 1, 2, 1, 0, 1, 2, 0, 0, -1, -3, -2, -1, -1, 1, 4, 1, 2, 1, -1, -2, -5, -3, -2, -2, 0, 2, 3, 2, 1, 1, 1, 0, 0, 0, -1, -3, -2, -2, -1, 1, 5, 2, 0, 0, 0, -1, -3, -2, -2, 0, 1, 2, 2, 1, 2, 1, 1, -1, 0, -2, -2, -4, -2, -1, -1, 3, 6, 0, 0, -1, 0, 0, -2, -2, 0, 0, 2, 2, 2, 2, 3, 2, 0, 0, -2, -1, -2, -2, -2, -2, -1, 3, 5, 1, 0, -1, 0, -1, -1, 0, 1, 4, 3, 3, 2, 1, 0, 1, 0, -1, -3, -4, -4, -4, -3, -1, -1, 1, 5, 0, 1, -1, -1, -2, 0, 2, 2, 3, 5, 2, 3, 0, 1, -1, -3, -3, -3, -3, -3, -3, -3, -3, -2, 0, 6, 0, 1, 0, 0, 0, 0, 2, 3, 3, 2, 2, 1, 0, 0, -2, -2, -4, -5, -4, -4, -4, -2, -3, -2, 2, 5, 0, 0, 1, 1, 1, 2, 2, 4, 2, 1, 1, 0, -1, -1, -2, -2, -2, -1, -3, -1, -2, 0, 0, 0, 3, 7, -4, -4, -1, 0, -1, -1, -3, -3, -4, -5, -6, -5, -5, -7, -5, -5, -3, -3, -2, -3, -2, -1, -2, 0, 0, 1, -4, -2, -1, -1, 0, -1, -2, -1, -2, -2, -2, -3, -3, -4, -3, -2, -3, -1, 0, -1, -1, -1, -1, -1, -1, 1, -2, -2, -1, 0, 0, 0, 0, 0, -1, -1, -2, 0, -1, -1, -1, -2, 0, 0, 0, -1, -2, -1, 0, -1, 0, 0, -3, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 1, -2, -1, 0, 0, 0, -1, 0, 0, 2, 2, 3, 3, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 3, -1, 0, 0, 0, 0, 0, 0, 1, 2, 3, 3, 3, 3, 2, 1, 2, 3, 1, 2, 0, 0, -1, -1, 1, 1, 2, -1, 0, -1, 0, -2, 0, -1, 1, 1, 1, 5, 3, 4, 4, 4, 1, 2, 1, 1, 0, 0, 1, 0, 0, 1, 2, 0, -1, 0, -1, -2, 0, 0, 2, 3, 4, 3, 3, 5, 3, 4, 3, 1, 0, 1, 0, 0, 0, 0, 0, 1, 2, -2, -2, 0, -1, 0, 0, 0, 2, 2, 4, 5, 4, 5, 5, 3, 3, 2, 0, 1, 0, 0, 0, 0, -1, 0, 0, -4, -2, 0, 0, 0, 1, 0, 2, 2, 2, 5, 6, 4, 6, 5, 2, 1, 1, 0, -1, -1, -1, -2, -2, -1, 0, -4, -3, 0, 0, 1, 0, 2, 1, 2, 2, 5, 4, 6, 6, 4, 1, 1, 0, 0, -1, -1, -1, -3, -3, -1, -1, -3, -3, -1, 0, 0, 1, 1, 3, 2, 3, 4, 6, 7, 7, 3, 3, 0, -1, -2, -2, -1, -2, -1, -1, -1, 0, -3, -2, 0, 0, 3, 1, 3, 2, 3, 4, 6, 8, 6, 6, 5, 3, 1, -1, 0, -2, -1, -3, -1, -2, -1, 0, -5, -1, 0, 2, 0, 1, 2, 3, 6, 6, 6, 6, 6, 6, 6, 2, 1, 0, 0, -2, -2, -3, -1, -1, 0, 0, -3, -1, 0, 2, 2, 0, 2, 3, 4, 6, 6, 6, 5, 5, 6, 5, 1, 0, -1, -1, -2, -3, -2, -3, 0, 0, -3, -1, 0, 1, 1, 2, 1, 3, 4, 3, 4, 4, 3, 5, 4, 3, 2, 1, 0, 0, -2, -2, -3, -2, 0, 0, -3, -1, 0, 1, 1, 1, 2, 2, 2, 3, 3, 4, 3, 4, 4, 3, 2, 1, 0, 0, -1, -1, -3, -3, -2, 0, -3, -1, 0, 0, 0, 2, 1, 0, 2, 3, 4, 4, 4, 4, 4, 4, 3, 1, 1, 1, 0, -2, -3, -3, 0, 0, -4, 0, 0, -1, -1, 0, 0, 0, 2, 3, 3, 3, 3, 3, 3, 3, 2, 1, 2, 1, 0, -1, -2, -2, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 2, 3, 2, 4, 1, 2, 2, 2, 2, 2, 2, 0, 0, -1, -2, -1, 0, 1, -4, -2, 0, -2, 0, 0, 0, 1, 0, 1, 3, 3, 2, 2, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, -3, -2, -1, -2, -1, 0, 0, 0, 1, 1, 3, 3, 3, 0, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 3, -4, -4, -1, -1, -1, 0, 1, 0, 2, 1, 1, 1, 2, 2, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 1, 2, -3, -3, -3, -3, -1, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, 3, -3, -2, -3, -3, -3, -1, -1, 0, -1, -2, -1, -1, -1, -3, -3, -1, -1, -1, -2, -2, -2, -4, -2, 0, 0, 2, -2, -2, -4, -2, -4, -3, -2, -2, -3, -3, -5, -4, -4, -6, -4, -4, -3, -2, -3, -3, -2, -3, -2, 0, 1, 1, -2, -1, -1, 0, 1, 0, 1, 0, 0, 0, -2, -1, -1, -1, -1, -1, -3, -2, -1, 0, 0, 0, 0, 2, 3, 4, 0, -1, -1, 0, -1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, -2, -1, -1, -1, 0, 1, 1, 1, 3, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 2, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 4, 0, 1, 0, 0, -1, -1, -1, -2, 0, 1, 2, 3, 3, 2, 1, 2, -1, -2, -1, 0, -1, 0, 0, 0, 2, 2, 0, 0, 1, -1, -2, -1, -1, -3, -2, 0, 2, 3, 3, 3, 3, 1, 0, 0, 0, 0, -1, -1, 0, 0, 2, 2, 2, 3, 0, -1, -2, -1, -4, -3, -2, 0, 0, 1, 2, 4, 1, 0, 0, -1, -2, -1, -1, -2, -1, 0, 0, 1, 0, 1, 0, 0, -2, -2, -3, -2, -2, 0, 2, 2, 2, 4, 2, 1, 0, 0, -1, -1, 0, 0, -2, -1, 0, 1, 0, 2, 2, -1, 0, 0, -2, -1, -1, 0, 0, 2, 2, 1, 2, 2, 0, 1, -1, -1, -1, 0, -2, -2, -1, 1, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 1, 2, 4, 2, 2, 2, 2, 0, 0, 0, 0, -1, -3, -2, -1, 1, 0, 0, 0, -1, -1, -2, -2, -1, 0, 1, 3, 3, 3, 3, 2, 2, 0, 0, 0, 0, 0, -1, -2, -2, -2, 0, -3, -2, -2, -1, -1, -1, -2, 0, -1, 0, 3, 5, 3, 3, 3, 0, 0, 0, -1, -2, -1, -2, -3, -1, 0, 0, -1, -2, -2, 0, 0, 0, 0, -1, -1, 1, 2, 3, 5, 4, 2, 0, 1, -1, -2, -2, -1, -1, -1, -2, -1, 0, -3, -1, -1, -1, 0, 0, 0, 0, 0, 1, 2, 4, 4, 2, 4, 1, 0, 0, -2, -3, -3, -1, -2, -2, -2, 1, -2, -1, 1, 0, 1, 0, 0, -1, 0, 0, 3, 3, 3, 4, 4, 1, 1, 0, 0, -1, -1, -1, -2, -1, -1, 0, -1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 2, 4, 3, 2, 2, 1, 0, 0, -1, -2, -1, -2, -3, -1, 0, -1, 0, 0, 2, 0, -1, 0, 0, 1, 0, 1, 1, 2, 4, 1, 0, 0, 1, 0, 0, -1, -3, -3, -2, -1, 1, -1, 0, 0, 0, 1, -1, 0, -1, 0, 0, 2, 2, 3, 3, 2, 0, 0, 0, 1, -1, 0, -3, -2, -1, 0, 1, 0, 0, 0, 0, 0, -2, -3, -2, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -2, -1, -1, -1, 0, 1, 0, 0, 0, 1, -1, 0, -3, -3, -2, -1, -1, 0, 1, 1, 0, 2, 1, 1, 0, 0, -2, -3, 0, 0, 0, 3, 0, 1, 1, 0, 0, -2, -3, -1, -1, 0, 0, 0, 1, 1, 1, 1, 1, 0, -1, 0, -2, -1, -2, 0, 0, 3, 0, 1, 0, 0, -2, 0, -3, -1, -1, 0, 1, 1, 1, 2, 1, 0, -1, 0, -1, -2, -2, -1, 0, 0, 2, 3, -1, -1, 0, 0, -1, -2, -2, -1, 0, 2, 0, 3, 2, 1, 0, 0, 0, -1, -2, -2, -2, -2, -1, 0, 2, 4, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 0, -3, -3, -3, -4, -2, -3, -1, 0, 0, 2, -1, -1, 0, 0, -1, -1, -1, 0, 0, 2, 1, 1, 2, 1, 0, -1, -2, -3, -5, -4, -4, -1, -3, -1, 0, 3, -1, -2, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, -2, -1, -1, -3, -2, -3, -2, -1, 0, 0, -1, 1, 4, -4, -1, -1, 0, 0, -1, 0, 1, 1, 1, 0, -1, 0, -1, -2, 0, -1, -2, 0, 1, 1, 2, 3, 3, 4, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, -1, 1, 0, 0, 0, 0, -1, 1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -2, 0, 0, -2, 0, -2, 0, 0, 0, -2, -1, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, -1, -1, 0, 1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 1, 0, 0, 0, 1, -1, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, -1, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, -2, -1, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, -1, 0, -1, -1, -1, 0, -2, 0, 0, -1, 0, -1, 0, -1, -2, -2, -2, 0, 0, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 2, 3, 2, 3, 2, 1, 0, 0, 0, -1, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 1, 0, 0, 1, 0, -1, -2, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, -1, 0, -1, 0, -2, -2, 0, 0, 0, -2, -1, 0, -2, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -2, 0, 1, 0, -1, -1, 0, -2, 0, 0, 0, 2, 0, 0, 1, 1, 0, 0, 0, -1, -2, -1, 0, -1, 0, -1, -2, 1, 0, 1, 0, -2, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, -1, -2, -2, -1, -1, 0, -1, -1, 1, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, 1, 1, 1, 0, 1, 0, 0, -1, -1, -1, 0, 0, -1, -2, -2, 0, 0, 0, -1, -1, -3, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, -2, -2, 0, -1, -1, -1, 0, -1, 2, 1, -1, -1, -1, -4, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -2, -1, -1, 0, 0, -2, -2, -3, -3, -3, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, -2, -2, -4, -4, -2, -2, -1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -2, -1, -2, -2, -2, -3, -3, -3, -3, -1, 1, 0, 0, 2, 0, -1, 0, -1, -1, 0, 0, -1, -1, 0, -2, -2, 0, -1, 0, -1, -3, -3, -4, -3, -3, -1, 0, 0, 0, 0, 1, -1, -1, 0, 0, -1, 0, -2, -1, -2, -2, -1, -1, 0, 0, -2, -2, -4, -5, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, -1, 0, -1, -2, -3, -5, -3, -3, -3, -2, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, -2, -2, -2, 0, 0, -1, -1, -2, -3, -5, -4, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, -2, 0, 0, 0, 0, -1, -2, -2, -3, -2, -2, -2, 0, 0, 1, 1, 0, 0, 0, 2, 2, 2, 1, -1, -2, 0, -1, -1, 0, 0, 0, -1, -1, -3, -2, -3, -1, -1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, -1, -2, -1, -1, -2, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -2, -2, -3, -2, -1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, -1, -1, -1, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, -2, -2, -1, -2, -1, -1, -2, 0, 0, 1, 1, 0, 1, 1, 1, 1, 2, 0, 0, 0, 0, -1, 0, -2, -2, -1, -3, -3, -4, -4, -3, -3, 0, 0, -1, -4, -4, 0, 0, 1, 3, 4, 6, 9, 7, 6, 3, 0, 1, 2, 1, 2, 2, 4, 7, 7, 6, 4, 0, 1, -1, -1, 0, 3, 2, 1, 2, 3, 4, 4, 5, 2, 1, 0, 2, 2, 1, 0, 0, 0, 1, 3, 0, -1, -5, 2, 1, 0, 1, 2, 0, 0, 1, 2, 3, 3, 1, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, 0, -2, -3, -6, 1, 1, 0, 0, 0, 0, 0, 1, 1, 2, 4, 2, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -2, -6, 0, 0, 0, -2, -1, -2, 0, 0, 0, 2, 2, 2, -1, -1, -1, -1, 0, 1, 0, 0, 0, 0, -1, 0, -2, -5, 0, 0, 0, -2, -2, -1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 2, 3, 1, 0, 0, 0, 0, -1, 0, -1, -3, 1, 2, 1, -2, -2, -1, -2, -1, -2, 0, 1, 2, 2, 2, 3, 2, 1, 0, 0, 0, 0, -1, 1, 0, 0, -3, 4, 4, 1, 1, 0, -1, -2, 0, 0, 0, 1, 3, 3, 4, 3, 0, -1, -2, -3, -2, 0, 0, 0, 1, 0, -3, 5, 5, 2, 0, 0, -2, -1, 0, -1, -1, 0, 1, 4, 3, 0, 0, -3, -2, -3, -2, 0, 1, 3, 3, 0, -3, 7, 4, 0, 0, 0, -3, -3, 0, -2, -1, 0, 0, 1, 4, 2, -1, 0, 0, 0, 1, 1, 3, 4, 3, 2, -1, 4, 2, 0, -2, -2, -2, -2, -1, -1, 0, 0, 0, 2, 5, 3, 2, 2, 1, 1, 3, 3, 5, 4, 4, 0, -1, 2, 0, -1, -4, -3, -4, -2, -3, -2, 0, 0, 2, 4, 7, 4, 2, 2, 1, 3, 3, 3, 3, 2, 3, 0, 0, 0, -1, -2, -2, -3, -3, -3, -4, -4, 0, 2, 5, 5, 6, 3, 0, -1, 0, 0, 2, 3, 1, 2, 2, 0, -1, -2, -4, -6, -4, -5, -4, -6, -5, -4, -2, 1, 5, 4, 5, 2, 0, -1, 0, 2, 3, 1, 3, 3, 4, 1, 0, -3, -5, -4, -2, -4, -6, -6, -3, -4, -2, 0, 4, 4, 4, 2, 0, 0, 2, 4, 3, 2, 4, 3, 5, 2, 0, -3, -4, -3, -1, -2, -3, -5, -3, -1, -1, 1, 5, 4, 3, 4, 1, 1, 2, 3, 5, 3, 4, 6, 5, 1, 0, -4, -3, -2, -1, -1, -4, -2, -2, -1, 0, 1, 5, 6, 7, 4, 3, 2, 2, 3, 3, 6, 5, 4, 2, 0, -2, -3, -2, 0, -1, -2, -4, -2, -3, -2, -1, 0, 5, 6, 6, 4, 0, 0, 2, 1, 3, 6, 6, 4, 0, 0, -3, -2, -2, -1, -2, -2, -1, 0, -1, -2, -1, 0, 4, 6, 5, 1, 1, 0, 2, 3, 4, 5, 5, 2, 1, 0, -3, -2, -1, 1, -1, 0, -3, 0, 0, -1, -2, 0, 5, 6, 5, 0, 0, 0, 1, 3, 4, 6, 5, 4, 2, 0, -3, 1, 2, 0, 1, 1, 0, -1, -2, -3, -2, 0, 2, 4, 2, 1, 1, 1, 3, 3, 4, 3, 5, 3, 1, -1, -4, 2, 0, 1, 0, 0, 0, 0, -2, -3, -2, 0, 0, 3, 2, 2, 2, 3, 4, 3, 2, 2, 4, 2, 0, -1, -5, 0, 0, 0, 0, 0, -1, 0, -2, -1, -2, 1, 0, 2, 1, 2, 2, 1, 1, 1, 1, 3, 3, 2, 0, -4, -4, 0, 0, 0, 0, 1, -1, -2, -1, 0, 0, 1, 2, 1, 2, 2, 2, 1, 2, 2, 2, 4, 3, 1, 0, -2, -4, 0, 0, 1, 2, 1, -1, 0, 0, 0, 2, 2, 1, 3, 2, 3, 5, 4, 3, 3, 1, 1, 3, 1, -1, -3, -5, 1, 1, 2, 0, 0, -1, 0, 0, 0, 1, 2, 3, 1, 0, 2, 3, 1, 0, 0, 0, -2, -2, -3, -4, -3, -6, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -1, 0, 1, 1, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, -1, 0, -2, -1, 0, 0, 0, 0, 1, 0, -1, -2, -2, -3, -5, -5, -5, -4, -4, -3, -2, 0, 0, 0, 1, 0, 2, 5, -3, -1, 0, -1, 0, 1, 0, 0, 0, -1, 0, -1, -2, -3, -3, -3, -3, -3, -2, -1, -1, 0, 0, 0, 1, 4, -2, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -2, -3, -1, -1, -1, 0, 0, 0, 1, 2, 3, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 2, 1, 2, 2, 0, 0, -1, -1, 0, 0, 0, 0, 1, 2, 2, 4, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 4, 2, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 2, 3, 0, 0, 1, 0, 0, 0, -3, -2, 0, 1, 3, 3, 3, 4, 3, 2, 1, 0, 0, 0, 0, 0, 0, 1, 2, 3, 1, 1, 1, 0, 0, -3, -3, -1, 0, 0, 3, 5, 4, 5, 2, 2, 2, 0, 0, 0, 0, -1, -1, 1, 0, 2, 1, 0, 0, -1, -2, -2, -1, -1, 0, 1, 2, 4, 3, 3, 4, 3, 2, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, -1, -1, 0, 0, 1, 2, 3, 4, 3, 4, 3, 2, 2, 0, 1, 0, -1, -1, -1, 0, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 1, 2, 4, 3, 4, 3, 3, 2, 2, 0, 0, -1, -1, -3, -2, -2, 0, -1, -1, 0, 0, 1, 1, -1, 0, 0, 2, 2, 3, 4, 4, 3, 4, 3, 0, 0, 0, -1, -2, -3, -3, -2, 0, -2, 0, 0, 0, 0, 0, 0, 0, 1, 2, 5, 5, 4, 4, 3, 1, 2, -1, 0, -2, -3, -4, -4, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 3, 5, 6, 4, 3, 1, 1, 1, 0, -1, -2, -3, -3, -4, -3, -3, 0, -1, -1, 0, 1, 1, 0, 0, 0, 1, 4, 5, 6, 5, 4, 3, 2, 1, -1, -2, -2, -2, -3, -4, -2, -2, -1, 0, -1, 0, 1, 0, 0, 0, 0, 1, 4, 5, 6, 5, 3, 3, 2, 2, 0, 0, 0, -2, -3, -4, -3, -3, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 2, 5, 6, 4, 3, 3, 3, 3, 0, 0, 0, -1, -3, -3, -4, -1, 0, -1, 1, 0, 2, 0, 0, -1, 0, 0, 2, 3, 4, 6, 4, 4, 3, 3, 1, 0, -1, -1, -1, -3, -3, -2, 1, -1, 0, 1, 1, 0, 0, -2, -2, 0, 0, 4, 5, 6, 3, 4, 1, 2, 1, 1, 0, 0, -1, -3, -2, 0, 1, 0, 0, 1, 0, 0, -2, -1, -1, -1, 0, 3, 4, 3, 4, 2, 3, 0, 0, 0, 0, 0, -3, -2, 0, 0, 3, 0, 0, 1, 0, -2, -1, -2, -3, -2, 0, 1, 3, 4, 3, 1, 3, 1, 0, 0, 0, -2, -2, 0, -1, 1, 3, 0, 1, 0, -1, -1, -1, -3, -2, -1, 0, 1, 2, 4, 3, 2, 3, 0, 0, -1, -2, -1, 0, 0, -1, 2, 3, -1, 0, 0, -2, -1, -2, -1, -2, 0, 0, 2, 2, 3, 1, 1, 0, -1, 0, -2, -1, -1, -2, 0, 0, 1, 4, 0, -1, -1, -2, -2, -2, -3, 0, 0, 0, 2, 3, 1, 1, 0, -1, -2, -3, -3, -1, -2, -3, -1, 0, 2, 5, -1, 0, -1, -1, -2, -3, -2, 0, 1, 1, 1, 2, 0, -1, 0, -2, -2, -4, -3, -3, -3, -1, -1, 0, 1, 4, -3, -1, -2, -1, -2, -2, -1, 0, 0, 1, 0, 0, 0, 0, -2, -3, -5, -3, -5, -2, -3, -3, -2, -2, 1, 4, -2, -2, -1, -1, -2, -2, -2, 0, 0, -1, -2, -1, -3, -4, -4, -4, -4, -4, -3, -2, -2, -1, -2, 0, 1, 4, 2, 2, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, -2, 0, 0, -2, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 1, 2, 2, 2, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 2, 1, 2, 0, 2, 1, 1, 2, 0, 2, 2, 1, 0, -1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 3, 4, 2, 3, 2, 4, 1, 3, 2, 1, 0, 0, -2, 2, 2, 1, 0, 0, -1, 0, 0, 0, 0, 1, 3, 2, 1, 3, 4, 3, 2, 3, 3, 1, 1, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 2, 2, 1, 1, 3, 5, 3, 3, 2, 3, 1, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 2, 1, 3, 3, 4, 4, 3, 3, 1, 0, 0, 0, -1, -2, 2, 0, 1, -1, -1, -2, 0, -1, 0, 1, 1, 2, 1, 2, 2, 2, 4, 3, 3, 1, 3, 2, 1, 0, 0, 0, 0, 1, 0, -1, 0, -1, -2, -1, -1, 0, 0, 2, 2, 2, 2, 3, 4, 2, 2, 1, 3, 2, 2, 0, 0, -2, 0, 1, 0, 0, -2, -3, -3, -2, -1, 0, 1, 1, 2, 2, 1, 2, 1, 2, 1, 2, 2, 1, 2, 0, 0, -2, 1, 1, -1, 0, -1, -3, -2, -4, -2, 0, 0, 1, 2, 2, 3, 2, 1, 2, 3, 3, 3, 1, 2, 0, 0, -2, 2, 0, -1, 0, -2, -3, -3, -3, -2, 0, 0, 2, 2, 2, 1, 1, 1, 1, 2, 1, 1, 1, 0, 0, 0, -1, 1, 0, 0, -1, -2, -1, -2, -3, 0, -1, 1, 2, 3, 3, 3, 1, 2, 3, 3, 3, 1, 1, 0, 0, 0, 0, 1, -1, -1, -1, -2, -4, -2, -1, -1, 1, 0, 1, 3, 4, 1, 2, 0, 2, 3, 2, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -2, -2, -2, -2, -1, 0, 1, 1, 3, 3, 1, 2, 1, 4, 2, 3, 3, 0, 0, -1, 0, 0, 0, 0, -1, -2, -1, -3, -3, -1, 0, 0, 0, 1, 2, 3, 3, 0, 2, 3, 2, 3, 2, 1, 0, 0, -1, -2, 0, 0, -2, -1, -1, -1, -2, -3, -2, 1, 2, 2, 3, 2, 3, 1, 1, 2, 4, 4, 3, 1, 1, -1, 0, 0, 0, 0, -1, -1, -1, -2, -1, -2, -1, 1, 1, 2, 4, 3, 3, 2, 4, 4, 3, 2, 2, 2, 0, 0, 0, -1, 1, 0, 0, -1, 0, -3, -1, -2, -1, 0, 3, 3, 6, 6, 3, 3, 3, 4, 3, 2, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, -3, -1, 1, 2, 4, 5, 5, 5, 3, 3, 2, 4, 3, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -2, -2, 0, 0, 4, 5, 5, 5, 4, 3, 2, 2, 2, 1, 0, 1, 0, -1, 0, 1, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 1, 3, 2, 1, 1, 2, 3, 2, 0, 1, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 3, 2, 3, 2, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 1, 0, 0, 0, 0, -1, -2, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, -2, 3, 4, 5, 4, 3, 3, 3, 3, 4, 2, 2, 0, 1, -1, -2, -4, -4, -3, -3, -3, -2, -3, 0, 2, 5, 7, 2, 2, 3, 2, 3, 3, 2, 2, 2, 3, 3, 2, 0, -2, -2, -5, -5, -5, -6, -5, -3, -2, 0, 0, 3, 7, 2, 2, 2, 1, 0, 0, -1, 0, 0, 3, 5, 3, 2, 0, -1, -3, -6, -6, -7, -4, -2, -3, 0, 1, 2, 5, 3, 1, 0, 0, -2, -2, -2, 0, 0, 2, 3, 2, 1, 0, 0, -3, -4, -6, -5, -5, -4, -1, 0, 0, 2, 5, 2, 3, 1, -1, -2, -4, -3, -4, -3, 0, 2, 1, 2, 1, 1, -1, -3, -5, -5, -4, -5, -2, 0, 1, 2, 4, 4, 2, 2, -1, -2, -3, -6, -6, -4, -1, 0, 1, 2, 1, 0, -1, -4, -4, -3, -3, -4, -2, -1, 0, 0, 4, 3, 1, 2, 0, -2, -3, -7, -6, -5, -2, 0, 1, 3, 1, 1, 0, 0, -3, -3, -2, -4, -5, -3, -1, 1, 2, 1, 2, 0, 0, -1, -3, -7, -6, -5, -4, 0, 0, 1, 0, 0, 0, 0, 1, 0, -2, -4, -4, -4, -2, 0, 2, 1, 1, 2, 0, -1, -4, -6, -6, -5, -2, -2, 0, 0, 1, 1, 3, 2, 2, 1, -1, -2, -3, -4, -4, -1, 2, 0, 0, 0, 0, -2, -5, -9, -8, -5, -3, -2, 1, 2, 1, 2, 2, 2, 1, 0, 0, -4, -4, -4, -5, 0, 0, -2, -2, -2, -1, -4, -7, -10, -9, -7, -4, 0, 1, 1, 1, 2, 3, 1, 0, 0, -4, -5, -4, -5, -3, -1, 0, -1, -1, -1, -2, -6, -7, -9, -9, -7, -5, -2, 1, 2, 3, 2, 0, 0, 0, -1, -3, -3, -5, -4, -4, -2, 0, -1, 0, 0, -1, -4, -8, -10, -10, -7, -5, -1, 0, 1, 3, 1, 0, 0, 0, -3, -3, -5, -5, -6, -6, -4, 0, 0, 1, 0, -2, -4, -7, -9, -8, -7, -4, 0, 1, 1, 1, 3, 1, 1, 0, -3, -3, -5, -6, -5, -5, -3, 0, 0, 0, 0, -2, -4, -6, -8, -8, -6, -2, 0, 1, 4, 3, 2, 2, 1, 0, -1, -2, -5, -7, -8, -4, -2, 0, 0, 1, 0, -1, -4, -5, -7, -7, -4, -3, -1, 2, 2, 3, 3, 2, 2, 0, -1, -2, -4, -5, -5, -3, -2, 0, 2, 1, 0, -2, -2, -5, -7, -7, -4, -4, 0, 1, 2, 2, 3, 4, 2, 0, -2, -2, -5, -5, -4, -2, 1, 2, 2, 3, 0, -1, -3, -6, -6, -6, -6, -4, 0, 2, 1, 1, 2, 1, 1, 0, -1, -2, -4, -3, -4, 0, 0, 4, 3, 3, 3, 0, -1, -4, -6, -5, -3, -1, -1, 2, 2, 3, 2, 2, 0, 0, -2, -2, -4, -4, -1, 1, 3, 6, 4, 5, 3, 2, 0, -4, -4, -3, -2, -2, 0, 2, 2, 1, 2, 1, 0, -1, -4, -2, -3, -4, -1, 0, 2, 6, 2, 3, 2, 2, -1, -4, -4, -3, -2, 0, 0, 1, 0, 0, 0, -2, -4, -4, -5, -5, -4, -4, 0, 0, 3, 6, 1, 1, 2, 0, -2, -3, -2, -3, 0, 0, 1, 1, 2, 0, -2, -3, -5, -7, -7, -5, -5, -4, -1, 0, 3, 5, 2, 1, 0, 0, -1, -1, -3, -1, 0, 0, 2, 1, 0, 0, -2, -7, -8, -8, -7, -6, -3, -3, -1, 0, 3, 6, 1, 1, 0, 0, -1, 0, 0, 1, 2, 2, 0, 1, 1, -1, -5, -7, -8, -9, -7, -6, -5, -3, -1, -1, 1, 5, 2, 1, 2, 1, 1, 1, 2, 3, 3, 1, 0, 0, 0, -2, -5, -7, -9, -9, -7, -3, -4, -1, 0, 1, 4, 7, 1, 1, 3, 3, 3, 3, 4, 3, 2, 1, 3, 2, 0, 0, -2, -3, -5, -5, -2, 0, 2, 3, 4, 6, 6, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, -1, 1, 0, 1, -2, -1, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -2, -3, -3, -4, -4, -4, -3, -3, -4, -2, 0, 0, 0, -3, -2, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, -1, -1, -3, -4, -2, -2, 0, 0, -1, 1, 3, 3, -3, -2, 0, -1, -1, 1, 2, 2, 2, 0, 1, -1, -2, -1, -1, -2, -2, -2, -1, 0, 1, 0, 1, 2, 3, 2, -4, -3, -2, -1, 0, 1, 4, 2, 2, 2, 1, -1, -1, -1, -1, -2, -2, -2, 0, 0, 0, 2, 0, 0, 1, 2, -4, -4, -1, 0, 0, 1, 4, 1, 3, 1, 0, 0, -2, -1, -2, -2, -1, 0, 0, 1, 1, 1, 0, 0, 1, 1, -2, -2, -2, 0, 0, 1, 4, 2, 2, 2, 2, 0, 0, -2, -3, -2, -2, 0, -1, 0, 1, 3, 2, 0, 0, 3, 0, -2, 0, 0, 0, 3, 4, 4, 4, 4, 2, 2, 0, -1, -2, 0, -2, 0, 0, 0, 1, 2, 2, 0, 0, 3, -1, -1, 0, 0, 1, 2, 5, 4, 4, 4, 3, 4, 1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, 2, 0, 0, 0, 1, 0, 4, 5, 5, 5, 5, 3, 3, 2, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, -2, 0, 3, 1, 1, 1, 2, 3, 4, 6, 6, 4, 4, 4, 4, 3, 2, -1, -1, -1, 0, 0, -2, -2, -1, 0, -1, 1, 3, 1, 2, 2, 3, 3, 4, 6, 7, 5, 5, 7, 4, 5, 0, -2, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 2, 2, 2, 2, 2, 3, 4, 6, 6, 7, 7, 8, 6, 4, 0, -3, -3, -1, 0, 0, -1, -2, -2, -3, -2, 0, 2, 2, 2, 1, 0, 1, 3, 4, 5, 7, 6, 8, 5, 3, 0, -3, -3, -1, 0, 0, 0, 0, -2, -1, -1, 0, 1, 2, 0, 1, 0, 1, 4, 4, 5, 6, 7, 7, 6, 2, 0, -3, -1, -1, 0, 0, 0, -2, -4, -1, 0, 0, 2, 2, 1, 0, 0, 0, 2, 4, 3, 4, 6, 6, 4, 3, 0, -2, -2, -1, -2, 0, -1, -1, 0, -1, -1, 0, 2, 1, 0, 0, 0, 1, 2, 3, 2, 1, 4, 5, 5, 0, 0, 0, -2, -3, -3, -2, 0, -1, -1, 0, -1, 0, 1, 0, 0, -1, 0, 1, 2, 1, 0, 2, 2, 5, 4, 0, 0, -1, -2, -4, -3, 0, 0, -1, -1, -1, 0, 0, 2, 1, -1, 0, 1, 2, 3, 1, 0, 2, 3, 6, 5, 1, 0, -1, -1, -2, -2, -1, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 3, 3, 1, 0, 0, 3, 4, 4, 2, 0, 0, -2, -1, -1, 0, 0, 0, 0, -1, -1, 1, 0, -2, 0, 1, 1, 3, 4, 3, 1, 2, 2, 4, 4, 0, 0, 0, -1, -3, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 2, 3, 2, 2, 3, 4, 3, 2, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, -2, -1, 0, -1, 2, 3, 3, 2, 1, 1, 2, 1, 1, -1, -1, 0, 0, 0, 2, 0, 0, 0, 0, 2, 2, 2, -2, -2, -1, 0, 0, 2, 2, 2, 0, 1, 1, 0, 0, -3, -1, 0, 0, 1, 1, 0, -1, -1, 1, 2, 3, 1, -2, -1, -2, -1, 0, 0, 1, 1, 1, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -2, -2, 0, 1, 4, 4, 2, -2, -2, -1, -2, -1, -1, 1, -1, 0, 0, 0, 1, 0, -2, -2, 0, 1, 1, -1, -2, 0, -1, 2, 4, 5, 2, -2, -3, -2, 0, -2, -2, 0, -1, 0, 1, 0, 2, 0, -1, -3, 0, 0, 0, -1, -2, -1, 0, 2, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 2, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 0, 1, 1, -1, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 2, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, -1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 2, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, 1, 2, 1, 1, 1, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 2, 2, 1, 0, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, 2, 0, 2, 0, 0, 2, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 1, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 1, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 1, 0, 1, 2, 0, 1, 1, 0, 0, 1, 0, 2, 1, 1, 0, 0, 1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 2, 0, 2, 1, 0, 1, 0, 0, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 2, 0, 2, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 2, 2, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -3, -2, -1, -1, -2, -1, -1, -2, -2, -3, -1, -2, -5, -4, -3, -3, -3, -2, -2, -1, 0, -1, 0, 0, 1, 1, -4, -3, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, -3, -3, 0, -1, 0, 0, 0, 1, 3, -3, -4, -4, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -2, -1, -2, 0, -1, 0, 1, 1, 1, 2, 2, -5, -3, -2, 0, 0, 0, 2, 1, 0, 2, 1, 1, 1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 1, 1, 3, -5, -4, -1, 0, -1, 1, 0, 2, 1, 3, 3, 4, 1, 0, 0, 1, 0, 0, 0, 1, 0, 2, 1, 2, 1, 4, -5, -4, -3, -2, 0, 0, 1, 0, 2, 2, 3, 4, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 5, -3, -2, -2, 0, -1, 0, 2, 2, 2, 2, 5, 5, 2, 3, 1, 1, 2, 0, 0, 0, 1, 0, 2, 0, 1, 2, -1, -2, -1, -1, 0, 1, 0, 2, 3, 3, 3, 6, 4, 3, 2, 2, 1, 0, 0, 0, 0, 0, 1, 0, 2, 2, -1, 0, -1, 0, 1, 0, 2, 2, 3, 4, 3, 6, 4, 2, 2, 1, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 4, 2, 3, 4, 4, 5, 4, 3, 2, 1, 0, 0, 0, -2, -1, -2, -1, -1, 0, 1, 0, 0, 0, 0, 1, 3, 3, 2, 4, 5, 6, 6, 3, 4, 1, 0, 0, 0, 0, -1, -2, -3, -3, -4, -2, 1, 0, 0, 0, 1, 1, 4, 3, 4, 4, 5, 8, 7, 5, 2, 0, 0, 0, 0, -1, -1, -2, -2, -4, -2, -2, 0, -1, 0, 1, 0, 2, 2, 3, 5, 4, 7, 6, 6, 5, 2, 1, 0, -1, 0, 0, -2, -1, -3, -3, -3, -2, 0, 0, 0, 0, 0, 1, 2, 2, 3, 5, 7, 8, 6, 3, 1, 1, 0, -1, 0, 0, -1, -2, -4, -3, -2, -2, 0, -2, -1, -1, 0, 0, 1, 2, 3, 3, 6, 8, 5, 3, 4, 1, 0, 0, 0, -1, -1, -2, -4, -3, -3, -2, 1, -2, -1, -1, 0, 0, 2, 1, 0, 3, 4, 6, 5, 4, 1, 0, 1, 1, 0, -1, -2, -2, -2, -2, -3, -1, 0, -1, -1, -1, 0, 1, 2, 0, 0, 3, 3, 6, 6, 5, 4, 2, 0, 0, 0, 0, -1, -2, -2, -2, -1, 0, 0, -2, -1, -1, 0, 0, 0, 1, 0, 2, 4, 6, 6, 4, 4, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 1, -2, -1, -1, 0, 0, 0, 0, -1, 0, 4, 6, 6, 4, 2, 2, 1, 0, 0, 0, 0, -2, -2, -1, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 1, 3, 5, 5, 3, 1, 2, 0, 0, 1, 1, -1, 0, -2, 0, 0, 1, 1, -4, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 3, 2, 1, 1, 0, 1, 0, 0, -2, 0, 0, 0, 0, 2, -2, -3, -2, -1, 0, -1, 0, -1, 0, 0, 2, 1, 2, 0, 1, 0, 0, 1, 0, -1, -2, 0, 0, 0, 2, 3, -2, -1, -3, -1, -2, 0, 0, -1, 0, -1, 0, 1, -1, -1, 0, 0, -1, 0, 0, -2, -1, 0, 0, 0, 2, 2, -2, -3, -2, -3, -1, -1, 0, 0, -2, 0, 0, 0, 0, -2, -1, -2, -3, -2, -1, -1, -2, -1, 0, 1, 3, 3, -5, -4, -4, -4, -4, -2, -2, -3, 0, 0, 0, -1, -2, -3, -4, -3, -3, -3, -1, -3, -3, -1, 1, 1, 1, 1, -5, -4, -5, -5, -3, -5, -3, -5, -1, -2, -1, 0, -1, -3, -3, -4, -3, -2, -2, -2, -3, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 4, 5, 6, 6, 5, 4, 5, 2, -1, 0, -1, -2, -2, -3, -1, -1, -2, -1, -1, 0, 2, 5, 8, 12, 0, 0, 2, 3, 2, 1, 2, 2, 3, 1, 0, 1, 0, 0, -1, -5, -3, -3, -3, -4, -4, -1, 0, 1, 5, 9, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 2, 2, 1, 0, -3, -5, -5, -5, -4, -3, -2, -1, 1, 3, 7, 1, 0, 1, 0, 0, -2, -3, -1, 2, 2, 2, 3, 4, 2, 0, -2, -3, -4, -6, -5, -5, -2, -1, 2, 3, 5, 2, 1, 0, 0, 0, -3, -5, -4, 0, 1, 1, 3, 4, 3, 0, -1, -5, -5, -4, -5, -4, -4, 0, 1, 3, 6, 3, 1, 0, 0, -3, -6, -6, -5, -1, 0, 1, 4, 5, 3, 1, -1, -3, -4, -5, -4, -4, -3, -1, 0, 1, 5, 3, 1, 1, -1, -3, -5, -7, -8, -4, -1, 0, 2, 2, 3, 1, -2, -2, -2, -4, -4, -5, -5, -3, -1, 0, 1, 3, 3, 0, 0, -3, -5, -8, -6, -5, -1, 0, 2, 2, 1, 1, 0, 0, -1, -3, -5, -5, -5, -3, -1, 0, 0, 3, 1, 0, 0, -2, -5, -8, -7, -5, -2, 0, 0, 1, 1, 2, 1, 2, 0, 0, -3, -4, -5, -4, -2, 0, 2, 0, 1, 0, -1, -2, -6, -9, -9, -7, -2, -1, 1, 0, 1, 2, 2, 1, 0, 0, -2, -3, -6, -5, -3, 0, 2, 0, 0, 0, 0, -4, -8, -10, -9, -6, -3, 0, 1, 0, 0, 0, 1, 0, 0, 0, -3, -3, -5, -4, -4, -2, 1, -2, -1, 0, 0, -5, -8, -11, -11, -7, -3, 0, 2, 1, 2, 0, 0, 0, -3, -3, -4, -5, -4, -3, -3, -3, 0, 0, 0, 0, -1, -4, -8, -11, -10, -6, -4, 0, 1, 3, 1, 1, 0, -1, -3, -5, -6, -5, -4, -3, -2, -3, 0, 0, 1, 1, 0, -6, -8, -10, -9, -6, -2, -1, 0, 2, 2, 0, 0, 0, -2, -4, -5, -6, -3, -5, -4, -2, 0, 1, 3, 1, 0, -4, -7, -9, -8, -4, -2, 1, 2, 2, 1, 0, 1, 0, -1, -5, -5, -6, -5, -6, -3, -2, 2, 2, 3, 2, 0, -3, -7, -7, -6, -5, -2, 0, 2, 2, 2, 2, 1, 0, -2, -2, -4, -4, -5, -5, -4, 0, 2, 3, 5, 1, -1, -2, -5, -7, -6, -5, -2, 0, 3, 4, 2, 0, 0, 0, -1, -2, -4, -4, -5, -5, -1, 0, 4, 4, 5, 1, 0, -4, -6, -6, -6, -4, -2, 0, 2, 2, 2, 1, 0, 0, -1, -3, -4, -5, -5, -3, -1, 2, 3, 4, 5, 2, 0, -4, -7, -5, -5, -3, 0, 1, 2, 1, 1, 0, 0, -1, -2, -1, -3, -5, -4, -3, 0, 3, 6, 5, 5, 3, 0, -2, -6, -6, -6, -3, -1, 0, 0, 2, 1, 0, -1, -2, -2, -4, -4, -5, -4, -1, 0, 3, 7, 5, 3, 2, 0, -3, -4, -5, -3, -3, 0, 2, 3, 1, 0, 0, -2, -4, -5, -5, -4, -3, -3, -1, 2, 5, 9, 1, 1, 1, 0, -2, -4, -3, -4, 0, 2, 3, 2, 1, 2, 0, -4, -5, -6, -5, -5, -3, -3, 0, 0, 3, 8, 0, 0, 0, -1, -3, -4, -2, -2, 2, 2, 3, 2, 2, 1, -3, -5, -6, -6, -5, -5, -4, -4, -1, 0, 3, 8, 1, 1, -1, -2, -1, -1, 0, 0, 3, 3, 3, 2, 2, -1, -3, -7, -7, -9, -8, -6, -3, -5, -2, -1, 2, 10, 3, 2, 1, 0, 0, 0, 1, 3, 5, 4, 3, 1, 0, 0, -3, -7, -9, -7, -7, -5, -3, -2, -2, 0, 4, 8, 3, 4, 2, 0, 1, 2, 3, 3, 4, 3, 2, 3, 2, 0, -1, -5, -4, -5, -3, -1, 0, 0, 0, 1, 6, 10, 2, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, -1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 2, 1, 0, 0, 0, 1, 2, 1, 1, -1, -1, 2, 1, 1, 0, 0, 0, 0, -1, 1, 0, 1, 2, 0, 0, 2, 1, 2, 3, 1, 2, 1, 0, 1, 0, -1, -2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 3, 3, 3, 2, 3, 2, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 2, 4, 3, 1, 1, 0, 1, 1, 0, -1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 2, 2, 2, 4, 3, 3, 3, 2, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 2, 1, 2, 2, 2, 2, 1, 1, 1, 0, 0, 2, 0, 0, -1, 0, 0, -1, -2, -1, 0, 1, 1, 1, 1, 2, 1, 2, 2, 1, 3, 1, 2, 2, 1, 0, 0, 1, 0, -1, 0, 0, -1, -2, -1, -1, -1, 0, 1, 2, 0, 1, 2, 1, 1, 2, 2, 1, 2, 1, 2, 0, 0, 1, 0, 0, -1, -1, -2, -2, -1, -1, 0, 0, 0, 1, 1, 1, 1, 0, 2, 3, 2, 2, 2, 2, 0, 0, -1, 1, 0, 0, 0, -1, -1, -2, -3, -1, -1, 0, 1, 2, 1, 1, 0, 1, 1, 1, 3, 1, 1, 1, 0, -1, -1, 0, 0, -1, -2, -1, -2, -2, -1, -2, 0, 1, 0, 2, 1, 2, 1, 0, 1, 2, 2, 3, 2, 1, 0, -1, 0, 1, 0, 0, 0, -2, -3, -2, -2, 0, 0, 1, 1, 2, 2, 2, 0, 0, 2, 2, 3, 2, 1, 1, 0, 0, 0, 0, 0, 0, -2, -2, -3, -2, -3, -2, 0, 1, 1, 2, 1, 2, 0, 1, 1, 3, 4, 1, 1, 1, -1, -1, 0, 0, -1, -1, -1, -2, -2, -2, -1, -1, 0, 0, 2, 1, 0, 0, 1, 1, 1, 2, 3, 1, 2, 0, 0, -1, 0, 0, 0, 0, -2, -2, -2, -1, -3, -1, 0, 1, 3, 2, 2, 2, 2, 2, 1, 2, 3, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, -2, -3, -1, -2, 0, 2, 2, 4, 4, 2, 3, 3, 3, 3, 3, 2, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, 1, 2, 4, 4, 4, 2, 4, 3, 3, 3, 3, 1, 1, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 2, 3, 4, 5, 4, 3, 4, 4, 2, 3, 3, 0, 0, 1, 0, 0, 2, 1, 1, -1, 0, 0, -2, 0, -1, 0, 1, 2, 2, 3, 2, 3, 3, 3, 3, 1, 1, 1, 1, 0, 0, 0, 2, 1, 0, 1, 1, -1, -1, 0, -1, 0, 0, 0, 2, 2, 3, 2, 2, 2, 2, 2, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 2, 1, 0, 0, 0, 0, 0, -2, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, -2, 1, 1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 2, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 1, 0, 1, 1, 0, 2, 1, -1, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, -1, 0, -2, -1, -1, 0, -1, -1, -1, 0, 0, 0, 1, 1, 3, 1, 3, 1, 1, 0, 0, 0, 0, 0, 1, 2, 2, 2, 1, 1, 0, 2, 0, -1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, -2, -4, 0, 1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, 1, 0, 0, -1, -1, 0, -2, -1, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, -1, -1, -2, -2, -1, 0, 0, 3, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -2, -1, -2, -1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, -2, -1, -1, -1, 0, 0, 0, 1, -1, 0, -2, -1, -1, 0, 0, 1, 1, 0, 0, -1, 2, 1, 0, -2, 0, -3, -2, 0, 0, -1, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 2, 0, 0, -3, -2, -3, -1, -2, -1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 1, 2, 0, 2, 0, 0, 1, -1, -2, -3, -3, -3, -2, -3, -2, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -2, -3, -3, -3, -3, -2, -3, -1, 0, 0, 1, 2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -2, -2, -3, -2, -3, -3, -2, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -2, -3, -3, -2, -3, -3, -3, 0, 0, 1, 1, 0, 0, 1, -1, 0, 1, 0, 1, 0, 0, 1, 2, 0, 0, 0, -2, -2, -2, -2, -3, -3, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 1, 0, 0, 0, -1, 0, -1, -3, -3, -2, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 1, 1, 0, 1, 0, 1, 0, 0, -1, -1, -2, -2, -2, -1, -2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, -1, -2, -2, 0, 0, -2, -2, -2, 0, -1, -1, 0, 2, 2, 1, 1, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, -2, 0, -1, -1, -1, 0, -2, -2, -2, -1, -1, 0, 1, 2, 0, 0, 0, -1, 0, -1, -1, 0, 1, 0, 1, 0, -1, 0, -1, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -1, 0, 0, 0, -1, -2, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, -2, -1, 0, 1, 1, 0, 0, -2, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 2, 1, 0, 0, 0, -1, 0, 1, 0, -1, -3, 1, 1, 0, 0, 1, 0, 1, 2, 1, 1, 2, 2, 1, 0, 1, 0, 0, 0, -2, -3, -1, -2, -2, 0, -3, -3, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 3, 0, 1, 1, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 2, 2, 1, 2, 2, 2, 2, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 1, 3, 2, 4, 2, 3, 2, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 2, 2, 2, 1, 3, 3, 2, 2, 1, 0, 1, 1, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, -1, 1, 1, 0, 1, 0, 2, 2, 2, 1, 1, 1, 2, 2, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 2, 1, 2, 0, 2, 2, 1, 2, 2, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 0, 1, 1, 3, 3, 1, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 2, 1, 2, 1, 2, 1, 0, 2, 1, 2, 0, 1, 1, 1, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 1, 0, 2, 2, 2, 2, 2, 2, 1, 1, 0, 2, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 2, 3, 2, 1, 0, 1, 2, 3, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 2, 0, 2, 2, 1, 0, 0, 1, 2, 2, 2, 1, 2, 1, 0, 0, -1, 0, 0, 0, -1, -1, -2, -2, -1, 0, 1, 3, 3, 1, 2, 1, 1, 2, 3, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 1, 1, 2, 2, 2, 0, 1, 1, 3, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 1, 2, 3, 2, 1, 1, 0, 0, 2, 3, 3, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 1, 2, 3, 4, 2, 2, 1, 0, 3, 1, 2, 1, 2, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 2, 2, 1, 2, 1, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 2, 2, 4, 4, 2, 2, 2, 3, 3, 2, 3, 2, 1, 0, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 1, 0, 2, 2, 1, 2, 3, 3, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 1, 0, 2, 3, 1, 2, 1, 1, 3, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 2, 0, 0, 1, 1, 2, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 2, 1, 1, 1, 0, 2, 2, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 1, 1, 1, 1, 0, 1, 0, 2, 4, 5, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 2, 1, 1, -1, 1, 0, 1, 0, 0, 0, 0, -1, 0, -2, -2, -1, -2, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, -1, -2, -1, -3, -1, 0, -1, -2, -2, -1, -2, -1, 0, 0, -2, 0, -1, 0, 0, -2, -1, 1, 0, 1, 1, 0, 0, -2, 0, -2, -1, -2, -3, -1, -1, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, -1, -2, -3, -2, -2, -3, -2, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -2, 0, -3, -2, -1, -2, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, -2, -3, -3, -2, 0, 0, 0, 0, 0, -1, -1, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -2, -2, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, -2, -1, -2, -2, -3, -2, 0, 0, 1, 1, 1, 1, 1, 1, 2, 0, 1, 1, 2, 1, 1, -1, 0, -1, 0, -1, -2, -3, -3, -1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 1, 1, 0, 0, -1, -1, -1, 0, -1, -2, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 1, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, -2, -2, -2, -2, -1, -2, -2, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, -1, 0, -2, -1, -1, -1, -1, -2, -1, -1, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -2, -2, -3, -3, -2, -2, 0, 0, -1, 1, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -2, -2, -2, -1, -1, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 2, 0, 0, 0, 0, 0, -1, -2, -1, -2, -4, -4, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, 0, 0, 1, 1, 1, 0, 0, -1, -2, -3, -4, -3, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, -2, -1, -1, -3, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 1, 1, 0, -1, -2, -2, -2, -2, -3, -2, -2, 0, 0, -1, 0, 0, 1, 0, 1, 1, 1, 0, 2, 1, 2, 2, 0, 1, -1, 0, 0, -2, -2, -3, -2, -3, -2, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 2, 2, 1, 2, 0, 0, 0, 0, 0, 0, -1, -3, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, -1, -1, -2, -1, -1, 0, -2, -1, -1, -2, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, 0, -1, -1, -1, -2, -3, -1, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 3, 3, 3, 4, 3, 3, 3, 4, 5, 5, 7, 5, 4, 1, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 1, 1, 2, 2, 1, 2, 1, 0, 1, 3, 2, 2, 2, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, -1, -2, 0, -1, 0, 1, 0, 1, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, -1, -1, 0, -1, -1, -2, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, 0, -3, -3, -3, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 2, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, -2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 2, 2, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -1, 0, 0, -1, -1, 0, 0, 1, 1, 2, 2, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -1, -2, -1, 0, -1, -1, 1, 0, 1, 3, 2, 1, 3, 1, 0, 2, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, 1, 0, 0, 1, 2, 1, 2, 2, 3, 2, 1, 0, 2, 0, -1, -1, 0, 1, -1, 0, 0, 0, -2, -1, -2, -1, 0, 0, 0, 0, 1, 0, 0, 2, 0, 1, 1, 1, 0, -1, 0, -2, 0, -1, -1, -2, -1, -1, -2, -1, 0, -1, -1, -2, 0, 1, 0, 2, 1, 2, 2, 0, 2, 1, 0, 0, -1, 0, 0, -1, 0, -1, -1, -2, -2, -2, 0, 0, -1, 0, 0, 0, 0, 1, 0, 2, 2, 0, 2, 1, 0, 0, 0, 0, 0, -1, 0, -2, -2, -3, -1, -1, 0, -1, 0, 0, 0, 1, 0, 2, 1, 2, 1, 2, 1, 0, 0, 0, 1, 1, 0, 0, -1, 0, -2, -3, -3, -2, -1, -1, 1, 1, 0, 2, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -3, -1, -2, -3, -2, -2, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -2, -3, -3, -2, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, -1, -1, -2, -3, -1, -2, -1, -1, 0, -2, 0, 0, 0, 1, 0, 0, 0, 0, 2, 1, 1, 1, 2, 1, 0, -1, -1, -1, -1, -3, -4, -2, -1, -1, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 0, 0, 1, 0, -1, -1, 0, -2, -2, -2, -2, -1, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 2, 1, 2, 0, 0, 0, -1, -1, -3, -1, -2, -2, -1, -1, -1, 0, -1, -2, 0, 0, 1, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -2, 0, -2, -2, -1, 0, -1, 0, 2, 3, 2, 1, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, -2, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, -3, -3, -2, -1, 0, -1, -3, -3, -1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -5, -4, -5, -3, -3, -3, 0, -1, -1, 0, 0, 2, 4, 6, -1, -1, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, -2, -2, -2, -3, -2, -2, -1, -2, 0, -1, 0, 0, 2, 4, -3, -1, -1, -1, 0, -2, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, 1, 4, 0, -1, 0, -1, 0, -1, -1, 0, 0, 1, 2, 2, 2, 1, 1, 1, -1, -2, -1, -2, -1, 0, 0, 1, 2, 4, 0, 1, 0, 0, 0, -2, -2, -2, -1, 1, 1, 3, 3, 3, 1, 1, 1, 0, 0, 0, -1, 0, 0, 1, 2, 4, 0, 1, 0, 0, 0, -4, -3, -2, 0, 2, 2, 2, 4, 3, 3, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 3, 0, 0, 0, 0, -3, -2, -5, -2, -1, 0, 2, 4, 5, 4, 4, 1, 2, 1, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, -3, -3, -2, -1, 2, 2, 2, 5, 5, 3, 3, 3, 3, 1, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -3, -1, -2, 0, 1, 3, 5, 5, 5, 3, 2, 3, 0, 1, 0, -1, -2, -2, -1, -2, 0, -2, 0, 0, 0, -1, 0, -2, 0, 0, 2, 3, 4, 5, 4, 4, 1, 1, 0, -1, -2, -2, -4, -4, -2, -1, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 2, 4, 4, 4, 5, 2, 2, 0, 0, 0, -2, -1, -2, -3, -3, -2, 0, -3, -2, -1, -1, 0, 0, 0, 0, 0, 3, 6, 5, 5, 4, 2, 2, 1, -1, -2, -2, -2, -2, -3, -2, -2, 0, -2, -1, 0, 0, 0, 0, 0, 0, 2, 3, 5, 5, 4, 5, 3, 3, 0, -1, -1, -2, -1, -3, -3, -4, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 2, 3, 5, 5, 5, 4, 4, 1, 1, 0, -1, -2, -1, -4, -3, -3, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 4, 4, 6, 6, 4, 4, 2, 1, 1, -1, -1, -1, -2, -4, -4, -2, 1, -1, 0, 1, 1, 0, 1, 1, 0, 0, 2, 4, 6, 6, 4, 3, 3, 1, 0, 0, -1, -2, -4, -4, -3, -1, 0, -1, 0, 1, 1, 1, 0, -1, -2, 0, 1, 4, 4, 5, 4, 3, 2, 0, 1, 0, 0, -2, -3, -2, -1, 0, 3, 0, 1, 0, 0, -1, 0, -2, -1, -1, 2, 3, 3, 4, 4, 1, 1, 2, 0, -1, -1, -1, -2, -3, -1, 0, 2, 0, 0, 0, 0, -2, -2, -3, -2, -1, 0, 4, 4, 3, 3, 2, 2, 0, 0, 0, 0, -2, -2, -1, -1, 1, 3, 0, 0, 0, 0, -1, -1, -3, -2, -1, 1, 4, 3, 3, 4, 1, 2, 0, 0, -1, 0, -1, -3, -1, 0, 3, 4, 0, 0, -1, 0, -2, -3, -3, 0, -1, 0, 3, 2, 1, 2, 1, 0, 0, -1, 0, -1, -2, -3, -2, 0, 2, 5, -1, 0, -1, -1, -2, -2, -2, 0, 0, 1, 1, 3, 2, 2, 0, 0, -1, -1, -3, -2, -2, -4, -2, 0, 2, 6, -1, -1, -1, -2, -3, -3, 0, 0, 1, 0, 1, 2, 0, 1, -1, -1, -2, -2, -4, -2, -4, -3, -1, -1, 3, 6, -1, -2, -1, -2, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -3, -4, -3, -2, -2, -3, -1, -1, 2, 5, -3, -3, -1, 0, -2, -2, 0, 0, 0, 0, 0, -1, -1, -2, -3, -2, -3, -3, -2, -3, -2, 0, 0, 0, 2, 7, -3, -3, -3, -2, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -3, -3, -3, 0, -1, 0, 1, 2, 1, 3, 5, 8, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -2, -3, -1, -1, 0, -1, 0, 0, -2, 0, -1, -2, -2, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, -1, -2, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, -1, -1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, -2, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 1, 1, -1, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -1, -2, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -1, -1, -1, 0, -2, 0, -1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -2, 0, -1, 0, -1, 0, -2, 0, 1, 0, -1, -1, -2, 0, 0, -1, -2, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, -1, -1, 0, -1, 0, -2, -1, 0, -1, -2, -1, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, -2, -1, -1, 0, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 1, 1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -2, -1, 0, -1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 1, 1, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, 0, 1, 0, 0, 0, -1, 0, -1, 0, -1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -2, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 1, 0, 0, 2, 2, 4, 3, 3, 4, 2, 2, 2, 0, 0, 0, -2, -3, -1, -1, -1, 0, -2, 0, 1, 2, 4, 1, 0, 0, 1, 0, 0, 2, 1, 2, 3, 3, 3, 2, 1, -1, -2, -3, -3, -2, -1, -2, -1, -1, 0, 0, 3, 2, 0, 0, 0, 1, 0, 0, 0, 2, 2, 3, 3, 1, 0, 0, 0, -1, -3, -4, -2, -1, -2, 0, 0, 1, 3, 1, 0, 0, -1, -1, -1, -1, -2, 0, 2, 3, 3, 2, 2, 0, 0, -1, -3, -4, -3, -3, -3, 0, 0, 0, 1, 1, 2, 0, 1, -2, -2, -2, -2, -2, -1, 1, 2, 2, 2, 0, 0, 0, -2, -2, -4, -2, -2, -1, -1, 0, 1, 4, 2, 1, 0, -1, -1, -3, -5, -4, -1, 1, 2, 1, 2, 3, 1, 0, -1, -2, -3, -2, -3, -1, 0, 0, 1, 3, 4, 2, 0, 0, -1, -4, -4, -2, -1, 1, 0, 1, 2, 1, 0, 0, 0, -1, -1, -3, -4, -3, -3, 0, 0, 3, 1, 2, 0, 0, 0, -3, -4, -4, -2, 0, 0, 2, 2, 1, 0, 0, 0, 0, -1, -2, -2, -1, -2, -2, 0, 1, 1, 0, 0, 0, -2, -4, -5, -3, -1, 0, 1, 2, 2, 1, 1, 1, 0, 0, 0, -2, -3, -4, -3, -1, 0, -1, 0, 0, -1, 0, -2, -4, -4, -4, -3, 0, 1, 2, 3, 1, 0, 1, 1, 0, 0, -1, -2, -4, -2, -1, 0, 0, -1, -2, -1, -1, -3, -6, -5, -4, -3, 0, 2, 2, 3, 0, 1, 1, 1, 0, -1, -3, -2, -3, -2, -2, 0, -2, -2, -1, -2, -2, -3, -6, -5, -6, -2, 0, 1, 4, 1, 2, 0, 0, 0, -2, -2, -1, -3, -4, -2, -1, 0, -2, -2, -1, -1, -1, -4, -5, -6, -6, -4, 0, 1, 4, 2, 2, 1, 0, 0, 0, -2, -3, -4, -3, -3, -2, 0, -1, -1, -1, 0, -2, -5, -7, -7, -4, -2, 0, 2, 2, 3, 1, 0, 0, 0, 0, -1, -3, -3, -2, -2, -2, -1, -1, 0, 1, 1, -2, -4, -4, -5, -4, -2, -1, 1, 2, 2, 2, 1, 0, 0, 0, -2, -4, -5, -3, -2, -3, 0, -1, 0, 0, 1, 0, -3, -4, -5, -5, -2, -1, 2, 2, 2, 2, 0, 1, 1, 0, 0, -3, -4, -5, -3, -1, 1, 0, 1, 1, 1, -1, -4, -4, -4, -3, -3, -1, 1, 2, 3, 2, 0, 0, 0, -1, -1, -1, -3, -3, -3, 0, 0, 1, 2, 2, 0, 0, -4, -3, -3, -3, -3, 0, 1, 2, 1, 1, 0, 0, 0, -1, -1, -2, -4, -3, -2, 0, 2, 2, 2, 2, 1, 0, -2, -3, -3, -4, -1, 0, 2, 2, 2, 0, 0, 1, -1, 0, -1, -2, -2, -2, 0, 0, 3, 3, 2, 2, 2, -1, -2, -4, -3, -2, -2, 0, 1, 2, 2, 0, 0, 0, -2, -1, -2, -1, -2, -2, 0, 1, 2, 1, 2, 3, 1, -1, -1, -1, -2, -3, -1, 0, 3, 2, 2, 0, 0, -2, -3, -4, -2, -3, -3, -1, 0, 1, 2, 0, 1, 2, 0, 0, -1, -1, -1, 0, 0, 1, 2, 2, 1, 0, -1, -2, -3, -4, -4, -4, -1, -3, -1, 0, 3, 1, 0, 1, 0, 0, -1, -2, -1, 0, 2, 2, 1, 1, 1, -1, -1, -3, -4, -5, -5, -2, -2, -2, -1, 0, 3, 0, 0, 1, 0, 0, -2, -1, 1, 2, 3, 2, 3, 1, 0, -1, -2, -5, -5, -5, -5, -3, -3, -1, -1, 0, 1, 0, 0, 1, 2, 1, 0, 0, 1, 3, 3, 3, 1, 1, 0, 0, -4, -5, -5, -6, -4, -2, -1, 0, -1, 0, 3, -1, 0, 0, 3, 1, 0, 2, 2, 3, 2, 1, 1, 2, 0, 0, -1, -3, -4, -3, -1, 0, 2, 3, 1, 3, 5, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, -1, 0, 1, 0, 0, 0, -2, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -2, 0, -2, -1, 0, 0, -1, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, -2, -1, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -2, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 2, 1, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 1, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, -1, -2, 0, -2, -1, -1, 0, 0, 1, 0, 0, 2, 1, 2, 1, 0, -1, 0, 0, 0, 0, -1, -2, 0, -1, -1, 0, -2, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 0, 0, -1, -1, 0, -1, -1, -2, 0, -2, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -2, 0, 1, 1, 1, 0, 0, 1, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, -1, -1, -1, -1, -2, 0, -1, 1, 0, 0, 2, 1, 0, 1, 0, -1, 0, -1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 2, 2, 3, 3, 3, 2, 2, 2, 1, 2, 2, 3, 0, 0, -1, -3, -2, -5, -1, -2, -1, -1, 0, 0, -2, -1, 1, 2, 3, 3, 3, 3, 2, 2, 2, 2, 4, 2, 0, -1, -2, -2, -2, -3, -4, -2, 0, -1, 0, 0, 0, -2, 2, 3, 2, 1, 1, 1, 2, 1, 1, 2, 1, 2, -1, 0, -2, -1, -3, -3, -3, -2, -1, -2, 0, -2, -2, -2, 2, 1, 2, 3, 2, 1, 0, 0, 1, 1, 0, 0, -2, -2, -1, -2, -3, -3, -3, -1, -1, 0, 0, -2, -2, -1, 0, 0, 2, 2, 2, 2, 2, 1, 1, 0, -1, -2, -2, -4, -2, -1, -2, 0, -2, -3, -2, -1, -1, -1, -2, -1, 2, 1, 1, 2, 2, 1, 2, 0, 0, 0, -1, -3, -4, -3, 0, -1, 0, -1, -1, -1, -2, -1, 0, -1, -1, 0, 2, 2, 1, 2, 3, 0, 2, 0, 0, 0, 0, -1, -3, -2, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -2, 0, 2, 2, 2, 3, 2, 1, 1, 1, 0, 0, -2, -3, -2, -2, 0, 0, 0, 0, 1, 0, -1, -3, -2, -2, -3, -1, 1, 2, 2, 2, 2, 1, 1, 0, 0, -1, -1, -3, -4, -2, 0, 0, 0, 0, 0, -1, -3, -4, -4, -3, -1, -1, 2, 2, 2, 2, 0, 2, 2, 0, 0, 0, -3, -3, -3, -2, -1, 0, 0, 1, 0, -1, -2, -3, -5, -4, -1, -3, 3, 1, 3, 3, 0, 0, 2, 0, 0, -1, -2, -3, -2, -3, -1, 0, 0, 0, 1, 0, -1, -3, -4, -3, -4, -4, 3, 1, 1, 2, 1, 1, 1, 0, -1, -1, -4, -3, -3, -2, -2, 0, 0, 1, 2, 1, -2, -4, -7, -6, -6, -4, 2, 1, 2, 1, 2, 1, 0, 0, -2, -1, -2, -2, -4, -3, -3, -2, 1, 0, 0, 0, -2, -5, -7, -6, -5, -6, 1, 0, 1, 0, 1, 0, 0, -1, -3, -2, -4, -2, -2, -2, -3, 0, 0, 1, 1, -1, -2, -5, -6, -5, -6, -6, 3, 1, 1, 0, 0, 0, -2, -3, -3, -3, -3, -3, -4, -4, -2, 0, 0, 0, 0, -1, -2, -5, -6, -6, -6, -5, 2, 1, 1, 1, 1, 0, -2, -1, -3, -4, -4, -4, -3, -3, -2, -1, 2, 2, 1, 0, -2, -3, -6, -6, -6, -6, 0, 1, 1, 1, 2, 1, 0, -1, -2, -2, -3, -4, -3, -1, -1, 0, 2, 2, 0, -1, -1, -3, -6, -4, -5, -6, 1, 0, 3, 3, 1, 0, 1, 0, -2, -3, -4, -2, -2, -2, -1, 1, 0, 0, 1, 0, 0, -3, -5, -5, -3, -5, 1, 2, 4, 5, 2, 1, 0, 0, -2, -3, -1, -2, -2, -2, 0, 0, 2, 0, 1, -1, -1, -3, -3, -4, -5, -5, 3, 3, 4, 3, 3, 3, 0, 0, -2, -3, -3, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -3, -3, -3, -5, -4, 3, 3, 3, 3, 3, 2, 1, 0, -1, -2, -1, -2, 0, -1, 0, 1, 0, -1, -1, -1, -1, -3, -3, -4, -4, -3, 0, 1, 2, 4, 2, 4, 3, 0, 0, -2, -3, -1, -2, -1, 0, 0, 0, -1, -2, -3, -2, -2, -4, -2, -4, -2, 0, 1, 2, 2, 3, 2, 2, 1, 0, 0, 0, -1, -2, 0, 0, -1, -1, -1, -3, -2, -2, -3, -3, -2, -2, -4, 0, 2, 2, 2, 1, 4, 3, 2, 1, 0, -1, -2, -4, -2, -3, -3, -3, -3, -3, -3, -2, 0, -1, -1, -4, -4, 0, 0, 1, 0, 2, 2, 3, 3, 3, 1, 2, -1, -2, -3, -4, -4, -4, -4, -4, -5, -1, 0, -1, -2, -2, -3, 0, 0, 1, 1, 1, 1, 0, 2, 2, 2, 2, 1, 0, -2, -4, -4, -5, -5, -5, -4, -3, -2, -3, -2, -3, -4, 3, 1, 2, 2, 1, 1, 0, 0, 2, 2, 2, 0, 1, 0, -3, -3, -3, -3, -3, -4, -2, -2, -3, -1, 0, 0, 2, 2, 1, 1, 0, 1, 0, 0, 2, 3, 2, 2, 0, 0, -2, -2, -3, -3, -3, -3, -2, -3, -1, -1, -2, -1, 1, 0, 0, 0, 0, -1, 0, 0, 2, 3, 3, 3, 1, 0, -1, -1, -3, -3, -3, -3, -2, -1, -1, 0, 0, -2, 2, 2, 0, 0, 0, -1, 0, 0, 1, 3, 2, 2, 2, 0, 0, 0, -2, -3, -3, -2, -2, -1, 0, -1, 0, -1, 1, 2, 0, 0, 1, 0, -1, -1, 0, 2, 1, 1, 0, 1, 1, 0, 0, -1, -2, -2, -2, -2, 0, -2, -1, 0, 2, 0, 1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, -2, -2, -2, -3, -1, -1, -2, -1, 2, 1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, -1, -1, -2, -2, -2, -3, -1, 0, 0, 0, 0, 0, -1, -2, -2, -1, 0, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, -1, -2, -3, -1, -1, -1, -1, 0, 0, 0, 0, -1, -2, -3, -2, 0, 0, 0, 1, 2, 2, 0, 1, 1, 1, -1, -1, -2, -2, -3, -3, -2, -2, -1, 0, 0, 0, -1, -3, -2, -3, -2, 0, 0, 3, 4, 2, 1, 1, 0, 1, 0, -1, 0, -2, -2, -3, -3, -3, -1, -1, 0, 0, -2, -4, -5, -4, -1, 0, 1, 3, 2, 1, 1, 1, 0, 1, -1, -1, -1, -3, -4, -3, -1, -1, 0, 0, 0, -1, -2, -4, -5, -5, -3, -1, 0, 3, 4, 2, 0, 1, 0, -1, -1, -2, -3, -3, -3, -4, -4, -2, -1, 0, -1, -2, -3, -6, -5, -4, -3, -1, 1, 3, 3, 1, 1, 0, 1, 0, 0, -2, -3, -3, -5, -4, -3, -2, 0, 0, -2, -2, -4, -5, -3, -5, -3, 0, 1, 3, 2, 2, 2, 1, 1, 0, -1, -2, -4, -3, -5, -3, -3, -1, 0, 0, -2, -3, -2, -3, -4, -3, -3, 0, 1, 1, 2, 1, 2, 1, 0, 0, -1, -1, -2, -5, -5, -5, -4, -2, 0, 0, -1, -2, -2, -4, -3, -2, -2, -1, 0, 3, 1, 2, 1, 1, 0, 0, 0, 0, -1, -4, -4, -3, -2, -1, 0, 0, 0, 0, -2, -3, -2, -2, -1, -1, 0, 2, 1, 2, 2, 0, 0, 0, 0, -1, -2, -4, -3, -1, -1, -1, 1, 1, 0, -1, 0, -2, -2, -1, 0, 0, 0, 3, 3, 3, 1, 0, 1, 1, 1, -2, -3, -3, -3, -2, -1, -1, 1, 2, 1, 1, 0, -1, -2, 0, 0, 1, 2, 2, 3, 2, 3, 0, 0, 1, 0, 0, -2, -1, -2, -1, 0, 0, 0, 2, 0, 1, 0, 0, 0, -1, 0, 1, 1, 4, 2, 3, 1, 0, 0, 0, 0, -2, -1, -2, -2, -1, -1, -1, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 2, 3, 2, 2, 0, -1, -1, 0, -2, -1, -3, -1, -3, -1, -3, -2, 0, -1, 0, -1, 0, 0, 0, 0, 2, 2, 2, 3, 1, 1, 0, -1, -2, -2, -2, -2, -1, -1, -4, -2, -3, -1, 0, -1, -1, 0, 0, 0, 0, 1, 3, 2, 2, 1, 0, -1, -1, -2, -3, -2, -3, -2, -3, -2, -3, -2, -3, -2, 0, 0, 0, 0, 0, 1, 1, 1, 3, 3, 2, 1, 0, -2, -3, -2, -3, -2, -2, -2, -2, -2, -2, -2, -3, -1, 0, 0, 0, 0, 1, 1, 2, 3, 2, 3, 2, 1, 0, 0, -2, -3, -3, -4, -3, -4, -2, -2, 0, -2, -1, 0, 1, 0, 0, 0, 1, 1, 2, 4, 2, 3, 1, 1, 0, 0, -3, -2, -4, -2, -2, -3, -1, 0, 0, 0, 0, 0, 1, 1, -2, -4, -2, 0, 0, 1, 2, 4, 5, 8, 5, 1, -1, -1, 0, 1, 0, 1, 4, 3, 2, 0, 0, 0, 0, 0, -1, -3, -1, 0, 2, 1, 4, 5, 7, 8, 6, 3, 2, 0, 1, 1, 2, 4, 5, 6, 2, 2, 0, -1, 1, -1, -2, -1, -1, 0, 0, 3, 3, 4, 8, 9, 5, 3, 4, 3, 2, 3, 2, 3, 5, 5, 5, 3, 1, 0, 2, 1, 0, -2, 0, 0, 2, 3, 3, 6, 7, 7, 5, 3, 3, 3, 2, 3, 2, 5, 5, 4, 3, 3, 3, -1, 0, 1, 0, 0, -1, 0, 0, 4, 3, 6, 7, 6, 5, 4, 2, 3, 2, 2, 1, 2, 5, 5, 4, 3, 2, 0, 1, 2, 0, -1, 0, 0, 2, 4, 3, 4, 8, 8, 6, 4, 4, 3, 3, 2, 3, 4, 5, 5, 4, 2, 1, -1, 0, 2, 1, 0, 0, 1, 3, 5, 5, 5, 7, 7, 6, 5, 5, 3, 3, 2, 4, 4, 5, 4, 3, 3, 3, -1, 1, 3, 0, 0, 0, 0, 3, 4, 5, 5, 6, 8, 7, 6, 7, 4, 3, 1, 2, 3, 5, 4, 5, 5, 2, 0, 0, 0, 0, 0, 0, 1, 4, 4, 4, 6, 8, 9, 7, 8, 6, 3, 1, 0, 0, 3, 4, 4, 5, 4, 4, 0, 0, 1, -2, -1, 0, 0, 3, 4, 5, 7, 8, 10, 9, 8, 5, 1, 1, 0, 0, 3, 3, 5, 6, 6, 3, 0, 0, 0, -1, 0, 0, 0, 2, 3, 5, 5, 8, 7, 10, 10, 5, 1, 2, 0, 0, 0, 2, 5, 7, 7, 5, 1, 0, -1, -1, 0, 0, 1, 2, 3, 5, 4, 5, 8, 9, 10, 6, 4, 2, 1, 0, 1, 0, 2, 5, 5, 5, 2, 0, 0, 0, 0, 2, 3, 2, 3, 2, 5, 5, 6, 11, 10, 6, 4, 3, 1, 3, 0, 1, 3, 4, 5, 5, 4, -1, -2, 0, 2, 3, 3, 4, 2, 2, 6, 7, 8, 10, 9, 6, 3, 3, 1, 2, 1, 1, 1, 4, 6, 6, 2, -2, -1, 0, 1, 4, 3, 4, 4, 4, 3, 4, 6, 9, 7, 5, 3, 0, 3, 2, 3, 3, 4, 6, 6, 6, 3, -1, -2, 0, 3, 3, 3, 3, 4, 5, 3, 4, 7, 8, 7, 3, 2, 0, 0, 2, 4, 3, 4, 5, 5, 5, 1, -3, 0, 1, 1, 1, 3, 3, 3, 3, 4, 3, 7, 4, 6, 3, 0, 0, 0, 1, 3, 4, 5, 5, 6, 4, 2, -1, 1, 1, 3, 0, 3, 5, 5, 3, 4, 4, 6, 5, 5, 5, 0, -1, 0, 0, 3, 3, 4, 4, 5, 2, 1, -2, 1, 2, 1, 1, 2, 4, 5, 5, 3, 4, 6, 8, 4, 3, 1, 0, -1, 0, 2, 3, 3, 2, 3, 2, 0, -2, 0, 1, 1, 2, 3, 4, 5, 6, 3, 6, 5, 6, 4, 1, 1, 1, 0, 0, 1, 5, 4, 2, 3, 0, -1, -1, 1, 2, 1, 1, 3, 4, 6, 4, 4, 4, 7, 6, 4, 1, 1, 1, 0, 0, 0, 3, 5, 3, 1, -1, -2, -1, 0, 1, 2, 0, 2, 3, 5, 3, 5, 5, 5, 4, 4, 1, 1, 2, 0, 0, 0, 3, 5, 3, 0, 0, -1, -1, 0, 1, 2, 1, 0, 1, 1, 4, 5, 6, 6, 5, 2, 3, 1, 1, 0, 0, 1, 3, 5, 4, 1, -2, -4, 0, 0, 1, 2, 1, 0, 0, 0, 2, 5, 7, 6, 4, 4, 3, 2, 2, 0, 0, 1, 3, 5, 2, 0, -1, -2, 0, -1, 1, 2, 1, -1, 0, 0, 2, 5, 5, 6, 5, 3, 1, 3, 2, 0, 2, 2, 4, 3, 1, 0, -3, -2, -2, 0, 0, 0, 0, 0, 0, 0, 3, 6, 5, 4, 5, 2, 2, 4, 3, 2, 1, 3, 2, 2, 2, 0, -2, -3, -1, 0, -1, -2, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 2, 0, 2, 2, 1, 2, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -2, -1, -2, -2, -1, -1, 0, -1, -2, 0, -1, -1, -1, -1, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, -2, -1, 0, -2, -2, -3, -2, -2, -1, -2, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, 0, -2, -3, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, -2, -1, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -2, -1, -2, -1, -1, 0, -1, 0, 1, 1, 0, 2, 1, 0, 1, 0, 0, -1, -1, -2, -1, 0, -1, -2, -1, -2, -2, -2, -2, 0, 0, 0, 0, 0, 1, 2, 0, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, 1, 0, 1, 1, 1, 2, 1, 2, 2, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 1, 1, 1, 0, 2, 2, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 0, 1, 1, 0, -1, -1, -1, -1, -1, -1, -1, -2, -1, 0, 0, 1, 1, 0, -1, -1, -1, 0, 0, -1, 1, 1, 1, 0, 0, 0, -2, -2, 0, -2, -2, 0, -2, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 2, 1, 1, 1, 1, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 3, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 1, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 1, 1, -1, -2, -1, 0, 0, 0, 1, 1, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, 0, -1, 0, -2, -2, 0, 0, 0, 0, 0, 1, 1, 2, 0, -1, 1, 1, 0, 1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, -2, -1, 0, 0, 1, 1, 1, 1, 0, 2, 0, -1, 1, 0, 1, 0, 0, 0, -1, -1, -1, -1, -2, -2, 0, -1, 0, 0, 0, 0, 1, 0, 1, 2, 0, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, -1, 0, 0, 0, 1, -1, 0, -1, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, 0, 1, 2, 1, 1, 2, 1, 1, 0, 2, 2, 2, 1, 0, 0, -2, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 1, 1, 3, 2, 2, 0, 0, 0, 0, 0, -1, -1, 0, -2, -2, 1, 3, 1, 2, 0, 1, 0, 0, 1, 0, 1, 0, -1, 0, -1, -3, -1, -2, 0, -1, 0, 0, 0, -1, -1, -1, 3, 2, 1, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -2, 2, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 3, 2, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, 2, 0, 2, 2, 2, 1, 2, 0, 0, 1, 0, 0, -2, -2, 1, 1, 0, 0, 0, 0, 0, -1, 1, 2, 2, 3, 2, 2, 2, 3, 3, 2, 1, 1, 1, 0, 0, 0, -2, -1, 2, 2, 0, 1, 0, 0, -1, 0, 1, 1, 1, 1, 2, 2, 1, 2, 3, 2, 1, 2, 1, 0, 0, -1, 0, -2, 1, 1, 1, 0, -1, -2, -1, 0, 0, 0, 0, 1, 0, 1, 3, 1, 1, 2, 3, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, -2, -2, 0, 0, 0, 0, 1, 3, 3, 2, 1, 3, 1, 2, 1, 1, 1, 0, 0, -1, -2, 1, 0, -1, -1, -2, -2, -3, -1, 0, 0, 1, 1, 3, 1, 1, 0, 2, 0, 2, 0, 2, 2, 1, 0, -1, -1, 2, -1, -1, 0, -1, -4, -3, -2, 0, 0, 1, 2, 3, 3, 3, 2, 1, 2, 1, 0, 2, 0, 0, 0, -2, -2, 1, 0, -2, -1, -2, -2, -4, -2, -1, -1, 1, 2, 1, 1, 0, 1, 1, 0, 0, 2, 0, 0, 1, 0, 0, -1, 1, 0, -1, -1, -3, -4, -4, -2, -1, 0, 0, 1, 1, 3, 1, 0, 1, 1, 2, 1, 0, 0, 0, 0, -1, -2, 0, 0, 0, -2, -2, -4, -3, -3, -1, 0, 0, 2, 2, 3, 1, 0, 1, 0, 3, 1, 0, 0, -2, -2, -1, -2, 0, 0, 0, -2, -3, -3, -4, -2, -1, 0, 2, 2, 2, 1, 2, 2, 1, 2, 2, 1, 0, 0, 0, -2, -1, -1, 0, 0, -2, -3, -4, -4, -2, -1, -1, 0, 0, 2, 3, 2, 1, 1, 1, 2, 2, 3, 0, 0, -1, -1, -2, 0, 1, 0, -2, -1, -3, -4, -3, -3, -1, 0, 0, 2, 1, 0, 0, 1, 2, 3, 3, 1, 1, 0, 0, 0, -2, -1, 1, 0, -1, -2, -3, -3, -2, -2, -2, 1, 2, 1, 3, 2, 0, 1, 2, 2, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -2, -1, 0, 1, 4, 3, 1, 2, 2, 2, 4, 3, 2, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 2, 4, 3, 4, 2, 2, 2, 3, 2, 2, 1, 1, -1, 0, -2, -2, 1, 0, 1, 0, 0, -1, -1, -1, -1, 1, 1, 3, 4, 4, 3, 2, 2, 1, 1, 1, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, -2, 0, -1, 0, 1, 3, 2, 4, 2, 2, 3, 3, 0, 1, 1, 0, -1, 0, -2, -3, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 2, 1, 1, 0, 1, 0, 0, -1, 0, -1, 0, -2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 1, 1, 0, 2, 0, 1, 0, 1, -1, 0, 1, 1, 0, 1, -1, 0, -2, -2, -2, -2, -1, -2, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -2, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, 2, 2, 2, 2, 2, 0, 0, 0, -2, -1, -1, 0, -1, -2, -1, -1, -1, 0, 0, 0, -1, -2, 0, 2, 4, 5, 4, 5, 4, 3, 0, -3, -3, -2, -2, -1, -1, 0, 0, 0, -1, 2, 2, 3, 8, 12, 15, 0, 0, 1, 1, 1, 3, 3, 2, 3, 2, 0, 0, 0, -1, -2, -2, -2, 0, -1, -1, 0, -1, 2, 3, 7, 13, -1, -1, 0, 0, 0, 0, 0, 3, 2, 3, 3, 2, 1, 0, 0, -2, -1, -1, -2, -3, -1, 0, 0, 2, 6, 10, 0, -1, 1, 0, -1, -1, 0, 0, 1, 3, 2, 5, 4, 2, 0, -1, -1, -1, -3, -3, -1, -2, 0, 0, 3, 8, 0, 0, 1, 0, -2, -3, -2, 0, 3, 2, 4, 5, 5, 4, 2, -1, -2, -1, -2, -1, -1, 0, 0, 0, 3, 8, 3, 1, 1, -2, -5, -5, -4, 0, 1, 2, 5, 6, 5, 5, 3, 0, -2, -2, -3, -3, -3, 0, 0, 0, 3, 5, 3, 1, 0, -1, -5, -6, -3, -1, 1, 3, 5, 7, 7, 5, 4, 0, 0, -1, -2, -4, -1, -2, -1, 0, 2, 4, 2, 1, -1, -2, -3, -4, -4, 0, 1, 3, 5, 5, 6, 4, 4, 1, 1, 0, -1, -4, -2, -2, 0, 0, 0, 3, 2, 1, -1, -2, -3, -3, -4, -1, 1, 4, 4, 5, 5, 6, 4, 3, 1, 0, 0, -3, -3, -2, 0, -1, 0, 1, 1, 0, 0, -2, -2, -2, -2, 0, 1, 5, 5, 6, 7, 6, 6, 4, 1, 0, -1, -3, -3, -4, -1, 0, 0, 2, -1, 0, -1, 0, -3, -3, -1, 0, 2, 7, 6, 7, 6, 7, 4, 4, 2, -1, 0, -4, -3, -2, -2, -1, 0, 2, -2, -1, 0, -1, -3, -3, -2, 0, 2, 6, 7, 9, 8, 6, 3, 3, 0, 0, -3, -4, -4, -2, -3, -3, -1, 2, 0, 0, -1, -2, -2, -2, -2, 0, 4, 7, 9, 9, 7, 6, 4, 1, 1, -1, -2, -2, -2, -4, -3, -3, 0, 2, 0, 1, 0, -2, -5, -4, -1, 0, 4, 6, 9, 9, 8, 6, 4, 2, 0, -3, -2, -2, -4, -4, -4, -1, 0, 3, 0, 1, 0, -1, -4, -2, -1, 0, 3, 5, 7, 8, 8, 4, 3, 4, 1, -2, -2, -3, -3, -3, -5, -1, 0, 5, 1, 1, 1, -2, -2, -4, -2, 0, 2, 4, 6, 8, 7, 5, 3, 2, 1, 0, -2, -3, -3, -3, -4, -1, 0, 5, 3, 2, 0, -1, -3, -4, -3, -1, 0, 3, 7, 6, 4, 3, 2, 2, 1, 0, -2, -2, -2, -2, -2, -1, 2, 6, 3, 2, 1, 0, -4, -4, -3, -2, 1, 2, 5, 5, 5, 1, 4, 3, 2, 1, -2, -3, -3, -1, -2, -1, 2, 7, 4, 3, 0, -1, -6, -5, -4, -2, 0, 3, 5, 6, 3, 2, 1, 3, 1, 0, 0, -2, -3, -2, -1, 0, 4, 10, 4, 2, 1, -2, -4, -7, -4, -4, 0, 3, 4, 5, 4, 3, 3, 3, 1, -1, -1, -3, -2, -1, -1, 2, 4, 10, 4, 1, -1, -3, -5, -5, -3, -2, 0, 4, 5, 6, 3, 3, 1, 1, 0, 0, -3, -1, -1, 0, 0, 1, 6, 12, 1, 1, -1, -2, -3, -4, -2, 0, 2, 3, 5, 5, 3, 4, 1, 0, -2, -3, -2, -2, -2, -1, -1, 2, 7, 13, 0, 0, -1, -2, -4, -2, -1, 0, 2, 5, 4, 3, 3, 1, 0, -2, -2, -2, -5, -3, -3, -3, -2, 1, 8, 12, 1, 0, -2, -2, -2, 0, 0, 2, 3, 4, 4, 2, 1, 0, -1, -3, -4, -5, -4, -2, -3, -4, -1, 2, 8, 13, 1, 0, 0, -1, -1, 1, 3, 4, 5, 4, 2, 1, 0, 0, -2, -5, -4, -4, -3, -2, -3, -4, -1, 3, 8, 14, 0, 0, 0, 0, 0, 1, 3, 3, 3, 3, 1, 0, 0, -2, -3, -5, -2, -2, 0, 0, 0, 0, 0, 6, 11, 17, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, -1, -1, -1, 0, 0, 1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 4, 4, 3, 3, 2, 1, -1, 0, 0, 0, -1, -2, 0, 0, -1, -1, -1, 0, 0, 1, 1, 2, 0, 0, 2, 1, 1, 1, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, -2, -2, -3, 0, 0, 0, 0, 1, 2, 0, 0, 2, 2, 1, 0, 0, 0, 1, 0, 2, 1, 0, 0, -1, 0, -1, 0, -1, -2, -2, 0, 0, 0, 1, 2, 0, 1, 2, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -2, -2, -1, -2, -1, 0, 0, 2, 3, 1, 0, 0, 0, 0, -2, -1, -1, 0, 1, 0, 1, 0, 0, -1, -1, 0, -3, -2, -3, -1, -1, 0, 0, 1, 2, 2, 2, 1, 1, 0, -2, -2, -1, 0, 0, 0, 0, 1, 0, 0, -1, -2, -1, -2, -1, -1, 0, 0, 0, 0, 1, 3, 0, 0, 0, -2, -2, -1, -2, 0, -1, 0, 1, 0, 0, 0, -1, -1, -2, -2, -2, -2, -2, -1, 0, 0, 1, 0, 2, 0, -1, -2, -2, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, -2, 0, 0, 0, 0, 1, 1, 1, 0, -2, -3, -3, -1, -2, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, -1, -2, -1, 1, 0, 0, 0, 0, 0, 0, 0, -2, -3, -2, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 1, 1, 0, -1, -1, -1, -2, -4, -4, -3, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, -2, -3, -3, -3, -4, -2, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -2, -3, -4, -2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, 0, -1, 0, -1, -1, 0, 1, 0, 0, 0, -1, -3, -5, -5, -3, -2, -1, 0, 0, 0, 0, -1, 0, 0, -2, 0, -1, -2, -1, 0, 0, 0, 1, 0, 0, 0, -1, -3, -5, -4, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 1, 0, 1, 0, 0, -1, -4, -3, -3, -3, -2, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, 1, 0, 1, 1, 2, -1, -1, -2, -4, -5, -3, 0, 0, 0, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, -2, 0, 0, 2, 2, 1, 1, 0, -2, -3, -5, -4, -2, -3, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 2, 3, 0, 0, -2, -4, -3, -4, -3, -1, -2, 1, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 4, 2, 1, 0, 0, -4, -4, -5, -3, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, -1, 0, 0, 0, 1, 0, 2, 3, 1, 0, -1, -1, -1, -4, -3, -1, 0, 0, 2, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 3, 0, 1, -1, -1, -1, -3, -2, 0, 0, 0, 2, 1, 1, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 2, 3, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 1, 1, 2, 1, 2, 1, 0, -1, 0, 0, 1, 1, 1, 2, 1, 0, 1, -1, -3, -1, -2, -3, -1, -1, 0, 0, 0, 0, 3, 0, 0, 1, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, -2, -3, -1, -3, -2, 0, 0, 0, 0, 0, 0, 3, 0, 1, 0, 1, 0, 1, 3, 2, 2, 1, 0, 0, -1, -1, -1, -3, -2, -2, 0, 0, 0, 0, 0, 1, 2, 5, 6, 7, 7, 6, 5, 3, 4, 5, 4, 5, 1, 0, -1, -1, -4, -4, -5, -5, -4, -2, -1, 0, 0, -1, -2, -4, 6, 5, 6, 6, 4, 2, 3, 3, 4, 1, 2, 1, 0, 0, -2, -2, -2, -3, -2, -1, 0, 2, 2, 2, -1, -3, 7, 6, 6, 6, 5, 4, 3, 3, 2, 2, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 1, 0, 1, -1, -3, 7, 5, 5, 4, 4, 2, 4, 2, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -2, -3, 6, 4, 5, 3, 3, 3, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, -1, -2, -2, 6, 5, 3, 3, 2, 1, 2, 1, 0, 0, 0, -2, -1, -2, 1, 1, 2, 1, 2, 3, 1, 1, 0, 0, -1, 0, 6, 4, 2, 2, 1, 0, 0, 0, 0, 0, -1, -2, -3, -1, 0, 1, 3, 2, 1, 3, 1, 1, -1, -1, 0, 0, 5, 3, 2, 1, 2, 0, 0, 0, -1, -1, -3, -1, -1, -1, 0, 2, 1, 2, 4, 1, 2, 1, 0, 0, -1, 0, 6, 2, 2, 0, 1, 1, 0, 0, -2, -2, -2, -3, -1, -2, 0, 0, 1, 2, 1, 3, 0, 1, -1, 0, 1, 0, 6, 2, 2, 1, 1, 1, 0, -1, -2, -2, -3, -3, -3, -2, -1, 1, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, 4, 3, 1, 1, 0, 0, -2, -1, -3, -2, -4, -2, -3, -1, -1, 0, 1, 1, 1, 3, 0, 0, -1, 0, 0, 0, 5, 3, 0, 0, 0, -1, -1, -3, -2, -5, -3, -2, -4, -1, -2, 0, 0, 2, 2, 2, 0, 0, 0, -1, -2, -1, 5, 4, 1, 0, -2, -1, -3, -3, -3, -4, -4, -4, -2, -2, 0, 0, 1, 2, 2, 1, -1, -2, -1, -2, -2, -2, 4, 2, 0, 0, -2, -2, -4, -5, -5, -5, -5, -2, 0, -1, -1, 0, 1, 2, 3, 2, -1, -2, -4, -4, -2, -3, 6, 2, 0, 0, -1, -4, -3, -5, -6, -5, -3, -3, -3, -3, -2, 0, 1, 1, 3, 1, 1, -2, -3, -1, -2, -3, 5, 2, 0, 0, -1, -3, -4, -4, -4, -5, -3, -3, -3, -2, -1, -1, 0, 3, 2, 1, 0, 0, -3, -2, -2, -2, 4, 3, 2, 0, -1, -2, -3, -4, -3, -3, -4, -2, -2, -2, -1, 0, 0, 3, 3, 2, 2, 0, -1, -2, 0, -1, 3, 3, 3, 1, 1, 0, -1, -1, -4, -4, -4, -2, 0, 0, 0, 0, 1, 2, 3, 1, 0, 0, -1, 0, -1, -3, 6, 4, 2, 3, 0, 0, -2, -3, -3, -3, -3, -2, 1, 2, 1, 2, 2, 3, 3, 0, -1, -1, 0, 0, -2, -1, 6, 3, 4, 2, 2, 0, -2, -1, -3, -3, -4, -1, 0, 1, 1, 4, 3, 3, 0, 0, -1, 0, 0, -1, -2, -2, 5, 3, 3, 3, 1, 0, -1, -3, -2, -3, -4, -1, 0, 2, 2, 3, 3, 1, 0, 0, -2, -1, -1, -1, -2, -2, 5, 2, 2, 3, 2, 1, 0, 0, -1, -4, -3, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, -1, 0, 0, -1, -3, 5, 4, 2, 2, 3, 3, 2, 0, 0, -3, -3, -3, -1, -1, 0, 1, 0, -1, -2, -3, -1, 0, 0, 0, -1, -3, 3, 3, 3, 3, 3, 3, 2, 3, 0, -1, -2, -4, -3, -2, -1, 0, -2, -3, -4, -2, -1, -2, 0, 0, 0, -3, 4, 3, 3, 4, 4, 5, 3, 3, 2, 0, 0, -2, -3, -3, -3, -4, -3, -5, -6, -3, -2, 0, -1, 0, 0, -2, 2, 3, 2, 5, 5, 3, 3, 3, 4, 3, 1, -1, -3, -3, -4, -4, -5, -5, -5, -5, -4, -1, -2, -2, -4, -3, 0, 2, 1, 2, 2, 1, 1, 1, 2, 2, 2, 1, 0, 0, -2, -2, -2, -2, -2, -1, -1, -1, -1, 0, 1, 0, 1, 0, 0, 1, 2, 0, 2, 3, 1, 3, 2, 1, 0, 0, -2, -3, -2, -1, -1, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 4, 4, 3, 2, 1, 0, -1, -2, -1, -2, -1, 0, 0, 0, 1, 0, 1, 0, 2, 1, 1, 0, 1, 0, 2, 3, 3, 3, 4, 2, 0, 0, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 3, 2, 3, 3, 2, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 1, 3, 2, 1, 2, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 1, 2, 3, 3, 2, 1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, -1, 0, 0, 2, 2, 1, 2, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, -1, 0, 1, 1, 2, 2, 1, 2, 2, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, -1, 0, 1, 2, 3, 1, 2, 3, 1, 0, 1, 0, 0, 0, -1, -1, -1, 1, 1, 0, 0, 2, 1, 0, -1, 0, 0, -1, 0, 0, 3, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, -1, -3, 0, -1, 1, 2, 2, 3, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, 0, 1, 2, 3, 2, 1, 0, 0, 0, 0, -1, -1, 0, -2, -1, 0, 0, 0, 1, 1, 0, -1, -1, -2, -3, 0, 0, 1, 3, 2, 3, 0, 0, 0, -1, 0, -1, -1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 1, 1, 3, 3, 3, 2, 1, 0, 0, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 2, 1, 3, 2, 1, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 2, 1, -1, 0, 0, 0, -1, 0, 1, 1, 2, 2, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 2, 2, 2, 1, 1, 2, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, 0, 0, 2, 3, 2, 4, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 1, 2, 2, 4, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 2, 2, 2, 3, 3, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 3, 3, 2, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 2, 1, 2, 2, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 1, 2, 2, 0, 1, 0, -2, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 3, 3, 1, 1, 0, 0, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 1, 2, 0, 1, 2, 1, 0, 0, -2, -1, 0, -1, -1, 0, -1, 0, -1, 0, 1, 0, -1, -2, -2, 0, 0, -1, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, -1, 0, 1, 0, 1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 1, 0, 1, 1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 2, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, 2, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 2, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -3, -2, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 2, -2, -1, 0, 0, 0, -1, 0, 0, 0, -2, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, -1, -2, -2, 0, 1, 0, 0, 1, 1, 3, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 2, 2, 2, 2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 2, 1, 1, 0, -1, 0, -1, 0, 0, 2, 1, 1, 0, 1, 1, 2, 1, 0, 1, 0, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 3, 2, 2, 0, 0, -1, -2, 0, -1, 0, 0, 0, 1, 0, -1, 0, -1, 0, 1, 2, 2, 2, 1, 3, 2, 3, 2, 2, 0, 1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 2, 3, 2, 2, 1, 2, 3, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 2, 3, 3, 1, 1, 2, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 2, 2, 4, 4, 4, 3, 3, 1, 1, 0, -1, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 2, 3, 3, 2, 3, 2, 1, 1, 2, 0, 0, -1, 0, -1, -2, -1, -1, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 1, 3, 2, 2, 2, 1, 1, 2, 1, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 2, 2, 2, 1, 2, 2, 1, 0, 0, 1, 0, 0, -1, -2, -1, -1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 2, 1, 2, 1, 2, 1, 0, 0, 0, -1, -2, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 3, 0, 2, 2, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 2, 0, 0, 1, 0, 0, 1, 1, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, -1, -1, 0, -1, -1, 0, 1, 1, 2, 2, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 3, 0, 0, 0, -1, 0, -2, -1, 0, 0, 1, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 3, 1, 1, -1, 0, 0, -1, 0, 0, 0, 2, 1, 1, 2, 1, 0, 1, -1, 0, -1, -1, 0, 0, 0, 0, 2, 4, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 2, -1, 0, -1, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, -1, -1, -1, 0, -1, -1, 0, -2, -2, 0, 1, 4, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -2, 0, 0, 3, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, -2, -1, 0, 0, 0, -1, 0, -2, 0, 0, 2, 4, 0, 0, -1, -1, 0, 2, 1, 1, 2, 3, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 5, 0, 0, 0, -1, 0, 1, 1, 0, 1, 1, 1, 1, 1, 0, 0, 0, -1, -2, -2, 0, -1, -1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, -2, -2, -1, 0, 0, -2, -2, 0, 0, 2, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, 2, 2, 0, 0, -1, 0, -2, -2, -1, -1, 0, -1, 0, 1, 1, 0, 1, 0, 0, -1, -1, -2, -1, 0, 1, 0, 2, 1, 0, 2, 0, 0, 0, -1, -2, 0, -2, -1, 0, 0, 1, 0, 2, 0, 0, 0, -1, -2, -1, -2, -1, 0, 1, 1, 1, 1, 1, 0, -1, -2, -2, -1, 0, 0, -1, 0, 0, 0, 2, 1, 0, 0, -2, -2, -2, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, -2, -3, -2, -2, -1, 0, 1, 1, 2, 0, 0, -1, 0, -3, -2, -3, 0, -1, 1, 2, 1, 2, 0, 0, 0, -1, -1, -2, -2, -2, -2, -1, 0, 1, 0, 1, 0, 0, 0, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -3, -1, 0, 0, 1, 0, 0, -1, 0, -3, -2, -2, -2, -1, 0, 2, 0, 2, 1, 1, 2, 0, 0, -1, -1, -3, -2, -1, 0, 0, 0, -1, -2, -1, -2, -3, -3, -3, -2, 0, 0, 1, 2, 0, 1, 0, 1, 1, 0, 0, -1, -1, -4, -1, -1, -1, -2, -2, -1, -1, -1, -2, -3, -3, -2, 0, 1, 1, 3, 2, 0, 1, 0, -1, -1, -1, -1, -3, -3, -1, -1, -1, -3, -2, 0, -2, -1, -3, -3, -4, -3, 0, 0, 1, 3, 1, 0, 1, -1, -1, -1, -2, -3, -3, -3, -2, 0, -1, 0, 0, 0, 0, -3, -3, -3, -2, -2, -1, 1, 1, 1, 1, 0, 1, 0, -1, -2, -2, -3, -4, -2, -2, 0, -1, 0, -1, 0, -1, -2, -3, -4, -2, -2, -1, 1, 2, 1, 3, 1, 0, 0, 0, -1, -1, -3, -3, -2, -1, 0, -2, 0, 0, 1, 0, -2, -3, -2, -2, -1, 0, 1, 1, 2, 1, 1, 0, 0, -1, 0, -2, -2, -3, -3, -1, -1, -1, 0, 0, 0, 0, -2, -1, -1, -2, -1, -1, 0, 1, 2, 1, 0, 1, 0, -1, -1, 0, -2, -3, -1, 0, 0, 0, 1, 1, 0, 0, -2, -2, -1, -1, -2, -1, 1, 2, 0, 1, 0, 1, 0, -1, 0, -1, -3, -3, -2, -1, 0, 0, 1, 2, 1, 0, -2, -3, -3, -3, -2, -1, 1, 1, 1, 0, 1, 0, 0, 0, -1, -2, -2, -3, -2, -1, 0, 0, 0, 1, 0, -1, -2, -1, -3, -2, -1, 0, 0, 1, 0, 0, -1, 0, -1, 0, -1, -2, -1, -1, -2, 0, 0, 1, 0, 1, 2, 0, -2, -2, -1, -1, -3, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, -2, -1, -2, -2, 0, 0, 0, 0, 0, 1, 0, -1, -3, -2, -2, -1, 0, 2, 1, 0, 1, 0, 0, -1, -1, -2, -2, -3, -2, -1, -1, 0, 0, 1, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 2, 1, 0, 0, -1, -1, -2, -3, -1, -1, -2, -1, -1, 0, 0, 0, 0, 1, -1, -2, -2, -1, 0, 0, 1, 2, 1, 0, 0, -1, -1, -3, -2, -2, -2, -1, -1, 0, -1, 1, 0, 0, 0, 1, 0, -1, 0, -1, 1, 2, 2, 0, 2, 0, 1, 0, -2, -2, -2, -2, -2, -2, -2, -2, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 1, 2, 1, 2, 0, 0, 0, -1, -2, -2, -2, -3, 0, -1, 0, 0, 0, 1, -3, 0, 0, 0, 0, 0, 0, -1, -2, -1, -3, -4, -2, -2, -4, -1, -2, -1, -1, 0, 0, 1, 1, 2, 3, 6, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -2, 0, -1, -1, -2, -2, 0, 0, 0, 0, 0, 1, 2, 4, -3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 3, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 1, 4, 0, 0, -1, 0, 0, 0, -1, 0, 0, 2, 2, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 5, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 5, 2, 2, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 2, 4, 0, -1, 0, 0, -1, 0, 0, 0, 1, 3, 3, 4, 3, 3, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 3, -1, 0, 0, 0, 0, -2, 0, 0, 1, 1, 2, 4, 4, 4, 3, 3, 2, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 4, 4, 2, 2, 3, 2, 0, 0, 0, 0, -1, -1, -1, -1, 2, -1, 0, 1, 0, 0, 0, 0, 1, 0, 2, 2, 3, 3, 4, 3, 2, 0, 0, 0, 0, -1, -2, -3, -2, -1, 0, -1, 0, 0, 2, 0, 1, 0, 0, 0, 2, 4, 3, 3, 3, 3, 2, 0, 0, -1, 0, -2, -4, -2, -3, -1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 2, 4, 4, 6, 3, 3, 1, 2, 1, 0, -1, -1, -2, -3, -2, -3, -1, -1, 0, 1, 1, 0, 2, 2, 1, 0, 3, 3, 4, 4, 4, 2, 2, 1, 0, 0, -2, -2, -3, -3, -4, -5, -4, -1, 0, 0, 2, 1, 0, 0, 1, 0, 2, 4, 5, 6, 3, 1, 2, 2, -1, -2, 0, -1, -2, -3, -4, -3, -3, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 3, 4, 5, 5, 2, 2, 1, 0, 0, 0, 0, -2, -3, -3, -4, -2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 2, 5, 5, 3, 3, 2, 2, 1, 0, -1, -1, -1, -2, -3, -2, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 4, 5, 6, 5, 2, 3, 3, 2, 0, 0, 0, -1, -1, -4, -3, 0, 1, 0, 0, 0, 1, 0, 1, 0, -1, 0, 2, 6, 6, 6, 4, 2, 2, 2, 0, 0, 0, -1, -3, -2, -1, 0, 3, 0, 0, 1, 0, 0, 0, -1, 0, 0, 3, 5, 5, 3, 4, 1, 1, 1, 0, 0, 0, 0, -2, -1, 0, 0, 2, 0, 0, 0, -1, 0, 0, -1, 0, 1, 3, 3, 4, 3, 2, 1, 1, 0, 0, -1, 0, -1, -1, -2, 0, 0, 3, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 3, 4, 3, 3, 2, 2, 0, 0, 0, 0, -2, -2, -1, 0, 2, 3, -1, -1, -1, -2, 0, -1, -2, 0, 0, 2, 2, 2, 2, 2, 1, 1, 0, 0, -1, -1, -2, -1, -1, 0, 1, 3, -1, -2, -1, -1, -2, 0, -1, 0, 0, 0, 0, 2, 1, 0, -1, -1, -1, -1, -2, -1, -1, -3, -2, 0, 3, 5, -1, -2, -1, -2, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, -2, -2, -4, -2, -2, -1, -2, -2, -1, 0, 3, 4, -2, -2, -1, -2, -1, -2, -2, -1, 0, 0, 0, 1, -1, -3, -4, -4, -4, -4, -1, -2, -2, -3, -1, 0, 2, 4, -3, -3, -2, -3, -3, -2, -1, -1, -1, 0, 0, 0, 0, -3, -3, -3, -3, -2, -2, -2, -1, -2, 0, 0, 4, 4, -8, -6, -5, -4, -4, -4, -4, -4, -4, -6, -4, -4, -6, -6, -8, -4, -4, -3, -2, -2, -2, -2, -2, -2, -1, -1, -7, -4, -2, -1, -2, 0, -2, -2, -3, -1, -1, -2, -1, -3, -4, -1, 0, -1, 0, 0, -2, 0, -1, -1, -1, -2, -5, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -3, -1, -1, -4, -1, -1, 0, 0, 0, 0, 2, 2, 2, 3, 2, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -2, -2, -2, -3, 0, 0, 0, 1, 1, 2, 2, 3, 3, 2, 2, 3, 2, 3, 2, 2, 0, 1, 0, 0, 1, 0, 0, -1, -3, -2, 0, 2, 0, 2, 2, 3, 5, 5, 5, 5, 3, 3, 3, 3, 3, 4, 1, 3, 0, 2, 0, 0, 0, 0, -3, 0, 0, 0, 0, 0, 2, 2, 4, 4, 5, 5, 6, 6, 4, 3, 3, 2, 1, 2, 2, 0, 1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 2, 4, 5, 4, 5, 5, 5, 7, 6, 4, 2, 1, 0, 1, 0, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 3, 5, 5, 5, 6, 6, 8, 6, 3, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 1, 2, 2, 3, 4, 5, 5, 6, 5, 7, 6, 5, 2, 1, 0, 1, 0, 1, 0, 0, 1, 0, -2, -2, -1, 0, 2, 1, 2, 4, 4, 6, 5, 5, 6, 8, 6, 5, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, 1, 3, 3, 4, 5, 6, 8, 7, 6, 7, 8, 6, 3, 1, 0, -2, -1, 0, 0, 0, 0, -1, -1, -3, -2, 0, 1, 2, 3, 6, 7, 7, 8, 8, 8, 7, 7, 7, 4, 2, 0, 0, -2, -3, -1, 0, 0, 0, -1, -3, -1, 1, 2, 3, 3, 5, 6, 6, 9, 8, 9, 8, 7, 7, 4, 2, 0, -2, -2, -2, 0, 0, 0, 0, -1, -4, -2, 0, 0, 1, 4, 3, 6, 5, 7, 6, 7, 7, 6, 7, 4, 2, 0, 0, 0, -1, 0, 0, 0, 0, -1, -4, -3, 0, 2, 2, 2, 4, 4, 5, 6, 7, 6, 7, 8, 6, 3, 3, 0, 0, 0, 0, 1, 0, -1, 0, -1, -6, -2, 0, 1, 3, 3, 3, 3, 5, 5, 4, 6, 7, 6, 6, 4, 2, 2, 1, 1, 0, 0, 0, 0, -1, -2, -5, -3, 0, 1, 1, 2, 3, 3, 6, 6, 4, 6, 7, 7, 7, 4, 2, 3, 2, 1, 0, 1, 0, -1, -1, -2, -5, -4, 0, 0, 2, 2, 2, 4, 5, 6, 5, 6, 6, 6, 5, 6, 3, 4, 2, 2, 2, 2, 0, -1, -3, -1, -6, -2, -1, 0, 2, 1, 1, 2, 4, 5, 6, 5, 7, 5, 4, 4, 4, 5, 3, 4, 3, 1, 0, -1, -2, -1, -5, -2, 0, 0, 2, 0, 0, 1, 2, 4, 5, 4, 4, 5, 3, 2, 3, 4, 4, 4, 2, 2, 0, 0, -2, -1, -5, -4, -2, 0, 0, 0, 1, 1, 2, 2, 2, 4, 3, 5, 5, 3, 4, 4, 4, 3, 4, 2, 0, -1, -3, -2, -5, -4, -2, 0, -1, 0, -1, 0, 0, 0, 0, 1, 2, 4, 3, 3, 3, 4, 2, 1, 2, 1, 0, -1, -3, -3, -5, -5, -2, -2, -1, -2, -2, -1, -1, 0, -1, 0, 0, 2, 0, 2, 0, 2, 0, 0, 2, 0, -2, -3, -3, -4, -5, -5, -3, -5, -5, -4, -5, -4, -4, -3, -3, -2, -2, -2, -1, -1, 0, 0, 0, 0, -1, -2, -3, -2, -3, -2, -6, -5, -5, -5, -6, -5, -6, -7, -7, -6, -5, -6, -5, -7, -4, -4, -4, -2, -2, -2, -3, -3, -3, -4, -3, -3, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 1, 0, 0, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 1, 2, 2, 1, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 3, 1, 1, 2, 2, 2, 2, 3, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, 1, 0, 0, 1, 2, 2, 2, 3, 3, 2, 1, 1, 2, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 3, 1, 3, 4, 3, 3, 1, 2, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, -1, 1, 0, 2, 2, 3, 3, 3, 3, 2, 2, 3, 2, 2, 1, 0, 0, 0, 0, -2, 1, -1, -1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 2, 4, 3, 2, 1, 2, 1, 0, 2, 0, 0, 0, -1, 0, 0, -1, -1, 0, -2, -1, 0, 0, 0, 1, 1, 3, 3, 3, 1, 0, 1, 2, 2, 1, 2, 0, 0, 0, 0, -2, 0, 0, -1, -1, 0, -1, -1, 0, 1, 1, 0, 3, 3, 4, 3, 2, 2, 1, 2, 1, 1, 0, 1, -1, 0, 0, -1, -1, -1, -1, -1, -1, -1, -1, 0, 2, 2, 2, 3, 2, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, 0, -2, -2, -2, 0, 1, 3, 4, 3, 2, 1, 0, 1, 2, 2, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -2, -1, 0, 0, 1, 2, 3, 3, 2, 1, 1, 0, 0, 2, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, -1, -2, -2, -2, 0, 0, 0, 1, 2, 3, 3, 2, 1, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -1, 0, 1, 1, 4, 3, 2, 3, 0, 1, 2, 3, 1, 1, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, -1, 0, -1, 1, 1, 2, 3, 2, 3, 1, 0, 2, 1, 1, 3, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, 2, 3, 4, 3, 2, 1, 1, 3, 2, 3, 2, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 4, 3, 4, 4, 3, 1, 1, 2, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 3, 5, 5, 4, 3, 3, 1, 3, 3, 1, 1, 1, 1, -1, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 3, 4, 3, 4, 3, 3, 3, 3, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 2, 2, 1, 2, 1, 1, 2, 2, 2, 1, 1, 0, -1, 0, -1, -1, -2, 0, 0, -1, -2, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, -1, -1, -1, -2, -1, -2, 0, 0, 0, -1, 0, 0, 1, 0, 1, 2, 1, 1, 1, 2, 0, 0, 1, 0, -1, -1, -1, -2, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -1, -1, -1, -2, -2, -2, -2, -3, -4, -5, -7, -8, -11, -12, -10, -8, -7, -8, -8, -9, -5, -5, -3, -3, -2, 0, -1, 0, 0, -1, -3, -1, -1, -1, -1, -2, -4, -6, -9, -8, -7, -7, -4, -5, -5, -4, -3, -1, 0, 0, 0, 0, 0, 2, 1, 1, -4, -3, -1, -1, -1, -2, -3, -5, -6, -5, -4, -3, -3, -4, -3, -2, -1, 0, 0, 0, 0, 0, 2, 1, 2, 0, -5, -2, -1, 0, 1, -1, -2, -4, -3, -3, -3, -2, -2, -2, -2, 0, 1, 1, 0, 0, 0, 1, 1, 2, 2, 0, -3, -3, -1, 0, 1, 0, -2, -2, -1, 0, -2, -1, -2, -3, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 1, 1, -3, -1, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 2, 3, 2, 0, 2, 2, 1, 4, 1, -3, -2, 0, 0, 1, 0, 0, 0, 0, 2, 2, 1, 0, 0, 0, 0, 1, 2, 3, 4, 2, 3, 2, 3, 4, 1, -4, -3, 0, -1, -1, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, 1, 2, 1, 4, 2, 3, 3, 2, 3, 3, 3, -3, -3, 0, 0, -1, 1, 0, -1, 1, 2, 3, 2, 1, 0, 0, 0, 1, 1, 1, 1, 2, 3, 1, 3, 3, 3, -3, -1, 1, 1, 1, 1, 0, 0, 2, 1, 2, 1, 1, 0, -1, -1, 0, 0, 2, 1, 2, 2, 3, 3, 3, 4, -1, 0, 0, 2, 1, 2, 0, 0, 2, 1, 1, 2, 0, 0, -1, -1, 0, 0, 0, 1, 2, 1, 2, 1, 4, 3, 0, 0, 0, 2, 2, 1, 1, 2, 3, 2, 1, 1, 1, 0, 0, -1, 0, 1, 0, 0, 0, 1, 2, 2, 3, 4, -2, 0, 1, 1, 3, 2, 1, 1, 4, 2, 2, 1, 0, -1, -1, 0, 0, 0, -1, -2, 0, 1, 3, 2, 2, 3, 0, 1, 2, 2, 1, 2, 2, 4, 3, 3, 2, 2, 0, 1, 1, -1, 0, -1, -2, -1, 0, 0, 3, 2, 2, 2, 0, 0, 0, 0, 1, 2, 2, 2, 3, 2, 3, 1, 0, 1, 0, 0, -2, -2, -3, -3, -1, 0, 1, 2, 3, 3, -1, 0, 0, 1, 2, 1, 1, 2, 2, 1, 3, 1, 0, 1, 1, -1, -3, -2, -1, -2, 0, 0, 1, 1, 2, 1, 0, 0, 1, 1, 2, 0, 1, 2, 3, 3, 1, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 2, 0, 0, -2, 0, 1, 1, 1, 0, 1, 2, 3, 4, 2, 1, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -2, -1, 0, 0, 1, 0, 0, 2, 2, 3, 2, 1, 1, 0, 2, 1, 1, 2, 0, 0, 0, 0, 1, 0, 0, -1, -3, -3, 0, 0, 0, 0, 0, 0, 3, 3, 1, 1, 1, 0, 1, 3, 2, 1, 2, 0, 1, 1, 1, 0, 0, -1, -2, -2, 0, 1, 0, -1, -1, 0, 0, 2, 0, 0, 0, 0, 1, 1, 2, 2, 2, 3, 3, 1, 2, 0, -1, -1, -4, -1, 0, 0, 0, 0, -2, -1, 0, 1, 0, 0, 0, 1, 2, 3, 3, 3, 3, 1, 3, 4, 3, 2, -1, -2, -4, -2, 0, 0, 0, -1, -4, -1, -2, 0, -2, -1, 0, 0, 0, 2, 2, 1, 1, 0, 2, 3, 2, 0, 0, -2, -2, -2, -1, -1, -2, -3, -5, -4, -4, -4, -3, -2, -2, 0, 0, 0, 1, 0, -1, -1, 1, 3, 1, 2, 0, -3, -2, -2, -2, -1, -2, -4, -5, -4, -5, -3, -5, -4, -5, -2, -2, -1, -3, -1, -1, -1, -1, 1, 0, 0, -3, -4, -2, -2, 0, -1, -2, -4, -5, -5, -5, -6, -6, -7, -6, -4, -4, -4, -5, -5, -6, -4, -2, -3, -3, -2, -5, -4, -1, -1, 0, 1, 3, 4, 3, 2, 3, 1, 0, 0, 0, 0, 0, -1, -1, -2, 0, -2, 0, 0, -1, 1, 2, 4, -1, 0, 0, 0, 1, 1, 1, 1, 2, 3, 2, 1, 1, 0, -1, 0, -1, -2, -2, -1, -3, -2, -2, 0, 1, 3, 0, 0, 0, 1, 0, 0, 0, 0, 2, 3, 2, 3, 3, 2, 1, 0, -1, -2, -2, -1, -3, -2, -1, 0, 1, 3, 0, -1, 0, -1, 0, 0, -2, -1, 0, 2, 1, 1, 2, 3, 0, 0, 0, -2, -1, -2, -1, -2, -1, 0, 0, 3, 1, 0, 0, -1, -2, -3, -3, -1, -1, 1, 1, 3, 3, 1, 1, 0, 0, 0, -3, -2, -4, -2, -3, 0, 0, 2, 3, 3, 1, 0, -2, -2, -4, -3, -1, 0, 0, 2, 4, 3, 1, 1, 0, -1, -1, -2, -4, -2, -4, -2, 0, 0, 4, 2, 1, -1, -2, -4, -4, -2, -3, 1, 1, 1, 3, 2, 0, 1, 0, 0, -2, -2, -3, -4, -4, -2, -1, 1, 2, 2, 1, 0, -1, -2, -4, -3, -2, 0, 2, 0, 1, 2, 1, 2, 0, 0, -2, -2, -2, -3, -3, -3, -1, 0, 2, 2, 0, -1, -1, -1, -4, -3, 0, -1, 1, 2, 1, 2, 0, 0, 0, 1, 1, -1, -3, -3, -4, -2, -2, 0, 0, 0, 0, -1, 0, -1, -4, -2, 0, 0, 2, 2, 2, 1, 2, 1, 2, 1, 1, 0, -1, -4, -4, -2, -2, 0, 0, -1, -2, -2, -2, -3, -2, -2, -1, 0, 2, 4, 2, 1, 0, 2, 1, -1, 0, -2, -2, -2, -4, -2, -2, 0, -1, -1, -2, -2, -2, -3, -3, -4, -1, 1, 2, 4, 3, 1, 0, 0, 0, -2, 0, -1, -2, -1, -3, -2, -2, -1, -2, 0, -2, -1, -1, -3, -4, -3, -2, 0, 2, 3, 2, 2, 1, 0, -1, 0, -3, -1, -3, -1, -3, -3, -3, 0, -1, -1, 0, -1, -3, -5, -5, -3, -1, 0, 2, 2, 4, 1, 0, 0, 0, -1, -1, -2, -2, -2, -2, -2, -2, 0, 0, 0, 0, -1, -2, -4, -5, -4, -1, 0, 0, 3, 2, 2, 1, 1, 0, -1, -1, -2, -1, -1, -4, -2, -1, 1, 0, 0, 0, 0, -2, -4, -4, -4, -2, 0, 0, 1, 3, 2, 0, 0, 0, 0, 0, -2, -1, -3, -2, -2, -2, 0, 0, 1, 0, -1, -1, -4, -5, -4, 0, 0, 1, 1, 2, 1, 1, 0, 0, 1, 1, -1, -1, -3, -2, -1, 0, 0, 2, 2, 1, 0, -3, -5, -5, -4, -1, 0, 0, 2, 0, 1, 0, 0, 1, 0, 0, 0, -2, -3, -1, -2, 0, 3, 1, 0, 0, 0, -3, -5, -5, -4, -2, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, -1, -2, -1, -1, 0, 0, 2, 0, 0, 1, 0, -3, -3, -6, -4, -3, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, -2, -2, 0, 0, 0, 2, 4, 2, 0, 0, 0, -3, -2, -2, -3, -1, 0, 1, 2, 1, 1, 1, 1, 0, 0, 0, -1, -1, -2, -1, 0, 1, 3, 1, 0, 1, -1, -2, -1, -1, -1, 0, 0, 2, 3, 1, 2, 0, 0, 0, -2, -2, -3, -2, 0, 0, 0, 0, 4, 0, 1, 0, 0, 0, -1, -1, 0, 1, 3, 2, 2, 2, 1, 0, 0, -2, -3, -1, -2, -1, -2, -1, 0, 0, 3, 0, 0, 0, -1, 0, -1, 1, 3, 4, 4, 3, 2, 1, 2, 0, 0, -3, -4, -3, -3, -1, -1, -2, -1, 0, 4, 0, 0, 1, 1, 1, 2, 1, 3, 4, 3, 2, 1, 2, 0, 0, -1, -3, -2, -3, -3, -2, -2, -2, -1, 1, 5, 0, 1, 0, 1, 0, 2, 4, 3, 3, 3, 3, 1, 1, 1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 3, 6, 1, 0, 2, 3, 1, 1, 2, 1, 3, 2, 4, 2, 1, 0, -2, -2, -3, -4, -4, -2, -1, 0, 0, 1, 1, 3, 0, 2, 0, 1, 0, 0, 2, 2, 4, 4, 3, 3, 0, 0, -3, -4, -5, -5, -4, -3, -1, 0, 0, 0, 2, 4, 1, 1, 0, 0, 0, 0, 2, 3, 4, 3, 4, 4, 1, -2, -2, -4, -4, -4, -3, -2, -1, 0, 0, 0, 1, 4, 1, 0, 0, 1, 0, 0, 0, 3, 2, 3, 4, 3, 0, -1, -2, -3, -4, -3, -3, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 3, 2, 0, 0, -2, -1, -4, -3, -3, -1, -1, -1, 0, 0, 0, 2, 0, 0, 1, 1, 0, 0, 0, 0, 1, 2, 2, 2, 0, 0, -1, -3, -3, -3, -1, -3, 0, 0, 0, -1, 0, 2, 0, 0, 2, 1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, -1, -2, 0, 0, -2, -1, -1, 0, 0, -1, 0, 1, 2, 3, 2, 2, 0, 0, 0, 0, 1, 1, 2, 2, 0, 1, 0, 0, 0, -1, 0, -2, 0, -1, 0, -1, -1, 2, 1, 2, 3, 1, 0, -1, -1, 0, 0, 3, 1, 1, 2, 1, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, -1, 2, 2, 1, 2, 0, -1, -1, -1, 0, 1, 2, 2, 3, 1, 0, 0, 1, 0, 0, 0, -2, -2, -3, -2, -2, 0, 1, 2, 1, 1, 0, 0, -1, 0, 0, 0, 2, 1, 2, 1, 2, 0, 0, -1, 0, -1, -1, -2, -2, -2, -3, 0, 0, 3, 1, 3, 1, 0, -1, -1, 0, 0, 0, 2, 2, 1, 0, 0, -1, 0, 0, 0, -1, -3, -2, -2, -1, 0, 1, 3, 3, 1, 0, 0, -2, -1, -1, 0, 2, 2, 2, 1, 1, 0, 0, -1, -1, 0, 0, -2, -2, -2, -4, -1, 0, 1, 1, 0, 0, 0, -1, 0, -1, -1, 0, 3, 2, 2, 2, 0, -2, 0, -2, -1, 0, -3, -3, -3, -3, -2, 0, 1, 1, 0, -1, -1, -1, -2, -1, 0, 0, 1, 4, 2, 1, 1, 0, -1, 0, -2, 0, -1, -4, -2, -3, 0, 0, 2, 1, 0, 0, -1, 0, 0, -2, -1, 0, 2, 3, 2, 1, 0, 0, -1, 0, -1, -2, -2, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 2, 2, 1, 1, 1, 0, 0, 0, -1, -2, -2, -1, -2, -2, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, -1, 0, 2, 4, 1, 1, 1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 1, 2, 1, 1, 1, 2, 1, 0, 0, 1, 1, 3, 4, 1, 1, 0, 0, 0, -2, 0, -2, 0, -1, -1, 0, 1, 0, 3, 3, 1, 1, 0, 0, 1, 0, 1, 2, 3, 3, 2, 0, -1, 0, -1, -3, -3, -1, -1, -1, -1, -1, 1, 0, 0, 0, 1, 1, 0, 1, 2, 1, 2, 1, 4, 3, 1, 0, 0, -1, -1, -2, -1, -2, -2, -1, -1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, 1, 1, 3, 2, 3, 1, 0, -1, -2, -3, -2, -1, -1, -1, 0, -1, 0, 1, 1, 0, -1, 0, 0, 0, 0, 1, 3, 2, 3, 3, 2, 1, -1, -3, -3, -2, -2, 0, -2, -1, -2, -1, 0, 1, 2, 0, -1, 0, 0, 1, 0, 2, 2, 2, 2, 2, 1, 0, -1, -4, -4, -3, -1, -2, -3, -2, -2, -1, 0, 1, 2, 0, 0, 0, 0, 1, 1, 2, 3, 2, 2, 2, 3, 1, 0, -3, -3, -2, -2, 0, -2, -1, -1, 0, 0, 2, 4, 1, 0, 0, 0, 1, 0, 0, 1, 1, 3, 3, 3, 2, 0, -2, -3, -2, -1, 1, 0, 1, 0, 2, 2, 2, 4, -6, -5, -2, -1, -1, -2, -3, -2, -3, -3, -4, -4, -4, -7, -8, -9, -7, -3, -4, -3, -2, -3, -2, -1, -1, 0, -6, -4, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, -2, -4, -5, -4, -3, -2, -3, -2, -1, -2, -2, -2, -3, 0, -2, -2, -1, 1, 0, 1, -1, -1, 0, 1, 1, 1, 0, -2, -3, -2, 0, 0, 0, 0, 0, -3, -2, -3, -1, -1, -3, 0, 0, 0, 0, 0, 0, -1, 2, 1, 3, 3, 3, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -1, 0, 0, 2, 2, 0, 0, 0, 0, 1, 4, 5, 5, 4, 3, 3, 2, 3, 1, 0, 0, 0, -2, -1, -2, -2, 0, 0, 0, 0, 2, 1, -1, 0, 0, 2, 4, 5, 4, 4, 3, 5, 4, 3, 1, 1, 0, 0, -1, -3, -1, -1, 0, 0, 3, 1, 1, -1, -1, 0, 0, 1, 4, 4, 5, 4, 5, 6, 5, 3, 3, 0, 1, 0, -1, -2, -2, -2, -1, 1, 2, 0, 0, -1, 0, 0, 1, 3, 6, 4, 6, 5, 5, 5, 6, 3, 1, 1, 0, 0, -2, -2, -1, -2, 0, 0, 0, 0, 0, 0, -1, 0, 2, 5, 6, 5, 5, 6, 7, 6, 5, 3, 1, 0, 0, 0, -1, -3, -4, -2, -3, 0, -1, 0, 1, 1, 0, 0, 3, 4, 5, 5, 6, 7, 7, 5, 5, 2, 0, 0, -1, -1, -2, -4, -4, -3, -3, -2, -1, 0, 0, 1, 0, 1, 3, 5, 7, 6, 7, 8, 7, 6, 2, 1, 0, -1, -1, -2, -3, -4, -3, -3, -3, -4, -2, 0, 2, 2, 3, 4, 3, 5, 5, 6, 8, 8, 6, 6, 3, 0, 0, -1, -1, -2, -3, -4, -4, -2, -3, -3, -1, 0, 0, 2, 2, 2, 5, 6, 6, 6, 8, 9, 8, 5, 3, 0, 0, -2, -1, -3, -3, -3, -3, -3, -2, -4, -1, 0, 1, 4, 3, 3, 4, 5, 6, 8, 8, 7, 6, 4, 3, 0, 0, -1, -1, -1, -2, -2, -4, -4, -1, -4, 0, 0, 2, 2, 3, 3, 3, 4, 6, 5, 5, 6, 5, 5, 4, 1, 0, 0, -1, -1, -2, -3, -3, -3, -2, -2, -1, 0, 3, 3, 2, 1, 3, 2, 2, 4, 3, 4, 5, 3, 2, 2, 2, 1, 0, -1, -1, -4, -3, -4, -3, -3, -2, 1, 2, 3, 0, 2, 1, 2, 3, 3, 4, 3, 5, 4, 2, 2, 3, 2, 0, 0, -1, -2, -4, -4, -2, -4, -1, 1, 1, 1, 1, 0, 0, 2, 3, 3, 3, 4, 4, 2, 2, 2, 2, 0, 1, 0, 0, -3, -3, -3, 0, -3, -1, 0, 2, 1, 1, 1, 2, 3, 3, 4, 4, 3, 4, 3, 2, 3, 3, 2, 2, 0, -2, -2, -3, -3, -1, -2, -1, 0, 2, 2, 0, 1, 0, 2, 3, 3, 4, 4, 2, 1, 2, 3, 3, 2, 1, -1, -2, -2, -3, -2, 0, -3, -2, 0, 2, 1, 0, 1, 0, 1, 2, 3, 5, 3, 2, 3, 2, 2, 2, 0, 0, 0, -1, -2, -2, -3, 0, -3, -2, 0, 1, 0, 0, 0, 0, 2, 2, 3, 3, 3, 2, 3, 1, 3, 0, 0, 0, 0, -2, -2, -3, -1, 0, -3, -2, -1, 0, 0, 0, 0, 0, 2, 2, 2, 3, 3, 3, 3, 3, 1, 0, 0, 0, 0, -2, -4, -3, -2, 0, -3, -3, -1, 0, -1, -1, -1, 1, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, -2, -2, 0, -3, -3, -4, -2, 0, -4, -3, -3, -2, -3, -4, -2, -2, -2, 0, -1, -3, -2, -2, -2, -3, -2, -2, -2, -1, -1, -3, -3, -2, -3, 0, -4, -3, -4, -4, -2, -5, -3, -4, -3, -2, -5, -4, -5, -5, -5, -6, -5, -4, -3, -3, -1, 0, -3, -1, -1, 1,
    -- filter=0 channel=2
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, -1, 0, -1, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, -1, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, 1, -1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 1, -1, 0, -1, -1, 1, 0, 1, -1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 1, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, -1, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, 1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, -1, -1, 0, 0, 0, -1, 0, 0, 1, 1, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, -2, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -2, -1, 0, -1, 0, 0, -2, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, -1, 0, 0, -2, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -2, -2, -2, 0, -1, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, -2, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, -1, 0, 1, 0, 1, 0, 0, -1, -1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 1, -1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 1, -1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, -1, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 1, 0, -1, 1, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -2, 0, 0, -2, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, -1, 1, 0, 0, 0, -1, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 1, 0, 0, 0, 0, 1, -1, 0, 1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -2, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -2, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 1, -1, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, 1, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, -1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, -1, -1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 1, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, -1, -1, 1, -1, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, -1, 1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 1, 0, 1, -1, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, -1, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, -1, 0, 1, 1, 1, 0, 0, 1, 0, 1, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, -1, -1, 0, -2, -2, -1, -1, -2, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -2, -1, -1, 0, -2, 0, 0, 0, -1, -1, -1, -1, -2, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, -2, 0, -2, -1, -2, -1, 0, -2, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, -1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, -1, -1, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, -1, -1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, -1, 0, 1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, -1, 1, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, -2, 0, -2, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, -2, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, -1, -1, -2, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, 0, -2, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -2, -2, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, 1, -1, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, -1, -1, -1, 1, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 1, 0, -1, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, -1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, -1, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, -1, 0, 1, -1, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 1, 0, 0, -1, 0, 1, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, 1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, -1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, -1, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, -1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 1, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 1, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, -1, 0, 1, 0, -1, -1, 0, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, -1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 1, 1, 1, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 1, -1, 0, 0, 1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 1, -1, 1, 1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, -1, 0, 0, 1, 0, 0, 1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, -1, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 1, 0, 0, 1, 0, 0, -1, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, -1, 1, 1, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 1, 0, -1, 1, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, -1, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, -1, -1, -1, -1, -1, -1, 0, -1, -1, 0, -1, -1, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, -2, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, -1, 1, 1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 1, 0, -1, 1, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, 0, -1, 0, 1, -1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, -1, 0, -1, 1, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, -1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 1, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, 1, -1, 0, -1, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 1, -1, 1, 0, 0, 0, -1, 0, 1, -1, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, -1, -1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, -1, -1, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, -2, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -2, -2, -1, 0, -1, -1, -1, -1, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, -1, -2, -1, -1, -2, 0, -1, -2, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -2, -1, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, -2, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -1, -1, -1, 0, -1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, -1, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 1, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 1, 1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, -1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, -1, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, -1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, -1, -1, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, -1, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, 1, 1, 0, 0, 0, 0, 1, -1, 0, -1, 0, -1, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, -1, 1, 0, 0, 0, -1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 1, 1, -1, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, -1, -1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, -1, 0, -1, 1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    -- filter=0 channel=3
    -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, 0, -1, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -2, -2, -1, -1, -1, -2, -2, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, -1, -1, -2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 1, -2, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -2, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, -2, -1, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 2, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 2, -1, 0, 2, 0, 2, 2, 3, 3, 5, 4, 3, 2, 3, 2, 3, 1, 2, 1, 2, 0, 2, 1, 2, 1, 1, 1, -1, -1, 0, 1, 3, 3, 3, 3, 2, 2, 3, 2, 2, 0, 2, 1, 1, 1, 2, 1, 2, 0, 1, 2, 2, 3, -3, 0, -1, 0, 0, 2, 0, 1, 0, 0, 2, 1, 0, 1, 0, 1, 0, 1, 0, 2, 0, 0, 0, 1, 0, 1, -2, 0, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, -1, 1, 0, 0, 1, 2, 1, 1, 0, 1, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, -2, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 1, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -2, 0, -1, -1, -1, 0, 0, 0, -1, -1, -1, 0, 1, -1, 0, -2, -1, 0, -1, 0, -1, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, -1, 0, 0, -1, 0, -1, -1, -2, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 2, -1, 0, 0, 0, -2, -3, -2, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 2, -1, 0, 0, -2, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 2, 1, 0, 1, 0, 3, 0, 0, -1, -1, -1, -2, -2, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 3, -1, 0, 0, -2, 0, -1, -2, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 4, -1, 0, 0, 0, -2, -1, -1, -2, -1, 0, -1, 1, 0, 0, 0, 0, 1, 2, 2, 0, 0, 2, 1, 2, 1, 3, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 1, 1, 3, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 0, 0, 1, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 2, 0, -1, 0, 0, 1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 2, 0, 2, 0, 0, 0, 0, 2, 2, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 3, 2, 2, 0, 0, 0, 1, 1, 2, 3, 3, 2, 3, 2, 0, 1, 1, 0, 1, 0, 0, 1, 2, 1, 2, 1, 1, 3, 2, 1, 2, 1, 1, 0, 0, -1, 0, -1, -1, -1, 0, 0, -2, -1, -2, -1, 0, 0, 0, -1, -1, -2, 0, 0, -1, 2, 3, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 2, 1, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, -1, 3, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 1, 0, 0, -2, -2, -2, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, -2, -2, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 1, 2, 1, 0, -1, -1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 1, 2, 2, 1, 1, 1, 1, 0, 2, 2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 1, 1, 2, 2, 3, 3, 1, 3, 1, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 2, 3, 2, 0, 2, 0, 1, 1, 1, 3, 2, 3, 2, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 3, 1, 1, 2, 2, 0, 0, 2, 2, 2, 3, 3, 0, 0, -1, -1, 1, 1, 1, 0, 0, 0, -1, 1, 0, 1, 0, 3, 2, 1, 2, 0, 1, 1, 2, 4, 3, 2, 1, 1, 0, 0, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 2, 2, 1, 1, 1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 1, 2, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 2, 1, 2, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 2, 2, 0, 0, 1, 0, -1, 2, 1, 1, 0, 1, 2, 1, 1, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, -1, 2, 2, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 3, 0, 0, 0, 0, 1, 1, 2, 2, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 2, 1, 3, 1, 0, 1, 3, 2, 1, 0, 0, 1, 1, 1, 0, 1, 1, -1, 0, 0, 0, 0, 2, 1, 2, 1, 2, 4, 2, 2, 2, 1, 1, 1, 2, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 4, 5, 3, 2, 1, 3, 1, 2, 0, 0, 0, 0, 2, 2, 0, 0, 0, 1, 1, 2, 0, 1, 1, 0, 1, 2, 4, 3, 4, 1, 0, 3, 1, 2, 0, -1, 0, 1, 1, 2, 0, 2, 1, 2, 3, 2, 0, 1, 0, 1, 1, 1, 3, 3, 3, 1, 0, 2, 3, 1, 0, -1, 0, 1, 1, 1, 2, 1, 2, 3, 1, 2, 1, 0, 0, 1, 1, 1, 0, 2, 0, 1, 0, 2, 1, 1, -1, -1, 0, 0, 0, 1, 0, 1, 3, 2, 2, 1, 2, 2, 1, 0, 1, 1, 1, 2, 0, 0, -1, 3, 2, 2, 0, 0, 0, -1, 0, 0, 0, 1, 2, 1, 1, 2, 2, 1, 1, 1, 0, 1, 0, 0, 0, -1, -3, 3, 1, 1, -1, -1, -2, -1, -1, 0, -1, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -2, -1, -2, 0, 0, 0, 0, 2, 1, 1, 2, 0, 0, 0, 1, 1, 0, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, 2, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 2, 0, 0, 1, 2, 2, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 2, 0, 0, 1, 1, 0, 2, 2, 1, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 2, 0, 2, 1, 2, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 2, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, -1, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 1, 1, -1, 0, 0, -1, -2, -2, -1, -2, 0, 1, 0, 0, -1, 0, -1, 0, 0, 1, 2, 1, 1, 0, 1, 0, 1, 0, 0, -1, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 2, 0, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 2, 2, 0, 1, 2, 2, 2, 2, 0, 0, 0, 1, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 2, 2, 1, 0, 1, 1, 2, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 1, 0, 2, 1, 1, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, -1, 0, -1, 0, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 2, 1, 1, 0, 1, -1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 2, 2, 0, 0, 1, 1, 0, 0, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 0, -1, 0, 1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 1, 0, 1, 0, 2, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 2, 1, 1, 2, 1, 2, 0, 1, 1, 0, 1, 2, 0, 0, 0, -1, 0, -2, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 2, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -2, 0, -1, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 2, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 0, 2, 1, 2, 0, 2, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 2, 0, 0, 2, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 2, 1, 1, 0, 1, 0, 2, 1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 2, 0, 1, 1, 1, 2, 1, 0, -1, 0, 0, 0, 0, 2, 1, 1, 1, 1, 3, 1, 1, 1, 0, 2, 0, 2, 2, 2, 1, 1, 2, 1, 0, 1, 0, -1, 0, 1, 1, 0, 0, 1, 0, 1, 2, 2, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 1, 1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 2, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 2, 1, 2, 2, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 2, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, -1, -1, 0, 0, 0, -1, 0, 1, 2, 1, 1, 1, 1, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 3, 2, 2, 3, 2, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 4, 3, 2, 1, 0, 2, 2, 1, 1, 0, 1, 2, 1, 2, 1, 1, 1, 2, 1, 0, 1, 0, 0, 0, 0, -1, 0, 2, 2, 1, 1, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 1, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -2, 0, -2, 0, 0, -1, 0, 0, -1, 2, 0, 1, 0, 0, 0, 0, 2, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, -3, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -1, 0, 0, 0, 0, 2, 0, -1, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 1, 0, 0, 1, 1, 1, 0, -1, -1, -1, -2, -1, -3, -2, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 2, 1, 0, 1, 2, 0, 0, -1, 0, -1, -3, -3, -1, -2, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 2, 0, 1, 1, 0, 0, -1, -2, -1, -3, -3, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 1, -1, -1, 0, -2, -1, -3, -1, -1, -1, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, -2, -2, -3, -1, -3, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, -2, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, -1, 0, -2, -3, -3, -2, 0, 0, -1, -1, -1, 0, 1, 1, 0, -1, 0, -1, -1, -1, 2, 0, -1, -2, -2, 0, 0, -2, 0, -2, -1, -2, -2, -2, -1, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, -2, 1, 0, -1, -2, -2, -1, -1, -2, -3, -2, -3, -2, -1, -2, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 2, 1, 0, -2, 0, 0, 0, -1, -2, -3, -1, -3, -3, -1, -3, -2, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 2, 0, 0, 1, 0, 0, 0, -1, 0, -1, -3, -2, -3, -1, -1, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, 3, 1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -3, -3, -2, -3, 0, -2, 0, -1, 0, -2, -2, -1, 0, 0, 3, 1, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, -2, -3, 0, -2, -1, 0, -2, -2, 0, -1, 3, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -2, 0, -1, -2, -1, -1, -1, -1, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, 0, -2, -1, -3, 0, -2, 2, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -2, -2, -2, -4, 2, 0, 1, 0, -1, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -2, -3, -3, 2, 2, 0, 0, 0, -1, -1, -1, -2, 0, -1, 0, 0, 1, 0, 0, 0, 0, 2, 0, 0, -1, -2, -4, -3, -6, 7, 4, 2, 1, 0, 0, -1, -2, -2, 0, 0, -1, -1, -4, -4, -5, -5, -3, -2, -3, -4, -6, -7, -7, -7, -9, 6, 3, 2, 1, 0, 0, 0, -2, -1, -1, 0, -2, -2, -2, -2, -3, -3, -2, -3, -2, -2, -4, -5, -4, -4, -8, 5, 3, 2, 1, 0, 1, 0, -1, 0, -1, 0, -1, -1, -1, -2, -2, 0, 0, 0, -1, 0, -2, -4, -4, -4, -5, 6, 2, 0, 0, 2, 2, 1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 1, -1, -1, -2, -1, -2, -3, 5, 2, 1, 0, 0, 3, 1, 0, 0, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 6, 3, 1, 0, 1, 3, 3, 0, 0, -1, 0, 1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 4, 2, 1, 0, 2, 5, 3, 2, 0, 0, 0, 1, 0, -1, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, -1, 0, 3, 3, 3, 3, 0, 0, 1, 1, 0, -1, -1, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 2, 1, 0, -2, 0, 3, 1, 3, 3, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 1, 1, -1, -2, -2, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 1, 0, 2, -1, -3, -1, -1, 2, 2, 3, 1, 2, 0, 0, -1, 1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 2, 0, 0, 1, -2, -4, -2, 0, 0, 1, 1, 2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, -1, -4, -3, 0, 1, 1, 2, 3, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 2, 3, 2, 3, 0, 0, -4, -5, -4, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, -1, -1, 0, 1, 0, 2, 1, 3, 1, 0, 1, 0, -3, -4, -3, 0, 0, 1, 1, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 3, 2, 0, 0, 0, 0, 1, -3, -4, -4, -1, 0, 1, 0, 0, 0, 1, 1, 0, 0, -2, -1, -2, -1, 0, 1, 2, 3, 2, 0, 0, -2, 1, 0, -2, -2, -2, 0, -1, 0, 0, 2, 0, 0, 0, 0, -2, -2, -1, 0, 1, 2, 1, 3, 0, 0, -1, -4, 2, 0, -2, 0, -1, -1, 0, 0, 0, 1, 0, 0, -1, -2, 0, 0, -1, 0, -1, 0, 2, 1, 1, -1, -1, -3, 2, 0, 0, 0, -1, 0, 0, 1, 0, 2, 1, -1, -2, -2, -3, -1, 0, 0, 0, 0, 0, 0, 1, 1, -1, -3, 3, 2, 2, 0, 0, 0, 1, 1, 3, 2, 2, -1, -2, -1, -3, -2, -2, 0, 0, 0, 0, 1, 0, 1, 0, -2, 3, 3, 2, 3, 0, 0, 0, 1, 2, 3, 2, 0, 0, -1, -1, 0, 0, -1, -1, 0, 1, 0, 0, 0, 1, -1, 4, 4, 3, 5, 3, 0, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 5, 6, 6, 5, 2, 1, 2, 2, 2, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, -3, 7, 6, 4, 3, 3, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, 0, -2, -3, 5, 4, 4, 3, 1, 0, -1, 0, 0, 0, -1, -2, -2, 0, 0, 0, 0, 0, 0, -2, -1, -4, -3, -2, -4, -4, 3, 3, 2, 2, 0, 0, 0, 0, -1, 0, 0, -3, -2, -2, -1, 0, 0, 0, 0, -1, -1, -1, -4, -3, -4, -7, -6, -3, -2, 0, 0, 2, 2, 5, 6, 6, 6, 5, 7, 4, 6, 5, 5, 4, 3, 4, 4, 5, 3, 3, 3, 0, -5, -4, -2, -2, 0, 1, 1, 2, 4, 5, 5, 4, 3, 3, 2, 2, 3, 1, 0, 0, 1, 3, 3, 1, 2, 3, -6, -4, -2, -1, -1, 0, 1, 1, 0, 1, 3, 1, 1, 1, 0, 0, 2, 1, 1, 1, 2, 1, 2, 0, 2, 3, -5, -3, -4, -2, -1, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, -5, -3, -3, 0, 0, 0, 1, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -4, -2, -1, -1, 0, 1, 2, 0, -1, -1, -2, -1, -3, 0, -2, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 1, -5, -4, -2, 0, 0, 2, 1, 0, -1, -2, -3, -2, -4, -2, -2, -2, -1, -2, -1, 0, -1, 0, 0, 0, -1, 1, -5, -4, -2, -1, 0, 0, 1, 0, -1, -3, -2, -4, -4, -2, -1, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 2, -6, -4, -3, -1, -1, 0, 0, 0, -1, -1, -2, -2, -4, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -3, -2, -4, -3, -2, -1, 0, -2, -1, -2, -1, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -5, -2, -2, -3, -1, -1, -1, -2, -1, -1, -2, 0, -1, 0, 0, 0, 0, 2, 3, 3, 2, 0, 0, -1, -1, 1, -3, -1, -2, -2, -2, -3, -1, -1, -2, -1, 0, 0, 2, 0, 0, 1, 0, 0, 2, 3, 3, 2, 0, 0, 0, 0, -2, -2, -1, -2, -2, -1, -1, -2, 0, 0, 1, 0, 1, 2, 0, 1, 1, 1, 2, 3, 1, 0, -2, -2, 0, 1, -1, 0, -2, -3, -3, -3, -3, -1, -2, -1, 0, 0, 1, 0, 2, 1, 0, 0, 0, 3, 2, 0, -1, -2, 0, 3, -1, -2, -2, -3, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 2, 0, 1, 0, -1, 1, 2, -1, 0, -1, -2, -2, -2, 0, -2, -1, 0, 0, 0, 1, 0, 0, 1, 1, 2, 2, 2, 1, 1, 0, 1, 3, 3, -2, 0, -2, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 2, 2, 1, 1, 1, 0, 0, 0, 1, 2, -2, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -2, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, -3, -3, -2, -2, -2, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 2, 0, 0, 0, 0, -3, -3, -2, -2, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 2, 3, 4, 2, 0, -1, 0, 0, -2, -4, -2, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 4, 4, 3, 2, 0, 0, 0, -4, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 1, 2, 1, 2, 1, 1, 1, 2, 1, 1, 1, -4, -2, -1, -1, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, -1, 0, 1, 2, 2, 1, 3, 2, 0, 1, 2, 1, -3, -2, 0, 0, 2, 2, 2, 2, 3, 3, 3, 3, 1, 1, 0, 0, 0, 0, 2, 2, 2, 1, 2, 2, 4, 2, -4, -2, 0, 2, 3, 2, 4, 5, 4, 4, 6, 4, 5, 3, 3, 2, 3, 4, 4, 2, 4, 2, 4, 5, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, -1, 0, -2, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 1, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 2, 2, 2, 1, 0, 1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -4, -1, 0, 2, 2, 4, 5, 7, 6, 9, 9, 7, 7, 6, 4, 5, 4, 4, 3, 3, 3, 4, 3, 1, 1, 1, -4, -1, -1, 0, 2, 2, 3, 5, 6, 7, 5, 5, 4, 4, 2, 1, 3, 2, 0, 3, 3, 4, 2, 2, 2, 2, -4, -3, 0, 0, 0, 2, 3, 3, 4, 3, 4, 2, 2, 2, 2, 1, 2, 1, 1, 2, 4, 2, 3, 1, 2, 2, -4, -2, -1, -1, 2, 1, 2, 0, 1, 2, 2, 0, -1, 0, -1, 0, 1, 1, 1, 3, 2, 2, 1, 0, 2, 3, -4, -2, 0, 0, 1, 1, 2, 1, 0, 0, 0, -1, -2, -1, 0, 0, 0, 2, 2, 3, 0, 2, 0, 0, 1, 3, -5, -1, 0, 0, 2, 3, 2, 1, 0, 0, -1, -3, -2, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 2, -5, -4, -1, 0, 0, 1, 1, 0, 0, 0, -1, -2, -3, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -5, -5, -2, -1, -1, 0, 0, 0, -1, -2, -1, -3, -2, -1, -1, -1, -1, -1, -2, -1, -1, -1, -1, 0, 0, 3, -6, -5, -4, -4, -2, 0, 0, -1, -2, -1, -1, -1, -2, -2, -2, 1, 0, 0, 0, 0, 0, -2, -2, -1, 1, 1, -5, -4, -4, -3, -3, -2, -2, -1, -3, -3, -1, -2, -1, -1, 0, 1, 2, 2, 2, 0, 0, 0, -1, 0, 0, 2, -4, -4, -4, -4, -4, -2, -3, -4, -2, -2, -2, -1, 0, 0, 2, 1, 3, 2, 3, 2, 0, 0, -1, 0, 0, 1, -4, -3, -3, -5, -6, -5, -2, -2, 0, 0, 1, 1, 1, 2, 1, 1, 2, 3, 2, 3, 2, 0, 0, 0, 0, 2, -3, -3, -4, -5, -4, -3, -5, -4, -1, 0, 1, 3, 3, 4, 3, 1, 2, 3, 4, 3, 3, 2, 0, 0, 0, 2, -3, -4, -3, -4, -4, -3, -3, -3, -1, 0, 1, 2, 2, 2, 2, 3, 2, 2, 3, 3, 1, 0, -1, 0, 0, 3, -3, -3, -4, -5, -4, -5, -2, -3, -2, 0, 0, 0, 1, 2, 2, 2, 0, 2, 2, 2, 1, 0, 0, 0, 2, 4, -2, -2, -1, -4, -3, -4, -3, -3, -1, -1, 1, 0, 0, 1, 0, 2, 1, 2, 1, 4, 2, 2, 2, 2, 2, 3, -3, -1, -1, -2, -3, -2, -1, -2, 0, 0, 2, 0, 1, 0, 1, 2, 2, 4, 2, 2, 1, 2, 1, 1, 1, 2, -3, -2, -2, -1, -2, -1, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, -2, -2, -2, -3, -2, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -2, -1, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 3, 3, 1, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 1, 2, 1, 2, 4, 4, 2, 0, 0, 2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 1, 1, 2, 3, 1, 0, 1, 1, 1, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 1, 2, 1, 2, 1, 2, 1, 1, 2, -2, 0, 0, 2, 2, 3, 2, 4, 4, 5, 4, 2, 0, 0, 0, 1, 0, 0, 1, 2, 2, 2, 1, 3, 3, 3, -3, 0, 0, 4, 6, 5, 6, 5, 6, 6, 6, 4, 3, 3, 1, 1, 2, 1, 2, 2, 2, 1, 4, 3, 4, 4, 0, 0, 1, 1, 1, 1, 1, 4, 3, 3, 5, 4, 3, 3, 5, 5, 3, 5, 5, 4, 5, 5, 4, 5, 2, 3, 0, 0, 0, 1, 1, 1, 2, 3, 4, 3, 2, 2, 4, 3, 2, 4, 4, 3, 3, 4, 4, 3, 4, 2, 4, 3, 1, 0, 0, 0, 0, 2, 1, 1, 3, 4, 3, 3, 3, 2, 4, 3, 3, 2, 1, 3, 3, 2, 2, 3, 2, 4, 0, 0, 0, 1, 1, 1, 1, 3, 4, 4, 3, 1, 2, 1, 2, 3, 2, 2, 0, 1, 1, 0, 2, 1, 1, 2, 1, 0, 1, 0, 1, 0, 0, 1, 1, 2, 2, 0, 0, 2, 1, 2, 1, 0, 0, 1, 2, 2, 2, 1, 1, 1, 0, 1, 0, 0, 0, 1, 1, 0, 2, 1, 1, 2, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 2, 0, 1, 0, 0, 1, 1, 2, 1, 2, 0, 0, 2, 0, 0, -1, 0, 0, 0, 1, 2, 2, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 2, 2, 2, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, 0, 1, 0, 0, 1, 2, 0, 1, 0, 0, 1, 0, 0, 0, 0, -2, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 2, 2, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, -1, 0, -1, 0, 1, 2, 1, 1, 1, 1, 2, 2, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, -2, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, -1, -1, 0, -1, -1, -1, 0, 1, 3, 2, 1, 0, 0, 1, 0, 3, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 2, 4, 2, 1, 0, 0, 0, 3, 3, 2, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 4, 4, 3, 2, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 3, 3, 2, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 2, 0, 0, 0, -1, -1, -1, 1, 1, 0, 1, 0, 1, 1, 2, 1, 2, 1, 1, 1, 0, 2, 1, 0, 1, 2, 2, 0, 0, 0, -1, 0, 0, 0, 2, 1, 2, 2, 1, 2, 2, 1, 0, 1, 1, 0, 0, 1, 1, 0, 2, 2, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 2, 2, 2, 1, 2, 0, 0, 0, 1, 0, 0, 1, 0, 1, 2, 0, 0, 1, 0, 1, 0, 1, 1, 1, 2, 0, 0, 3, 3, 3, 1, 1, 2, 3, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 2, 0, 0, 2, 2, 2, 2, 2, 1, 1, 3, 3, 1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 2, 0, 2, 2, 1, 2, 1, 2, 1, 3, 3, 3, 2, 2, 3, 2, 0, 1, 0, 0, 2, 1, 1, 2, 4, 2, 2, 3, 3, 2, 3, 2, 2, 3, 3, 2, 2, 4, 2, 3, 2, 1, 2, 1, 1, 1, 1, 1, 3, 2, 3, 2, 2, 2, 3, 2, 3, 4, 4, 4, 3, 3, 2, 4, 1, 3, 3, 3, 1, 0, 1, 2, 1, 2, 0, 2, 3, 4, 5, 4, 4, 4, 3, 5, 5, 3, 5, 5, 5, 4, 3, 4, 5, -1, 0, 0, 0, 1, 2, 2, 1, 2, 3, 3, 2, 2, 0, 0, 0, 0, -1, -1, 0, 1, 1, 0, 0, -1, -2, -1, 0, 0, 1, 2, 2, 3, 2, 2, 0, 0, 2, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 1, 2, 1, 3, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, 3, 1, 3, 2, 3, 2, 1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 1, 0, -1, -1, -1, 1, 1, 2, 1, 3, 2, 1, 3, 2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 1, 1, 3, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -4, -2, -1, 0, 1, 1, 2, 2, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -2, -3, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, -2, -1, 0, 0, -2, -2, -3, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -2, -4, -3, -2, -3, -3, -2, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -4, -3, -3, -2, -3, -2, -2, -1, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 1, 1, 1, -2, -3, -3, -3, -3, -3, -2, -2, -2, -1, 0, -1, -1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 2, 1, -3, -2, -4, -3, -4, -3, -4, -2, -3, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -2, -3, -2, -4, -3, -5, -4, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 1, 2, -1, -2, -1, -3, -3, -3, -2, -3, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 2, 1, 2, 1, 1, 1, 2, -2, 0, -2, -2, -2, -1, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 2, 1, 1, 1, 0, -1, 0, 0, -1, -2, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, -2, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 2, 1, 0, 0, 0, 1, 0, 0, -2, -1, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, -3, -1, 0, 0, 1, 2, 2, 2, 1, 1, 0, 2, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 1, 0, 1, 1, 2, 2, 1, 2, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -2, -1, -2, -1, 0, 1, 0, 1, 1, 0, 0, 2, 1, 1, 2, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, 0, -1, 0, 1, 0, 1, 1, 0, 0, 0, 2, 2, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 1, 1, 1, 2, 1, 2, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 2, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 2, 1, 2, 1, 1, 0, 1, 0, 0, 0, -1, 0, 1, 0, 2, 2, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 1, 2, 1, 0, 0, 0, -2, -1, -3, -1, -1, 1, 0, 1, 2, 1, 3, 2, 0, 0, -1, 0, 0, -1, -1, 0, 1, 0, 1, 1, 0, -1, -1, -2, -3, -2, -1, 0, 0, 1, 0, 1, 2, 1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, -1, 0, -2, -2, -1, -1, 0, -1, 0, 1, 0, 1, 0, 1, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, -1, -1, 1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -3, -2, -3, -2, 0, -2, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -3, -3, -3, -3, -3, -2, -1, -3, -1, 0, -2, 0, 0, -1, 0, 0, -1, -1, 0, 0, 1, 1, 0, 2, 0, 0, -2, -3, -2, -2, -2, -1, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 1, -3, -2, -3, -3, -2, -3, -1, -2, -1, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, -1, -3, -3, -3, -4, -2, -2, -2, -3, -1, -1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 2, 2, 2, 0, 0, 1, -3, -2, -2, -2, -1, -2, -2, -2, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 0, 1, 0, -1, -2, -2, 0, -2, -3, -1, -1, -2, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 2, 2, 2, 0, 1, 0, -2, -1, -2, 0, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, -1, -1, 0, 1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, -2, -1, -1, -1, -2, 0, -1, -1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, -1, 1, -2, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, 0, 0, 1, 1, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -4, -1, 1, 1, 4, 4, 5, 5, 7, 6, 7, 5, 6, 6, 4, 4, 3, 3, 3, 3, 4, 5, 5, 4, 4, 4, -4, -3, -1, 0, 1, 3, 2, 4, 3, 5, 4, 3, 4, 3, 2, 2, 3, 2, 3, 2, 4, 3, 3, 2, 2, 4, -3, -2, 0, 1, 1, 1, 0, 0, 2, 2, 2, 0, 0, 0, 1, 1, 2, 1, 2, 1, 1, 1, 3, 2, 2, 4, -4, -3, -1, 0, 2, 1, 0, 2, 2, 1, 1, 0, -1, -1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 3, 2, -4, -3, 0, 0, 0, 0, 1, 2, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 3, -4, -3, 0, 1, 2, 2, 1, 0, 0, -1, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, -4, -1, -1, 0, 0, 1, 0, 0, 0, -2, -3, -1, -2, -3, -2, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, -4, -2, 0, 0, 0, 0, 0, 0, -1, -2, -3, -2, -2, -2, -2, -1, 0, 0, 0, 2, 1, 0, 0, 0, 1, 3, -2, -2, -2, 0, -1, -1, 0, -1, -1, -1, -3, -2, -2, -2, -1, 0, 0, 2, 2, 0, 1, 1, 0, 1, 0, 2, -2, -1, -2, -1, -2, -2, -2, -1, -1, -2, -3, -2, 0, -1, 0, 0, 0, 0, 2, 3, 2, 2, 1, 2, 3, 3, -2, 0, 0, -2, -1, -1, -1, -3, -3, -3, -1, -2, -1, -2, 0, 0, 0, 2, 4, 4, 4, 1, 1, 1, 1, 2, -1, 0, 0, -2, -1, -3, -2, -3, -2, -1, 0, -1, 0, 0, -1, 0, 0, 2, 2, 3, 3, 0, 1, 0, 2, 4, 0, -1, -1, -1, -2, -2, -2, -1, -2, -3, -1, -1, 0, -2, 0, -1, 1, 2, 2, 2, 3, 2, 1, 1, 4, 5, 0, -2, 0, -2, -4, -3, -3, -3, -3, -3, -2, -1, 0, -1, -2, -2, -1, 0, 2, 3, 1, 0, 1, 2, 3, 6, -3, 0, -1, -1, -3, -2, -2, -3, -3, -1, -2, 0, -1, -1, 0, -1, 0, 2, 1, 1, 1, 1, 2, 2, 3, 5, -1, -1, 0, -2, -1, -3, -2, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 1, 1, 2, 2, 2, 1, 2, 3, 6, -3, -1, -2, -1, -1, -2, -2, -1, -2, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 2, 3, 2, 4, -2, -2, -2, -2, -2, 0, -3, -1, -2, -1, -2, 0, 0, -1, 0, -2, -1, 0, 0, 0, 0, -1, 1, 0, 1, 2, -3, -2, -2, -1, -1, -1, -1, -1, -1, -1, -2, -1, 0, 0, -2, -1, -1, -1, -1, 0, 0, 0, -1, 0, 2, 2, -2, -2, -1, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 1, -4, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, -5, -2, -1, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -3, -4, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, -5, -2, -1, 0, 1, 0, 1, 2, 3, 3, 1, 0, 1, -1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 2, 1, 1, -5, -2, -1, 0, 1, 2, 3, 4, 4, 4, 3, 4, 2, 0, 0, 1, 2, 1, 1, 1, 2, 3, 2, 3, 3, 3, -3, 0, 0, 2, 4, 4, 4, 6, 4, 4, 4, 6, 4, 4, 3, 4, 4, 1, 2, 2, 3, 3, 2, 2, 3, 2, -1, 0, 1, 1, 1, 1, 1, 2, 3, 3, 4, 3, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 0, 1, 2, 3, 3, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, -1, -1, 1, 1, 1, 2, 3, 2, 0, 0, 2, 2, 0, 0, -1, -1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 3, 4, 2, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 1, 2, 1, 2, 1, 1, 0, 1, -1, 0, 1, 2, 3, 3, 4, 3, 2, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 2, 2, 1, 1, 1, 0, 0, -2, 0, 0, 2, 1, 3, 4, 3, 2, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 2, 1, 1, 0, 1, 1, -3, -2, 0, 0, 2, 3, 1, 2, 0, 0, 0, -1, 0, 0, 0, -1, -1, -2, -1, 0, 0, 2, 1, 0, 0, 1, -2, -3, -2, -1, 1, 0, 0, 0, 0, 0, -2, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 2, -4, -3, -1, 0, 0, 0, 0, 0, -2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, -2, -1, -2, -2, -1, -2, -2, -2, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, -4, -3, -3, -2, -2, -1, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 2, 1, 1, 0, 2, 0, 0, 2, 2, -3, -2, -2, -2, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 1, 1, 0, 2, 2, -3, -3, -3, -3, -3, -2, -1, 0, 0, 0, 1, 0, 1, 2, 0, 2, 1, 0, 1, 1, 2, 2, 0, 0, 0, 1, -3, -3, -4, -3, -4, -2, 0, -1, 0, 0, 0, 1, 1, 0, 0, 2, 2, 0, 0, 3, 1, 1, 0, 1, 2, 2, -1, -1, -1, -3, -2, -2, -2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 2, 2, 2, 2, 1, 1, 3, 0, 0, -1, -2, -2, 0, -1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 1, 1, 2, -2, 0, -2, -2, -2, 0, -2, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 1, 1, 1, -2, -1, -2, -2, -2, -1, -1, 0, -1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 2, 0, 0, 0, -2, 0, 0, 0, 0, 1, 0, 1, 2, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 2, 2, 2, 0, 2, 2, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 3, 2, 1, 1, 2, 1, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 3, 1, 2, 2, 3, 1, 2, 1, 1, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 3, 1, 2, 1, 3, 2, 3, 2, 1, 1, 0, 0, 1, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 1, 1, 1, 2, 2, 3, 4, 2, 1, 2, 2, 2, 2, 1, 1, 0, 0, 1, 0, -1, 0, 0, 1, 1, 3, 4, 3, 3, 4, 5, 4, 5, 4, 3, 2, 3, 2, 2, 2, 3, 4, 3, 4, 3, 1, 2, 2, -1, 0, 1, 1, 1, 2, 3, 3, 3, 3, 1, 1, 2, 2, 2, 1, 1, 0, 2, 3, 2, 3, 2, 2, 2, 1, -2, -1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, 1, 2, 2, 2, 0, 0, 0, 0, 3, -3, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, -1, -1, -2, -1, -1, 1, 0, 0, 1, 1, 0, 0, 0, 1, 1, -2, -2, 0, 0, -1, 0, -1, -2, 0, -1, -1, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 2, -3, -1, 0, 0, -1, -2, -2, -2, -2, -1, -3, -1, -2, -1, -2, -1, -1, 0, 0, 0, -1, 0, 0, -1, 1, 1, -2, 0, -1, 0, -1, -2, -3, -1, -1, -4, -2, -3, -2, -2, -3, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, -3, -1, 0, -2, -2, -2, -3, -2, -2, -1, -2, -3, -3, -2, -2, -3, -1, 0, 0, -1, -1, 0, 0, 0, 0, 2, -1, -1, -1, -2, -2, -3, -1, -2, -2, -3, -2, -2, -2, -4, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 3, 0, 0, -1, -1, -1, -2, -1, -3, -1, -3, -2, -4, -3, -3, -2, -1, -2, -1, 0, -1, 0, 0, 0, 1, 1, 2, 0, 0, -1, -2, -1, -2, -1, -3, -3, -1, -4, -3, -2, -3, -4, -1, -2, -2, 0, -1, 0, 0, 0, 0, 1, 2, 0, -1, -1, -2, -1, -3, -2, -1, -2, -3, -3, -4, -4, -3, -4, -2, -1, 0, -1, 0, 0, 0, 0, 1, 0, 3, 0, -1, -1, -1, -2, -3, -3, -3, -2, -2, -3, -2, -2, -4, -3, -1, -2, -1, 0, 0, 0, 0, 0, 1, 2, 3, 0, -2, 0, -1, -3, -3, -4, -3, -3, -3, -3, -1, -3, -2, -2, -3, -2, -1, -1, 0, -1, 0, 0, 0, 0, 2, -1, 0, -2, 0, -1, -1, -4, -2, -4, -2, -2, -4, -2, -3, -2, -2, -1, -2, 0, 0, 0, 0, 1, 1, 1, 2, -1, -1, -2, -1, -2, -3, -4, -3, -2, -2, -2, -3, -3, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 2, 1, 2, -2, -2, -1, -2, -1, -3, -3, -3, -3, -3, -1, -1, -2, -1, -1, -1, -2, 0, -1, 0, 0, 0, 1, 0, 1, 2, -3, 0, -2, -1, -1, -3, -2, -1, -2, -1, -1, -2, -1, -1, -3, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, -2, -1, -1, -2, -1, 0, 0, -1, -1, -2, -3, -2, -2, -2, -2, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -2, -2, -1, -1, -2, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, -2, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, -3, -1, -2, -1, 0, 0, 0, 0, 0, -2, -1, -2, -2, 0, 0, -1, -1, 0, 0, 0, -1, 0, -2, -1, -2, -1, -3, -3, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, -2, 0, 0, -3, -1, 0, 0, 0, 1, 1, 1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, -2, -2, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, -2, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 2, 2, 0, 0, 1, 1, 1, 2, 2, 1, 0, 0, 1, 1, 0, -3, -1, 0, 0, 0, 2, 2, 1, 2, 2, 3, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 3, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 1, 1, 2, 3, 2, 2, 1, 0, 1, 0, 0, 0, 1, 0, 1, 2, 2, 2, 1, 1, 0, -1, 0, 0, 0, 2, 3, 1, 2, 2, 2, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 2, 0, 2, 0, 1, 0, 0, -1, -1, 0, 1, 2, 3, 3, 3, 1, 2, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -3, 0, 0, 0, 3, 2, 2, 3, 1, 2, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 2, 0, 0, 0, 1, -2, -2, 0, 0, 1, 1, 2, 3, 2, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, -1, 0, 1, -3, -1, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -4, -1, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -2, -2, -2, -2, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 2, 1, 1, 0, 1, 0, 0, -4, -1, -3, -2, -2, -1, -1, 0, -1, 1, 0, 2, 0, 2, 0, 0, 0, 0, 2, 3, 3, 2, 2, 0, 1, 0, -2, -2, -2, -3, -4, -3, -1, -2, 0, 0, 2, 1, 0, 2, 1, 0, 0, 1, 2, 2, 2, 1, 1, 0, 0, 2, -3, -1, -3, -2, -3, -3, -1, -2, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 1, 2, 2, 1, 2, 0, 2, 1, -3, -2, -2, -2, -3, -2, -3, -1, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 2, 2, 1, 1, 2, 2, 1, 2, -1, -1, -2, 0, -3, -2, -1, -2, -1, 0, 1, 1, 0, 1, 1, 0, 1, 0, 2, 3, 2, 1, 1, 2, 0, 3, -1, 0, -1, 0, 0, -2, -2, -1, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 2, 2, 2, 1, 2, 1, 2, -2, -2, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 1, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 1, 0, 0, 0, 1, 0, 1, 2, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 2, 2, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 3, 2, 2, 0, 1, 0, 1, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 3, 3, 3, 2, 3, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 2, 2, 3, 3, 2, 3, 2, 3, 2, 2, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 2, -2, 0, 0, 0, 1, 4, 2, 2, 2, 3, 2, 3, 3, 2, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, -1, -1, 1, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 1, -1, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 3, 1, 3, 2, 1, 2, 2, 2, 2, 3, 3, 1, 2, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 1, 0, 0, 1, 1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, -1, 1, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 2, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, -2, 0, -1, -1, -1, -1, -1, 0, 0, -1, 0, 1, 0, 0, 2, 0, 0, 0, 0, 2, 0, 0, 0, -2, -1, -1, -2, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, -2, -1, -2, -2, -2, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, -2, -1, -1, -2, 0, 0, 0, 0, 1, 0, 2, 1, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 1, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, -2, -2, -1, -1, 0, 0, 0, 0, -1, -1, -1, -2, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, -1, -2, 0, -2, 0, -1, 0, 0, 0, 0, 0, -1, -1, -2, 0, 2, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -2, -2, -3, -2, -1, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -3, -2, -1, -3, -2, -2, -2, 0, 0, -2, 0, 0, -2, 0, 0, 2, 0, 0, 0, -1, -1, 0, 0, -1, -1, -2, -3, -1, -2, -3, -3, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -2, -3, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, -1, -3, -2, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 2, 1, 1, 0, 0, 0, 0, -1, -1, 0, -2, -1, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 1, 2, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 1, 0, 1, 0, 1, 1, 1, 2, 3, 1, 1, 1, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 3, 3, 2, 3, 3, 2, 0, 0, 0, 2, 2, 1, 1, 1, 1, 1, 1, 2, 3, 2, 1, 3, 0, 0, 0, 2, 1, 2, 1, 2, 3, 2, 1, 0, 1, 0, 1, 0, -1, -2, -2, -1, -1, 0, 0, 2, 1, 2, -1, -1, 1, 1, 1, 1, 2, 1, 3, 1, 0, 0, 1, 0, 0, -1, -3, -3, -5, -4, -3, -1, 0, 0, 1, 3, -1, -1, 1, 0, -1, 0, 0, 0, 1, -1, 0, 0, 0, 0, -1, -1, -4, -3, -3, -3, -2, -1, 0, 2, 1, 2, 1, 0, 0, 0, 0, -1, -1, 0, -1, -2, 0, 0, 1, -1, -2, -3, -4, -4, -3, 0, 1, 1, 1, 1, 0, 2, 3, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -3, -3, -3, -2, 0, 1, 1, 0, 0, 0, -1, 1, 2, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -3, -2, 0, 0, 0, 0, 0, 0, 0, -2, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -3, -2, -4, -2, -1, -3, -3, 0, 0, 1, 2, 3, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -2, -3, -2, -4, -4, -3, -3, -2, -2, -2, -2, -1, 0, 2, 3, 2, 3, 1, 2, 0, 0, 0, 0, 0, -2, -2, -5, -4, -3, -3, -3, -4, -3, -3, -3, -2, -3, 0, 1, 2, 3, 4, 3, 2, 1, 0, -2, -1, -1, -3, -3, -5, -4, -4, -4, -4, -3, -1, -2, -1, 0, 0, -1, 0, 0, 2, 3, 3, 1, 0, 0, -1, -2, -3, -4, -5, -5, -4, -5, -3, -3, -3, -2, 0, 0, 0, 0, 0, 0, 0, 1, 5, 4, 1, 0, -1, -2, -1, 0, -1, -3, -4, -3, -5, -5, -3, -2, 0, 0, 1, 2, 2, 1, 0, -2, 0, 2, 6, 6, 2, 0, -2, 0, -1, 0, -1, -2, -2, -3, -3, -5, -2, -1, -1, 0, 0, 1, 1, 1, 0, 0, 0, 3, 4, 4, 0, 0, 0, 0, 0, 0, -2, -2, -4, -4, -2, -3, -3, -1, -1, -3, 0, 0, 1, -1, -1, -1, 1, 2, 3, 3, 0, 1, 0, 0, 0, -1, -3, -3, -3, -5, -4, -3, -2, -1, -1, -3, -1, 0, -1, -1, -1, -2, 0, 4, 4, 0, 0, 0, 0, -1, -3, -3, -6, -6, -4, -3, -3, -3, -3, -2, -2, 0, 1, 1, -1, -1, -1, 0, 1, 2, 3, 3, 1, 0, 1, 0, -1, -3, -3, -6, -4, -3, -2, -3, -1, 0, 0, 0, 2, 0, -1, -3, -3, 0, 2, 3, 4, 4, 2, 3, 2, 0, 0, -2, -2, -5, -3, -2, -2, -2, -2, -1, -1, 0, 0, -1, -2, -3, -2, 1, 4, 2, 3, 2, 3, 2, 0, -1, -2, -3, -4, -5, -3, -4, -4, -2, -4, -4, -3, -2, -2, -1, -3, -1, 0, 2, 4, 4, 4, 4, 3, 1, 0, -1, -2, -4, -4, -2, -2, -3, -5, -4, -4, -4, -4, -2, -2, -1, -2, 0, 0, 3, 4, 5, 6, 5, 4, 4, 0, -1, -1, -2, 0, -1, -2, -4, -4, -4, -6, -5, -4, -1, 0, 0, -1, 0, 1, 4, 4, 5, 5, 6, 4, 3, 0, -1, 0, 0, 0, -1, 0, -2, -2, 0, -2, -2, -2, -2, -1, -2, -1, 0, 1, 2, 4, 5, 3, 4, 3, 3, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -2, 0, 3, 3, 4, 4, 4, 5, 4, 2, 0, 1, 0, 0, 0, 0, 2, 1, 1, 1, 0, 2, 1, 0, 0, -2, 0, 1, 3, 5, 6, 5, 7, 6, 6, 4, 1, 1, 0, 0, 1, 2, 3, 2, 1, 3, 3, 3, 3, 1, 2, 0, 0, 1, 4, 7, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 1, 1, 2, 1, 1, 3, 1, 4, 4, 4, 4, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -3, -1, 0, 1, 0, 1, 3, 1, 2, 2, 2, 3, 1, 2, 0, 0, 0, 0, 0, 2, 2, 2, 1, 1, 0, -1, -1, 0, 0, 1, 1, 2, 3, 3, 2, 1, 1, 1, 2, 0, 0, 0, 0, 1, 1, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, 1, 2, 2, 1, 3, 2, 2, 2, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 2, 0, 1, 0, -1, -1, -1, 0, 1, 0, 2, 2, 2, 2, 2, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, -1, -1, -2, 0, 0, 0, 2, 1, 3, 4, 2, 1, 0, 0, -1, 0, -2, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, -1, -3, -1, 0, 0, 1, 3, 3, 2, 3, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -3, -1, -1, 0, 0, 0, 1, 2, 1, 1, 1, 1, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -2, -2, -2, -1, -1, 0, 1, 1, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -2, -3, -3, -3, -2, -1, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, -2, -4, -4, -4, -4, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, -3, -2, -4, -4, -4, -1, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, -1, -3, -2, -3, -4, -2, -3, -3, -1, -1, -1, -2, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 2, 0, 1, 1, 0, -1, -4, -3, -3, -2, -3, -3, -2, -2, -1, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, -1, -2, -3, -3, -3, -4, -2, -2, -3, -2, -1, -1, -1, -1, 0, 0, -1, 0, 1, 0, 2, 1, 1, 2, 1, 1, -1, -1, -2, -1, -3, -2, -2, -2, -1, -1, 0, 0, 0, 0, -1, -2, -1, 0, 0, 1, 1, 1, 1, 2, 2, 1, -2, -2, -1, 0, -2, -2, -3, -2, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 2, 0, 1, 2, 2, 1, 1, 1, -1, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 2, 1, 2, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 2, 2, 1, 0, -1, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 2, 0, 1, 1, 1, 0, -1, -1, 0, -2, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, -1, -1, 0, 0, 1, 1, 1, 0, -1, 0, -1, -1, -1, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -2, -1, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -3, -1, -1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 1, 3, 2, 2, 4, 2, 2, 3, 4, 2, 2, 1, 2, 2, 2, 0, 2, 0, 0, 0, 3, 1, 0, -1, 0, 0, 1, 2, 1, 2, 2, 2, 3, 1, 3, 3, 1, 1, 0, 0, 0, 0, 2, 0, 0, 0, 2, 0, 0, 0, -1, 0, 0, 1, 1, 0, 2, 1, 0, 0, 1, 0, 1, -1, -1, -1, -1, 0, 0, 0, 0, 1, 2, 0, -1, 0, 0, 0, 1, 0, 2, 2, 1, 0, 1, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -2, -1, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -2, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, -1, 0, -2, -1, -1, -2, -2, -2, 0, -1, 0, -1, 0, -1, 0, -2, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, -2, -1, -3, -1, -2, -1, -2, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 2, 0, 2, 1, 0, 0, -1, -1, -1, -2, -3, -2, -1, -2, -1, 0, 0, 0, 0, -2, -1, 0, 0, -1, 1, 0, 0, 2, 2, 0, 0, -1, 0, -1, -2, -1, -2, -2, -3, -2, -1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 1, 0, 2, 1, 0, 0, 0, -1, 0, -2, -2, -1, -3, -2, -1, -1, -2, -1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, -2, -1, -2, -2, -3, -1, -1, 0, 0, 0, 0, -1, -2, -1, -2, 0, -1, 2, 1, 0, 0, 0, -1, 0, 0, -2, -1, -2, -3, -2, -2, -2, -2, -1, -1, -1, 0, -2, -1, -2, -2, -1, -1, 2, 1, 0, 0, 0, 0, 0, 0, -1, -3, -4, -3, -3, -1, -1, 0, 0, -2, -2, -1, 0, 0, -2, -2, -1, 0, 2, 0, 0, -1, -1, 0, 0, -2, -1, -2, -2, -2, -1, -3, -1, -3, -1, -1, 0, -2, -2, -2, -2, -1, 0, 0, 2, 1, 0, -1, -1, 0, 0, -2, -3, -3, -4, -3, -3, -3, -1, -1, -2, -2, -1, -1, -2, -2, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, -2, -3, -3, -3, -3, -1, -1, -1, -3, -2, -3, 0, 0, 0, -3, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, -2, -3, -2, -3, -3, -2, -1, -1, 0, -1, -1, -1, 0, 1, 2, 1, 0, 0, 0, -2, -1, -1, -2, 0, -2, -1, -2, 0, -2, -2, -1, -2, -1, -2, 0, -1, -2, 0, -1, 0, 2, 0, 0, -1, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, -2, -1, 0, -2, -1, 0, 0, -1, 0, -1, 0, -1, 2, 1, 0, 0, 0, -1, -2, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -2, -1, 0, 3, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 1, 1, 1, 2, 1, 1, 0, 0, -1, -1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 0, 1, 2, 1, 0, 0, 0, 0, -1, -1, 3, 3, 2, 1, -1, 0, -1, -1, 0, 1, 0, -1, 0, -3, -4, -2, -2, -3, -1, -1, 0, -2, -3, -5, -6, -9, 4, 3, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -3, -3, -1, 0, 1, 1, 0, 0, -1, -3, -4, -6, 5, 4, 2, 2, 1, 1, 2, 0, 2, 1, 0, 0, -1, -1, -2, 0, 1, 2, 3, 2, 1, 0, -1, -1, -1, -5, 4, 4, 2, 1, 0, 1, 3, 3, 1, 1, 1, 0, 0, 0, 0, 0, 1, 3, 2, 4, 3, 2, 1, -1, -1, -4, 3, 2, 0, 0, 0, 3, 4, 3, 3, 2, 1, 1, 0, 0, 0, 0, 0, 1, 2, 1, 2, 1, 0, 0, 0, -2, 0, 0, 0, 0, 1, 4, 3, 5, 2, 3, 2, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, -1, -2, -3, -1, -1, 0, 1, 5, 3, 2, 2, 0, 2, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -2, -3, -2, 0, 1, 3, 1, 1, 2, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -3, -2, -4, -3, -2, -1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 1, 1, 0, 1, -2, -3, -4, -4, -2, -1, 0, 1, 1, 2, 0, 0, 1, 2, 2, 1, 0, 1, 1, 2, 0, 1, 2, 0, 1, 0, -1, -4, -4, -4, -4, -2, 0, 1, 3, 2, 3, 2, 0, 1, 0, 2, 0, 0, 0, 0, 0, 1, 3, 1, 1, -1, -3, -4, -5, -6, -5, -2, 0, 0, 3, 2, 3, 2, 3, 2, 2, 0, 0, 0, -1, 0, 0, 2, 2, 3, 1, 0, -2, -5, -5, -6, -5, -1, 0, 0, 1, 0, 1, 2, 3, 2, 1, 2, 0, 0, 0, 0, 2, 3, 2, 2, 0, 0, -2, -5, -7, -7, -4, -1, 0, 0, 0, 0, 1, 0, 0, 2, 2, 1, 1, 0, 0, 1, 1, 2, 2, 0, 0, -1, 0, -3, -5, -3, -2, -2, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, -1, -1, 0, 2, 3, 2, 2, 0, 0, 0, 0, -2, -3, -2, -2, -1, -1, 0, 0, 0, 1, 2, 1, 1, 0, -2, -1, 0, 1, 3, 3, 3, 2, 0, -2, -3, 0, -1, -3, -1, -2, -2, 0, 0, -1, 1, 1, 2, 1, 1, -1, -1, -2, -1, 0, 2, 4, 3, 2, 0, -2, -3, 2, 0, -2, 0, 0, -1, 0, 0, 2, 0, 3, 3, 1, 0, 0, -1, 0, 0, 2, 2, 3, 2, 0, -1, -2, -1, 1, 1, 0, 1, 0, 1, 0, 2, 2, 4, 4, 2, 0, 0, 0, 0, 1, 2, 1, 3, 4, 2, 2, 1, 0, -2, 4, 2, 2, 0, 1, 0, 1, 3, 3, 3, 4, 0, 0, -1, 0, 1, 1, 2, 3, 1, 2, 3, 1, 0, 0, -1, 4, 4, 3, 3, 3, 3, 1, 2, 2, 2, 2, 0, -1, 0, 0, 1, 1, 2, 2, 0, 1, 1, 2, 0, 0, -1, 5, 5, 3, 4, 3, 2, 4, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, -1, 0, -1, 4, 4, 4, 4, 4, 3, 4, 4, 3, 1, 1, 0, 1, 1, 0, 1, 2, 1, 0, 0, -1, -1, 0, -2, 0, -2, 3, 4, 2, 2, 3, 2, 3, 2, 2, 0, 0, 0, 1, 0, 0, 0, 1, 2, 2, 0, 0, -2, -1, -3, -2, -3, 1, 1, 2, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, -2, -2, -3, -4, -2, -6, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, -2, -2, -2, -2, -3, -2, -1, -1, -2, -3, -2, -5, -4, -7, -8, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, -1, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -1, -3, -3, -4, -4, -2, -1, 0, 0, 0, 0, 0, 4, 2, 3, 2, 0, 1, 1, 0, -2, 0, -1, -2, -1, 0, 0, -3, -2, -3, -2, 0, 1, 0, 0, 0, 0, 1, 3, 3, 3, 0, 0, 0, 1, 0, -2, 0, -1, -2, -1, -2, -2, -1, -3, -2, -1, 1, 0, 0, 1, 0, 1, 0, 2, 3, 1, 1, 0, 0, 0, 0, -2, -2, -2, -3, -4, -1, -2, -1, -3, -2, -1, 0, 2, 1, 1, 1, 1, 2, 2, 2, 0, 0, 0, -1, -1, -2, -3, -3, -5, -4, -3, -1, 0, -1, -1, -1, 0, 0, 1, 2, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, -1, -2, -3, -4, -5, -2, -1, 0, 0, -2, -2, 0, 2, 2, 1, 1, 0, 1, 2, 0, 0, -1, -1, -2, -1, 0, 0, 0, -1, -3, -2, -2, -1, 0, 0, 0, 0, 0, 2, 3, 0, 1, 0, 3, 3, 1, 0, 0, 0, 0, 0, 1, 1, 1, -1, -3, -1, 0, 0, 0, 1, 1, 0, 3, 4, 2, 0, 0, 2, 2, 0, 2, 0, 1, 1, -1, 0, 1, 1, 2, -1, -3, -1, 0, 0, 0, 1, 1, 1, 3, 3, 2, 2, 1, 2, 0, 1, 1, 1, 0, 0, 0, 0, 2, 1, 0, -1, -1, -2, 0, 0, 0, 2, 3, 3, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -2, -2, -2, -3, 0, 2, 1, 3, 3, 3, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, -1, 0, 0, 1, 2, 1, 3, 2, 2, 1, 0, 1, 3, 2, 2, 1, 0, -1, 0, -2, 0, 0, 0, -2, -1, -3, -1, 0, 0, 1, 2, 3, 3, 1, 1, 2, 1, 0, 1, 3, 1, 2, 2, 0, -1, 0, -1, 0, -1, -2, -1, -3, -2, -1, 0, 1, 2, 2, 1, 0, 1, 0, 0, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -3, 0, 0, 0, 1, 2, 3, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -3, -4, 1, 0, 0, 3, 4, 1, 1, 2, 0, 2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 2, 0, 1, 0, -2, -3, 0, 0, 0, 2, 3, 3, 3, 2, 3, 1, 1, 0, 0, 1, 0, 1, 1, 1, 1, 0, 1, 2, 1, 0, -2, -4, 0, -1, 0, 1, 1, 1, 2, 2, 3, 2, 1, 1, 0, 0, 1, 2, 1, 2, 2, 2, 1, 3, 2, 1, -1, -2, 0, 0, -1, 0, -1, 0, 0, 2, 2, 1, 1, 0, 0, 1, 0, 1, 2, 3, 1, 2, 1, 2, 5, 4, 0, -2, -2, -1, -2, -2, -1, 0, -1, 2, 3, 2, 0, 0, 1, 1, 0, 1, 1, 4, 2, 3, 2, 4, 5, 3, 2, 0, -3, -3, -4, -4, -5, -1, -1, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 4, 5, 4, 0, -2, -3, -2, -2, -5, -5, -4, 0, 0, 0, 0, 0, 2, 0, 1, -1, 0, 0, 1, 0, 1, 2, 2, 2, 3, 0, -1, -3, -3, -3, -5, -3, -3, 0, -1, 0, 0, 0, 1, 2, 0, 0, 0, 1, 0, 1, 0, 1, 1, 2, 1, 0, -1, -2, -3, -4, -4, -4, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 2, 1, 1, 2, 0, -3, -3, -2, -4, -5, -6, -3, -1, -2, -2, 0, -2, -2, -2, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, -4, -2, -2, -3, -6, -6, -5, -3, -2, -2, -2, -2, -4, -5, -3, -2, -1, 0, -1, -1, 0, 0, 1, 0, 1, 0, -3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, -1, 1, 1, 0, 0, -1, 0, 0, 0, -1, 0, -2, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, -1, 0, 0, 0, -2, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, -1, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, 1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 1, -1, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, -1, -3, -4, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -4, -1, -2, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 2, 1, 1, -1, -1, -1, -1, -3, -2, -2, -3, -2, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, -1, -1, -1, 1, 0, 0, 0, -1, -1, -1, -2, -2, -3, -4, -2, -1, 0, -1, -1, -2, 0, -1, 0, 0, 0, -2, -1, 0, -1, -1, 0, 0, -1, -2, -1, -3, -3, -4, -3, -4, -3, -3, -1, 0, 0, 0, 0, 0, -1, -1, -1, -3, -2, 0, -1, 0, 0, -1, -1, -1, -2, -2, -1, -3, -2, -4, -4, -1, 0, 0, -1, 0, 0, -1, 1, -1, -1, -2, -2, 0, -1, 0, -1, -1, -2, -3, -2, 0, -1, -2, -3, -4, -3, -3, -2, -1, -1, 0, -1, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, -1, 0, -2, -2, 0, 0, -1, -3, -5, -4, -2, -3, -3, -1, 0, 0, -1, -2, -1, -2, 0, -1, -1, -1, -1, 0, -2, -1, 0, -1, 0, -1, -2, -3, -4, -4, -3, -1, -2, -1, -2, -1, -1, -1, -2, -2, -2, -1, -2, -2, -2, -1, -2, -1, -1, 0, 0, -2, -3, -2, -2, -4, -3, -2, -2, -2, -1, -3, -2, -3, -4, -1, -1, -1, -2, -2, 0, -2, -3, -2, -1, -1, 0, -1, -2, -1, -2, -2, -2, -3, -3, -2, -3, -4, -2, -3, -3, -2, -3, -1, -2, -2, -2, -2, -2, -3, -1, -2, -1, 0, -2, -2, -3, -2, -2, -1, -2, -4, -4, -3, -3, -3, -5, -3, -4, -3, -1, -2, -1, -2, -1, -3, -1, 0, -1, -1, -2, -1, -2, -2, -3, -2, -2, -2, -3, -3, -3, -4, -4, -4, -4, -1, -2, -3, -1, -1, -1, -1, -2, -2, -1, -3, -4, -2, -3, -1, -1, -1, -1, -3, -3, -3, -4, -3, -3, -2, -3, -2, -3, -1, 0, 0, -1, -1, 0, 0, -1, -2, -4, -1, -1, -2, -2, -1, -3, -2, -2, -4, -4, -3, -2, -3, -4, -2, -1, -1, -2, 0, 0, 0, 0, 0, -2, -3, -4, -1, -2, -1, 0, -2, -2, -1, -4, -2, -2, -2, -2, -4, -3, -3, -2, -1, 0, -1, 0, 0, 0, 0, -2, -2, -3, -2, -1, -2, -2, -1, -2, -1, -3, -1, -1, -1, -3, -4, -1, -3, 0, -1, 0, 0, -1, 0, 0, 0, 0, -2, -3, -1, -1, -3, -3, -2, -1, -1, -2, -1, -1, -1, -3, -2, -1, -3, -1, -1, 0, 0, -1, -1, 0, 1, 0, -1, -4, -3, -4, -3, -4, -2, -3, -3, -3, 0, -1, -2, -3, -2, -1, -3, -3, -3, -3, -2, -1, -1, 0, 0, 0, 0, -2, -2, -5, -5, -5, -3, -3, -2, 0, -1, -1, -2, -2, -3, -3, -3, -4, -3, -2, -2, -1, 0, 0, 0, 0, -2, -4, -2, -3, -3, -4, -4, -2, -2, 0, -1, -2, 0, -2, -2, -1, -4, -4, -4, -1, 0, 0, -1, 0, -1, 0, 0, -3, -5, -3, -3, -4, -3, -3, -3, -1, -3, -3, -2, -3, 0, -2, -4, -4, -1, -2, 0, -1, 0, -1, -1, -1, -1, -3, -4, -5, -3, -4, -5, -2, -3, -2, -1, -4, -2, -3, -3, -2, -2, -3, -2, -1, 0, 0, -2, -1, 0, 0, -2, -2, -3, -5, -5, -4, -4, -2, -3, -2, -4, -4, -3, -3, -5, -3, -3, -1, 0, -2, 0, -1, -1, -1, -1, 0, -1, -4, -4, -4, -5, -5, -5, -2, -2, -3, -3, -2, -4, -4, -4, -4, -4, 0, -2, -2, 0, -1, -1, -1, 0, -3, -3, -4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, -1, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, -1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, -1, 0, -2, -2, -2, 0, 0, -3, -4, -5, -5, -5, 2, 1, 0, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 2, -1, -2, -4, -4, -2, 4, 2, 1, 2, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 2, 0, 0, -2, -2, -1, 3, 4, 2, 1, 1, 3, 4, 2, 0, 1, 0, 0, 0, 0, 1, 0, 0, 2, 3, 4, 3, 2, 0, -1, 0, 1, 2, 3, 3, 0, 3, 4, 5, 3, 3, 0, 1, 0, -1, 1, 0, 0, 0, 0, 2, 2, 0, 2, 0, -1, 0, 0, 1, 3, 2, 1, 3, 6, 5, 5, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 3, 3, 6, 4, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 0, -2, -2, -2, 1, 2, 3, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, -1, -3, -3, -3, -1, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 2, -1, -3, -4, -4, -2, 0, 0, 2, 1, 1, 0, 1, 0, 1, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, -1, -3, -4, -4, -4, -1, 0, 1, 3, 4, 2, 0, 0, 2, 2, 0, 0, 1, 2, 1, 0, 0, 1, 0, 1, 1, -2, -2, -5, -5, -5, 0, 0, 2, 4, 5, 3, 3, 2, 4, 0, 2, 1, 1, 2, 1, 0, 0, 0, 2, 1, 2, -1, -5, -6, -4, -4, -1, 0, 2, 2, 4, 4, 3, 2, 2, 2, 1, 1, 0, 0, 1, 1, 1, 0, 1, 2, 0, -2, -4, -5, -4, -4, -1, 0, 1, 2, 4, 2, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 2, -2, -3, -4, -3, -4, -1, 1, 2, 2, 2, 1, 2, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 1, -1, -2, -2, -3, -3, -1, 0, 0, 2, 1, 1, 0, 1, 0, 1, 0, 0, -2, 0, 1, 0, 2, 1, 0, 0, -1, 0, -1, -1, -2, -1, -1, 0, 0, 1, 2, 3, 0, 1, 0, 0, 0, 0, -1, 0, 0, 2, 2, 2, 2, 0, -2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 3, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, -2, 2, 1, 0, 0, 0, 0, 2, 1, 3, 4, 3, 1, 0, -1, -2, 0, 0, 1, 0, 0, 0, 1, 2, 1, -1, 0, 1, 0, 0, 1, 0, 0, 3, 3, 3, 4, 4, 0, -1, -1, -2, 0, 0, 0, 0, 1, 1, 1, 1, 1, -1, -1, 2, 2, 1, 3, 3, 3, 4, 3, 4, 3, 2, 1, -1, -2, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, -1, 4, 3, 3, 4, 4, 2, 2, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 1, 0, -1, -1, 2, 4, 4, 4, 3, 3, 1, 2, 0, 0, -1, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -2, 3, 4, 3, 4, 3, 1, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, -2, -1, 0, 0, -2, 2, 1, 4, 3, 3, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, -1, -1, -2, -2, -1, -2, -2, 1, 1, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -2, -1, 0, -1, -2, -2, -2, -3, -4, -6, 0, -1, 0, 0, 1, 3, 3, 4, 2, 1, 3, 2, 2, 1, 3, 3, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 2, 3, 2, 1, 1, 2, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 2, 1, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 2, 0, 0, 0, 0, -1, 0, -1, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -2, -2, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -2, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, -2, -2, -2, -2, -1, -2, -2, 0, 0, 0, -1, -2, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, -2, -2, 0, 0, 0, -1, -1, 0, 0, 0, 1, 2, 1, 0, 0, 1, 2, 1, 0, 0, -2, 0, -1, -1, -3, -1, -2, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 2, 0, 0, 1, -1, 0, 0, -2, -2, -3, -3, -2, -2, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -2, -2, -2, -3, -1, -2, -3, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 2, 1, 2, 1, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 2, 0, 1, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, -2, -1, -2, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 2, 0, 1, 0, 0, -1, 0, -1, -1, -1, -3, -1, -3, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, -2, -3, -2, -3, -3, -2, -1, 0, -2, -1, -1, 0, 0, 0, 0, -1, 0, -1, 1, 0, 1, 0, -1, 0, 0, -1, -2, -3, -2, -3, -3, -2, -3, -1, -3, 0, -1, 0, -1, -1, 0, -1, 0, 0, 2, 0, 0, -1, 0, 0, -1, -1, -2, -2, -1, -1, 0, -3, -2, -1, -1, -2, -2, 0, 0, 0, -1, -1, 0, 1, 2, 0, 0, 0, -1, 0, 0, 0, -1, -1, -2, -2, -1, -2, -1, -2, -2, -1, -2, 0, 0, -1, 0, 0, 1, 1, 1, 2, 0, 0, 0, -2, -1, 0, 0, 0, 0, -2, -1, -2, 0, -1, 0, -1, -2, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 0, 0, 0, 2, 2, 2, 1, 1, 0, 0, 0, 1, 2, 1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 2, 0, 1, 1, 1, 3, 3, 1, 0, 2, 1, 0, 0, 0, 2, 2, 0, 1, 2, 2, 2, 3, 2, 3, 2, 0, 2, 2, 2, 0, 1, 0, 1, 1, 1, 0, 2, 3, 1, 3, 1, 1, 2, 1, 0, 0, 1, 2, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 2, 1, 0, 1, 0, 0, 1, 0, 3, 1, 1, 1, 0, 0, 1, 0, -1, -1, -1, -1, -1, 0, 0, 1, 1, 1, 1, 0, 1, 2, 0, 0, 0, 0, 1, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 2, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, -1, 0, 1, 0, 0, 2, 0, 0, 1, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, -1, -2, 0, 0, 1, 0, 0, -1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 1, 1, 1, 3, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -2, -2, -3, -2, -2, 0, -1, 0, 0, 0, 0, 1, 1, 0, 2, 0, 0, 0, 0, -1, -1, -2, -1, -2, -1, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, -1, 1, 1, 2, 1, 0, 0, -1, 0, 0, -2, -2, -2, -2, -2, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 3, 2, 2, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 0, -1, 0, 0, 1, -1, 0, 0, 0, -1, -1, 0, 0, -1, -1, -2, 0, 0, -1, -1, -1, -1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, -2, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 1, 1, 1, 1, 1, 0, 0, -2, -2, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 2, 1, 2, 1, 1, 2, 0, 0, -1, 0, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 3, 2, 2, 1, 1, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -2, -2, 0, -2, -2, 0, -1, 0, -1, -1, 0, 0, 1, 2, 1, 2, 1, 2, 2, 0, 0, 0, -1, -1, 0, -1, -1, -3, -2, -3, -1, -1, 0, -1, 0, 0, 0, 0, 2, 2, 4, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -2, -2, -1, -1, 0, 0, 1, 0, 1, 2, 2, 4, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, -1, 1, 0, 0, 1, 1, 2, 2, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 3, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 1, 1, 3, 3, 2, 2, 1, 1, 2, 1, 1, 1, 0, 0, 1, 1, 1, 2, 1, 0, 2, 1, 0, 1, 0, 1, 1, 3, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 1, 2, 2, 2, 1, 0, 1, 0, 0, 1, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 1, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, -2, 0, 0, 0, -1, -1, -1, -2, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -2, 0, 0, -2, 0, -1, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, -2, -1, -1, -3, -1, -2, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, -1, -2, -2, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -2, -2, -1, -2, -2, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -2, 0, -1, -1, -1, 0, -1, 0, -1, 0, -1, 0, -1, 1, 1, 0, 0, 0, 0, -1, 0, -1, -1, -2, -1, 0, -2, -1, 0, -1, 0, -1, -1, 0, 0, -1, -1, 0, -1, 1, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, -1, 0, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, -2, -1, -2, 0, -2, -2, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -2, 0, 0, -2, 0, -1, 0, -1, -1, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 3, 0, 0, 0, 1, 0, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 2, 0, 1, 2, 1, 0, 0, 0, 1, 2, 0, 2, 2, 3, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 0, 1, 1, 0, 1, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 1, 2, 1, 1, -1, 0, 0, -1, 0, 0, 0, 1, 1, 2, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 1, 1, 1, 0, 2, 1, 1, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 0, 2, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 0, 0, 2, 0, 2, 2, 1, 0, 0, -1, -1, -1, -1, -2, 0, -1, -1, 0, 0, 1, 0, 0, 1, 1, 2, 0, 1, 2, 0, 1, 1, 1, 1, 0, 0, 0, -1, 0, -1, -1, -2, -1, -1, 0, 0, 1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -2, -2, -2, -1, 0, 0, 0, 1, 0, 1, 0, -1, -1, 0, 2, 1, 1, 1, 0, 1, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 2, 0, 2, 2, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 3, 2, 2, 1, 0, 1, 2, 1, 1, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 1, 1, 1, -1, 1, 1, 1, 1, 0, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, -1, 1, 1, 1, 0, 1, 0, 2, 2, 1, 1, 0, 0, 2, 0, 0, 0, 1, 1, 2, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 1, 0, 1, 2, 1, 2, 1, 2, 1, 0, 0, 2, 3, 2, 1, 0, -1, -1, 2, 1, 0, 0, 0, 2, 2, 0, 1, 2, 0, 0, 2, 1, 1, 1, 1, 0, 2, 3, 3, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 2, 1, 2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 1, 2, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 1, 2, 1, 0, 0, 0, 1, 2, 0, 0, 1, 1, 1, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 2, 1, 1, 1, 1, 3, 0, 2, 0, 0, 1, 1, 0, 1, 0, 1, 3, 1, 2, 0, 1, 1, 1, 0, 1, 0, 1, 2, 1, 1, 1, 3, 0, 1, 1, 0, 1, 0, 0, 0, 1, 1, 0, 2, 1, 2, 0, 1, 0, 0, 1, 0, 0, 0, 1, 2, 1, 3, 2, 1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 2, 1, 0, 1, 0, 0, 2, 0, 2, 0, 3, 2, 2, 3, 2, 1, 0, 0, 0, 1, 1, 2, 2, 0, 1, 1, 0, 0, 0, 1, 1, 2, 2, 2, 2, 4, 3, 1, 3, 2, 1, 1, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 3, 2, 2, 3, 2, 2, 0, 1, 1, 0, 1, 1, 2, 1, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 2, 1, 0, 1, 1, 0, 2, 2, 2, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 2, 0, 0, 1, 0, 0, 0, 2, 1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 2, 1, 2, 2, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 2, 3, 1, 2, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 1, 2, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, -1, 0, -1, -1, -1, -2, 0, -1, 0, 1, 2, 2, 0, 0, 2, 0, 0, 1, 0, 1, 1, 2, 1, 0, 0, 0, -1, -1, -3, -2, -3, -1, -1, -1, 1, 0, 1, 0, 0, 0, 0, 1, 2, 2, 2, 0, 1, 2, 2, 2, 1, -1, 0, -1, -1, -3, -2, -3, -1, -2, -1, 0, 1, 1, 0, 1, 0, 2, 0, 0, 2, 2, 0, 1, 0, 1, 1, 0, 1, 0, 0, -1, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 2, 0, 0, 0, 1, 1, 0, -1, 0, -1, -1, 0, -1, 0, -1, 1, 1, 1, 3, 2, 1, 0, 2, 3, 3, 4, 2, 2, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 2, 1, 1, 3, 3, 1, 3, 3, 1, 2, 2, 2, 0, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 3, 1, 1, 1, 2, 2, 1, 1, 2, 1, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 2, 2, 1, 3, 3, 1, 1, 1, 2, 1, 3, 3, 1, 1, 1, 2, 2, 0, 2, 0, 0, 1, 0, 0, 1, 1, 0, 1, 2, 1, 3, 3, 2, 2, 2, 2, 1, 2, 2, 3, 2, 3, 2, 1, 2, 2, 1, 1, 0, 0, 2, 1, 0, 2, 1, 2, 4, 4, 3, 2, 1, 1, 2, 2, 2, 3, 3, 2, 3, 3, 2, 2, 1, 1, 1, 0, 0, 0, 1, 0, 1, 1, 2, 2, 3, 2, 2, 1, 1, 2, 3, 2, 2, 1, 2, 0, 0, 3, 3, 2, 0, 0, 0, -1, 0, -1, 0, 1, 1, 1, 1, 0, 0, 1, 2, 2, 0, 0, 1, 2, 1, 2, 2, 1, 2, 1, 2, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 2, 2, 2, 1, 2, 2, 0, 1, 1, 0, 1, 2, 1, 1, 3, 3, 2, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 2, 1, 3, 1, 1, 1, 0, 0, 0, 1, 1, 2, 3, 1, 2, 2, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 2, 1, 2, 3, 3, 3, 1, 0, 0, 1, 3, 3, 2, 2, 3, 3, 2, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 2, 1, 3, 2, 1, 2, 1, 1, 1, 1, 4, 2, 3, 4, 2, 2, 0, 0, 0, 2, 0, 0, 0, 1, 0, 2, 0, 2, 3, 1, 2, 0, 0, 2, 3, 2, 4, 3, 3, 3, 0, 0, 0, 2, 2, 1, 4, 2, 4, 2, 3, 3, 2, 0, 0, 1, 1, 1, 2, 0, 1, 0, 0, 0, 0, -1, 0, 1, 2, 2, 1, 2, 3, 3, 3, 3, 2, 1, 0, 0, 0, 0, 1, 0, 2, 2, 3, 1, 2, 1, 0, 0, 0, 0, 0, 2, 1, 3, 4, 3, 2, 1, 3, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 1, 3, 3, 3, 3, 2, 3, 2, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 1, 0, 0, -2, -1, 0, 0, 2, 4, 2, 2, 3, 1, 1, 0, 0, 0, -2, -1, 0, 0, 0, 2, 1, 0, 1, 0, 0, 0, -2, 0, 0, 2, 1, 2, 2, 3, 2, 0, 0, 1, -1, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, -3, -2, -1, 0, 0, 0, 3, 2, 2, 0, 0, 0, 0, -1, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -4, -3, -3, -1, -1, -1, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, -4, -4, -3, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, -4, -4, -5, -4, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 2, 1, 1, -4, -3, -3, -3, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, -3, -2, -5, -3, -4, -2, -2, -3, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 1, 0, 1, 2, 2, 2, -3, -3, -2, -4, -3, -4, -3, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 2, 2, 2, 2, 3, -1, -3, -2, -4, -3, -3, -2, -2, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 1, 2, 2, 1, 3, 2, 3, 3, -2, -3, -3, -3, -3, -2, -3, -2, -1, -2, 0, 0, 1, 0, -1, 0, -1, 1, 0, 1, 3, 1, 2, 3, 1, 1, -1, -1, -3, -2, -2, -3, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 1, 2, 3, 1, 2, 0, 0, 0, -2, -1, -2, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 1, 3, 1, 1, 0, 0, -1, -1, -2, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 1, 1, 0, 1, 2, 1, 2, 1, 0, -2, -1, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, -2, -1, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 2, 2, 2, 1, 0, 0, 1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 2, 2, 2, 2, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, 0, -1, 0, 0, 1, 2, 1, 2, 2, 1, 0, 0, 0, -2, 0, -1, -1, 0, -1, -1, -1, -1, -2, -2, -3, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, -1, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 2, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 1, 0, 2, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, -2, 0, -1, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, -1, -1, -1, 0, 0, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, -2, -1, -2, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, 0, 1, 1, 0, -1, -1, -1, 0, 0, -1, 0, -2, 0, -1, 0, 1, 1, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, -1, -3, -2, -4, 1, 1, 3, 0, 2, 0, 1, 1, 0, -1, -1, 0, 0, 0, 0, -2, -1, 0, 1, 0, 0, 1, -1, 0, -2, -2, 1, 2, 2, 1, 1, 0, 1, 2, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 2, 0, 2, 0, 0, 0, 0, 0, 2, 1, 2, 1, 0, 1, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 1, 0, -1, 0, 1, 1, 2, 1, 0, 0, 3, 3, 2, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 2, 0, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 4, 2, 2, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 2, 2, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 1, -2, -1, -2, -1, 0, 0, 1, 3, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, -1, -2, -2, -2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -2, -1, -2, -3, -2, -1, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -2, -2, -1, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -2, -2, -3, -3, -3, -3, -1, 0, 0, 0, 2, 0, 1, 1, 2, 1, 0, -1, -1, 1, 0, 1, 0, 0, 0, 1, 0, -1, -3, -2, -3, -3, -1, 0, 1, 2, 2, 2, 0, 1, 0, 1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 1, 0, -3, -3, -3, -2, -2, 0, -1, 0, 0, 2, 1, 1, 1, 0, 0, 1, -1, -1, 0, 1, 2, 2, 0, 0, 1, -1, -2, -2, -2, -2, 0, -2, -1, 0, 0, 2, 0, 0, 0, 0, -1, 0, -1, -1, 0, 1, 1, 1, 0, -1, 0, -1, -2, 0, -1, -3, -1, -1, 0, 0, 0, 0, 2, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 2, 0, 0, -1, 0, 0, -1, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, -1, -2, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -2, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 2, 0, 1, 2, 2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 4, 3, 1, 1, 1, 1, 0, 2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 2, 2, 2, 1, 2, 1, 1, 2, 2, 2, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 2, 2, 3, 1, 3, 2, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 2, 1, 3, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 2, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -2, -2, -2, -1, -2, 0, 0, 1, 2, 2, 0, 2, 0, 0, 0, 2, 2, 2, 2, 1, 1, 0, 0, 0, 1, 0, 2, 1, 1, 2, 3, 0, 0, 0, 1, 2, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 1, 1, 1, 2, 0, 2, 0, 0, 0, 2, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 2, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 2, 1, 0, 1, 0, 2, 1, 0, 0, -2, -1, -3, -1, -2, -2, 0, 0, 0, 0, -1, 0, -1, 1, -1, 0, 0, -1, 0, -1, -4, -4, 3, 1, 0, -1, -1, -1, -2, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -2, 0, -1, 0, 0, -1, -2, -4, 2, 0, -1, -3, -3, -2, -2, -1, 1, 0, 2, 1, 1, 1, 0, -1, -2, -1, -2, -2, -1, 0, -1, -2, -3, -5, 0, 0, -2, -2, -2, 0, -2, 0, 1, 0, 1, 1, 2, 0, 1, -1, 0, -2, -1, -2, 0, 0, 0, -1, -2, -3, 1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 1, 2, 2, 2, 1, 0, -2, -2, 0, -1, -1, 0, 0, -1, -3, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 2, 1, 1, 1, 0, 0, -1, 1, 0, 1, -1, -2, 1, 1, 0, 1, 2, 1, 1, 2, 1, 0, 0, 0, 2, 1, 0, 2, 2, 2, 2, 1, 0, 3, 2, 0, 1, -2, 2, 1, 1, 0, 1, 2, 3, 4, 1, 1, 2, 0, 0, 1, 2, 3, 3, 5, 2, 3, 2, 3, 2, 1, 2, 0, 4, 3, 2, 3, 2, 3, 4, 4, 3, 0, 1, 0, 1, 0, 0, 1, 2, 3, 1, 1, 2, 3, 1, 2, 0, 0, 4, 2, 2, 2, 4, 6, 5, 5, 3, 1, 0, 1, 2, 1, 2, 1, 1, 0, 0, 0, 1, 2, 2, 0, 0, -2, 5, 1, 0, 2, 4, 6, 6, 5, 1, 1, 1, 1, 2, 2, 2, 2, 0, 0, 0, 0, 0, 1, 1, 0, -1, -1, 2, 1, 0, 2, 3, 4, 4, 4, 3, 0, 0, 2, 1, 2, 2, 3, 1, 2, 0, -1, 0, -2, -2, -1, 0, -1, 1, 0, 0, 0, 1, 4, 3, 2, 0, 0, 1, 1, 1, 3, 3, 3, 3, 1, 0, 0, -1, -2, -3, -2, -1, -4, 2, 0, 0, 0, 2, 2, 1, 1, 0, 0, 0, 0, 1, 1, 2, 2, 2, 0, 1, 0, 0, -1, -2, -2, -2, -4, 2, 1, 2, 0, 2, 3, 4, 2, 0, 0, 0, 0, 1, 2, 2, 0, 1, 0, 0, 1, 0, 0, -1, -2, -1, -3, 4, 2, 0, 2, 3, 3, 2, 1, 1, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -4, -3, 4, 3, 0, 0, 3, 3, 2, 0, 1, 1, 0, 0, 0, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, -1, -3, -2, 4, 1, 0, 1, 1, 2, 1, 1, 1, 0, 1, 1, 2, 0, 2, 1, 2, 1, 0, 0, 1, 3, 0, 0, -1, -3, 3, 3, 1, 0, 1, 1, 1, 1, 1, 0, 1, 1, 1, 2, 2, 1, 0, 1, 0, 2, 3, 4, 2, 1, -1, -2, 4, 3, 1, 1, 2, 2, 3, 1, 1, 2, 2, 2, 1, 0, 0, 1, 1, 0, 3, 4, 4, 5, 4, 0, 0, -2, 3, 1, 0, 0, 1, 2, 2, 1, 1, 1, 2, 3, 1, 1, 0, 1, 1, 1, 2, 2, 5, 3, 3, 1, 1, -1, 1, 1, 0, 1, 0, 1, 3, 1, 1, 3, 4, 3, 4, 1, 1, 1, 0, 1, 1, 2, 2, 1, 1, 0, 1, 0, 2, 0, 1, 0, 0, 1, 0, 2, 3, 2, 3, 3, 3, 2, 1, 0, 0, 0, 1, 2, 1, 2, 1, 0, 0, 0, 1, 0, -1, 0, 0, -1, 1, 1, 1, 2, 2, 2, 2, 1, 1, 0, 0, 1, 2, 2, 1, 0, 0, 0, -1, -2, 1, 0, -1, -2, -2, -2, 0, 0, 1, 1, 2, 2, 1, 0, 2, 1, 1, 2, 2, 2, 2, 1, 0, 0, -1, -3, 0, 1, -1, -1, -2, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 1, 1, 1, 2, 1, 0, -2, -3, -4, 4, 4, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -2, -1, -3, -2, 4, 3, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, -2, -1, 3, 2, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 3, 2, 2, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, 1, 0, -1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, -1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 2, 0, -1, 0, 0, 1, 2, 1, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 1, 0, 2, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 2, 1, 1, 2, 0, 0, -1, 0, 1, 0, 0, 1, 0, -1, 0, -1, -2, -1, 0, 0, 0, 0, 1, 1, 2, 1, 2, 0, -1, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, -1, 1, 0, -1, 0, -1, 1, 0, 2, 1, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 1, 0, 2, 1, 1, 0, 0, 1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -2, 1, 0, -2, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, -1, -3, 2, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 1, -1, -1, -2, -2, 2, 0, 0, 0, -2, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -2, 0, -1, 0, 0, 0, 0, -1, -2, -1, 2, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, -2, -2, -2, -1, -2, 0, 0, 0, 0, -1, 0, -1, 0, 3, 3, 1, 0, 1, 0, 0, 1, 0, 0, 0, -2, -1, -2, -2, -2, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 4, 3, 2, 3, 1, 1, 1, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, -1, -1, -1, 1, 0, 0, 0, 0, 0, 5, 4, 3, 2, 3, 1, 1, 2, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, -1, 5, 4, 3, 3, 3, 1, 2, 2, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -1, 0, -2, -1, 4, 3, 3, 4, 2, 2, 2, 0, 2, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -2, -2, 0, -3, 4, 4, 2, 1, 1, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, -1, -1, -2, -1, -3, -4, 4, 3, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, -2, -4, -4, -4, 1, 0, 0, 0, 0, -1, -2, -1, -2, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, -3, -5, -6, -6, -6, -2, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 1, 1, 1, 3, 3, 1, -1, -1, 1, 1, 0, 0, -1, 0, 0, 0, -3, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 2, 1, -2, 0, 0, 1, 0, 0, 0, 0, 0, -1, -4, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 1, -1, -1, 0, 1, 0, -2, -2, -1, -1, -3, -4, -3, -1, 0, 0, 0, -1, 0, 0, -2, 0, 0, 0, 0, 1, 3, -2, -1, 1, 0, -1, -1, -2, 0, 0, -3, -3, -3, -1, -1, -1, -1, -1, -2, 0, -1, -1, 0, 0, 0, 0, 1, -2, -1, 0, 2, -1, -3, -2, -1, -1, 0, -2, -2, -2, -3, -4, -4, -2, -1, 0, 0, 0, -1, -1, -1, -1, 1, -2, 0, 0, 0, -1, -2, -2, -2, 0, -1, -1, -1, -3, -3, -4, -5, -4, -2, 0, 0, -1, 0, -2, -1, -1, 0, -3, -2, 1, 1, -2, -3, -1, -2, 0, -2, -2, -1, -3, -2, -2, -4, -3, -2, -1, 0, 0, 1, 0, 0, 0, 0, -2, -1, 0, 0, 0, -2, -1, -1, -2, -2, -2, -1, -1, -1, -4, -3, -3, -4, -1, 0, 0, 0, 0, 0, -1, 0, -4, -1, 0, 1, 0, 0, -2, -3, -2, -2, -1, 0, -1, -3, -2, -4, -5, -2, -3, 0, 0, 2, 2, 0, 0, 0, -3, 0, 1, 2, 0, -1, -2, -1, -3, -2, -3, -1, -2, -3, -4, -3, -3, -4, -3, -1, 0, 2, 3, 0, -1, 0, -3, 0, 1, 2, 0, 0, 0, 0, -2, -2, -2, -2, -2, -5, -3, -3, -4, -3, -2, -1, 1, 3, 2, 0, 0, 0, -1, 1, 2, 1, 0, 0, 0, 1, 0, -2, -1, -1, -3, -4, -4, -4, -4, -4, -4, -3, 0, 1, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -3, -2, -3, -2, -2, -2, 0, 2, 2, 0, 0, 0, 0, 2, 2, 0, -1, 0, 1, 2, 1, -1, -1, 0, -2, -2, -4, -2, -3, -3, -3, -3, 0, 2, 0, 0, 1, 1, -1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, -1, -2, -2, -4, -3, -3, -1, -2, -1, 0, 0, 0, 0, 2, 1, -2, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -2, -4, -3, -2, -1, -2, -2, 0, 0, -1, 0, 1, 1, -1, 1, 1, 0, -1, 0, 0, -1, -1, -1, 0, 0, -1, -2, -1, -2, -1, -1, -1, -1, -1, 0, -2, -1, 0, 3, -2, 0, 0, 0, -2, -1, -2, 0, -1, -2, -1, -1, 0, -1, -2, -3, -2, -1, -1, -1, -1, -3, -3, -1, 0, 3, -1, 1, 0, 0, 0, -1, 0, -3, -3, -1, -1, -2, -2, -3, -3, -2, -4, -1, -2, -2, -2, -4, -2, 0, 1, 3, -2, -1, 0, 0, 0, 0, -2, -2, -2, 0, -2, -1, -2, -2, -3, -4, -4, -1, -1, -2, -1, -4, -1, 0, 1, 3, 0, 0, -1, 0, 0, -1, -1, -3, -3, -2, 0, -1, -1, -1, -2, -3, -3, -2, 0, 0, -1, -2, -2, 0, 2, 3, -1, -2, -1, 0, 0, -1, -2, -1, -1, 0, -1, 0, -2, 0, -1, -2, -3, -2, 0, 0, -1, -1, -1, 1, 2, 4, -2, -3, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 4, 5, -3, -2, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 2, 4, 5, -2, -4, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 4, 4, 7, 2, 2, 1, 2, 1, 2, 1, 0, 1, 1, 2, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 2, 1, 0, 1, 1, 1, 1, 1, 1, 1, 0, 1, 2, 2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, -1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 1, 0, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 2, 1, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 2, 2, 2, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 1, 1, 2, 2, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 2, 1, 1, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 1, 1, 2, 0, 1, 1, 0, 0, 1, -1, 0, -1, -2, 0, 0, -1, 0, -1, 1, 0, 1, 0, 1, 0, 0, 0, 1, 2, 0, 1, 2, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 2, 2, 2, 1, 1, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 1, 2, 2, 3, 0, 0, 0, 1, 2, 1, 1, 2, 2, 2, 2, 0, 0, 0, 1, 0, 2, 1, 2, 0, 0, 1, 2, 2, 1, 0, 1, 0, 2, 0, 2, 1, 2, 1, 2, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 0, 0, 1, 2, 2, 0, 0, 1, 1, 2, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 2, 1, 1, 1, 1, 0, 2, 2, 2, 2, 2, 1, 2, 1, 2, 3, 1, 2, 0, -1, 1, 1, 1, 2, 2, 1, 1, 1, 3, 1, 2, 1, 1, 0, 0, 1, 2, 3, 3, 3, 3, 3, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 3, 1, 1, 2, 1, 1, 1, 2, 2, 1, 1, 0, 2, 0, 2, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 1, 0, 2, 2, 0, 0, 2, 1, 1, 2, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 2, 1, 2, 1, 2, 1, 1, 1, 1, 1, 0, 1, 1, 1, 2, 0, 0, 1, 1, 0, 0, 1, 1, 2, 1, 1, 1, 1, 3, 3, 2, 2, 2, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 2, 1, 1, 3, 1, 0, 0, 1, 2, 0, 1, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 2, 3, 2, 2, 2, 2, 2, 2, 2, 0, 0, 0, -1, -1, 0, 1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 1, 2, 3, 2, 3, 2, 3, 3, 2, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 2, 1, 2, 3, 4, 0, 0, 1, 1, 2, 2, 3, 4, 4, 2, 4, 2, 2, 2, 3, 4, 1, 3, 3, 2, 1, 2, 2, 1, 1, 1, 2, 1, 1, 1, 1, 2, 2, 2, 2, 1, 2, 1, 2, 2, 2, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 2, 1, 0, 0, 1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, -2, -1, -1, -1, -1, 1, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, -1, 0, 0, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 1, -1, -1, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, -2, -2, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 2, 2, 2, 1, 0, 0, 0, -2, -1, 0, -2, -1, -2, 0, -1, 0, 0, -1, 0, 1, 1, 0, -1, 1, 1, 2, 2, 3, 1, 1, 0, -1, -1, 0, -2, 0, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 2, 1, 0, 2, 1, 2, 1, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 2, 1, 1, 1, 2, 1, 0, 0, -1, -2, -2, -1, -1, -2, 0, -1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, -1, 0, -3, -1, -1, 0, -1, -1, -1, 0, 0, 1, 0, -1, -1, 0, -1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -2, -1, 0, 0, 0, 1, 0, -2, -1, 0, 0, -1, 0, 2, 1, 0, 1, 0, 0, 1, -1, -1, -2, -1, -1, -2, -2, 0, -1, 0, -1, 0, 0, 0, -2, -2, -2, -1, 0, 1, 1, 1, 0, 0, 0, 0, -1, -1, -2, -1, -2, -2, -2, -2, -1, 0, 0, 0, -1, -1, -2, -1, -1, -1, -1, 2, 0, 0, 0, 0, 0, 0, -1, -3, -1, -2, -1, -2, -3, -2, -1, 0, 0, -1, -2, -1, -1, 0, -1, -1, 0, 3, 1, 0, 0, 0, -1, 0, 0, -2, -2, -2, -4, -3, -1, -2, -1, -2, -2, -1, -1, -1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, -3, -3, 0, 0, -1, -1, -2, -1, 0, -1, 0, 0, -2, 0, 0, 0, 2, 1, 0, 1, -1, -1, 0, -1, 0, -1, 0, 0, 0, -2, 0, -1, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, 4, 2, 0, -1, -2, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, -2, -2, -1, -2, 0, 0, -1, -1, -1, 0, 0, 3, 2, 1, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, 0, -1, 0, 0, 0, 3, 2, 0, 0, 0, -1, 0, -1, 0, 1, 0, 1, 0, 2, 1, 1, 0, 0, 0, 1, 1, 0, -1, -2, 0, 0, 3, 0, 0, -1, 0, -1, -2, 0, 1, 0, 0, 1, 0, 2, 0, 2, 2, 1, 2, 1, 0, 0, -1, -2, -1, -2, 2, 1, 0, 0, -1, 0, 0, -1, 0, 1, 2, 2, 1, 2, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0, -1, -1, -2, 0, 0, 2, 1, 3, 2, 3, 4, 3, 2, 1, 2, 2, 0, -1, 0, 0, 0, 2, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 3, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 1, 0, -2, 0, -1, 0, -1, 0, 0, 1, 3, 3, 2, 0, 1, 0, 0, 1, 0, -2, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 2, -1, 0, 0, 1, 3, 3, 3, 0, 1, 0, 0, 0, 0, -2, 0, -1, 0, 0, 2, 1, 2, 0, 0, 0, 2, 3, -1, 1, 0, 2, 2, 4, 2, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 2, 2, 0, -1, 0, 2, 3, 4, 2, 0, 0, -1, 0, -2, 0, 0, -1, 0, -1, -2, 0, 0, 1, 0, 0, 0, 1, 3, -2, 0, -1, 1, 2, 3, 2, 1, 0, -1, -1, -1, -1, -2, -2, -2, 0, 0, -2, 0, -1, 0, -1, 0, 1, 3, -4, -3, -1, 0, 0, 0, 0, -1, -2, -2, -1, -1, -2, -2, -1, -1, -2, -1, -2, -2, -1, 0, 0, 0, 2, 5, -4, -5, -3, -2, 0, 0, -1, -3, -2, -2, 0, 0, -2, -2, -2, -2, 0, -1, 0, -2, -2, 0, 0, 0, 0, 4, -4, -6, -4, -5, -2, -2, -2, -2, -2, -2, -2, -1, -1, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 4, -4, -6, -5, -4, -3, -3, -2, -1, -1, -1, -1, -1, 0, 0, 0, -1, 1, 0, 0, 1, 0, -1, 0, 0, 1, 2, -3, -5, -5, -7, -4, -2, -2, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 3, 4, -4, -4, -6, -5, -5, -3, -2, -1, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 5, -5, -5, -5, -6, -3, -2, -1, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 1, 2, 5, -5, -3, -4, -4, -2, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 2, 2, 3, 6, -2, -3, -3, -3, -2, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 2, 0, 0, 1, 1, 3, 4, -2, -3, -2, -2, -2, -1, -1, -1, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -3, -3, -2, -2, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, -1, -2, -1, 0, 0, 0, -1, 1, 1, 0, 0, 0, -3, -2, -1, 0, 0, 0, 1, 0, 1, 2, 2, 0, 0, -1, -2, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 2, 3, 0, 0, -2, -1, -2, -2, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 2, 2, 1, 0, -2, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 3, 1, 2, 1, 1, 1, 0, 0, -2, -2, -2, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 2, 1, 0, 1, 1, 3, 2, 2, 1, 0, 1, 0, 0, 0, -1, -1, 0, 1, 1, 0, 0, 0, 0, 1, 2, 2, 2, 1, 1, 0, 2, 3, 3, 1, 1, 3, 2, 1, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 0, -1, 2, 2, 3, 3, 2, 3, 2, 2, 3, 2, 2, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, -1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 2, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 2, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, -1, -2, 0, 0, -2, -1, 0, 1, 1, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 2, 1, 0, 1, 1, 1, 0, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 1, 1, 2, 0, 0, 2, 0, 0, 0, 0, 1, 0, -1, -2, -1, 0, -1, 0, 0, 0, -1, -2, -1, 1, 0, 1, 3, 1, 1, 0, 0, 0, 2, 0, 1, 1, 1, 0, 0, 0, -2, -2, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -2, 0, -1, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, 1, 0, -1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 1, 1, 0, 0, -2, -1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 0, 1, 1, 0, -1, -2, -1, -1, 0, 1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 1, 1, 1, 2, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 2, 2, 3, 1, 1, 2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 2, 2, 3, 2, 2, 0, 1, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 2, 1, 3, 5, 3, 5, 6, 6, 6, 6, 6, 5, 5, 4, 4, 5, 5, 5, 2, 3, 2, 1, 0, 0, -1, 0, 0, 0, 1, 2, 4, 4, 4, 3, 4, 5, 5, 4, 1, 1, 1, 3, 4, 4, 1, 2, 2, 1, 0, -3, -1, -1, 0, 0, 2, 3, 5, 5, 5, 3, 3, 3, 3, 2, -1, 0, 0, 1, 2, 2, 2, 2, 1, 0, -2, -3, -2, 0, 0, 0, 0, 1, 4, 3, 2, 3, 2, 3, 3, 1, 0, 0, -1, -1, 0, 0, 2, 0, 0, 0, -2, -2, -2, -1, 0, 0, 2, 3, 2, 4, 4, 4, 5, 5, 2, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 2, 3, 2, 4, 2, 1, 1, 0, 0, 0, 0, 1, 2, 1, 1, -1, 3, 0, 0, 0, 1, 3, 2, 2, 2, 1, 1, 2, 1, 3, 2, 3, 2, 0, 2, 2, 2, 2, 3, 1, 0, -1, 2, 0, 0, 0, 2, 1, 3, 3, 3, 3, 3, 1, 0, 1, 2, 2, 1, 1, 1, 2, 1, 2, 2, 2, 1, -1, 1, 2, 0, 1, 4, 4, 4, 4, 4, 3, 0, 0, 1, 1, 3, 1, 2, 3, 2, 2, 0, 0, 2, 3, 1, -1, 2, 1, 2, 3, 3, 5, 5, 2, 2, 1, 0, 0, 1, 1, 2, 3, 1, 2, 1, 0, 0, 1, 1, 0, 0, -3, 1, 0, 1, 2, 4, 4, 5, 3, 3, 1, 2, 1, 3, 1, 2, 1, 2, 2, 1, 0, 1, 0, 0, -1, -1, -2, 3, 2, 2, 3, 4, 4, 5, 3, 2, 2, 2, 2, 3, 1, 2, 2, 3, 1, 3, 0, 0, 0, 0, 0, 0, -1, 2, 3, 1, 1, 3, 5, 5, 2, 3, 2, 0, 0, 1, 2, 2, 3, 1, 3, 3, 2, 1, -1, -2, -2, -2, -1, 4, 2, 1, 3, 2, 3, 2, 3, 2, 2, 0, 0, 1, 2, 1, 1, 1, 3, 1, 1, 0, -1, -2, -2, -3, -1, 5, 4, 3, 2, 3, 1, 1, 2, 2, 2, 0, 0, 0, 0, 1, 0, 3, 2, 3, 1, 0, 0, -1, -1, -3, -1, 7, 3, 4, 3, 3, 1, 3, 2, 2, 1, 0, 0, -1, 0, 0, 2, 3, 2, 2, 0, 0, 0, -1, -1, -1, -3, 5, 3, 2, 2, 2, 1, 3, 1, 2, 1, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, -1, 0, -1, 0, -3, -2, 6, 4, 0, 2, 0, 2, 1, 1, 0, -2, -1, 0, 0, 0, 1, 0, 2, 1, 2, 0, 2, 1, 0, 1, 0, 0, 6, 1, 0, 1, 2, 2, 2, 1, 0, 0, 0, -1, 0, 0, 2, 0, 2, 0, 3, 2, 3, 3, 1, 1, 1, 0, 5, 3, 0, 1, 1, 3, 1, 1, 0, 0, 0, 0, 1, 0, 0, 2, 1, 0, 1, 4, 5, 3, 3, 1, 2, 1, 5, 3, 1, 1, 1, 2, 1, 1, 1, 0, 2, 2, 1, 2, 2, 0, 0, 1, 1, 3, 6, 3, 2, 0, 3, 1, 5, 2, 0, 0, 0, 0, 0, 2, 1, 2, 2, 1, 4, 2, 2, 2, 0, 2, 1, 5, 5, 4, 2, 1, 3, 3, 3, 3, 1, 0, 0, 0, 0, 2, 2, 2, 3, 3, 3, 4, 2, 2, 1, 2, 3, 5, 5, 4, 2, 3, 2, 2, 5, 3, 2, 0, 0, 0, 0, 0, 4, 5, 3, 5, 4, 4, 4, 3, 3, 3, 4, 5, 4, 4, 2, 2, 2, 0, 4, 3, 1, 0, 0, 0, 2, 1, 3, 4, 4, 4, 4, 4, 5, 4, 5, 3, 4, 5, 4, 3, 3, 1, 1, 0, 6, 2, 0, 1, 0, 0, 0, 1, 0, 2, 4, 5, 5, 6, 4, 5, 4, 5, 5, 7, 5, 3, 2, 3, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -3, -3, -3, 3, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -2, -2, 1, 2, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, -1, -2, -1, -2, -3, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, -1, -2, -2, 2, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 1, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 2, 1, 1, 0, 0, 1, 0, 2, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 1, 2, 2, 2, 1, 1, 0, 2, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, -1, -2, -2, 0, 0, -1, -1, 1, 1, 0, 1, 2, 2, 0, 1, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, 1, 0, 1, 1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 1, 1, 0, 0, -1, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 2, 1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, -1, 0, -2, -1, 0, 1, 2, 1, 0, 0, 0, 0, -2, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -2, 0, 2, 0, 1, 0, 0, 0, 0, 1, 1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 1, 1, 0, 0, 0, 0, 2, 1, 0, 0, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 3, 2, 1, 1, 1, 0, 0, 0, 1, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 1, 2, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 3, 2, 2, 2, 2, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, 1, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, -1, 0, -1, 0, -2, -2, -2, -2, -3, 1, 1, 0, -1, -2, -1, -2, -1, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -3, -2, -3, -5, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, -1, -1, 1, 1, 2, 0, 1, 2, 1, 2, 2, 0, 1, 2, 2, 1, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, -2, 0, -1, 1, 1, 0, 0, 1, 0, 2, 1, 1, 1, 1, 0, 1, 0, -1, 0, 2, 1, 1, 0, 0, 2, 2, -2, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 1, 0, 2, -2, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 2, -1, 0, 0, 0, 1, 0, -1, -1, 0, -1, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -2, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -2, 0, 0, 0, 0, 0, 0, -2, -1, -1, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 2, -1, -2, 0, 0, -1, 0, -2, -2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, -1, -2, -1, 0, -1, 0, 0, -2, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, -1, -1, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 2, 1, 0, -1, -1, 0, -2, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, -2, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 2, 1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -2, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 2, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 2, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -2, -2, 0, -1, -1, -1, -2, -2, 0, 0, 0, 0, 1, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 2, 0, 0, 0, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 1, 1, 2, 1, 2, 0, 1, 1, 2, 0, 1, 0, 0, 0, -1, -1, 0, 1, 1, 1, 2, 2, 2, 1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 3, 1, 2, 0, 1, 0, 0, 0, -1, 0, 1, 0, 1, 1, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 2, 3, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, 0, 0, 1, 1, 2, 2, 2, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, -2, 0, 0, -1, -1, -2, 0, -1, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 2, 0, 1, 1, 0, -3, -2, -1, -1, -2, -2, 0, 0, -1, 0, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, 2, 2, 2, 1, 0, 0, -1, -2, -1, -1, -3, -1, -1, -1, 0, 1, 1, 2, 1, 2, 1, 1, 0, 1, 0, 1, 0, 2, 1, 1, 0, 0, 0, -1, -2, -1, -2, -1, 0, 0, 0, 0, 1, 1, 3, 1, 0, 2, 2, 0, -1, 0, 0, 1, 1, 0, 1, 0, -2, -1, -1, -1, -3, -1, 0, -1, 0, 0, 1, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, -2, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, -1, 0, -1, 0, 2, 1, 0, 1, 0, 0, -2, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 1, 0, 0, 2, 2, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 0, 1, 0, 1, 0, 0, 2, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 2, 0, 2, 2, 1, 0, 1, 2, 1, 0, 2, 0, 1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 1, -1, -1, 0, 1, 0, 0, -1, -1, -2, -1, -1, -1, 0, 0, 0, 2, 0, 1, 0, 1, 2, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 1, 0, 2, 1, 3, 2, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -3, -4, 0, 1, 1, 0, 2, 1, 3, 2, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 0, 2, 1, 0, 0, 0, 0, 1, 2, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, -1, 0, 1, 2, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 2, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 3, 1, 0, 0, 1, 0, 0, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -2, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -2, -4, -2, -2, -2, 0, 0, 0, 0, 0, -1, -2, -2, 0, -2, -2, 0, 0, 0, 0, -1, -1, 0, 0, 2, 0, 0, -3, -3, -2, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, -1, -1, -2, -2, -2, -1, -2, -2, -2, -2, -1, -1, 0, 0, -2, 0, -1, -1, -1, 0, -1, 0, 0, 2, 1, 1, 0, -2, -1, -3, -1, -2, -2, -1, -1, -1, -1, -2, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 1, 0, -2, -3, -3, -2, -2, -3, -3, -2, -1, -2, -1, -1, -2, -1, -1, -2, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, -2, -3, -2, -2, -1, -2, -2, -2, -2, -2, -1, -2, -1, -1, -2, -2, -1, 0, 1, 0, 1, 2, 2, 1, 1, 0, -1, 0, -1, -2, -3, -2, -2, -1, -1, -2, -1, -2, -2, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -3, -2, -2, 0, -1, -2, 0, 0, -2, -2, -1, 0, 1, 1, 2, 0, 2, 1, 1, 0, -1, -1, -1, 0, -2, -1, 0, -1, -2, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 1, 3, 2, 1, 1, -1, -2, -1, -1, -1, -2, -1, -2, -2, 0, 0, -1, 0, -1, -2, -2, -1, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, -1, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, -1, 0, 0, 0, 1, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 1, 1, 1, 0, 0, 0, -1, -2, 0, -1, -2, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 1, 0, 0, -2, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -3, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, -2, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, -3, -3, -2, -2, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 2, 2, 4, 3, 4, 4, 5, 6, 6, 5, 3, 4, 4, 5, 5, 4, 6, 5, 5, 5, 5, 2, 3, 3, 3, -1, 1, 2, 2, 3, 3, 2, 2, 2, 5, 4, 2, 3, 4, 3, 3, 4, 3, 4, 2, 2, 4, 1, 2, 2, 2, -3, 0, 1, 1, 1, 1, 2, 1, 2, 3, 0, 2, 2, 2, 3, 2, 1, 2, 2, 2, 1, 2, 0, 0, 1, 4, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 2, -4, -2, -2, -1, 0, -1, -2, 0, -1, 0, -2, -2, 0, -2, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, -3, -3, -3, -2, -1, -2, -2, -1, -3, -2, -2, -1, -2, -2, -2, -1, -1, -2, -2, 0, -1, 0, -1, 0, 0, 2, -4, -3, -1, -2, -3, -2, -2, -2, -2, -4, -3, -3, -2, -3, -3, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 3, -3, -3, -3, -1, -3, -2, -4, -3, -4, -2, -3, -2, -3, -2, -3, -3, -1, -1, 0, 0, 1, 1, 1, 0, 0, 2, -3, -1, -2, -2, -1, -4, -3, -2, -3, -4, -4, -3, -4, -2, -2, -3, -2, -1, 0, 0, 1, 0, 1, 1, 1, 3, -2, -1, -1, -3, -2, -3, -4, -3, -4, -3, -3, -5, -4, -3, -3, -3, 0, 0, 0, 1, 1, 1, 2, 2, 2, 3, 0, 0, 0, -2, -2, -4, -3, -3, -3, -4, -5, -5, -5, -3, -3, -2, -1, -1, 0, 1, 1, 0, 1, 0, 1, 3, -1, 0, -1, -1, -2, -3, -4, -2, -3, -5, -4, -5, -3, -3, -4, -3, -2, -1, 0, 0, 2, 0, 1, 0, 1, 3, 0, 0, 0, -2, -3, -3, -4, -4, -4, -5, -3, -4, -4, -4, -4, -3, -2, -1, 1, 0, 2, 0, 0, 1, 1, 3, -1, 1, -2, -2, -3, -4, -2, -3, -3, -5, -4, -3, -3, -5, -4, -3, -1, 0, 0, 2, 1, 2, 0, 0, 2, 4, 0, 0, -2, -1, -2, -2, -3, -4, -3, -5, -3, -4, -3, -4, -3, -3, 0, 0, 0, 1, 0, 1, 1, 0, 1, 4, 0, -2, -2, -1, -1, -2, -2, -3, -2, -2, -3, -4, -4, -2, -3, -1, -1, 1, 0, 1, 1, 2, 0, 0, 1, 4, -3, -1, -1, -1, -3, -1, -3, -3, -4, -3, -2, -4, -3, -3, -1, 0, -1, 0, 1, 1, 0, 2, 1, 1, 1, 2, -2, -2, -2, -3, 0, -2, -1, -1, -3, -3, -1, -2, -2, -1, 0, -1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 2, -3, -2, -1, -1, -1, -1, 0, -1, -2, -3, -2, -1, 0, 0, -1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -4, -3, -2, 0, 0, -1, -1, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, -1, -1, -2, -2, -1, 2, -4, -3, -3, -1, -1, 0, 0, 0, -1, -2, 0, 0, -1, 0, 1, 0, 0, 0, 1, 1, 0, -1, -3, -1, -1, 0, -5, -4, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, -1, -3, -1, -1, 0, -4, -4, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 1, 0, 2, 2, 0, 0, 0, 0, 0, -1, -2, 0, -4, -3, -1, -1, 0, 2, 1, 0, 1, 0, 1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -4, -3, -2, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 0, 1, 2, 0, 0, 1, 1, 1, 1, 0, 0, 1, 1, -3, -1, 0, 0, 1, 1, 3, 2, 1, 1, 1, 1, 2, 3, 3, 1, 1, 3, 3, 1, 2, 2, 2, 1, 1, 3, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 1, 1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 1, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 2, 0, 0, 1, 0, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 1, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, -1, -1, 0, -2, -1, -1, -1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -2, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, -2, -1, -2, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, -1, -1, -1, -2, -3, -1, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, -1, 0, -1, -1, -2, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -2, -2, -1, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, -2, 0, -1, -1, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -2, 0, 0, -1, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -2, -3, -3, -1, 0, -1, -2, 0, 0, 0, -1, 0, 0, 0, 2, 0, 1, 1, 0, -1, -1, -1, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, -1, -2, 0, -1, -1, -1, 0, -1, 0, 1, 0, 0, 1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -2, 0, 2, 2, 2, 1, 1, 2, 0, 1, 3, 3, 2, 3, 3, 5, 6, 7, 6, 6, 6, 6, 5, 4, 1, 3, 2, 0, 1, 2, 2, 2, 2, 1, 3, 2, 3, 3, 3, 2, 2, 3, 5, 6, 5, 6, 4, 4, 5, 4, 2, 1, 3, -2, 0, 0, 1, 0, 0, 0, 1, 2, 4, 3, 2, 2, 3, 2, 3, 4, 4, 5, 5, 2, 3, 0, 0, 2, 2, -2, -2, 0, 0, 0, 0, 1, 2, 2, 3, 4, 3, 4, 2, 2, 3, 4, 4, 3, 1, 1, 0, 0, 0, 0, 0, -3, -2, -1, 0, 0, -1, 0, 0, 1, 1, 4, 2, 1, 1, 2, 3, 3, 1, 3, 0, 0, 0, 0, 0, 0, 0, -4, -3, -1, 0, -1, 0, 0, -1, 0, 2, 1, 3, 1, 2, 2, 1, 2, 2, 0, 1, 1, 0, 0, 0, 1, 0, -4, -3, 0, 0, -1, -1, 0, 0, 1, 1, 2, 1, 1, 0, 1, 2, 0, -1, 0, -1, 0, 1, 0, -1, 0, 0, -3, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -3, -3, 0, 0, -1, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, -2, -1, -1, 0, 1, 2, 1, 0, 0, -3, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, 2, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, -1, -1, -2, -2, -2, -2, 1, 1, 2, 1, 2, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -3, -1, -3, 2, 3, 3, 4, 1, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -2, -3, -2, 1, 1, 3, 2, 3, 1, 1, 0, 1, 2, 0, 2, 1, 0, 2, 1, 1, 1, 0, 0, 0, 0, -1, -1, -2, -1, -1, 2, 2, 2, 2, 0, 1, 2, 2, 1, 2, 0, 1, 2, 1, 4, 1, 1, 2, 1, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 2, 1, 1, 1, 4, 4, 4, 2, 2, 3, 2, 2, 1, 0, 0, -1, -2, -2, -2, -1, 1, 1, 2, 0, 2, 1, 1, 4, 2, 3, 3, 3, 3, 3, 5, 4, 4, 3, 2, 0, 0, 0, -5, -4, -2, -1, 0, 0, 2, 1, 0, 0, 1, 2, 2, 1, 3, 2, 4, 3, 4, 5, 4, 3, 2, 0, -2, 0, -4, -5, -4, -2, -1, 0, 3, 2, 0, 1, 1, 3, 2, 1, 4, 3, 2, 4, 4, 4, 2, 2, 1, 0, 0, -1, -5, -6, -5, -2, -1, 1, 2, 0, 0, 1, 1, 2, 2, 1, 3, 2, 3, 2, 3, 4, 2, 2, 1, 0, -1, -1, -5, -6, -6, -3, 0, 0, 1, 1, 0, 2, 1, 1, 3, 3, 2, 2, 3, 2, 2, 3, 2, 2, 0, -1, -1, -2, -6, -5, -5, -2, 0, 0, 1, 0, 0, 1, 0, 3, 2, 3, 2, 3, 3, 2, 2, 4, 4, 3, 1, 0, 0, -1, -6, -6, -6, -3, -1, -1, 2, 0, 1, 1, 1, 3, 2, 1, 2, 2, 2, 2, 3, 2, 4, 3, 2, 0, -1, 0, -6, -5, -5, -3, -2, -1, 1, 2, 0, 0, 1, 2, 3, 4, 4, 3, 4, 3, 4, 4, 3, 4, 3, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 1, 1, 1, 1, 3, 2, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 2, 3, 1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 2, 0, 1, 0, 2, 0, 0, 0, 0, -1, 0, 1, 1, 2, 2, 3, 2, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -2, 0, 1, 2, 0, 3, 2, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -2, 0, 0, 0, 0, 2, 2, 2, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -3, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, 1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, -2, -2, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, -2, -1, -2, -2, -3, -3, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -2, -1, -1, -3, -2, -3, -2, 0, 0, 1, 2, 0, 2, 1, 1, 2, 0, 0, 2, 2, 2, 0, -1, -1, 0, 1, 0, -1, -2, -3, -2, -3, -1, 0, 0, 1, 0, 1, 3, 1, 0, 1, 0, 1, 1, 1, 0, 1, -1, -1, 0, 0, -1, 0, -2, -4, -2, -1, 0, -1, 1, 2, 1, 0, 0, 1, 2, 2, 1, 2, 1, 1, 1, 0, 0, -2, 0, 1, -1, 0, -1, -4, -2, -2, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -2, -2, -1, -2, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 2, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -2, -2, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, -1, -2, -1, -1, -1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, -1, -2, -2, -1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 3, 2, 3, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 2, 0, 1, 2, 3, 3, 2, 0, 0, 1, 0, 2, 1, 1, 0, 2, 1, 1, 2, 1, 0, 1, 0, 0, 1, 2, 2, 0, 0, 2, 3, 2, 1, 2, 1, 1, 2, 2, 2, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 3, 1, 1, 0, -2, 0, -2, -2, -3, -2, -2, 0, -2, -3, -2, -2, -2, -1, -1, -1, -2, -3, -4, -2, -5, -5, 4, 1, 1, 0, -1, -2, -2, -3, -1, 0, 0, 0, 0, -2, -1, 0, -1, 0, 0, -1, 0, -1, -2, -2, -3, -5, 4, 2, 1, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, -4, 3, 2, -1, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, 3, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, 1, 0, -1, 0, 1, 0, 1, 1, 1, 1, 2, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 2, 0, 0, 0, 0, 2, 1, 2, 0, 1, 2, 2, 2, 1, 0, 2, 2, 0, 0, 1, 1, 0, 0, 0, 0, -1, 2, 0, -1, 0, 0, 2, 1, 2, 1, 1, 3, 3, 2, 1, 1, 1, 1, 0, 1, 1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 1, 2, 1, 1, 3, 2, 3, 1, 0, 1, 1, 2, 2, 0, 2, 0, 0, 1, 2, 1, 1, 1, 0, -1, 0, 1, 0, 2, 3, 2, 3, 1, 1, 2, 1, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, -1, 0, 1, 1, 3, 5, 1, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, -2, -3, -1, 1, 1, 3, 4, 1, 0, 1, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 1, 0, -2, 0, -1, -1, -1, 0, 1, 1, 3, 3, 2, 2, 0, 2, 2, 2, 0, 2, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -3, -3, -1, -1, 0, 2, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 2, 1, 1, 0, 0, -4, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 0, 1, 0, 0, 0, 2, 2, 2, 2, 1, -1, 0, -2, 3, 2, 0, 0, 0, 0, 0, 1, 1, 0, 2, 2, 1, 0, 0, 0, 1, 1, 0, 2, 2, 1, 1, -1, -1, -3, 3, 2, 1, 1, 1, 1, 1, 1, 2, 1, 3, 0, 0, 0, 0, 0, 2, 2, 0, 1, 1, 0, 2, 0, -2, -2, 2, 2, 1, 0, 1, 2, 0, 2, 2, 4, 2, 0, -1, -1, 0, 0, 0, 1, 1, 2, 1, 2, 4, 3, 1, 0, 3, 3, 1, 1, 2, 0, 1, 2, 3, 3, 1, 0, 0, 0, 1, 2, 0, 1, 1, 2, 2, 2, 3, 2, 1, -1, 2, 3, 3, 3, 2, 1, 2, 1, 2, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 2, 1, 0, -1, 3, 3, 3, 2, 1, 2, 1, 2, 3, 1, 1, 2, 3, 2, 1, 0, 1, 0, 1, 0, 0, 1, 1, 1, -1, -1, 4, 4, 3, 2, 1, 1, 2, 2, 0, 1, 1, 1, 2, 1, 0, 1, 0, 1, 1, -1, -1, 0, 0, 0, 0, -1, 2, 3, 1, 2, 0, 0, 1, 1, 0, 0, 0, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -2, 2, 1, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -2, -4, 2, 2, 0, 0, 0, -2, -3, -2, -1, -2, -2, -2, -2, -2, -3, 0, -2, -2, -1, -1, -1, -2, -1, -3, -5, -8, -3, 0, 1, 2, 3, 3, 4, 5, 7, 5, 4, 6, 6, 5, 3, 4, 3, 2, 4, 3, 4, 4, 3, 3, 2, 1, -4, -1, 1, 2, 2, 3, 2, 2, 3, 4, 4, 4, 4, 2, 2, 1, 1, 0, 1, 1, 2, 4, 2, 0, 3, 1, -3, -2, -1, 0, 1, 2, 1, 2, 2, 1, 1, 2, 2, 1, 1, 1, 0, 1, 0, 0, 0, 1, 2, 0, 0, 2, -4, -3, -2, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 1, -4, -4, -2, 0, 1, 0, 0, -1, 0, 0, -2, 0, 0, -2, -1, -2, -1, -1, 0, 0, -1, -1, -1, 0, 1, 3, -4, -4, -1, 0, -1, -2, -1, 0, -2, -1, -1, -1, -1, 0, -2, -1, -2, -1, 0, 0, 0, 0, -1, 0, 1, 1, -4, -4, -1, 0, -1, -1, -1, -1, -3, -2, -3, -2, -3, -2, -3, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -5, -3, -2, -1, -1, -2, 0, -2, -3, -2, -3, -2, -3, -3, -3, -2, -2, 0, -1, 0, 0, 0, 0, 0, 1, 2, -3, -3, -1, -1, -1, -2, -2, -3, -2, -3, -2, -3, -3, -2, -3, -3, -1, -2, 0, 0, 0, 2, 0, 1, 1, 1, -2, -1, -1, -2, -3, -1, -1, -2, -3, -2, -2, -4, -2, -3, -2, -2, -1, 0, 0, 1, 1, 2, 1, 0, 1, 1, -3, -3, -3, -2, -2, -2, -2, -3, -4, -2, -3, -3, -2, -2, -2, -2, -3, 0, 0, 1, 3, 1, 0, 1, 2, 3, -3, -2, -4, -3, -2, -4, -3, -3, -3, -3, -3, -3, -3, -2, -2, -2, -2, -1, 0, 1, 3, 2, 1, 1, 2, 4, -2, -2, -3, -4, -3, -3, -2, -2, -2, -4, -2, -2, -2, -2, -3, -2, -3, 0, 0, 1, 1, 0, 1, 0, 1, 3, -2, -2, -2, -3, -2, -3, -4, -3, -4, -2, -2, -3, -2, -2, -1, -1, -1, -2, 0, 1, 1, 0, 0, 2, 1, 3, -3, -3, -2, -2, -3, -4, -4, -4, -3, -2, -1, -2, -2, -2, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 3, 2, -3, -2, -1, -3, -2, -4, -3, -4, -2, -3, -3, -2, -2, -2, -1, 0, -1, 0, -1, 1, 1, 1, 1, 1, 3, 4, -2, -3, -2, -3, -2, -2, -2, -3, -3, -2, -2, 0, -1, -1, -2, -1, 0, -1, 0, 0, 1, 0, 0, 0, 2, 3, -3, -2, -2, -1, -2, -2, -2, -2, -3, -2, -2, -1, -1, 0, 0, -1, -2, -2, -1, -1, 1, 0, 0, 1, 1, 1, -2, -1, -2, -1, -2, -2, -1, -1, 0, 0, -2, -2, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -3, -2, -2, -1, 0, 0, 0, 0, -1, -1, 0, -2, -1, -1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 1, -5, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, -1, -2, 0, 1, -4, -2, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 1, 1, 2, 1, 0, 1, 0, 0, -2, 0, 0, -5, -3, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -5, -4, -1, 0, 1, 1, 2, 0, 1, 1, 1, 1, 0, 1, 1, 1, 0, 1, 1, 0, 1, 0, 0, 2, 0, 0, -4, -3, -2, 0, 0, 1, 1, 2, 2, 3, 3, 2, 1, 2, 2, 2, 1, 2, 1, 1, 2, 0, 2, 1, 3, 1, -4, -1, -2, 0, 3, 3, 2, 3, 4, 2, 4, 3, 3, 2, 4, 2, 2, 2, 3, 3, 2, 3, 3, 3, 1, 2,
    -- filter=0 channel=4
    -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -2, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -2, -1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, -2, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, -1, -2, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -2, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -4, -2, -3, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, -3, -2, -2, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, -1, -1, 0, -2, 0, -1, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -2, -1, -2, -2, -3, -1, -2, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -3, -4, -1, -2, -2, 0, -1, -1, 0, 0, 1, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, -2, -1, -1, -4, -2, -2, -3, -1, -2, -2, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -4, -3, -5, -4, -3, -2, -1, -1, 0, -1, -1, -1, 0, 1, 0, 0, 0, -1, 0, 1, 0, -1, -1, 0, -1, -2, -3, -3, -4, -4, -4, -1, -1, -2, -1, -2, 0, 0, 0, 0, 1, 0, 0, -2, 0, 0, 0, -1, 0, -3, -2, -3, -4, -5, -3, -3, -2, -1, -3, -2, -3, -2, -2, 0, 0, 0, 1, 1, 0, -2, -1, 0, 0, -1, -2, -3, -2, -2, -2, -3, -3, -4, -3, -3, -2, -1, -3, -2, -2, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, -3, -2, -3, -4, -2, -2, -3, -2, -2, -3, -3, -2, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -2, -2, -3, -4, -3, -3, -4, -2, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -4, -3, -4, -3, -3, -2, -1, -3, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -2, -2, -3, -2, -4, -2, -1, -2, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, -1, -3, -1, -3, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, 0, 1, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 1, 0, -1, -1, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -2, 0, 1, 1, 0, -1, -1, 0, 0, -1, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -3, -1, -1, 0, 0, -1, 0, 0, -1, 0, -1, -2, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, -1, -1, 0, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 4, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 3, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 4, 3, 1, 1, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 1, 2, 4, 2, 0, 1, -1, 0, -1, 0, -1, 0, 1, 0, 0, -1, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 4, 3, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, -1, 1, 2, 0, 1, 1, 1, 0, 0, 0, 0, 0, 2, 2, 3, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 2, 2, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 2, 3, 2, 4, 0, 0, 0, -1, -1, 0, -1, 1, 0, 0, 1, 2, 1, 0, 1, 2, 1, 0, 0, -1, 0, 2, 2, 3, 3, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 3, 0, 1, 0, 0, 1, 1, 0, 2, 2, 1, 2, 3, 0, -1, 0, 0, 1, 0, 1, 2, 2, 0, 1, 3, 3, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 3, 2, 1, 0, 0, 0, 1, 2, 2, 2, 2, 1, 1, 2, 3, 2, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 0, 0, 0, 1, 1, 1, 2, 2, 2, 2, 2, 3, 2, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 1, 1, 1, 1, 2, 3, 2, 1, 1, 3, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 3, 2, 1, 0, 1, 0, 0, 1, 1, 2, 1, 3, 2, 1, 2, 0, 0, 1, 0, -1, 0, 0, -2, 0, 0, 0, 3, 2, 1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 2, 1, 0, 0, 0, 0, -1, 0, 1, 2, 1, 1, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, -1, -1, 1, 3, 2, 0, 0, 1, 0, 0, 0, 1, 2, 1, 2, 2, 1, 3, 1, 1, 0, 0, 0, -1, 0, -1, -2, 0, 0, 1, 2, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 1, 0, 2, 1, 1, 0, -1, 0, -1, -1, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, -1, 0, 0, -1, 0, 0, 1, 1, 3, 3, 2, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, -1, -1, 0, 0, 0, 0, 1, 1, 3, 3, 2, 0, 0, -1, -1, -1, -1, 0, -1, -2, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 1, 1, 2, 3, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, 0, 0, 2, 1, 2, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 2, 2, 1, 0, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, -2, 0, -1, -1, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, -1, 0, -2, -1, -2, -1, 0, -1, 0, -1, -1, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 1, 1, 0, 1, 1, 2, 2, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 1, 0, 2, 2, 0, 1, 2, 0, 1, 1, 1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 2, 1, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -2, 0, 0, -1, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -2, -2, 0, -2, 0, -2, -1, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, -2, -1, 0, 0, -1, -1, -1, 0, -2, -1, -1, -1, 0, -1, 0, -1, -2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, 0, 0, -1, -2, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, -2, -1, -1, -1, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -2, -3, -1, -2, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, -2, 0, -1, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, -1, -1, -1, -2, -2, -3, -2, -1, 0, -1, -1, -1, -1, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -2, -2, 0, -2, -1, -3, -3, -3, -2, -1, -2, -1, -1, -2, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -2, -1, -1, -2, 0, -3, -1, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -2, 0, -2, -3, -2, -2, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, -1, 0, 0, 0, -2, 0, -1, -2, 0, -1, -3, -2, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -2, -2, 0, 0, -2, 0, -2, -2, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -3, -2, -2, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 1, 2, 2, 3, 4, 3, 0, 1, 1, 0, 2, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 3, 2, 2, 4, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 3, 4, 3, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 2, 1, 2, 2, 1, 2, 3, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 2, 1, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 2, 0, 2, 0, 2, 1, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 0, 2, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 2, 0, 0, 0, 0, -1, 0, 0, -2, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 3, 0, 0, 0, -1, -1, 0, -1, -2, -1, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 3, 1, 0, 0, -1, 0, -1, -1, -2, -2, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 2, 0, 0, 0, -1, -1, 0, 0, -1, -2, -1, -2, -1, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 2, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, 1, 1, 0, 0, 1, 0, 1, 0, 1, 0, 2, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, -2, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, -1, 0, 0, -1, -2, -1, -1, -1, -1, -1, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, -1, -2, -1, -1, -2, 0, -1, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, -2, -2, -1, -3, -2, -1, -1, -1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -2, -1, -1, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, -1, -2, -1, 0, 0, 2, 1, 1, 2, 1, 1, 0, 0, -1, -2, -1, -3, -3, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 2, 1, 1, 2, 1, 1, 0, 0, -1, -3, -3, -2, -2, -2, -1, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 1, 2, 3, 1, 2, 2, 2, 1, 0, 0, -2, -1, -3, -1, -2, 0, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, 1, 0, 3, 0, 2, 1, 0, 1, 0, 1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, 3, 0, 1, 0, 0, 1, 1, 2, 0, 1, 1, 0, 0, 0, 2, 2, 2, 2, 2, 1, 0, 1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 2, 1, 2, 1, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 2, 1, 2, 3, 3, 2, 2, 1, 2, 3, 1, 1, 0, 0, 0, 0, 0, -1, 1, 0, 2, -1, -1, 0, 0, -1, 1, 0, 0, 2, 1, 1, 1, 2, 2, 3, 5, 3, 1, 0, 2, 1, 0, 0, 0, 0, 1, -1, -1, 0, 1, 1, 1, 0, 0, 1, 3, 2, 1, 1, 3, 4, 4, 2, 4, 2, 0, 1, 2, 1, 1, 1, 3, -1, 0, 0, 2, 2, 0, 0, 0, 1, 1, 1, 2, 3, 2, 3, 3, 2, 3, 1, 3, 2, 3, 2, 1, 1, 3, -1, -1, 1, 0, 2, 2, 1, 1, 1, 0, 1, 0, 0, 0, 1, 1, 1, 2, 3, 3, 3, 0, 2, 1, 2, 3, 0, 0, 0, 0, 2, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 3, 1, 1, 1, 2, 3, 3, 0, 0, 1, 1, 1, 2, 0, 1, 2, 0, 0, 0, -1, -1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 1, 3, 5, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, -1, -1, 0, 0, 0, 1, 0, 1, 2, 2, 2, 0, 1, 2, 3, 5, 1, 1, 0, 1, 1, 0, 0, 0, 2, 0, 0, -2, -1, 0, 0, 0, 0, 0, 1, 2, 2, 0, 1, 3, 3, 7, 1, 2, 0, 0, 1, 0, 1, 0, 1, -1, -1, -2, -2, 0, -1, 0, -1, 0, 0, 0, 1, 2, 2, 4, 4, 5, 1, 2, 0, 0, 0, 1, 0, 0, -1, -2, -2, -3, -3, -3, -1, -2, -2, -2, -1, 0, 1, 1, 4, 5, 5, 6, 1, 2, 1, 0, 0, 0, 0, 0, -1, -2, -5, -4, -5, -5, -5, -5, -2, -4, -4, -2, 0, 0, 1, 2, 4, 4, 2, 0, 0, 0, 1, 1, 1, 0, -1, -3, -4, -4, -5, -6, -5, -5, -6, -4, -3, -2, -1, 0, 1, 2, 3, 6, 1, 2, 2, 2, 2, 3, 3, 3, 1, -2, -4, -5, -5, -5, -6, -6, -5, -5, -4, -3, -1, -1, 1, 2, 2, 3, 1, 1, 2, 3, 3, 4, 2, 4, 3, 0, -3, -5, -6, -4, -4, -5, -4, -3, -4, -3, -3, -2, 0, 2, 4, 3, 1, 2, 2, 2, 3, 3, 2, 2, 1, 1, -2, -2, -4, -4, -4, -3, -3, -3, -3, -1, -1, -1, 0, 1, 4, 3, 2, 2, 2, 2, 2, 1, 1, 3, 2, 0, -2, -2, -2, -2, -2, -3, 0, -2, -2, -1, -2, 0, 0, 1, 4, 3, 2, 1, 0, 0, 2, 1, 0, 1, 0, 0, -2, -2, -3, 0, 0, -1, -1, -1, 0, 0, 1, 0, 1, 3, 1, 4, 3, 0, 0, 0, 0, 0, 0, 1, 0, -2, -1, -2, -1, -1, 0, 0, 0, 0, 1, 2, 2, 2, 2, 3, 4, 3, 4, 2, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, 1, 0, 1, 0, 0, 0, 1, 0, 1, 3, 2, 4, 3, 4, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -2, 0, 0, 1, 0, 0, 0, -1, 0, 0, 2, 1, 1, 4, 5, 4, 2, 1, 0, -1, -1, -1, -2, -1, -2, 0, 0, -1, 1, 1, 1, 0, -1, -1, 0, 1, 0, 2, 3, 2, 4, 3, 4, 1, 1, 0, -1, 0, -2, -2, -3, 0, 0, 0, 1, 1, 3, 1, 1, 0, 0, 0, 1, 2, 1, 3, 3, 2, 2, 2, 0, 0, 0, 0, -2, -2, -3, -3, 0, 0, 0, 1, 3, 4, 3, 1, 1, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 1, 1, 2, 4, 3, 2, 1, 2, 1, 0, 1, 1, 1, 1, 0, -1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 2, 1, 3, 3, 3, 4, 2, 3, 1, 0, -1, 0, 0, 1, 0, 0, -1, -2, -1, -1, 0, 1, 1, 1, 1, 1, 3, 1, 1, 2, 2, 3, 1, 0, 0, 0, -2, -1, -1, 0, 0, -7, -5, -4, -3, -3, -2, -2, 0, -2, -3, -4, -2, -2, -2, -3, -2, -1, -1, 0, 0, 0, 0, -2, -3, -2, -4, -5, -4, -4, -4, -3, -2, -2, -2, -2, -3, -2, -2, -1, -2, -1, 0, 0, 0, 1, 0, 1, 0, 0, -1, -2, -3, -5, -4, -2, -2, -3, -3, -2, -3, -1, -1, -4, -2, -2, -3, -1, -2, -1, 0, 0, 0, 1, -1, -1, -2, -1, -3, -5, -4, -4, -3, -3, -2, -3, -1, -1, -2, -4, -2, -3, -2, -2, -2, 0, -1, 1, 0, 1, 0, -1, -1, -2, -3, -6, -4, -3, -2, -1, -1, -1, -1, -1, -3, -2, -2, -3, -2, -3, -2, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -5, -3, -3, -3, -3, -2, -2, -3, -3, -3, -3, -3, -3, -4, -3, -1, -2, 0, 0, 0, 1, 0, 0, 0, -1, -2, -3, -1, -1, -3, -3, -1, -2, -3, -3, -3, -3, -4, -5, -4, -4, -2, -1, 0, 0, 0, 0, 0, 0, -2, -2, -2, -3, -2, 0, -2, -2, -2, -1, -2, -3, -2, -5, -6, -6, -4, -3, -4, -1, -1, 0, 0, 1, 0, 0, 0, -1, -2, -2, -1, -2, -1, -3, -2, -3, -2, -2, -5, -5, -6, -5, -5, -4, -3, -3, -1, -1, 1, 1, 0, 0, 0, -2, -3, -2, 0, 0, -1, -1, -3, -3, -3, -3, -5, -4, -4, -4, -4, -3, -3, -4, -2, -2, -1, 0, 0, 0, 0, -1, -3, -4, -2, -2, -2, -2, -2, -4, -3, -4, -5, -5, -4, -5, -4, -3, -3, -4, -4, -2, -2, -1, -1, 0, -1, 0, -2, -5, -3, -1, -3, -2, -3, -3, -4, -3, -4, -5, -6, -4, -4, -4, -3, -3, -4, -4, -3, -2, 0, 0, 1, -1, -1, -4, -2, -1, -1, -4, -4, -4, -5, -4, -4, -6, -6, -4, -3, -4, -2, -3, -3, -4, -2, -3, 0, 0, 0, 0, 0, -4, -3, -3, -3, -4, -4, -3, -5, -6, -5, -6, -4, -5, -4, -4, -2, -3, -3, -4, -2, -1, -2, -1, 0, 0, -2, -3, -2, -1, -2, -3, -3, -4, -3, -4, -5, -4, -6, -4, -3, -2, -4, -4, -3, -4, -1, -1, -2, 0, -1, -2, -1, -3, -2, -2, -1, -2, -3, -2, -4, -5, -7, -6, -6, -4, -2, -2, -4, -2, -3, -2, -3, -2, -1, -2, -3, -2, -1, -3, -2, -2, -2, -1, -1, -1, -2, -4, -5, -6, -4, -3, -3, -3, -2, -3, -4, -4, -3, -2, -1, 0, 0, -1, -3, -3, -1, -1, -2, -1, -3, -3, -2, -3, -4, -4, -3, -4, -3, -3, -4, -4, -3, -3, -3, -1, 0, -1, -1, 0, -1, -4, -3, -2, -2, -1, 0, -2, -2, -5, -4, -4, -3, -3, -4, -2, -3, -1, -3, -2, -1, 0, 0, 0, -1, 0, -2, -3, -3, -3, -1, -1, -2, -2, -2, -2, -3, -2, -3, -4, -4, -2, -2, -2, -3, -3, -2, -2, -1, 0, 0, -1, -1, -5, -2, -3, -2, 0, -1, -1, -3, -3, -3, -2, -3, -3, -3, -3, -2, -3, -3, -4, -3, -1, 0, -1, 0, -1, -2, -4, -3, -3, -1, -2, -1, -1, -2, -3, -2, -2, -3, -2, -4, -4, -4, -3, -2, -3, -3, -1, 0, -1, 0, 0, 0, -4, -1, -3, -1, -1, -2, -3, -2, -2, -3, -3, -2, -3, -5, -4, -3, -1, -3, -1, -2, 0, 0, -1, 0, 0, -2, -4, -2, -3, -2, -2, -2, -1, -3, -2, -2, -2, -4, -4, -4, -4, -2, -2, -2, -1, -1, -1, 0, 0, -1, 0, -3, -7, -4, -3, -3, -4, -2, -2, -1, -2, -4, -4, -2, -2, -3, -2, -2, -2, -2, -1, -1, 0, 0, -1, -2, -3, -2, -7, -5, -3, -4, -3, -4, -2, -2, -3, -4, -3, -2, -4, -3, -3, -2, -2, -2, -1, 0, 0, 0, 0, -2, -4, -4, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -3, -2, -2, -1, 0, 0, -1, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, -1, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, -2, -2, -1, -1, 0, -2, 0, -1, -1, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -2, -1, -1, 0, -1, -2, -1, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -12, -10, -7, -6, -5, -2, -2, -1, -3, -2, -4, -4, -3, -3, -1, 0, 0, 0, 0, 1, 0, -1, -1, -3, -4, -5, -9, -5, -5, -3, -4, -1, -2, -2, -3, -3, -3, -4, -3, -2, -1, 0, 0, 1, 1, 2, 0, 1, -1, -2, -4, -4, -8, -5, -5, -3, -1, -2, 0, 0, -3, -4, -3, -4, -3, -2, -1, 0, 1, 0, 0, 1, 1, 1, 0, 0, -4, -4, -8, -6, -3, -4, -3, -2, -1, -2, -1, -4, -2, -2, -2, -2, -1, -1, 0, 0, 2, 0, 1, 0, 0, -1, -3, -4, -8, -4, -2, -3, -1, -2, -2, -2, 0, -3, -3, -3, -3, -4, -2, 0, 0, 1, 2, 1, 1, 1, 0, 0, -3, -3, -5, -3, -2, -1, -2, -1, -1, 0, -2, -2, -2, -3, -2, -3, -2, -2, -1, 0, 2, 1, 0, 0, 0, -2, -1, -3, -5, -2, -2, -3, -1, -2, 0, -2, -3, -4, -3, -4, -4, -3, -3, -2, -1, 0, 0, 1, 1, 1, 0, -1, -3, -2, -3, -2, -1, -2, -2, -2, -1, -1, -2, -3, -5, -4, -5, -5, -3, -1, -1, -1, -1, 1, 1, 0, 1, -1, -1, -1, -3, -1, 0, -2, -2, -2, -1, -1, -2, -5, -5, -6, -6, -5, -4, -4, -2, -1, 0, 0, 1, 2, 0, 0, -2, -2, -4, -2, 0, 0, -2, -1, -1, -1, -3, -4, -8, -7, -8, -7, -3, -4, -2, -1, -2, -1, 0, 0, 1, 0, -1, 0, -4, -3, -2, -1, -3, -2, -2, -4, -4, -6, -7, -7, -6, -7, -5, -5, -4, -4, -2, -1, -1, 0, 2, 0, -1, 0, -4, -4, -2, -2, -3, -4, -4, -5, -6, -6, -6, -7, -6, -5, -5, -4, -5, -5, -6, -2, -2, 0, 1, 0, 0, -1, -6, -3, -1, -1, -2, -4, -5, -5, -6, -7, -6, -8, -7, -5, -4, -4, -7, -6, -5, -4, -1, 0, 2, 1, 0, -1, -5, -4, -2, -3, -3, -3, -4, -6, -6, -6, -6, -5, -6, -5, -4, -5, -6, -7, -5, -4, -3, -1, 1, 0, 0, 0, -6, -3, -1, -1, -3, -3, -3, -5, -6, -6, -7, -7, -6, -4, -4, -5, -6, -6, -5, -4, -4, -2, 0, 0, -1, -1, -5, -3, -3, -3, -3, -3, -3, -4, -5, -6, -6, -7, -5, -5, -4, -3, -5, -5, -4, -3, -1, -2, -1, -1, -2, -1, -5, -4, -3, 0, -2, -1, -2, -4, -5, -6, -6, -7, -5, -4, -4, -4, -5, -4, -3, -2, 0, -1, -1, 0, -2, -2, -5, -2, -1, -2, -1, -3, -3, -3, -4, -5, -6, -5, -5, -4, -2, -3, -3, -5, -3, -2, -1, 0, 0, -1, -2, -2, -3, -3, -2, -2, -1, -2, -4, -3, -4, -5, -5, -3, -5, -4, -4, -3, -3, -3, -3, 0, 0, 1, 1, 0, 0, -2, -4, -1, -2, -1, -1, -3, -3, -2, -4, -2, -2, -3, -2, -3, -4, -3, -2, -3, -3, 0, 0, 0, 1, 0, -1, -1, -5, -3, 0, -2, -2, -1, -2, -3, -2, -1, -2, -2, -1, -3, -2, -4, -3, -1, -2, -1, 0, 0, 0, -1, 0, -3, -6, -3, -2, -1, 0, -1, -1, -1, -3, -2, -2, -3, -2, -3, -2, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, -3, -6, -4, -2, -2, -1, -1, -1, -1, -2, -2, -3, -4, -2, -4, -2, -3, -1, -2, -2, -1, 0, 0, 1, -1, -2, -3, -7, -4, -1, -2, 0, 0, -2, -2, -2, -2, -4, -2, -3, -5, -2, -3, 0, -1, -1, -1, 0, 1, 0, 0, -1, -2, -8, -6, -5, -3, -3, -3, -1, -2, -3, -3, -3, -5, -3, -4, -3, -3, -2, -1, 0, 0, 0, -1, -1, -2, -2, -4, -11, -7, -7, -6, -4, -3, -3, -4, -3, -4, -3, -4, -4, -5, -2, -2, -2, 0, -1, -1, -2, -1, -2, -2, -3, -6, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -3, -2, -3, -2, -3, -1, -2, -1, -3, -1, -3, -3, -3, 0, 1, 1, 0, 0, -1, 0, 1, 0, -1, -2, -2, -2, -3, -3, -3, -1, -1, 0, -2, -2, -1, -2, -2, -3, -3, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -2, -3, -3, -3, -3, -1, 0, 0, -1, -1, -2, -2, -4, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, -2, -2, 0, -1, -2, -2, -2, -2, -3, -3, 0, 1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, -2, 0, 0, 0, -1, 0, -2, -1, -1, -2, -4, -3, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -2, -1, 0, 0, 0, -1, -2, -2, -1, -3, 0, 0, -1, 0, -1, -2, -1, -1, 0, -1, 0, 0, -1, -1, 0, -2, -1, -2, -1, 0, -1, 0, 0, -2, -1, -1, 0, 0, 0, 0, -1, -1, -2, -2, 0, 0, -1, 0, 0, -1, -1, -2, -1, -1, -1, -1, -1, -1, 0, -2, -2, -2, 0, 0, 0, 0, -1, -1, -1, -2, -1, -2, 0, -1, 0, 0, 0, -1, -1, -2, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 1, 1, 1, -1, 0, -2, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, 1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 1, 2, 1, 2, 0, -1, 0, 1, 0, 1, 1, 0, 0, -1, 0, 1, 0, 0, 0, -1, -2, -1, -1, -2, 0, 0, 1, 2, 2, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -2, -1, -3, -2, 0, -1, 1, 0, 2, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, -2, -2, -1, -1, -2, 0, 1, 2, 2, 2, 0, 1, 1, 0, 0, 1, 0, 0, -1, 0, -1, 0, -1, 0, 0, -2, -2, -1, -1, -2, -3, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, -1, 0, 0, -1, -2, 0, -1, -1, -1, 2, 1, 1, 0, 0, -1, 0, 0, 0, -1, -1, -2, 0, -2, 0, 0, 0, -1, 0, -1, -2, -2, -1, 0, 0, 0, 1, 2, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, -1, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, -1, -1, -2, 0, -2, -1, 0, -2, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, -2, 0, -1, 0, 0, 0, -1, -1, 0, -2, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, 0, -1, -1, 0, -1, -1, -1, -1, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, -1, -2, -2, -2, -2, -1, -1, -1, 0, -1, -2, -1, -1, -2, -1, -1, 0, 0, -1, -1, 0, 0, 2, 0, 0, 0, 0, 0, -1, -2, -3, -2, -1, 0, 0, -1, -2, -2, -3, -2, -2, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, -1, 0, -2, -3, -3, -3, -2, -2, 0, -1, -2, -1, -2, -1, -2, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, -1, -2, 0, -1, -2, -2, -2, -2, -2, -2, -1, -1, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, -3, -1, -2, -2, -3, -2, -1, -1, -2, -1, -1, -1, -8, -4, -3, -1, -1, 0, 0, 1, 1, 2, 2, 1, 3, 3, 3, 2, 2, 1, 2, 1, 1, 3, 0, 1, -1, -1, -7, -4, -3, -2, -1, -1, 0, 0, 0, 1, 2, 1, 2, 2, 2, 2, 1, 2, 1, 3, 2, 2, 0, 1, 0, 0, -6, -4, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 1, 1, 1, 1, 2, 1, 2, 2, 1, 0, 0, -5, -2, -2, 0, 1, 0, 1, 1, 2, 1, 1, 0, 2, 0, 1, 1, 0, 2, 1, 1, 1, 1, 0, 0, 1, 0, -3, -1, 0, -1, 0, 1, 0, 0, 2, 1, 1, 1, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 2, 0, 1, 1, -4, -1, 0, 1, 0, 1, 0, 2, 2, 2, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 2, 2, 0, 0, 1, 1, -2, 0, 0, 1, 0, 0, 1, 1, 2, 1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 2, -2, -1, 0, 1, 1, 1, 2, 0, 1, 0, 0, -1, -1, -2, -1, -2, 0, -1, 0, 2, 1, 1, 1, 1, 1, 2, 0, -1, 1, 0, 1, 1, 2, 1, 0, 0, -2, -3, -4, -3, -4, -2, -2, -1, 0, 0, 0, 3, 3, 1, 3, 3, -1, -1, 0, 0, 1, 0, 0, 1, 0, 0, -3, -2, -5, -3, -4, -3, -2, -3, -4, 0, 0, 0, 1, 3, 3, 4, -3, -1, 0, 0, 0, 0, 1, 1, 0, -2, -3, -4, -5, -6, -6, -5, -5, -5, -5, -2, -2, 0, 2, 1, 2, 1, -1, -1, 1, 1, 2, 0, 0, 0, 0, -2, -3, -4, -6, -5, -6, -7, -5, -5, -6, -4, -2, 0, 1, 2, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, -1, -4, -4, -3, -4, -6, -4, -7, -5, -6, -5, -3, -2, -1, 0, 0, 1, -1, 0, 1, 2, 2, 1, 0, 0, -1, 0, -3, -3, -4, -4, -3, -4, -5, -5, -5, -3, -3, -2, -2, 1, 1, 1, 0, 0, 0, 1, 3, 0, 1, 1, -1, -1, -2, -3, -5, -5, -4, -3, -4, -4, -4, -4, -3, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 2, 1, 1, 0, -2, -3, -4, -5, -4, -4, -2, -4, -3, -2, -1, -1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, -1, -1, -3, -3, -4, -1, -2, -1, -1, -1, 0, 1, 1, 2, 3, 2, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -1, -1, 0, -1, -1, 0, 0, 1, 1, 1, 1, 2, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, 3, 1, 2, 3, -1, 0, 0, 0, 0, 2, 2, 2, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 2, 0, 1, -3, 0, 1, 0, 0, 0, 1, 2, 2, 0, 0, 1, 2, 0, 1, 0, 1, 1, 1, 2, 1, 0, 0, 1, 0, 1, -3, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 2, 2, 1, 0, 2, 1, 1, 1, 1, 0, -4, -2, 0, 0, -1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 3, 2, 2, 3, 1, 1, 1, 0, -6, -4, -4, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 3, 1, 1, 1, 1, 1, 0, 0, -7, -5, -2, -3, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 3, 1, 0, 1, 0, -1, 0, 0, -2, -7, -6, -5, -2, -2, -3, -1, -2, 0, -1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -2, -3, -3, -2, -1, -8, -7, -6, -4, -2, -1, -1, -1, 0, 0, 0, 1, 2, 0, 2, 2, 1, 2, 1, 1, 1, 0, 0, 0, -1, -2, -6, -5, -4, -1, -1, 0, 0, 0, 1, 1, 0, 2, 2, 3, 3, 1, 2, 1, 0, 1, 2, 2, 1, 1, -1, 0, -6, -4, -3, -3, -2, 0, 1, 0, 1, 0, 0, 2, 1, 2, 0, 1, 1, 1, 1, 1, 0, 1, 0, 0, 1, -1, -4, -4, -3, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 2, 2, 0, 1, 2, 1, 1, 1, 0, -5, -2, -1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 0, 1, 0, 0, -4, -1, -1, 0, 1, 1, 0, 1, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 1, 2, 1, 1, 1, 1, -4, -1, -1, 0, 0, 0, 1, 2, 0, 1, 2, 1, -1, -1, -1, -1, 0, 0, 0, 1, 2, 1, 0, 1, 1, 1, -3, -2, 1, 0, 2, 1, 2, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 2, 1, 2, 0, 0, 2, -1, 0, 0, 2, 2, 1, 1, 1, 1, 1, 1, -1, -2, -2, -1, -2, -2, 0, 0, 0, 1, 1, 1, 2, 0, 1, -3, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -3, -4, -3, -3, -2, -2, -1, 0, -1, 0, 2, 0, 2, 1, -2, 0, 0, 0, 0, 0, 0, 1, 0, -1, -2, -2, -3, -4, -3, -2, -2, -3, -2, -2, -2, -1, 0, 0, 1, 1, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, -5, -5, -5, -4, -3, -4, -5, -4, -3, -2, 0, 0, 1, 1, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, -2, -3, -4, -4, -5, -4, -4, -4, -5, -4, -4, -2, 0, 0, 1, 1, 2, -2, 0, 0, 1, 1, 0, 1, 1, 0, -1, -2, -3, -5, -4, -4, -5, -5, -4, -5, -5, -2, -2, -1, 0, 1, 2, -1, -1, 0, 0, 1, 1, 1, 1, 1, 0, -3, -4, -4, -5, -5, -4, -5, -5, -4, -4, -4, 0, 0, 1, 0, 1, -3, 0, 0, 0, 1, 2, 0, 1, 0, 0, -2, -2, -4, -4, -3, -3, -3, -2, -3, -3, -1, 0, 0, 1, 1, 2, -2, -2, 0, 0, 1, 2, 0, 2, 0, 0, 0, -3, -2, -2, -2, -3, -2, -2, -2, -1, -1, 0, 2, 1, 2, 1, -3, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -3, -2, -1, 0, -1, -1, -1, 0, 0, 0, 3, 2, 1, 0, -2, -1, 0, 0, 0, 1, 0, 1, 0, 1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 1, 2, 1, 1, 2, 2, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 1, 1, 3, 3, 3, 0, -2, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 3, 1, 1, -3, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 1, 2, 1, 1, 0, -3, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 2, 3, 2, 1, 1, -4, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 2, 2, 2, 2, 1, 2, 1, 0, 0, -6, -5, -4, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 1, 1, 2, 1, 0, 1, 0, 0, 0, -5, -4, -5, -2, -2, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 2, 2, 1, 0, 0, 0, -2, -1, -6, -4, -3, -2, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, -1, 0, -1, -4, -3, -1, -1, -1, -1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 1, 0, 0, -1, -4, -1, -2, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, -3, 0, -1, 0, 0, -1, 0, 0, -1, -2, 0, -1, -1, -1, -1, 0, 1, 1, 0, 1, 0, 2, 1, 0, 0, 0, -2, 0, 0, 0, 0, 0, -1, 0, -2, -1, -1, -2, -2, -1, -2, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -2, -3, -2, -3, -2, -1, -1, 0, 0, 1, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -3, -4, -3, -2, -3, -2, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 1, 0, -2, -2, -3, -3, -4, -4, -3, -4, -2, -1, 0, -1, 0, 0, 1, 1, 1, 0, 0, -1, -2, 0, 1, 1, 0, -1, -1, -2, -3, -4, -4, -3, -3, -2, -3, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, -2, -1, -2, -5, -4, -4, -3, -2, -2, -3, -1, -1, -1, 0, 0, 0, 0, 0, -1, -2, 0, 1, 0, -1, -1, -2, -1, -3, -3, -4, -6, -6, -3, -4, -4, -3, -3, -2, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -3, -2, -3, -3, -5, -4, -5, -5, -5, -4, -3, -2, -3, -3, -2, 0, 1, 0, 1, 0, -2, -2, 0, 0, 0, -3, -3, -3, -4, -3, -5, -6, -5, -4, -5, -4, -4, -3, -4, -2, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -2, -1, -2, -4, -3, -4, -7, -6, -4, -4, -3, -2, -4, -3, -2, -3, -2, -1, 0, 0, -1, -1, -2, 0, 1, 0, -1, -1, 0, -3, -4, -4, -6, -5, -6, -5, -3, -3, -2, -3, -3, -2, -1, 0, -1, -1, -1, -1, -1, 1, 0, 0, 0, 0, 0, -1, -3, -4, -6, -5, -5, -3, -4, -1, -3, -3, -1, -2, 0, 0, 0, 0, -2, -1, -1, 1, 1, 0, 1, 0, 0, -2, -4, -5, -6, -4, -4, -4, -3, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, -1, -2, 0, 1, 0, 0, 0, -1, -2, -2, -4, -4, -4, -5, -2, -2, -3, -1, 0, -1, 0, 0, 0, 1, 0, 0, -1, -2, 0, 0, 2, 1, 0, 0, -2, -2, -4, -3, -2, -2, -2, -3, -1, -1, -1, -1, -1, 1, 1, 1, 1, 0, 0, -1, -1, 0, 1, 0, 0, 0, -1, -2, -3, -2, -3, -2, -2, -2, -2, -1, -2, 0, 0, 1, 0, 2, 1, 0, -1, -3, 0, 0, 0, 1, 1, 0, -1, -1, -2, -2, -1, -2, -1, -3, -2, -2, -1, 0, -1, 0, 1, 1, 1, 0, -1, -2, 0, 0, 0, 0, 0, -1, -2, -2, -1, 0, -2, -2, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -2, -1, -1, -1, 0, 0, 1, 1, 1, 1, 2, 0, 0, 0, -4, -1, -1, 0, 0, 0, 0, -1, -2, -1, -2, -1, -1, -1, 0, 0, -1, 1, 0, 0, 0, 1, 1, 0, 0, 0, -4, -3, -2, 0, -1, -1, 0, 0, 0, -2, -1, -1, 0, -1, 0, 0, 1, 0, 1, 0, 1, 2, 0, 0, -1, -1, -7, -4, -2, -3, -2, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 1, 1, 1, 0, 0, -2, -2, -5, -4, -2, -3, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, 1, 2, 1, 2, 2, 3, 2, 2, 0, -1, -1, -1, -6, -3, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 3, 3, 1, 3, 1, 3, 1, 1, 0, 0, -4, -2, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 2, 2, 2, 1, 3, 2, 2, 1, 0, 0, 0, -3, -2, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 1, 1, 0, 0, 0, 0, -4, 0, -1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 2, 1, 2, 0, 1, 0, 0, 1, -2, -1, 0, 0, 0, 1, 1, 2, 2, 0, 0, -1, 0, 0, 0, 0, 1, 2, 3, 1, 2, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 2, 1, 1, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, 1, 0, -1, 0, -1, -1, -2, 0, 0, 0, 1, 2, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, -2, -1, -1, -2, 0, 0, -1, 0, 0, 1, 2, 2, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, -4, -2, -4, -3, -1, -2, 0, -1, 0, 0, 1, 2, 1, 2, 1, 2, -1, 0, -1, 0, 0, 0, 0, -1, -2, -3, -4, -4, -4, -2, -1, -1, -1, -1, -1, 0, 0, 2, 1, 3, 1, 1, -2, -1, -1, 0, 0, 0, -2, 0, 0, -1, -4, -3, -2, -3, 0, -1, -3, -2, -1, 0, 0, 1, 2, 2, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, -2, -1, -3, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, -1, 0, -1, 1, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 1, 1, 2, 1, -3, 0, -1, 1, 0, -1, 0, 0, -1, -1, -3, -1, 0, 0, 0, 0, -2, -1, -2, 0, 0, 0, 1, 1, 1, 1, -2, -1, 0, 0, 0, 0, 0, 0, -2, -3, -1, -2, -1, -1, 0, 0, -1, -2, -2, 0, 0, 0, 2, 0, 1, 0, -1, -1, 0, -1, 0, 0, -1, -1, -3, -3, -2, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 1, 0, -1, -2, 0, -1, -1, 0, 0, -2, -2, -2, -1, 0, -1, 0, 0, 0, 1, 1, 0, 1, 1, 3, 1, 3, 2, 2, 0, -2, 0, 0, -1, 0, 0, -1, 0, -2, -1, 0, -1, 0, 0, 2, 1, 1, 0, 0, 2, 1, 2, 4, 1, 1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 2, 2, 1, 1, 0, -1, 1, 1, 1, 2, 1, 2, 1, -2, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 1, 1, 3, 0, 1, 0, -2, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 1, 0, 3, 2, 3, 1, 1, 0, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 3, 1, 3, 3, 3, 2, 2, 1, 0, -5, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 2, 2, 2, 1, 2, 3, 1, 1, 2, 0, -1, -6, -3, -2, -2, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 1, 1, 1, 2, 0, 0, 1, -1, 0, -3, -8, -5, -2, -4, -2, -2, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 2, 1, 0, 1, -1, -1, -1, -1, -3, -3, -1, -1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 2, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 2, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 1, 0, 1, 1, 1, 1, 2, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 2, 0, 0, 1, 1, 0, 0, 1, 0, -1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 2, 1, 2, 2, 1, 1, 0, 0, -1, 0, 1, 0, 1, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 0, 1, 2, 1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 1, 0, 1, 0, 2, 1, 0, 0, 0, 0, 2, 1, 2, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 2, 1, 0, 1, 1, 1, 3, 1, 2, 0, 1, 0, 0, 0, -2, -1, -2, 0, 0, 0, -1, -1, -1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, -2, -1, -2, -1, -2, -1, -1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, -1, -2, -3, -2, -3, -2, -2, 0, 0, -1, 0, -1, 1, 1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, -2, -3, -2, -1, -2, -2, -1, 0, -2, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, -2, -2, -2, -4, -2, -1, -1, -2, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, -2, -3, -3, -3, -2, -1, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 3, 2, 0, 0, 0, -1, -2, -1, -1, -3, -2, -1, -1, -2, -1, -1, 0, 1, 0, 0, 0, 0, -1, -1, 1, 0, 2, 2, 1, 1, 0, 0, 0, -1, -2, -2, -1, -2, -1, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 1, 3, 1, 2, 1, 1, 0, -1, -1, -1, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 2, 2, 2, 2, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 1, 0, 1, 1, 0, 2, 0, 0, 1, 0, 0, 2, 1, 3, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 0, 1, 0, 0, 2, 3, 3, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 2, 2, 3, 1, 2, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 2, 1, 0, 0, 1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 2, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 2, 0, 1, 1, 2, 1, 2, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -7, -4, -2, -3, -1, -2, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 2, 1, 2, 2, 1, 0, 0, 0, 0, -2, -5, -4, -2, -2, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 2, 1, 3, 2, 1, 1, 0, 2, 1, -1, 0, -5, -3, -2, 0, -1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 1, 2, 2, 3, 2, 1, 2, 0, 1, -1, -1, -5, -4, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 0, 0, 2, 2, 1, 0, 1, -1, 0, -4, -2, 0, 0, 0, 1, 1, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -3, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, -1, -3, 0, 2, 2, 1, 1, 0, 2, 1, 0, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -2, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -3, -3, -3, 0, -1, 0, 0, 0, 0, 1, 2, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, -3, -3, -3, -1, -1, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, -2, -1, 1, 0, 0, 1, 0, 0, 0, -1, -2, -3, -3, -3, -2, -1, 0, -1, 0, -1, 0, 1, 1, 1, 2, 2, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, -2, -3, -4, -4, -2, -2, -2, -2, -3, -1, -1, 0, 0, 1, 2, 1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -3, -4, -4, -2, -3, -2, -3, -2, -2, 0, 0, 1, 2, 2, 2, -2, -1, 0, 0, 0, 0, 0, -1, 0, -2, -1, -2, -2, -2, -1, -2, -3, -2, -3, -3, -2, -1, 1, 1, 1, 0, -2, -2, 0, 1, 0, 0, 1, -1, -2, -3, -1, -2, -2, -1, -2, -3, -3, -3, -4, -3, 0, -1, 0, 1, 1, 1, -1, -1, 0, 1, 0, 0, 0, -1, 0, -2, -2, -3, -3, -2, -2, -3, -3, -4, -2, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, -1, 0, -2, -2, -2, -3, -1, 0, 0, -1, -2, -2, 0, 0, 2, 2, 1, 1, 0, -2, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, -1, -2, -1, -1, -1, 0, -1, 0, 0, 1, 3, 2, 0, 1, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 3, 1, 1, 1, 1, -3, -1, 1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 2, 1, 0, -4, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 1, -3, -1, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, -3, -1, -1, 0, 0, 0, 0, 0, 2, 0, 1, 1, 1, 1, 0, 1, 0, 2, 1, 1, 0, 1, 2, 2, 0, -1, -5, -3, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 2, 1, 2, 1, 1, 0, 0, -6, -4, -1, -2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 2, 2, 2, 2, 2, 0, -1, -1, -8, -4, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -2, -1, -8, -5, -5, -2, -1, -1, -2, -1, -2, -1, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, -1, -2, -4, -3, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, -1, 1, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, -1, -1, 1, 1, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, -1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 1, -1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 2, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 2, 0, 2, 2, 1, 0, -1, -1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -2, -2, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 1, 2, 0, 0, 1, 1, 0, 0, -1, 0, -1, -2, -2, -2, -3, -1, -1, 0, 0, 0, -1, 0, 1, 0, 2, 2, 2, 2, 3, 2, 0, 0, 1, 0, 0, 0, 0, -2, -3, -1, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 2, 0, 2, 1, 2, 1, 1, 0, 0, 1, -1, 0, 0, -2, -1, -3, -2, -1, -2, 0, -1, 1, 0, 1, 2, 1, 2, 0, 3, 1, 3, 0, 2, 0, 1, 0, -1, 0, -2, -2, -3, -1, -2, 0, -1, -1, 0, 0, 2, 1, 1, 1, 1, 2, 1, 1, 3, 2, 1, 0, 0, 0, -1, 0, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 1, 3, 1, 2, 0, 2, 1, 2, 2, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 2, 1, 1, 3, 2, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 2, 1, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 2, 1, 2, 2, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, -2, 0, 0, 0, 1, 0, 2, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 2, 2, 2, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, -3, -2, -1, -2, -3, -3, -1, 0, 0, 0, -3, -4, -3, -2, -3, -1, -2, 0, -1, -1, 0, -1, 0, 0, 0, -1, -4, -3, -1, -3, -2, -3, -1, -1, 0, -2, -3, -4, -3, -3, -1, -3, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, -4, -4, -3, -2, -3, -3, -1, -2, 0, -2, -3, -1, -1, -2, -2, -2, 0, 0, 1, 1, 0, 2, 1, 2, 0, 0, -4, -2, -2, -1, -1, -1, -2, -1, -2, -2, -1, -2, -2, -1, -1, -1, 0, 1, 0, 0, 2, 2, 1, 1, 2, 0, -3, -2, -1, -1, -2, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 2, 1, 2, 1, 1, 0, -3, -3, -2, -2, -3, -3, -1, -2, -1, 0, 0, 1, 0, 0, -2, -2, 0, 0, -1, -1, 1, 2, 1, 0, 0, 0, -3, -2, -2, -3, -2, -3, -2, -1, -1, 0, 0, 0, -1, 0, 0, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -3, -4, -2, -1, -2, -2, -2, -2, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 1, 0, -1, -1, 0, -4, -3, -3, -1, -1, -2, -2, -1, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -4, -2, -2, -1, 0, -2, -1, -2, 0, 0, 0, 1, 2, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -2, -2, -2, -2, -2, -4, -2, -3, -1, 1, 2, 2, 2, 0, 2, 0, 2, 2, 2, 2, 2, 0, 0, 0, 0, 1, -1, -3, -3, -2, -4, -4, -6, -3, -2, 0, 1, 2, 0, 0, 1, 0, 1, 2, 2, 3, 1, 0, 1, 1, 0, 0, -3, -1, 0, -4, -5, -5, -5, -5, -1, 0, 2, 1, 0, 1, 1, 0, 1, 2, 3, 1, 0, 0, 0, 0, 0, 0, -1, 0, -3, -2, -3, -4, -5, -4, -1, 1, 2, 3, 1, 1, 0, 0, 2, 1, 1, 0, 1, 0, 0, 0, -2, -1, -2, -2, -2, -3, -3, -3, -4, -2, 0, 1, 1, 3, 2, 1, 2, 0, 0, 1, 1, 0, 0, 0, -1, -2, 0, 0, -2, 0, -1, -1, -3, -3, -3, 0, 0, 1, 3, 2, 1, 0, 0, 0, 1, 2, 2, 0, -1, 0, -1, 0, -1, 0, -1, -1, -1, -2, -2, 0, 0, 0, 2, 2, 1, 2, 1, -1, -2, -1, 0, 0, 0, 0, 0, -2, -2, -1, 0, -2, -2, -1, -2, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, -2, -1, 1, 1, 1, 0, -1, -1, -2, -1, -2, -1, -2, -1, -1, 0, -1, 1, 1, 0, 0, 1, 0, 0, -1, -1, 0, 0, 2, 1, 0, 0, -1, -1, -3, -1, -1, -2, 0, -2, -1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -3, -1, -1, 0, 0, 0, 0, 0, -1, -3, -3, -3, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -2, 0, 0, 0, 1, 0, -2, -1, -2, -2, -4, -2, -1, -1, -2, -1, -1, 1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 2, 0, -1, -1, -2, -4, -5, -4, -2, -2, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -2, -1, 0, 0, 1, 0, 0, -2, -1, -2, -2, -3, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, -2, -1, -3, -2, -2, -1, -1, -2, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -2, -3, -1, -1, -3, -2, -3, -3, -2, -2, -1, 0, -1, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, -2, -2, -1, -2, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -8, -6, -4, -4, -1, 0, 0, 1, 1, 1, 1, 3, 2, 3, 3, 3, 3, 3, 1, 2, 0, 0, 0, -1, -1, -1, -7, -5, -3, -3, -1, 0, 0, 0, 0, 2, 1, 3, 2, 2, 3, 2, 3, 3, 1, 1, 1, 1, 1, 0, 0, -1, -6, -3, -3, -1, 0, 0, 0, 1, 0, 0, 1, 1, 3, 1, 1, 3, 2, 2, 2, 2, 2, 1, 0, 0, 0, 0, -6, -3, -2, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 2, 2, 1, 1, 2, 1, 3, 1, 2, 2, 0, 0, 0, -5, -2, 0, -1, 0, 1, 1, 0, 2, 0, 2, 1, 0, 0, 0, 1, 1, 1, 1, 2, 1, 2, 1, 1, 1, 1, -4, -2, 0, 0, 0, 0, 0, 2, 1, 3, 2, 0, 0, 0, 0, 0, 0, 0, 1, 2, 4, 3, 3, 2, 2, 2, -2, 0, 0, 1, 1, 1, 0, 2, 1, 2, 2, 0, 0, -1, 0, -1, -1, 1, 1, 2, 3, 2, 2, 2, 3, 1, -3, -1, 0, 0, 1, 1, 0, 0, 2, 1, 1, 0, -1, 0, -1, -1, 0, 0, 1, 2, 3, 4, 3, 1, 1, 2, -2, 0, 0, 2, 1, 2, 1, 1, 0, 1, 0, -2, -1, -2, -3, -1, -1, 0, 0, 1, 3, 3, 3, 3, 2, 3, -1, 0, 0, 2, 2, 1, 2, 1, 1, 0, -1, -4, -5, -5, -3, -4, -2, -4, -2, 0, 1, 0, 1, 1, 2, 3, -1, 0, 1, 0, 1, 1, 0, 0, -1, 0, -2, -4, -5, -6, -5, -6, -4, -4, -3, -4, -1, 0, 2, 1, 3, 0, -2, 0, 0, 1, 1, 1, 0, 0, 0, -3, -5, -5, -5, -7, -6, -5, -7, -5, -6, -4, -4, 0, 0, 1, 2, 0, 0, 0, 1, 2, 2, 1, 1, 1, 0, -2, -3, -5, -7, -7, -7, -6, -6, -7, -5, -6, -2, -2, 0, 0, 2, 1, 0, 0, 2, 1, 2, 2, 1, 1, 0, -2, -5, -6, -8, -8, -8, -7, -7, -8, -5, -5, -2, -1, 0, 0, 0, 1, -1, 1, 1, 2, 2, 2, 2, 2, 0, -2, -3, -4, -6, -6, -6, -6, -5, -5, -6, -4, -3, -2, -1, 0, 1, 0, 0, 1, 1, 2, 2, 3, 1, 2, 0, -2, -2, -4, -5, -5, -5, -5, -4, -3, -4, -3, -3, -1, 0, 2, 2, 2, -1, 0, 0, 3, 2, 3, 1, 1, 0, -1, -1, -3, -5, -4, -4, -2, -2, -2, -3, 0, 0, 0, 1, 2, 3, 2, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, -2, -1, -2, -2, -1, 0, -1, 0, 0, 0, 1, 0, 3, 3, 2, 1, -2, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, -1, 1, 0, 1, 2, 2, 3, 1, -2, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 2, 2, 1, 3, -2, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 2, -3, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 1, 1, 1, 1, 0, 2, 2, 0, 2, 0, 0, -3, 0, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 3, 2, 2, 2, 3, 1, 1, 2, 0, 0, -3, -2, -3, 0, -1, 0, 1, 0, 1, 0, 1, 0, 1, 1, 2, 0, 2, 3, 3, 3, 3, 2, 1, 1, 0, 0, -6, -4, -3, -3, -1, -1, 0, 1, 0, 1, 0, 0, 1, 0, 1, 1, 3, 2, 3, 1, 1, 1, 1, 1, 0, 0, -6, -5, -3, -2, -1, 0, 0, 0, 2, 0, 1, 0, 0, 2, 2, 3, 3, 3, 2, 1, 1, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -2, -2, -1, 0, -1, -1, 1, 0, 0, 0, 1, 1, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, -2, 0, -2, -2, 0, -2, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -2, -1, -1, 0, -1, -2, -2, -1, -1, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, -1, -2, -1, 0, -1, -1, 0, 0, 0, 0, -1, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -2, -2, -1, 0, 0, -1, -1, 0, -1, -1, 0, -1, -1, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, -2, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, -2, 0, 0, -1, -2, 0, 0, -2, -1, 0, 0, -2, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, -2, -1, -2, -2, -2, -1, 0, -2, 0, -1, 0, 0, 0, 0, -1, 0, -1, -2, 0, -1, -1, -1, 1, 0, 0, 0, -2, -2, -2, -1, 0, -1, -1, -2, -2, -2, -2, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -2, -3, -1, -3, -2, 0, -2, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -3, -2, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, 0, -2, -1, -1, -2, -2, -2, -2, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, -2, 0, -2, 0, -1, -2, -2, -1, -3, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -2, -3, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -2, 0, 0, -2, -3, -2, -1, -1, -2, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -3, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, -1, -1, -1, 0, 0, -1, 1, 0, -1, -1, -2, 0, 0, -2, -1, -2, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, -2, -1, -1, -1, 0, 0, 0, 1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, -1, 0, -2, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -7, -6, -2, -1, -1, 0, 1, 2, 2, 2, 3, 2, 4, 5, 4, 6, 6, 5, 3, 3, 2, 3, 2, 2, 1, 1, -6, -5, -3, 0, 1, 2, 1, 1, 3, 3, 3, 5, 5, 4, 3, 5, 4, 5, 4, 2, 2, 3, 3, 3, 1, 0, -5, -4, -2, 0, 1, 0, 2, 1, 2, 3, 3, 2, 2, 3, 4, 2, 3, 3, 3, 3, 4, 3, 2, 2, 1, 0, -5, -2, 0, 1, 1, 2, 2, 1, 2, 4, 3, 2, 2, 1, 2, 2, 1, 1, 1, 2, 2, 2, 1, 1, 2, 0, -3, 0, 0, 1, 2, 2, 3, 2, 3, 4, 4, 2, 0, 1, 0, 0, 1, 1, 2, 3, 1, 2, 0, 1, 1, 0, -1, 0, 2, 1, 1, 1, 3, 4, 4, 3, 3, 2, 0, 0, 0, 0, 2, 3, 2, 3, 2, 2, 1, 1, 1, 1, -3, 0, 1, 1, 2, 1, 2, 2, 3, 1, 2, 0, 0, 0, 0, 0, 0, 2, 3, 3, 2, 2, 2, 1, 4, 4, 0, 0, 1, 2, 3, 3, 1, 1, 2, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 2, 3, 2, 3, 4, 4, 5, 0, 0, 1, 1, 2, 1, 2, 1, 0, 0, 0, -4, -4, -4, -3, -2, 0, 0, 0, 1, 3, 3, 4, 6, 4, 5, -1, 1, 0, 0, 0, 0, 1, 0, -1, -1, -4, -4, -7, -5, -4, -4, -3, -1, -2, -2, 0, 3, 3, 6, 5, 5, 0, 1, 0, 2, 2, 1, 0, 1, 0, -2, -3, -5, -6, -6, -6, -5, -5, -4, -5, -2, 0, 2, 3, 3, 5, 4, 1, 1, 0, 1, 1, 3, 3, 2, 1, 0, -3, -4, -5, -6, -5, -5, -4, -4, -5, -4, -2, 0, 1, 2, 4, 3, 0, 0, 2, 4, 4, 5, 4, 2, 2, 0, -3, -4, -6, -6, -6, -5, -4, -4, -4, -3, -3, -2, 0, 2, 2, 3, 0, 1, 2, 3, 4, 3, 3, 3, 1, 0, -3, -4, -5, -5, -3, -4, -3, -3, -5, -4, -2, 0, 0, 2, 3, 3, 0, 0, 1, 3, 3, 3, 2, 1, 0, -1, -2, -4, -5, -3, -4, -3, -2, -3, -5, -3, -1, 0, 0, 2, 2, 2, 0, 1, 0, 1, 1, 2, 0, 0, 1, 0, -2, -2, -3, -3, -2, 0, 0, -1, -1, 0, 0, 1, 2, 2, 2, 3, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, -3, -1, -1, 0, 0, 0, 0, 0, 1, 0, 3, 3, 4, 3, 2, 0, 1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 1, 1, 2, 2, 1, 1, 1, 3, 4, 3, 3, 5, 1, 0, 0, 1, 0, -1, 0, 1, 2, 2, 2, 2, 1, 1, 1, 2, 2, 1, 0, 0, 0, 2, 3, 5, 5, 5, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 2, 2, 2, 2, 0, 0, 0, 0, 2, 2, 3, 4, 4, -1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 2, 2, 3, 4, 4, 1, 2, 1, 2, 2, 4, 4, 3, 4, -1, 0, 0, 0, 0, 1, 0, 2, 0, -1, 0, 1, 1, 3, 2, 3, 3, 3, 3, 3, 4, 3, 3, 3, 3, 1, -3, -3, 0, 0, 0, 2, 2, 2, 0, 0, 0, 0, 1, 2, 1, 3, 3, 4, 4, 3, 3, 3, 3, 3, 3, 0, -5, -5, -2, -2, 0, 1, 0, 0, 0, 0, 1, 0, 0, 3, 1, 2, 3, 4, 5, 4, 1, 2, 1, 0, 1, 0, -7, -5, -4, -3, -2, 0, 0, 2, 0, 0, 0, 2, 2, 1, 3, 3, 2, 4, 2, 3, 0, 0, -1, 0, -2, -2, -8, -5, -6, -3, -2, -2, -1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 2, 0, -1, -3, -5, -4, -5, -2, -2, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 3, 2, 1, 1, 1, 2, 1, 0, 1, 2, 3, 3, 4, 6, 6, 4, 2, 0, 0, 0, 0, 0, -2, -1, -1, 0, 3, 1, 1, 0, 0, 0, 0, 0, 2, 2, 2, 3, 3, 4, 5, 3, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, 3, 0, 1, 1, 0, -1, -1, -1, 1, 2, 2, 1, 1, 2, 3, 1, 2, 0, 0, 0, 0, -1, -2, -1, -1, 0, 3, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 2, 0, 2, 1, 0, 0, 0, -2, -1, -1, 0, 0, 2, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, -1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 1, 0, 1, 2, 0, 0, 0, 2, 1, -1, 0, 0, 0, -1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 1, 2, 2, 0, 0, -1, -1, 0, 0, 0, 2, 1, 1, 3, 2, 1, 0, -1, 0, 0, -1, -2, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, -1, 0, 1, 2, 3, 2, 3, 3, 0, 1, 0, 0, 0, 0, -1, -2, 0, 0, 2, 3, 1, 1, -2, -2, -3, -2, -2, 0, 1, 2, 2, 1, 2, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 0, -1, -1, -2, -2, -2, -2, -1, 0, -1, 1, 1, 0, 2, 3, 2, 0, 1, 3, 1, 0, 1, 0, 0, 1, 0, 0, -1, -1, -2, -1, -2, -1, -1, -1, 0, -1, 0, 0, 0, 1, 1, 2, 4, 3, 3, 2, 3, 0, 1, 0, 0, -1, -2, -3, -3, -3, -2, -2, -4, -2, -3, -3, -1, 0, 0, 3, 2, 3, 3, 4, 4, 4, 3, 1, 0, 0, -2, -1, -4, -3, -3, -2, -3, -3, -4, -3, -4, -4, -2, 0, 0, 4, 4, 5, 5, 3, 2, 4, 4, 3, 0, 0, -1, -3, -5, -4, -2, -1, -3, -4, -3, -4, -2, -3, -1, 0, 1, 3, 2, 3, 3, 3, 1, 3, 4, 3, 1, -1, -1, -2, -4, -4, -1, -1, -1, -2, -1, -1, -3, -2, 0, 0, 0, 3, 2, 3, 3, 3, 2, 3, 3, 3, 1, 0, -1, -1, -3, -2, -2, -1, -1, -2, 0, 0, -1, 0, 0, 0, 0, 2, 2, 1, 1, 2, 1, 3, 3, 3, 2, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 2, 3, 1, 0, 0, 0, 2, 2, 3, 4, 5, 2, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 2, 3, 0, 0, -1, 1, 1, 0, 2, 3, 4, 3, 1, 2, 1, 0, 0, -2, 0, 0, 0, 0, 0, -1, 0, 1, 2, 2, 2, 0, -1, 0, 0, 0, 1, 1, 1, 2, 3, 2, 2, 1, 1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 2, 1, 1, 0, -1, 0, -1, 0, 1, 2, 1, 2, 0, 0, 0, 1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 2, 2, 1, 2, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 4, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 3, 0, 0, 0, 0, -1, 0, 1, 1, 1, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, -1, -2, -2, 0, 0, 0, 2, 1, 0, -1, -1, -1, 0, 1, 0, 2, 2, 3, 1, 1, 2, 1, 0, 0, 1, 0, -1, -1, -1, 0, 0, 1, 3, 1, 0, 0, -1, 0, 2, 1, 2, 2, 3, 2, 3, 2, 0, 1, 0, 0, 0, 0, -2, -1, -2, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, -1, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, -2, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, -1, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, 1, -4, -3, -1, 0, -2, 0, -1, 1, 0, 1, 4, 5, 5, 5, 5, 5, 4, 3, 1, 0, -1, -1, -2, -3, -2, -1, -3, -3, -1, -2, -1, -1, -1, 0, 0, 2, 3, 4, 4, 4, 4, 5, 4, 1, 0, 1, -1, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 3, 2, 4, 4, 4, 2, 2, 2, 0, 0, 0, -1, 0, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 3, 3, 3, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 2, 2, 1, 1, 0, 1, 1, 1, 2, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 2, 1, 4, 3, 1, 1, 3, 0, 1, 0, -1, 0, 2, 1, 1, 0, 1, 1, 0, 2, 3, 2, 1, 0, 0, 0, 0, 2, 1, 4, 4, 2, 3, 3, 3, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 3, 3, 1, 0, -1, -1, 0, 0, 0, 2, 3, 3, 4, 5, 3, 1, 1, 1, 0, 2, 2, 0, 0, -1, 0, 1, 1, 0, 0, 0, -1, -3, -2, -1, 0, 0, 1, 3, 3, 2, 1, 2, 0, 0, 1, 2, 2, 2, 1, 0, 0, 1, 1, -1, -2, -3, -2, -3, -3, -2, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 2, 2, 2, 0, 0, 0, 0, -1, -2, -3, -3, -3, -3, -1, -2, -3, -1, -1, 0, 0, 0, -1, 0, 1, 1, 2, 4, 2, 2, 2, 0, -1, -1, -4, -3, -5, -6, -4, -4, -2, -3, -3, -2, -1, -3, 0, -1, -1, 1, 3, 2, 4, 3, 3, 2, 4, 1, -1, -2, -3, -6, -5, -5, -6, -4, -2, -3, -3, -3, -2, -1, -1, -2, 0, 1, 1, 3, 2, 3, 4, 3, 3, 2, 1, -3, -5, -5, -7, -6, -4, -4, -3, -3, -4, -3, -2, -2, -1, -1, 0, 2, 2, 3, 3, 4, 2, 2, 2, 1, 1, -1, -2, -4, -5, -4, -3, -3, -2, -4, -4, -4, -2, -2, 0, 0, 0, 1, 1, 3, 2, 3, 4, 3, 3, 2, 0, 0, -1, -3, -5, -4, -3, -2, -1, -2, -2, 0, -1, 0, 0, 0, 2, 1, 0, 2, 2, 4, 3, 4, 3, 3, 1, 0, -1, -1, -2, -1, -2, 0, -1, -2, 0, 0, 0, 0, 2, 2, 2, 0, 1, 0, 1, 1, 2, 4, 4, 3, 1, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 1, 0, 2, 2, 4, 2, 3, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 1, 0, 0, 0, 0, 1, 0, 1, 3, 2, 2, 3, 3, 2, 0, 1, 0, 0, 1, 0, 0, 2, 1, 2, 3, 1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 2, 1, 3, 1, 1, 0, 2, 2, 0, 0, 1, 0, 0, 2, 0, 1, 0, 0, 0, 0, 1, 1, 1, 2, 2, 0, 0, 2, 1, 2, 2, 2, 1, 2, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 3, 2, 2, 3, 3, 2, 0, 1, 1, 0, 0, 0, 0, -1, -2, -2, -1, 1, 2, 2, 1, 1, 2, 1, 3, 1, 2, 2, 3, 3, 2, 1, 0, 0, 0, 1, 0, -1, 0, 0, -3, -2, -1, 0, 1, 1, 1, 2, 2, 2, 3, 4, 3, 2, 2, 3, 1, 1, 1, -1, 0, 0, 0, 0, 0, -1, -3, -2, -1, 0, 0, 2, 3, 4, 4, 4, 3, 4, 3, 4, 5, 2, 1, 0, -2, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 1, 1, 0, 0, 1, 0, 1, 0, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, -7, -3, -3, -1, 0, 1, 1, 1, 2, 3, 1, 3, 2, 2, 3, 3, 3, 3, 3, 2, 2, 1, 1, 0, -2, -2, -5, -3, 0, -1, 0, 1, 2, 1, 2, 1, 2, 2, 2, 1, 1, 2, 3, 3, 4, 2, 2, 2, 2, 2, 0, 0, -5, -3, 0, 0, 1, 2, 1, 1, 2, 1, 2, 2, 1, 1, 2, 2, 2, 2, 2, 3, 2, 1, 1, 1, 0, 0, -4, -2, -1, 1, 0, 1, 2, 2, 1, 2, 1, 2, 1, 1, 2, 1, 2, 3, 2, 2, 2, 2, 2, 1, 0, 0, -3, 0, 0, 0, 1, 2, 1, 2, 3, 2, 2, 1, 0, 0, 0, 1, 0, 3, 3, 2, 2, 0, 1, 1, 0, 0, -1, 0, 2, 1, 2, 2, 2, 4, 4, 3, 0, 0, 0, 0, 0, 0, 2, 2, 3, 2, 3, 1, -1, 0, 0, 0, 0, 0, 2, 2, 0, 2, 1, 3, 2, 1, 0, 0, -1, 0, 0, 0, 0, 3, 3, 3, 2, 1, 0, 0, 0, 0, 0, 1, 3, 1, 1, 2, 0, 0, 1, 0, 0, -3, -2, -2, 0, 0, 1, 3, 2, 4, 2, 2, 0, 0, 2, 1, 1, 2, 2, 2, 1, 1, 0, 0, 0, -1, -3, -4, -3, -4, -2, -1, 0, 0, 1, 3, 2, 2, 1, 1, 2, 3, 0, 3, 2, 2, 0, 0, 0, 0, 0, -2, -7, -6, -6, -4, -2, -1, -1, -1, 0, 0, 2, 2, 2, 2, 2, 2, 0, 1, 1, 1, 1, 1, 0, 0, -2, -4, -7, -7, -5, -5, -4, -2, -2, -2, -1, 0, 1, 1, 4, 4, 4, 4, 0, 2, 1, 0, 2, 1, 1, 0, -1, -3, -5, -6, -6, -3, -4, -4, -3, -3, -3, -1, 0, 2, 2, 2, 3, 4, 0, 0, 1, 2, 3, 1, 2, 0, -1, -3, -5, -4, -4, -3, -3, -3, -4, -4, -4, -2, 1, 2, 2, 1, 1, 3, 0, 0, 2, 1, 2, 2, 0, -1, -1, -1, -2, -3, -2, -2, -1, -1, -2, -3, -3, -1, 0, 0, 0, 3, 1, 1, 0, 0, 1, 3, 2, 2, 0, 0, -3, -3, -4, -3, -2, -1, 0, 0, -2, -1, -2, 0, 1, 0, 0, 0, 1, 0, 0, 1, 2, 2, 2, 1, -1, 0, -2, -3, -4, -3, -1, 0, 0, 0, -1, -1, 0, 1, 1, 3, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -3, -4, -2, -2, 1, 0, 0, 1, 0, 0, 1, 4, 2, 3, 1, 1, 0, 0, 1, 0, 0, -1, -2, -2, 0, -2, -2, -3, -2, -1, 0, 1, 2, 1, 2, 1, 1, 4, 4, 2, 2, 1, 2, 1, 1, 0, 0, 0, -1, -2, -2, 0, -1, -2, 0, 0, 1, 3, 3, 1, 0, 0, 1, 4, 3, 4, 2, 3, 3, 0, 2, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 2, 2, 3, 2, 2, 1, 2, 0, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 3, 3, 1, 1, 2, 4, 2, 2, 3, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 0, 1, 1, 0, 1, 2, 3, 2, 1, 2, 3, 3, 3, 3, 2, 1, 0, -3, 0, 0, 0, 0, 1, 1, 2, 2, 1, 1, 1, 0, 1, 3, 2, 4, 3, 4, 4, 3, 3, 4, 1, 0, 0, -3, -1, -1, 0, 2, 0, 1, 2, 0, 0, 0, 0, 0, 0, 1, 2, 4, 3, 3, 4, 4, 3, 1, 1, 0, -2, -6, -4, -1, 0, 0, 0, 0, 1, 1, 1, 0, 2, 0, 2, 1, 2, 2, 3, 1, 1, 2, 1, 0, -1, -1, -1, -7, -4, -3, -2, -2, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 2, 0, 2, 0, -1, 0, -2, -3, -4, -4, -3, -1, 0, 0, 0, -1, -1, -2, 0, -1, -1, -1, -2, -2, -1, -2, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, -2, -1, 0, 0, 0, 0, -1, -2, -2, -1, 0, -1, 0, -2, -1, 0, 0, -1, 0, 0, 0, 0, -1, -2, -2, -2, -2, 0, -1, -1, 0, 0, 0, -2, 0, -2, -1, 0, -1, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, -2, 0, -2, 0, 0, -1, -1, 0, -1, -1, -1, -1, -2, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, -1, -2, -2, 0, -1, -1, 0, -2, 0, -2, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -2, -1, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, -2, -2, -1, -1, -1, 0, 0, 0, 1, 0, -1, 0, 0, -2, 0, -2, -1, 0, -1, 0, 0, 0, -1, -1, -1, -2, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -2, -2, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, -1, -2, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -1, -1, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -2, -3, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, -1, -2, 0, 0, -2, -2, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -1, -1, -3, -2, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, -2, -2, -1, -1, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -2, 0, -1, 0, -2, -2, -1, -2, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, -2, -1, -2, -1, -2, -1, 0, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, -2, -2, -2, -1, -1, 0, 1, 1, 1, 0, 0, -1, -1, 0, -1, -1, -1, 0, -1, -2, 0, 0, -1, -1, 0, 0, -1, 0, -2, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -2, -1, 0, 0, -2, -1, 0, 0, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, -2, -1, -1, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, -2, 0, 0, -1, 1, 1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, 0, 0, 0, 0, -1, 0, -2, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, -2, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, -1, -2, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -2, -2, -3, -2, -2, -2, -2, -1, 0, 0, -1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -2, -1, -2, -1, -1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 1, 0, 1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -2, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 2, 2, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, -1, 0, -1, -1, 0, -2, -1, -3, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -2, -3, -2, -2, -3, 0, 0, 0, 0, 1, 2, 1, 1, 0, 2, 1, 0, 1, 0, 0, 0, 1, 0, -1, -1, -1, -1, -3, -2, -1, -1, -1, 0, 0, 0, 2, 2, 1, 2, 2, 1, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -2, 0, -2, -3, 0, -1, 0, 0, 1, 2, 1, 2, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -2, -2, 0, 0, 0, 1, 1, 2, 2, 0, 1, 1, 0, 0, 1, 0, 0, -1, 0, 1, -1, 0, 0, -1, 0, 0, -2, -2, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, -2, -1, 0, -2, -1, -2, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, -2, 0, 0, -1, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 1, -1, 0, 1, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, -1, -2, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, -1, 0, -1, 0, -1, -1, -2, -2, 0, -2, -1, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, -2, -1, 0, -2, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, -1, 1, 0, 1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, -1, 0, -1, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, -2, -2, -1, -2, -1, 0, 0, -2, -2, -2, -2, -2, -1, -3, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, -2, -2, 0, 0, -2, -1, 0, -1, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, -2, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, -1, 0, -1, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, -1, -2, 0, -1, -2, -2, 0, 0, 0, -1, 0, -2, 0, 1, 0, 0, 0, 0, -2, -1, -2, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, 0, -1, 0, 0, -2, -2, 0, 1, 0, 0, 0, -1, -2, 0, -2, -2, -1, 0, 0, -1, 0, 0, 0, 0, -1, -2, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -2, -1, -1, -1, -1, -2, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -2, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 2, 2, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, 0, 0, 0, 1, 0, 1, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, -1, 0, 0, 1, 0, -1, 0, -2, -2, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, -1, 0, -1, -2, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -2, 0, -1, -2, -1, -1, -2, 0, 0, 0, 0, 1, 0, -1, 0, 1, 1, 1, 0, 0, -1, 0, -1, -1, -1, -3, -2, -2, -2, 0, -1, -2, -1, 0, -1, -2, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -2, -1, -2, -1, -2, -2, -1, -1, -1, -2, -2, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -2, -2, -1, -1, -2, -2, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -2, -3, -2, -3, -3, -1, -2, -3, -2, -1, -2, -2, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, -1, -2, -2, -1, -2, -1, -2, -1, -1, -1, -1, -2, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, -2, -1, -3, -2, -2, -3, 0, -1, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -2, -3, -3, -1, -3, -1, -1, -2, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, -2, -2, -2, -3, -1, -3, -1, -3, 0, -1, -1, -1, -1, -2, 0, 1, 0, 0, 0, 0, 1, 0, 0, -2, -1, -1, -1, -2, -2, 0, 0, -3, -2, -2, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, -1, -2, -3, -3, -1, -2, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -2, -1, -1, -2, -3, -1, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, 0, -2, 1, 0, 0, 1, 0, -1, -1, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, -1, 0, -2, 0, -1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -2, -2, 0, -2, 0, -1, -1, -2, -2, 1, 1, 0, 0, -1, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, -1, 0, -2, -2, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -1, -1, -2, 0, 0, 2, 0, 0, -2, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, -1, -2, -1, -1, -1, 1, 0, -1, 0, -2, -1, 0, -2, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 1, 2, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 2, 1, 2, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -3, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, -1, 0, 0, -2, -1, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, -2, -3, -1, -1, -2, -1, -1, -1, -2, -2, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, -1, -3, -2, -2, -3, -1, -2, -1, -2, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -2, -1, -2, -2, -4, -2, -1, -2, -1, -1, -1, -1, -1, 0, 1, 1, 0, -1, 0, 0, 0, -1, 0, -1, -1, -2, -2, -1, -2, -3, -2, -1, -2, -3, -2, -2, -2, 0, -2, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -2, -2, -3, -3, -2, -2, -2, -1, -1, -2, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -2, -2, -1, -2, -2, -3, -2, -3, -1, -1, -1, -1, -1, -3, 0, 0, 0, 0, -1, 0, -1, -1, 0, 1, 0, 0, 0, -2, -2, -3, -2, -3, -3, -3, -1, -1, -2, -2, -2, -2, 2, 1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -2, -1, -2, -2, -3, -1, -2, -2, -2, -1, 0, 2, 0, 0, 1, -1, -1, -1, 0, -2, 0, 1, 0, 0, -2, -1, -2, -3, -2, -3, -3, -1, -1, -1, -2, -1, 0, 1, 1, 0, 0, 0, 0, 0, -2, 0, 0, -1, 0, 0, 0, -2, -3, -1, -3, -2, -1, -1, 0, -1, 0, 0, -1, 2, 1, 0, 1, 0, 0, -1, -1, -2, -2, -2, -2, 0, -2, -2, -1, -1, -1, -2, -1, 0, 0, 0, 0, -1, 0, -7, -5, -4, -2, -3, -1, 0, 1, 0, 1, 0, 3, 1, 2, 2, 3, 3, 2, 2, 2, 2, 0, 0, 0, 0, -1, -6, -5, -3, -2, -1, -1, 0, 0, 2, 1, 2, 2, 2, 1, 3, 2, 2, 1, 3, 2, 3, 0, 1, 0, 0, -2, -6, -4, -2, -1, 0, 1, 0, 1, 0, 2, 0, 0, 2, 1, 1, 1, 1, 2, 1, 2, 1, 1, 2, 0, 0, -1, -4, -3, -2, 0, 0, 0, 1, 1, 0, 2, 1, 0, 0, 0, 1, 1, 2, 1, 3, 1, 2, 2, 1, 0, 0, -1, -3, -1, -1, 0, 0, 1, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 3, 2, 1, 0, 0, 0, -3, 0, 0, 1, 1, 0, 1, 3, 1, 2, 0, 0, 0, 0, 0, 0, 1, 1, 2, 3, 3, 1, 0, 0, 1, 1, -2, -1, 0, 1, 1, 0, 1, 2, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 3, 3, 1, 2, 2, 1, 0, -2, 0, 1, 1, 2, 1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 1, 3, 1, 1, 1, 2, -1, 0, 0, 1, 2, 0, 0, 0, 0, 0, -2, -3, -4, -2, -2, -2, -1, -1, 0, 1, 0, 1, 2, 3, 2, 1, -2, 0, 0, 0, 2, 1, 0, 1, 0, -2, -2, -3, -3, -5, -3, -3, -3, -2, -2, -2, 0, 0, 2, 3, 1, 0, -1, 0, 0, 0, 0, 1, 1, 0, -1, -3, -4, -5, -5, -4, -6, -5, -6, -4, -4, -2, 0, 1, 2, 0, 0, 0, -1, 0, 0, 0, 0, 2, 0, 0, -2, -2, -3, -4, -4, -6, -5, -5, -5, -6, -4, -2, -2, 0, 0, 0, 0, 1, -2, 0, 0, 1, 2, 0, 1, 0, 0, -2, -5, -5, -4, -5, -5, -6, -7, -6, -6, -4, -2, 0, -1, 0, 0, 0, -1, 0, 1, 1, 2, 1, 0, 1, -1, -2, -3, -4, -5, -5, -5, -6, -5, -6, -5, -3, -3, -1, 0, 0, 1, 0, -2, 0, 1, 3, 2, 0, 1, 0, -1, -1, -3, -4, -6, -4, -5, -5, -4, -3, -3, -3, -1, 0, 0, 0, 0, 0, -1, 1, 0, 2, 0, 0, 1, 0, 0, 0, -2, -3, -4, -3, -3, -2, -4, -2, -3, -1, -1, 0, 0, 1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, -1, -1, -2, -3, -2, -2, -1, 0, 0, -1, 0, 1, 3, 2, 1, 1, -2, 0, 0, 0, 0, 0, 0, 1, 2, 0, -1, -1, -1, -1, -1, -1, 0, -1, 0, 0, 2, 1, 3, 3, 2, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 3, 1, 2, 2, 2, -2, 0, 0, 1, 0, 0, 0, 1, 2, 1, 1, 2, 0, 0, 1, 0, 0, 1, 0, 0, 0, 3, 1, 3, 2, 1, -1, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 2, 0, 2, 2, 2, 1, 1, 0, -2, -1, -1, 0, 0, 0, 2, 0, 0, 0, 0, 1, 0, 0, 2, 1, 2, 1, 1, 1, 2, 2, 2, 1, 0, 0, -3, -3, -2, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 2, 1, 1, 2, 3, 3, 2, 2, 2, 0, 0, 0, -6, -3, -3, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 1, 1, 4, 2, 3, 1, 2, 1, 0, -1, -2, -7, -5, -3, -3, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 3, 3, 1, 1, 0, 0, 0, 0, 0, -1, -7, -5, -4, -3, -4, -2, -1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 0, 0, 0, 0, -2, -1, -1, -3, -4, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -6, -3, -3, -1, 0, -1, 0, 0, 1, 0, 0, 0, 2, 2, 1, 1, 2, 1, 1, 3, 3, 3, 2, 1, 0, 0, -5, -4, -1, -2, 0, -1, 0, 0, 1, 0, 0, 1, 2, 2, 0, 1, 2, 2, 2, 2, 1, 3, 1, 2, 1, 0, -5, -3, -2, 0, 0, 0, 0, 2, 2, 1, 1, 1, 2, 0, 1, 1, 2, 2, 3, 2, 2, 2, 1, 0, 0, 0, -3, -1, 0, -1, 0, 1, 0, 2, 1, 1, 0, 1, 1, 0, 0, 0, 0, 2, 0, 1, 2, 2, 0, 1, 1, 0, -2, -1, 0, 1, 1, 0, 1, 0, 2, 2, 2, 2, 1, 0, 0, 0, 0, 0, 1, 0, 2, 2, 0, 0, 1, 1, -2, -1, 1, 2, 0, 0, 1, 1, 2, 2, 2, 1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, -3, 0, 1, 3, 1, 2, 0, 1, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 3, 2, 1, 0, 1, 1, -1, 0, 0, 3, 1, 2, 0, 1, 1, 0, 1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 2, 2, 1, 0, 1, 2, -1, 1, 1, 2, 1, 0, 2, 1, 0, 0, 0, -2, -2, -1, -2, 0, 0, -1, 0, 1, 0, 0, 2, 1, 3, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, -3, -2, -2, -1, -1, 0, 0, -1, -1, 0, 2, 1, 2, 2, -1, 0, 2, 1, 0, 0, 0, 2, 0, 1, 0, -3, -3, -3, -3, -3, -1, -2, -1, -2, 0, 1, 0, 1, 3, 4, -1, 0, 0, 1, 0, 2, 1, 1, 1, 1, 0, -3, -2, -3, -1, -1, -3, -2, -2, -2, -1, 0, 0, 3, 2, 2, -1, 0, 1, 1, 0, 3, 1, 2, 1, 0, -1, -2, -2, -3, -2, -3, -1, -2, -4, -4, -1, -1, 0, 0, 2, 1, -2, 0, 1, 2, 1, 2, 3, 2, 2, 0, -1, -1, -3, -1, 0, -2, -1, -1, -3, -4, -2, 0, 0, 0, 1, 2, -1, 0, 0, 2, 1, 2, 1, 1, 1, 0, 0, 0, -2, -2, 0, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, 1, -1, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, -1, -1, 0, 0, 1, 2, 2, 0, 1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, -2, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 3, 2, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 1, 2, 0, 1, 0, 1, 1, 2, 3, 2, 1, 1, 0, 1, 0, 1, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 1, 1, 2, 1, 1, -2, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 2, 0, 1, 0, 1, 2, 1, 2, 0, 2, -2, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 2, 2, 2, 1, 2, 2, 0, 1, 0, 0, 1, 2, 1, 0, -2, 0, 0, 1, 0, 0, 0, 2, 0, 0, 1, 1, 2, 1, 1, 2, 1, 2, 1, 2, 3, 1, 3, 2, 1, 0, -4, -2, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 2, 0, 2, 2, 1, 3, 1, 1, 1, 1, 1, 1, 1, 0, -5, -2, -2, -1, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 1, 2, 1, 1, 3, 1, 2, 1, 1, 1, 0, 0, -5, -4, -2, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 2, 2, 1, 1, 0, 0, -1, 0, -1, 0, -7, -4, -4, -3, -2, -2, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 1, 1, 0, 0, -1, -2, -2, -2, -1, -3, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -2, -1, 0, 0, -2, -1, -1, -1, -1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, -1, 0, -1, 0, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 1, 0, 0, -1, 0, -1, -2, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -2, -2, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, -2, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 2, 2, 1, 1, -1, 0, -1, 0, 0, 1, 2, 5, 6, 0, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, 2, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 2, 5, 3, -1, -2, -2, 0, -1, -1, -2, -1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 2, 4, 3, 0, -2, -2, 0, -2, -1, -1, -2, 0, -1, 0, 1, 0, 0, 0, 0, 0, 2, 0, 0, 1, 1, 3, 3, 3, 5, 0, 0, -1, 0, 0, -2, -2, -2, -1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 4, 5, 0, 0, -1, 0, -1, 0, -2, -2, -1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 3, 4, -1, -1, 0, -1, -1, 0, -2, -1, 0, 0, 0, 2, 2, 0, 0, -1, 0, -1, 0, 0, 2, 2, 2, 4, 5, 4, 0, -2, 0, 0, 0, -2, -1, -1, 0, 2, 2, 2, 0, 0, -1, 0, 0, -1, -1, 1, 1, 3, 3, 4, 5, 6, -1, 0, -1, -1, -2, -1, 0, 0, 2, 2, 3, 4, 2, 0, 0, -1, -2, 0, -1, 0, 2, 2, 2, 3, 5, 5, 0, 0, 0, 0, 0, 0, 1, 2, 3, 5, 6, 4, 3, 2, 0, -1, -1, -1, -2, 0, 0, 0, 1, 4, 3, 5, 0, 0, 1, 0, 2, 1, 4, 2, 4, 6, 6, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 3, 0, 1, 2, 1, 1, 2, 3, 5, 4, 4, 4, 4, 2, 0, -1, -1, -1, 0, 0, -2, -1, -2, 0, 2, 3, 5, 2, 2, 3, 3, 2, 2, 4, 4, 7, 4, 3, 1, 1, -1, -2, -1, 0, 0, 0, -2, -3, -3, 0, 1, 1, 4, 2, 2, 2, 3, 1, 3, 4, 5, 6, 4, 4, 0, 0, 0, -2, -1, 0, 0, -1, -2, -3, -2, -2, 0, 2, 3, 1, 2, 0, 1, 3, 2, 3, 5, 5, 4, 3, 1, 0, -1, -2, 0, 0, -1, 0, -2, -4, -3, -2, 1, 3, 3, 1, 0, 1, 2, 1, 2, 2, 4, 4, 2, 1, 0, 0, 0, -2, -1, 0, -1, -1, -2, -4, -3, -2, 0, 4, 4, 0, 1, 0, 0, 1, 2, 2, 2, 3, 2, 1, 1, 0, 0, -1, 0, -1, -1, -3, -2, -3, -2, -1, 0, 3, 4, 0, 0, 0, 2, 1, 1, 1, 1, 2, 1, 2, 1, 0, 0, 0, 0, -1, 0, -1, -1, -4, -2, -1, 1, 4, 6, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 0, 0, -2, -1, -1, -1, -1, -1, -2, -2, 0, 1, 5, 5, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, -1, 0, -1, 0, 0, -1, -1, 0, 1, 3, 3, 4, 3, 1, 0, 0, 0, -1, 0, -2, 0, 0, -1, -2, -3, -2, -2, -2, -2, 0, -1, 0, -2, 0, 0, 1, 3, 5, 2, 1, 0, -1, 0, 0, -1, -2, 0, -2, -1, -2, -2, -1, -2, -1, -1, -1, 0, -2, 0, 0, 0, 0, 1, 3, 2, 1, 0, -1, -2, 0, -1, 0, -1, -1, -1, 0, 0, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 2, 4, 2, 0, -1, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 2, 3, 3, 0, -1, -2, -1, -2, 0, 0, 1, 2, 2, 1, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 2, 3, 3, 4, 0, -1, -1, -2, -1, 0, 0, 1, 3, 3, 2, 3, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, 2, 2, 4, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 2, 2, 1, 3, 2, 2, -1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 1, 2, 2, 1, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 1, -1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 3, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 2, 2, 3, 0, 0, 0, 0, 1, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 2, -1, 0, 0, 0, 1, 0, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 2, 2, 3, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 2, 3, 2, 1, 1, 1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 3, 3, 4, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, -2, -1, 0, 0, -1, 0, 0, 0, 0, 2, 1, 3, 4, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -2, 0, 0, 0, -1, 0, 0, 0, 2, 1, 2, 3, 2, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 0, -1, -1, 0, -1, 0, 0, 0, 1, -1, 0, 0, 1, 2, 3, 3, 0, 1, 0, 1, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 2, 1, 3, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 3, 2, 0, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 0, 0, 0, 1, 0, 1, 3, 3, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 0, 0, 0, 0, 1, 2, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 0, 0, 0, 2, 1, 2, 1, 0, 0, 0, 0, -1, 0, -2, -1, 0, 0, 0, 0, 2, 1, 1, 2, 1, 0, 0, 1, 0, 0, 0, 1, 2, 1, 1, 1, 2, 1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 2, 2, 2, 2, 0, -1, 0, -1, 1, 1, 1, 2, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 2, 1, 2, 2, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 2, 1, 1, 1, 1, 1, 1, 0, 1, 0, 2, 2, 3, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 0, 2, 1, 1, 1, 1, 2, 2, -1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, -1, 1, 1, 2, 1, 2, 1, 0, 2, 1, 2, 1, 2, 0, 2, 0, -1, -1, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 3, 0, 2, 1, 3, 0, 0, 0, 0, 1, 1, 1, -1, 0, -1, -1, 0, 0, 0, 2, 2, 1, 2, 1, 2, 2, 1, 2, 2, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, -2, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, -2, 0, -1, 0, 0, -2, -1, -1, 0, -1, -1, 0, -3, -1, -1, 0, -1, -2, 0, -1, 0, -1, -2, -1, 0, -1, -1, -2, -1, 0, -2, -1, -1, -1, 0, -1, -1, -2, -1, -2, -1, -2, -2, -1, -1, 0, -1, -3, -1, 0, 0, 0, -2, -2, -1, 0, 0, -2, 0, 0, -1, 0, -1, -1, 0, -2, -2, -1, -2, -2, -1, 0, -1, -1, -1, -1, -2, -1, -3, -2, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, -1, -3, -1, -2, -1, -1, -1, -1, -1, -1, -2, -2, -1, -2, -2, 0, 0, -2, -1, -1, -1, -1, -2, 0, -1, 0, -1, -1, -2, -1, -1, -1, 0, -1, -1, -1, -1, -1, -2, -3, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, -2, -1, -2, -1, 0, 0, -1, 0, -2, -2, -2, -2, -1, -4, -3, -1, 0, -1, -1, 0, -2, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -2, -2, -1, -3, -1, -2, -1, 0, -3, -3, -2, -3, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, -1, 0, -3, -1, -1, -2, -1, -2, -2, -2, -3, -3, -4, -3, -1, -1, -2, 0, 0, 0, 1, 0, -1, -2, -3, -1, 0, -2, -2, -2, -1, -2, -2, -1, -1, -1, -5, -4, -3, -3, -2, -2, -3, 0, 1, 0, 1, -1, 0, -2, -2, -1, -1, 0, -3, -2, -3, -2, -4, -3, -2, -1, -4, -4, -2, -1, -3, -3, -2, 0, -1, 0, 1, 0, -1, -1, -2, -1, -2, -1, 0, -2, -2, -2, -2, -1, -2, -1, -3, -3, -2, -2, -2, -2, -2, -1, 0, 0, 1, 1, 1, -1, -2, -2, -1, -1, -1, -1, -2, -1, -3, -2, -1, 0, -3, -2, -3, -2, -3, -3, -2, -2, 0, 0, 1, 1, 0, -1, -1, -2, -1, 0, 0, -1, -2, -1, -2, -2, -2, -1, -2, -3, -2, -3, -4, -3, -4, -1, 0, 1, 0, 0, 0, -1, -2, -2, -2, -3, 0, -1, -2, -1, -3, -1, -1, -1, -4, -2, -2, -4, -2, -3, -3, 0, 0, 0, 1, 1, 0, -1, -1, -2, -3, -2, 0, -2, -2, 0, -3, -2, -2, 0, -2, -2, -3, -4, -2, -2, -2, -1, -1, 0, 1, 0, 0, -1, -2, -2, -1, -3, -2, -1, -1, -2, -2, -2, -1, -1, -2, -2, -1, -3, -2, -2, -1, -2, 0, 0, 0, 0, 0, -1, -2, -3, -1, -2, -1, -3, -2, -2, -3, -1, -1, -1, -3, -3, -3, -2, -1, -1, -3, -1, -1, 0, 2, 0, 0, -2, -3, 0, 0, -3, -1, -1, -1, -2, -2, 0, -1, -1, -3, -2, -1, -3, -2, -3, -2, 0, -2, -1, 1, 0, 0, -2, -1, 0, 0, -2, -2, -3, -1, -1, -2, -3, -1, -2, -2, -2, -1, -2, -2, -3, -3, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -3, -3, -2, -1, -1, -2, -3, -1, -2, -2, -1, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -2, -2, -2, -2, 0, -3, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -3, -1, 0, 0, 0, -2, -1, -2, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, -1, -3, -1, -1, 0, -1, -3, -2, -1, -1, 0, 0, 0, -1, -1, -1, -2, -3, -1, -1, -1, -1, -2, 0, 0, -1, -2, -1, -2, 0, -1, 0, -1, -2, -1, 0, -2, -2, -1, 0, -1, -2, -3, -2, -1, -3, -3, -1, -1, -1, 0, 0, -1, 0, 0, -2, -1, 0, -4, -1, -1, -1, -1, -1, 0, -1, -1, 0, -2, -2, -1, -1, -2, -2, -2, 0, 0, 0, -1, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 1, -1, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, 0, -1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -2, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 1, 0, 0, -2, 0, -2, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, -2, 0, -2, -2, 0, 0, -1, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, 0, -2, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -1, -1, -2, -3, 0, 0, -2, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -3, -1, -1, -1, -1, -1, -2, 0, -2, -1, -2, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -3, -2, -2, -2, -1, -2, -1, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, -2, -2, -2, -2, -1, -2, 0, -1, -1, -1, 1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, -1, -2, -2, -1, -2, -1, -1, -1, -1, -2, -1, -2, -1, -1, 0, 1, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, -1, -2, -1, 0, -2, -1, -2, -2, -2, -2, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -3, 0, -3, -3, -2, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, -1, -2, -3, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -2, -1, -1, -2, 0, -2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -3, -2, -1, -1, -2, 0, -1, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, -2, -1, -1, -1, -1, 0, 0, -1, -2, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 2, -1, -1, -1, -1, -1, -2, -1, 0, -1, 0, -1, 0, -2, 0, 0, -1, -1, 0, 1, 0, 0, 2, 0, 1, 2, 2, -1, -1, -1, -1, -1, 0, -1, 0, 0, -1, 0, -1, -1, -2, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 2, -1, 0, -1, -1, -1, -1, -1, 0, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 1, 0, 1, 1, 0, 1, 2, 0, 0, -2, -1, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 2, 1, 1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 2, 2, 0, 0, -1, 0, 0, -1, -2, 0, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, -2, -2, -2, -2, 0, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, 0, 0, -1, -1, -1, -3, -1, -1, -1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, -1, -1, 0, 0, -2, -3, -1, -2, 0, 0, -1, 0, 0, 1, 2, 1, 1, 0, 2, 0, 1, 1, 0, 0, 0, 0, -2, 0, -2, -1, -2, -1, -2, -2, 0, -1, 0, 1, 0, 1, 2, 0, 1, 2, 3, 2, 1, 0, 2, 1, 1, 1, 0, 0, -1, -3, -3, -2, -1, -2, -1, 0, -1, 0, 0, 1, 1, 2, 2, 1, 3, 0, 1, 0, 1, 1, 1, 0, -1, 0, -1, -2, -2, -1, -2, -2, -2, -1, 0, 1, 1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 1, 1, 1, 0, -2, 0, -1, -3, -2, -4, -2, -1, -1, -1, 0, 0, 2, 1, 2, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -3, -3, -1, -1, -1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, -1, -1, -1, 0, -2, -3, -1, -1, -2, 0, 0, 0, 0, 2, 1, 1, 1, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, -1, -2, -1, 0, -2, -1, -2, -1, -1, 0, 1, 2, 2, 0, 0, 1, 0, -1, -1, -2, -2, -1, 0, 0, 2, 0, -1, -2, -1, 0, -1, -2, -1, 0, -2, -1, 0, 1, 1, 1, 2, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, -1, 0, -1, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, -1, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 2, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 2, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 2, -8, -7, -5, -4, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 1, 2, 2, 2, 2, 2, 1, 0, -1, -3, -3, -4, -7, -4, -3, -2, 0, 0, 1, 0, 0, -1, 0, -1, 1, 0, 1, 3, 3, 2, 3, 3, 2, 1, -1, -1, -2, -3, -6, -2, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 2, 3, 4, 3, 3, 0, 0, 0, -1, -1, -5, -1, -2, -1, 1, 1, 2, 2, 1, 0, -1, 0, 0, 0, 0, 0, 2, 3, 1, 2, 1, 2, 0, 0, 0, -2, -4, -2, -1, 0, 0, 1, 1, 2, 2, 1, 0, 0, -1, 0, 0, 1, 2, 1, 3, 2, 1, 0, 0, -1, -1, -1, -2, 0, -1, -1, 1, 2, 2, 1, 2, 1, 0, -1, -2, 0, 0, 0, 0, 2, 3, 1, 1, 0, 0, 0, 0, -1, -2, 0, -1, 1, 1, 0, 2, 3, 0, 0, 0, -1, -1, 0, 0, 0, 2, 3, 2, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, -1, -2, -2, -1, 0, 0, 0, 1, 0, 2, 2, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -3, -5, -3, -3, -2, -1, 0, 0, 1, 0, 1, 2, 0, 1, 0, 1, 0, -1, 0, 0, -1, -1, -1, -1, 0, -2, -4, -4, -5, -3, -3, -3, -2, -1, 0, -1, 0, 0, 2, 2, 2, 2, 1, -1, -1, -2, 0, -1, -1, -1, -1, -2, -5, -6, -4, -5, -3, -2, -2, -2, -3, -3, -1, 1, 2, 1, 2, 2, 1, -1, 0, -1, -2, 0, -1, -1, -2, -4, -6, -6, -5, -3, -3, -4, -5, -4, -4, -4, -2, 0, 1, 2, 1, 1, 0, -3, -1, -1, -1, 0, 0, 0, -1, -3, -6, -5, -4, -3, -4, -4, -5, -4, -6, -4, -1, 0, 0, 3, 3, 0, 0, -2, -1, -1, -1, 0, -1, 0, -2, -2, -4, -4, -2, -1, -2, -3, -4, -6, -5, -3, -2, 0, 0, 0, 1, 0, 0, -3, -1, 0, 0, 1, 0, -1, -2, -4, -4, -4, -2, -3, -1, -3, -4, -3, -5, -4, -2, 0, 0, 1, 2, 0, 0, -2, -1, 0, 0, 0, -1, -2, -3, -2, -3, -3, -2, -3, -3, -4, -3, -3, -3, -2, 0, 1, 1, 1, 1, 0, 0, -1, 0, -1, 0, -1, -1, -1, -3, -3, -4, -4, -2, -1, -1, -1, -2, -3, -2, 0, 0, 1, 2, 2, 1, 0, 0, -2, -1, 0, 0, -1, -2, -1, 0, -1, -2, -2, -1, 0, 0, -1, 0, -1, 0, 1, 0, 3, 1, 2, 0, 0, 0, -2, -1, -1, -1, -2, -2, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 1, 2, 0, 0, 0, -1, 0, 0, 0, 0, -2, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 2, 1, 2, 3, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 3, 3, 0, 0, 0, -3, -2, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 2, 2, 3, 3, 1, 1, 0, -2, -3, -2, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 2, 3, 3, 3, 0, -1, -2, -4, -4, -1, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, 0, 1, 1, 2, 2, 1, 4, 3, 2, 1, -1, -2, -4, -7, -5, -3, -2, -1, 0, 0, 0, -2, -1, -3, -1, 0, 0, 0, 0, 1, 2, 1, 2, 1, 0, 0, -1, -2, -5, -8, -6, -5, -4, -1, 0, -2, -1, -1, -3, -3, -3, -1, -1, 0, 0, 1, 0, 0, 0, -1, -1, -2, -4, -4, -6, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, -2, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, -2, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, -1, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 1, 1, 0, 0, 0, 0, -1, 1, 0, 0, 1, 1, 0, 0, 0, -2, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, -1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, 1, -1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 1, 1, 2, 0, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, -1, 0, -2, -1, 0, 0, 0, 0, 1, 0, 0, 2, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 2, 1, 1, -1, 0, 0, -1, -1, 0, 0, -1, 0, -2, 0, 0, -1, -1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, -1, -2, -1, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, -2, 0, -2, 0, 0, -1, 1, 0, -1, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -2, -1, -2, -1, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, -3, -2, 0, -1, -1, 0, -1, -2, -1, -3, -2, -2, -2, 3, 4, 2, 1, 0, 0, -1, 0, 0, 0, -2, -2, -2, -2, -1, -1, -1, -2, -1, -2, 0, 1, 1, 4, 3, 4, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, -2, -1, -1, -1, 0, -1, 0, 1, 1, 1, 3, 4, 1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -2, -2, -1, -1, 0, 1, 0, 0, 1, 1, 1, 2, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -1, 0, 0, 1, 1, 1, 0, 1, 2, 2, 1, 0, 0, 0, -2, -2, 0, -2, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 1, 0, 0, 1, 2, 1, 3, 2, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 3, 2, 1, 2, 0, -1, 0, -1, -2, -2, -3, -2, -1, 0, 0, 1, 0, -1, -1, -1, 0, -1, -1, -2, 0, 0, 1, 2, 1, 3, -1, -1, -2, -2, -1, -3, -2, -2, -1, 0, 1, 0, 2, 1, 0, -1, 0, -2, -1, -1, -1, 0, 1, 2, 2, 2, 0, -2, -1, -1, -2, -1, -1, 0, 0, 0, 2, 1, 1, 1, 0, -1, -2, -2, -1, -1, 0, 0, 0, 1, 1, 0, -1, -1, -1, -1, -2, 0, 0, 0, 0, 3, 2, 3, 2, 1, 1, 0, -2, -2, -2, 0, -1, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 3, 3, 3, 2, 2, 0, -1, 0, 0, 0, -1, 0, 1, 0, 2, 1, -1, -1, 0, 0, -1, 0, 0, 2, 3, 3, 4, 4, 4, 3, 2, 2, 0, 0, 0, 0, -1, 0, 0, 2, 1, 2, 0, -1, -1, -1, -1, 0, 0, 1, 2, 4, 3, 3, 2, 3, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, -1, -2, -1, -1, -2, 0, -1, 0, 3, 3, 4, 2, 4, 3, 2, 2, 1, 0, -1, 0, -1, 0, 0, 0, 3, 3, 0, -2, -1, -3, -3, -2, 0, 0, 0, 2, 1, 3, 3, 4, 3, 1, 0, 0, 0, -2, -2, -2, -1, -1, 1, 2, 0, -1, -2, -2, -3, -2, -2, 1, 0, 1, 1, 3, 3, 4, 3, 1, -1, -1, -2, -1, -2, -3, -3, 0, 0, 0, 0, -1, -3, -3, -2, -2, 0, -1, 0, 0, 1, 3, 2, 4, 2, 0, -2, -2, -3, -4, -4, -3, -3, -1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 1, 0, 3, 2, 0, 0, 0, -2, -2, -2, -5, -4, -5, -3, 0, 0, 3, 0, 0, -2, 0, 0, 0, -1, -3, -1, 0, 0, 0, 0, 1, 0, -2, -1, 0, -2, -4, -4, -4, -1, 0, 2, 2, 0, 0, -1, 0, 0, -1, 0, -2, -3, -1, -1, 0, 0, -1, -1, -2, -1, 0, -1, -2, -2, -2, -1, 0, 1, 2, 0, 0, -1, 0, 0, 0, -1, -1, -2, -3, -3, -2, -3, -2, -2, -2, 0, -2, -1, -1, -1, 0, 0, 1, 3, 3, 0, -1, 0, 0, -1, -2, -1, -1, -2, -1, -1, -2, -1, 0, -1, 0, 0, 0, -2, -1, -1, -2, 0, 1, 2, 4, 0, 1, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, -1, -2, 0, -1, 0, 1, 2, 3, 2, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, -1, -2, -1, -1, -1, -1, 0, 0, 1, 3, 2, 2, 0, 0, -1, 0, 1, 2, 2, 2, 2, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 2, 3, 3, 0, 0, 0, 0, 0, 0, 3, 4, 4, 4, 3, 1, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 2, 1, 3, 1, 0, 1, 1, 0, 0, 2, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 1, 0, 1, 1, 2, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 2, 1, 1, 1, 1, 0, 0, 1, 2, 1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 1, 0, 2, 0, 0, 2, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 1, 0, 1, 2, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, -1, 0, 0, 2, 2, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, 0, 1, 2, 2, 0, 2, 1, 1, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 3, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 2, 0, 1, 1, 0, 0, 0, -1, -1, 0, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, 1, 0, -2, -2, -1, -2, -1, -1, -2, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, 0, -2, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -2, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, 0, -1, -1, 0, 0, 1, 2, 1, 2, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 2, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, -1, 1, 1, 2, 2, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 2, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 0, 0, 1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 2, 1, 0, 1, 0, 1, 0, 0, 0, 0, 2, 1, 0, 1, 0, 1, 0, 1, 0, -2, 0, 0, 0, 1, 0, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 0, 1, 1, 2, 0, 1, 2, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 2, 2, 2, 2, 2, 1, 1, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, -1, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -2, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -2, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -2, -1, -2, 0, -2, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, -1, -2, -2, -2, 0, -1, -1, -1, -1, 0, -2, -2, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -2, -1, -2, -2, -1, -1, 0, -2, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, -2, -2, -2, -2, -2, -1, 0, 0, 0, -2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -2, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -7, -5, -4, -2, -4, -2, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 2, 1, 2, 0, 0, 2, 1, 0, 1, 0, -6, -5, -3, -2, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 2, 2, 2, 2, 1, 1, 1, 1, 3, 1, 2, 0, -6, -5, -3, -1, 0, -1, 0, 0, 1, 0, 1, 1, 2, 1, 0, 0, 1, 1, 2, 1, 2, 2, 1, 1, 1, 2, -6, -4, -1, -1, 0, -1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 2, 0, 0, 0, 1, 1, 1, 1, 0, -5, -4, -1, 0, 0, 1, 0, 2, 0, 2, 2, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, -3, -3, 0, 0, 0, 1, 0, 1, 2, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 2, 0, 0, 1, 1, -2, -2, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, -1, 1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, -4, 0, 0, 1, 0, 0, 1, 1, 2, 2, 1, 1, 0, -1, 0, -1, 0, 0, 0, 1, 2, 2, 0, 0, 0, 1, -3, 0, 0, 0, 0, 1, 0, 2, 1, 0, 2, 0, -1, -1, -1, -1, 0, 0, 0, 1, 2, 1, 2, 1, 2, 2, -1, -1, 0, 0, 1, 0, 1, 1, 2, 1, 1, -1, -3, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, -3, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -2, -1, -3, -2, -1, -1, -1, 0, 1, 0, 2, 2, 1, -2, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, -1, -3, -1, -3, -1, -3, -3, -2, -2, -2, -1, 0, 1, 0, 2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -2, -2, -1, -2, -3, -1, -3, -2, -4, -2, -1, 0, 1, 1, 1, -2, -1, 0, 0, 1, 1, 1, 2, 2, 1, 0, -1, -2, -1, -2, -1, -2, -2, -4, -3, -2, 0, 0, 0, 0, 2, -1, 0, 0, 1, 2, 1, 2, 2, 1, 1, 0, 0, 0, -1, -1, -2, 0, -2, -1, -1, -2, -1, 0, 1, 2, 2, -2, 0, 0, 1, 2, 1, 0, 0, 0, 0, -1, -1, 0, -1, -2, 0, -2, -1, -2, -1, 0, 0, 0, 0, 0, 1, -3, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, -1, 0, -1, -2, 0, -1, 0, 0, -2, 0, 0, 0, 2, 1, 1, -3, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 2, 2, 1, 0, -3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 3, 2, 2, 0, -3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 2, 0, 0, -1, 1, 2, 2, 1, 0, 0, -3, -1, 1, 0, 0, -1, 1, 1, 0, 0, 0, 1, 1, 2, 1, 1, 1, 0, 0, 0, 0, 1, 0, 2, 2, 0, -3, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 1, 1, 1, 1, 2, 1, 0, 1, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 1, 1, 0, 1, 2, 2, 2, 2, 3, -5, -2, -2, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 2, 1, 2, 0, 2, 2, 2, 1, -6, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 2, 2, 2, 0, 1, 0, 0, 1, -6, -3, -2, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 0, 1, 0, 0, 0, -5, -4, -4, -2, -1, -1, 0, 0, 0, 1, 1, 2, 2, 4, 4, 3, 2, 3, 2, 0, 0, 0, -2, -1, -1, -1, -4, -2, -3, -1, 0, 0, 0, 0, 2, 0, 3, 3, 3, 3, 2, 3, 2, 2, 0, 1, 0, 1, 0, 0, -1, 0, -4, -1, -1, -1, 1, 0, -1, 0, 1, 2, 1, 1, 2, 2, 1, 3, 3, 2, 2, 0, 2, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 2, 0, 1, 2, 1, 1, 1, 1, 3, 2, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 2, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, 2, 2, 2, 3, 2, 2, 1, 0, 0, 0, -2, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 2, 3, 1, 2, 2, 2, 1, 1, -1, 0, 0, 1, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 3, 3, 3, 2, 3, 2, 1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 2, 2, 2, 1, 2, 3, 2, 3, 0, 0, 2, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, -2, -2, -3, 0, -1, 0, 0, 1, 1, 1, 3, 2, 3, 0, 0, 1, 2, 1, 0, 1, 1, 0, 0, -2, -1, -2, -4, -4, -3, -3, -3, -1, 0, 0, 1, 2, 2, 2, 1, -1, 0, 1, 1, 1, 1, 1, 0, 0, -2, -2, -3, -4, -4, -4, -3, -3, -3, -2, -2, -1, 0, 0, 0, 1, 1, -1, 1, 1, 1, 1, 2, 1, 0, 0, -3, -4, -4, -6, -5, -7, -5, -5, -4, -4, -2, -3, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 1, 1, -1, -1, -5, -5, -6, -7, -6, -5, -4, -4, -5, -3, -3, 0, 0, -1, 0, 0, 0, 0, 0, 3, 3, 1, 1, 1, 0, -1, -4, -5, -6, -7, -7, -6, -6, -4, -5, -5, -3, -1, 0, 0, 0, 0, 0, 1, 1, 2, 3, 0, 2, 0, 0, -2, -3, -6, -5, -7, -6, -4, -4, -3, -4, -3, -2, -1, 0, 0, 0, 1, 0, 1, 1, 2, 3, 1, 2, 1, 0, 0, -3, -4, -4, -5, -5, -5, -3, -3, -3, -2, -2, 0, 0, 1, 2, 0, 0, 1, 1, 2, 1, 2, 1, 0, 1, 0, -1, -4, -5, -4, -3, -2, -3, -2, 0, -2, 0, 0, 1, 0, 0, 2, 0, 1, 1, 2, 2, 0, 0, 1, 0, -1, 0, -1, -3, -2, -2, -1, 0, -1, -1, -1, 0, 1, 0, 2, 1, 1, 0, 0, 0, 1, 0, 0, 0, 2, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 2, 2, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 3, 1, 2, 0, -1, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 2, 1, 0, -1, -1, -1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 2, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 2, 3, 3, 2, 0, 0, 0, 0, 1, 0, -1, -3, -1, -1, -2, -1, -1, 0, 0, 1, 0, 0, 2, 1, 2, 1, 3, 3, 3, 2, 0, 1, 0, 0, 0, 0, -1, -2, -2, -2, -2, -2, -1, 0, 0, 0, 1, 1, 2, 2, 1, 3, 3, 3, 2, 2, 1, 0, -2, -1, -2, -1, 0, 0, 0, 0, 1, 0, 2, 2, 3, 2, 0, 2, 1, 0, 0, 0, 0, 0, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 3, 2, 2, 1, 2, 2, 2, 1, 2, 0, 2, 1, 2, 1, 0, 0, 0, 0, 1, 0, 1, 1, 2, 0, 0, 2, 3, 2, 1, 0, 0, 1, 2, 1, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 2, 0, 1, 0, 1, 3, 2, 0, 2, 1, 2, 2, 0, 2, 0, 1, 2, 2, 2, 0, 1, 0, 1, 0, 0, 1, 1, 1, 1, 1, 1, 3, 1, 0, 1, 2, 2, 1, 0, 0, 0, 0, 0, 1, 2, 2, 1, 2, 1, 2, 0, 1, 1, 2, 2, 1, 2, 1, 3, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 3, 1, 1, 2, 0, 0, 3, 1, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 2, 3, 1, 2, 2, 2, 3, 3, 1, 1, 0, 1, 0, 1, 1, 0, -1, -1, 0, -1, 0, 0, 0, 1, 0, 1, 2, 0, 2, 2, 0, 1, 2, 2, 3, 3, 1, 1, 0, -1, -1, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 2, 1, 2, 2, 1, 1, 1, 0, -2, -3, -1, -2, -2, -1, -1, 0, 0, 1, 0, 0, 1, 0, 0, 2, 0, 0, 1, 1, 3, 1, 2, 0, 0, -1, 0, -2, -2, -3, -1, -2, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 2, 1, 0, 1, 0, -1, -2, -1, -3, -2, -2, -4, -2, -2, -2, 0, 0, -1, 0, 1, 0, 1, 1, 0, 0, 1, 3, 3, 0, 0, 0, -1, -1, -2, -3, -4, -4, -4, -2, -2, -1, -2, 0, -1, -1, 0, 0, 0, 1, 0, 0, 2, 1, 1, 1, 0, 0, 0, -2, -3, -3, -4, -5, -4, -3, -3, -2, 0, -1, 0, -1, 0, 0, 0, 1, 0, 1, 1, 2, 1, 2, 0, 0, -2, -2, -2, -4, -3, -5, -2, -3, -1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 3, 1, 2, 0, 0, 0, 0, -2, -2, -2, -4, -2, -2, -2, -1, -2, -2, -1, -1, 1, 0, 0, 0, 0, 0, 2, 2, 3, 3, 3, 1, 0, 0, 0, -1, -3, -1, -2, -3, 0, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 2, 3, 2, 2, 0, 0, 0, -1, -2, -3, -1, -2, 0, -1, -1, 0, 0, 1, 0, 2, 2, 1, 0, 0, 2, 3, 3, 4, 3, 2, 0, 0, -1, -1, -2, -1, -2, -1, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 1, 0, 2, 3, 4, 3, 4, 1, 0, 1, 0, -1, 0, -2, 0, -1, 0, 1, 0, 0, 1, 1, 0, 2, 0, 0, 1, 1, 0, 1, 4, 2, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 1, 0, 2, 3, 1, 2, 1, 3, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 0, 1, 1, 2, 2, 1, 0, 0, 2, 1, 2, 3, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 1, 0, 1, 1, 1, 1, 1, 2, 2, 1, 2, 2, 2, 1, 1, 0, 1, 0, 1, 0, 3, 1, 1, 2, 1, 0, 1, 3, 0, 0, 0, 0, 0, 2, 2, 2, 1, 1, 2, 2, 0, 1, 1, 2, 2, 1, 1, 1, 1, 2, 2, 2, 1, 2, 2, 0, 0, 0, 1, 0, 2, 3, 2, 1, 3, 1, 2, 2, 1, 2, 2, 2, 3, 3, 2, 1, 2, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, -1, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, -1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, -1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 1, 1, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 2, 2, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 2, 1, 0, -1, -1, -1, -1, 0, -1, -1, -1, -1, -2, -1, 0, 0, 0, 1, 0, 0, 1, 1, 2, 1, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 2, 2, 1, 2, 2, 1, 1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 2, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, 1, 0, 0, 0, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 3, 2, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, -1, 0, 1, 0, 2, 2, 2, 2, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 3, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, -1, 1, 0, 0, 0, 2, 1, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 3, 1, 3, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 1, 1, 0, 0, 1, 0, -1, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 3, 4, 4, 4, 4, 4, 5, 4, 4, 5, 5, 2, 3, 1, 2, 0, 0, 0, 0, -2, -1, 2, 0, 2, 1, 3, 4, 3, 4, 4, 4, 3, 3, 6, 5, 6, 3, 2, 2, 0, 0, 2, 0, -1, -1, 0, -1, 2, 0, 0, 2, 2, 2, 2, 5, 4, 2, 4, 4, 6, 6, 4, 4, 2, 1, 2, 0, 0, 1, 0, 0, -1, -1, 2, 1, 0, 2, 0, 2, 3, 5, 4, 3, 4, 4, 6, 6, 3, 3, 3, 0, 0, 0, 1, 1, 1, 0, 0, 0, 3, 1, 1, 0, 0, 2, 2, 4, 3, 4, 2, 5, 5, 4, 3, 1, 1, 1, 0, 0, 1, 0, 0, 2, 1, 0, 2, 2, 1, 1, 2, 1, 1, 4, 2, 4, 3, 4, 3, 3, 2, 1, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 2, 2, 0, 1, 1, 1, 1, 2, 3, 4, 3, 5, 5, 3, 2, 0, 0, 1, 0, 0, 1, 1, 2, 2, 1, 1, 2, 1, 2, 1, 0, 0, 1, 1, 1, 2, 3, 3, 4, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 1, 1, 4, 3, 2, 1, 0, 0, 2, 2, 1, 1, 1, 2, 2, 3, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 2, 0, 4, 1, 1, 2, 1, 0, 1, 1, 0, 1, 0, 2, 1, 1, 1, -1, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 3, 4, 2, 3, 3, 1, 2, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 3, 2, 2, 1, 1, 3, 2, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -2, -1, -1, 0, 0, 0, 0, -1, 0, 2, 3, 3, 1, 1, 2, 2, 1, -1, 0, -2, 0, 0, 0, 0, 0, -2, -1, -2, -2, -1, 0, 0, -1, -1, -1, 3, 2, 2, 1, 2, 1, 2, 0, 0, -1, -1, -2, -1, 0, 0, 0, -2, -2, -1, -1, -2, -1, 0, 0, 0, 0, 2, 3, 2, 1, 1, 1, 2, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, -2, -1, -1, -1, -1, 0, -1, 0, -1, 1, 2, 1, 2, 2, 2, 2, 0, 0, 0, -2, 0, 0, -1, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 3, 1, 2, 1, 2, 2, 3, 2, 2, 0, -1, 0, 0, 1, 1, 0, 0, -2, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 1, 2, 4, 3, 1, 1, 0, 0, 1, 1, 0, 0, -1, -2, 0, 0, 1, 1, 1, 0, 0, 0, 2, 1, 2, 2, 3, 1, 3, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 0, 0, 0, 1, 1, 2, 3, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 2, 1, 2, 2, 2, 1, 0, 1, 0, 0, 1, 0, 3, 3, 2, 1, 2, 0, 1, 2, 1, 0, 0, 1, 1, 0, 2, 1, 1, 1, 2, 0, 0, 1, 2, 0, 1, 0, 1, 2, 2, 4, 2, 1, 0, 1, 0, 0, 1, 1, 2, 1, 2, 3, 3, 4, 1, 1, 0, 0, 0, 1, 0, 2, 1, 3, 4, 3, 3, 2, 1, 2, 2, 3, 2, 2, 0, 1, 2, 2, 2, 3, 2, 2, 1, 2, 1, 0, 0, 2, 1, 4, 5, 3, 3, 2, 3, 3, 3, 2, 1, 3, 1, 1, 2, 2, 2, 3, 3, 1, 1, 1, 1, 0, 0, 2, 1, 2, 3, 4, 4, 2, 3, 4, 3, 2, 1, 2, 1, 1, 2, 2, 2, 2, 2, 3, 1, 1, 2, 2, 0, 2, 3, 3, 4, 5, 4, 4, 4, 4, 3, 2, 2, 3, 2, 2, 3, 3, 3, 3, 3, 2, 2, -4, -3, -3, -3, -1, 0, 0, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, -2, -5, -3, -1, -2, -1, -1, -1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 1, 1, 2, 0, 0, 1, 0, -1, -1, -2, -4, -4, -2, 0, 0, -1, 0, -1, -2, 0, -2, -1, 0, -1, 0, 0, 1, 2, 0, 0, 1, 0, 0, 0, 0, -2, -3, -2, -2, 0, -1, -2, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 2, 1, 1, 1, 0, 0, 0, -2, -4, -2, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 2, 0, 0, 0, -1, -2, 0, -2, -1, 0, -1, -1, 0, -1, 0, 1, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, 2, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, 0, -2, 0, 1, 1, 0, 0, -1, 0, 0, -1, -2, -1, -2, -2, 0, -1, 0, 1, 1, 0, 1, 0, 0, -1, -1, -2, 0, 0, 0, -1, 0, 0, 0, -1, -1, -2, -2, -3, -2, -2, 0, -2, 0, 0, 0, 0, 1, 1, 0, 0, -1, -2, -2, -1, -1, 0, 0, -1, -1, -2, -1, -2, -2, -2, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -2, 0, 0, -2, -1, -1, 0, -2, 0, -2, -2, -2, -1, 0, -1, 0, 0, -1, -2, -2, 0, 0, 0, 0, 0, -1, -3, 0, 0, 0, 0, 0, 0, -2, 0, -2, -1, 0, 0, 0, -1, 0, -1, 0, -2, -1, 0, 1, 1, 1, 1, 0, -3, -3, -2, 0, 0, -1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, -2, -2, -2, -1, -1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, -2, -2, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, -1, -1, 0, -3, -2, -2, -2, 0, 0, -1, -1, -1, -1, -2, -1, 1, 0, 0, 1, 0, 0, 0, 0, 2, 1, 0, 0, 0, -1, -3, 0, -1, 0, -2, -1, 0, -1, -2, -1, -2, -2, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 2, 0, 0, -2, -2, -1, -1, -1, -2, -2, -1, -2, -3, -1, -2, 0, 0, 0, 0, 2, 1, 2, 2, 0, 1, 2, 2, 0, 0, 0, -1, -2, -1, 0, -2, -1, 0, 0, -1, 0, 0, 1, 0, 1, 2, 2, 1, 0, 1, 1, 1, 0, 0, 0, -1, 0, -1, -2, 0, 0, -1, 0, -1, 0, -1, -1, 0, 2, 1, 1, 0, 1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, -2, -1, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, -2, -1, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 2, 2, 1, 1, 0, 0, 0, 3, 0, 1, 0, 0, -4, -1, -1, -1, -1, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 2, 0, -2, -1, -5, -3, -2, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 2, 1, 1, 0, 0, -3, -6, -3, -2, -2, -1, 0, 0, -1, 0, -1, -2, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -2, -3, -2, -3, -6, -4, -3, -4, -1, -1, -2, -2, -3, -1, -2, -2, -3, -3, -3, -1, 0, 0, -1, -1, 0, -2, -3, -3, -5, -5, 0, -1, 0, 0, 0, 0, 1, 0, 0, 2, 2, 3, 2, 3, 4, 3, 2, 2, 1, 0, 0, 1, 0, 0, 2, 3, -1, -1, 0, -1, 0, 0, -1, -1, 0, 1, 1, 2, 1, 2, 2, 2, 3, 0, 1, 0, 1, 0, 1, 0, 2, 3, 0, -1, 0, -1, 1, 0, -1, 0, 0, 1, 1, 2, 0, 1, 2, 2, 1, 0, 1, -1, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 2, 1, 0, 0, 2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 2, 1, 1, 1, 1, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 1, 1, 1, 4, 1, 0, 0, 1, 2, 0, 1, 0, 1, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 2, 4, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, -1, 1, 1, 0, 0, 0, -1, 0, 1, 0, 0, 2, 3, 4, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 2, 2, 4, 5, 5, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -2, -1, 0, 0, 0, 3, 3, 6, 5, 2, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -2, -2, -3, -3, -3, -3, 0, 0, 1, 1, 4, 4, 4, 2, 1, 1, 0, 3, 3, 0, 2, 1, 0, 0, -1, -2, -1, -2, -3, -2, -5, -4, -3, -1, 0, 2, 1, 4, 4, 3, 1, 1, 1, 2, 3, 2, 2, 2, 0, 0, 0, -1, -2, -3, -4, -3, -3, -4, -3, -2, -1, 0, 1, 1, 3, 1, 2, 3, 3, 3, 5, 2, 4, 3, 1, 0, 0, -1, -3, -4, -4, -4, -4, -3, -3, -1, -1, 0, 0, 2, 3, 3, 4, 2, 2, 3, 5, 2, 4, 3, 2, 1, -2, -1, -4, -3, -5, -3, -2, -2, -3, -2, -2, -1, 0, 1, 3, 3, 2, 3, 3, 3, 2, 2, 3, 3, 1, 0, 0, -1, -4, -3, -3, -4, -3, -2, -2, -2, -1, -1, 1, 3, 2, 2, 0, 1, 2, 2, 1, 1, 2, 3, 2, 0, -1, -1, -2, -1, -1, -2, -1, -2, -1, -1, 0, 0, 1, 1, 2, 2, 0, 1, 2, 1, 2, 1, 1, 3, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, 3, 2, 3, 0, 1, 1, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 4, 4, 2, 0, 0, 0, 1, 0, 0, 3, 3, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 4, 4, 3, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 2, 3, 4, 3, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 3, 4, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 2, 1, 0, 1, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, -1, -1, 1, 1, 1, 2, 1, 0, 2, 2, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 2, 1, 2, 0, 1, 0, -2, -2, -2, 0, 0, 0, 0, 0, -1, -3, -2, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, -1, -3, -2, -3, -1, 1, 1, -4, -4, -2, -1, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -2, -3, -2, 0, -2, -1, -1, -1, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, 1, 1, 0, 1, -1, 0, 0, -1, -1, -3, 0, 0, 0, 0, -1, -1, 0, 0, -2, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -1, -2, -1, -2, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -3, -2, -2, -2, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, -1, 1, 0, 0, 0, 0, -2, -2, 0, -1, -3, -1, -3, -2, -1, -2, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -2, -4, -3, -2, -1, -3, -1, -1, 0, -2, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, -3, -2, -1, -2, -3, -3, -4, -4, -1, -1, -2, -1, -1, -1, -2, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, -2, -2, -1, -3, -2, -3, -2, -2, -3, -3, -3, -1, -3, -1, -3, -1, 0, 0, 0, -1, -2, -2, 1, 1, 1, 0, 0, 0, -3, -1, -3, -3, -3, -1, -2, -1, -2, -1, -2, -1, -1, 0, -1, 0, -1, 0, -1, 0, 1, 0, 1, 1, 0, 0, -2, -3, -3, -2, -3, -1, -1, -1, -2, -1, -2, -2, -1, 0, -1, 0, -1, 0, -2, 0, 0, 2, 1, 1, 0, 0, -1, -1, -2, -2, -3, -1, -2, 0, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 1, 2, 1, 0, 0, -1, -1, -1, -1, -1, -2, -2, 0, -1, -2, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 2, 1, 2, 1, 0, -1, 0, -1, -3, -1, -2, -1, 0, -1, -1, 0, -1, 0, 0, 1, 0, 1, -1, -1, -2, 0, 1, 1, 2, 0, 0, -1, 0, -2, -1, -1, -1, -2, 0, -2, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 2, 0, 0, 0, 0, -2, -1, -2, -2, -1, -2, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, -1, 0, -3, 0, 1, 2, 0, 0, 0, 0, 0, -1, -3, -1, -2, -1, -2, 0, -1, 0, 0, -1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -3, -2, 0, 0, -1, 0, -1, -1, -1, -2, -2, 0, 0, -1, -1, -1, 0, 0, -1, 0, 1, 1, -1, 0, 0, 0, -4, -2, -1, 0, 0, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, -1, -1, -5, -4, -1, -1, 0, -1, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -2, -1,
    -- filter=0 channel=5
    -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, -2, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -2, 0, 1, 0, 0, 0, 0, -1, -1, -2, 0, -1, -1, -1, 0, 0, -1, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, -1, -2, 0, -1, -1, -1, 0, -1, -2, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -2, -1, -1, -1, 0, 0, -1, -2, -2, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, -1, -1, -2, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -2, 0, 0, -2, -2, -1, -1, -1, 0, 0, 0, 0, -1, 1, 1, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -2, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, -2, 0, 0, 0, -1, -1, 0, 0, 0, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, -1, -1, 0, 0, -2, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, -2, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -2, 0, -2, -1, -2, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, -1, -1, -1, 0, -1, -1, 0, -2, 0, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, -2, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, 0, -2, 0, 0, 0, -2, 0, -1, -2, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, 0, -1, 0, -2, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, -2, -1, 0, 0, 0, 0, -2, 0, 0, 0, 0, -1, 0, -1, -1, -1, -2, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, -1, -2, 0, -1, -1, 0, 0, -1, -1, -1, -2, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -2, -2, -2, -1, 0, 0, 1, -3, -2, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -4, -2, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, -3, -2, 0, 1, 2, 1, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, -2, -1, -1, 0, 0, 1, 2, 1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 1, 1, -2, -1, 0, 1, 1, 2, 1, 1, 0, 1, 0, 1, -1, 0, 0, 0, 1, 2, 1, 0, 1, 0, 1, 1, 1, 1, -1, 0, 1, 0, 1, 0, 0, 2, 0, 0, 1, 0, 1, 0, 0, 0, 1, 2, 2, 1, 1, 0, 1, 3, 2, 2, -2, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 2, 2, 1, 1, 1, 0, 0, 1, 1, 1, 3, 1, -1, 0, 2, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 2, 2, 2, 0, 1, 2, 2, 0, 2, 2, 0, 0, 1, 1, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 1, 0, 2, 1, 1, -1, 0, 0, 2, 0, 2, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, -2, 0, 0, 0, 2, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 1, -1, -1, -2, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 2, 1, 1, 2, 1, 0, 0, 1, 0, 0, 2, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 1, 2, 1, 1, 1, 0, 0, 1, 0, 0, 2, 0, 1, 1, 1, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 2, 1, 1, 2, 1, 1, -1, 1, 2, 1, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 2, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 1, -2, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 1, 0, -2, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 2, 0, 0, 2, 0, 0, -2, -2, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 0, 1, 1, 0, 0, -1, -2, -3, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, 0, 0, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, -2, -3, -2, 1, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -2, 1, 0, 0, 0, 0, 1, 1, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 2, 1, 2, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -1, 2, 0, 0, 1, 0, 2, 0, 1, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -2, -1, 1, 1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, -1, 2, 0, 2, 2, 2, 1, 1, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, -1, -1, 0, 0, -1, -3, 1, 2, 0, 0, 2, 0, 2, 1, 0, 0, 2, 3, 1, 3, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 1, 1, 2, 0, 0, 0, 0, 0, 1, 0, 2, 2, 1, 1, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -2, 1, 1, 2, 1, 0, -1, 0, 0, 0, 1, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 1, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 1, 0, 0, 1, 0, 1, 1, 0, 1, 1, 1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, -2, -1, -2, 0, 0, 1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 1, 0, 0, -1, -1, 0, -2, -1, 0, -3, -2, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 4, 2, 1, 0, 0, 1, 1, 0, -1, -1, -2, 0, -1, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 2, 2, 0, 1, 2, 1, 1, 1, 2, 1, 0, 1, 1, 1, 2, 1, 0, 1, 0, 1, 1, 0, 0, 0, -3, 1, 0, 0, 1, 0, 1, 1, 3, 1, 2, 1, 0, 2, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -2, -1, 1, 2, 0, 0, -1, -1, 0, 2, 3, 2, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 3, 1, 2, 0, -1, -1, 0, 1, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 1, 0, 0, -1, -1, -2, -2, 2, 2, 1, 2, -1, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 2, 2, 2, 0, 0, 1, 0, 0, 0, 0, -1, 0, -2, 0, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, -2, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, 0, 0, 2, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 2, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 2, 1, 1, 1, 0, 1, 0, 2, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 1, 0, 1, 0, 2, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 2, 1, 2, 1, 1, 2, 2, 1, 1, 1, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 1, 0, 2, 2, 1, 0, 0, 1, 1, 2, 1, 1, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 2, 1, 1, 2, 0, 0, 1, 0, 1, 1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 2, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 2, 0, 0, 1, 0, 2, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 2, 1, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 2, 0, 1, 0, 1, 0, 2, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 2, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 1, 0, 2, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 2, 1, 0, 1, 0, -1, -1, 0, 1, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 1, 1, 1, 1, 2, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, -1, -1, -1, -1, -1, 0, 1, 0, 1, 2, 2, 1, 0, 1, 1, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 3, 2, 2, 2, 3, 2, 1, 1, 1, 0, 0, 0, 2, 0, 1, 1, 0, 0, 1, 0, 1, 0, -1, -1, 0, 0, 2, 2, 3, 2, 3, 2, 0, 1, 1, 0, 0, 1, 1, 1, 1, 0, 1, -1, 0, 1, 0, 0, 1, 0, 0, 0, 3, 3, 4, 2, 2, 1, 3, 1, 1, 0, 1, 2, 0, 1, 1, 0, 0, 0, 0, 1, 2, 1, 2, 0, 2, 2, 1, 3, 2, 2, 2, 2, 1, 2, 1, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 2, 2, 2, 1, 1, 1, 1, 1, 2, 1, 2, 2, 1, 2, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 2, 1, 0, 0, 0, 3, 2, 2, 1, 1, 2, 3, 3, 2, 1, 1, 0, 2, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 0, 0, 1, 3, 2, 2, 2, 3, 3, 2, 1, 2, 0, 1, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 2, 0, 2, 1, 4, 2, 3, 2, 2, 1, 3, 1, 1, 3, 2, 1, 0, 1, 1, 0, 1, 0, 1, 0, 1, 0, 1, 1, 1, 2, 3, 2, 2, 3, 1, 1, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 1, 2, 2, 1, 0, 0, 1, 3, 1, 3, 3, 1, 2, 2, 2, 2, 2, 1, 1, 1, 0, -1, -2, -1, -1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 1, 1, 0, 2, 2, 1, 2, 1, 0, 0, 0, 0, -1, -1, -2, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 1, 2, 1, 2, 2, 1, 2, 1, 2, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 2, 1, 3, 1, 2, 2, 1, 2, 2, 2, 2, 1, 1, 1, 1, 1, 0, 2, 0, 0, 0, 1, 2, 2, 1, 1, 2, 1, 2, 2, 2, 2, 2, 1, 3, 2, 1, 1, 0, 1, 1, 1, 3, 1, 2, 0, 0, 0, 1, 2, 2, 0, 1, 2, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 2, 0, 0, 1, 1, 2, 1, 2, 3, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 2, 0, 1, 1, 2, -1, 0, 1, 0, 1, 3, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 2, 0, 2, 0, 0, -1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 2, 0, 2, 1, 1, 1, 1, 1, 0, 2, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, -1, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, 1, 0, 0, 1, 1, 0, 1, 2, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 1, 1, 2, 0, 2, 1, 0, 0, 1, 1, 2, 0, 2, 1, 2, 1, 0, 0, 0, 0, -2, -1, -1, -1, -2, 0, 0, -1, -1, -1, -1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 2, 1, 2, 0, 0, -2, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 0, -1, -2, 0, -2, 0, -2, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 2, 1, 0, 0, -1, -2, -1, -3, -1, -2, -2, -3, -3, -1, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, -3, -2, -3, -3, -3, -4, -3, -3, -2, -2, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, -2, -1, -4, -4, -5, -4, -4, -3, -1, -1, -1, -2, -1, 0, 0, -1, 1, 1, 0, -1, 1, 1, 2, 0, 0, 0, -1, -3, -3, -5, -3, -3, -4, -3, -1, -2, -1, -1, 0, 0, 0, 1, 2, 2, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -2, -4, -5, -4, -2, -3, -1, 0, -1, 0, 0, 0, 1, 0, 1, 1, -1, 0, 0, 1, 0, 0, 1, 0, -1, -1, -2, -3, -4, -2, -3, -1, 0, -1, 0, 0, -1, 0, 1, 2, 2, 2, -2, -2, -1, 0, 0, 1, 0, 0, 0, -1, -2, -1, -1, -2, -3, -1, 0, -1, -1, 0, 0, 0, 0, 1, 2, 3, -1, -2, -1, 0, 0, 0, 1, 0, 0, -1, -2, -1, -2, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 2, 1, 1, -2, -2, -1, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 2, 1, 0, 1, 1, 1, 3, -3, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 0, 2, 1, 0, 2, 2, 3, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 2, 1, 2, 0, 2, 0, 1, 2, 2, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 2, 1, 0, 1, 1, 1, 0, -1, -1, -1, -1, 0, 1, 0, 0, 2, 2, 1, -1, -1, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, 0, 2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -2, 0, -2, -2, -1, -2, -1, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -2, -1, -1, -3, -1, -2, -2, -2, -2, 0, -1, 0, 0, 1, -1, -3, -1, -2, 0, -1, 0, 0, -2, -2, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -3, -5, -4, -6, -8, -10, 0, -1, -2, 0, 0, 0, -1, -1, 0, -1, 0, 1, 0, 0, 2, 0, 1, 0, 0, 0, -1, -2, -4, -4, -5, -7, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, -3, -5, -5, 2, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -2, -3, -6, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -3, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, -2, -2, 3, 3, 2, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 1, 1, -1, 0, -1, 0, -1, -1, -2, 0, 1, -1, -2, 5, 3, 1, 0, -1, -1, -1, -2, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 2, -1, 3, 3, 4, 2, 0, -1, -2, -3, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 6, 5, 3, 3, 1, -1, -4, -5, -4, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 7, 4, 5, 5, 2, -2, -4, -4, -4, -3, -1, 0, 0, 1, 0, -2, -1, 0, 1, 2, 2, 1, 1, 0, 1, 1, 7, 7, 6, 3, 3, 1, -1, -3, -4, -4, -1, 0, 0, -1, 0, -2, -3, -1, 0, 1, 0, 1, 0, 2, 2, 0, 8, 7, 6, 5, 3, 0, 0, 0, -3, -3, -2, -1, 0, 0, -2, -1, -1, -2, -1, -1, 0, 0, -1, 0, 0, -1, 9, 8, 6, 3, 2, -1, 0, 0, -2, -4, -2, -2, -1, -2, -2, -3, -2, -3, -1, -1, 0, -1, -1, 0, -1, -2, 7, 5, 4, 4, 1, 0, 0, -2, -3, -3, -3, -1, -1, -1, -2, -2, -2, 0, 0, 0, 0, -1, 0, 1, 0, -2, 6, 4, 4, 3, 4, 0, 0, -1, -3, -2, -3, -2, -1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, -2, 3, 5, 3, 2, 1, 2, 0, -2, -3, -2, -3, -3, -1, 0, 2, 1, 0, 0, 0, -1, 0, 1, 2, 1, 1, -1, 4, 2, 3, 3, 3, 2, 0, -2, -2, -1, -3, -2, -1, 0, 2, 0, 0, 0, -1, 0, 0, 1, 1, 2, 2, 0, 2, 3, 3, 3, 3, 0, 0, -2, -2, -2, -1, -2, 0, 0, 1, 2, 1, 0, 0, -1, 0, 0, 0, 2, 1, 0, 2, 1, 3, 2, 3, 2, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 0, 0, -1, 0, 0, 1, 0, -1, 0, 2, 3, 3, 1, 1, 0, 0, 1, 1, 1, 1, 1, 1, 3, 2, 0, 0, 2, 3, 2, 2, 2, 1, 0, -2, 0, 2, 4, 3, 0, 0, 0, 1, 0, 2, 2, 1, 1, 1, 2, 2, 0, 1, 2, 3, 3, 2, 0, 0, -1, -1, -1, 1, 2, 3, 1, 0, 0, 1, 0, 2, 2, 1, 1, 3, 2, 1, 1, 1, 1, 3, 4, 3, 0, 0, -1, -1, -1, 0, 4, 2, 1, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 1, 0, 1, 3, 3, 4, 1, 0, 0, -1, 0, 0, 1, 3, 2, 1, 1, 1, 1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 2, 3, 1, 2, 2, 0, -3, -7, -4, -3, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -3, -3, -2, -3, -1, -2, -1, -6, -4, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -2, 0, -1, -1, -5, -4, -2, -1, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, -1, -5, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, 1, 2, 1, 1, 1, 2, 1, 2, 2, 0, -5, -1, -1, 1, 1, 1, 2, 0, 2, 1, 0, 1, 0, 0, 0, 1, 1, 2, 1, 1, 1, 1, 2, 1, 2, 0, -3, -1, 0, 0, 0, 0, 1, 1, 1, 3, 4, 1, 0, 1, 0, 1, 1, 1, 3, 3, 1, 2, 3, 3, 3, 2, -2, 0, 1, 0, 0, 2, 2, 1, 2, 3, 4, 4, 2, 2, 3, 1, 3, 3, 2, 0, 0, 0, 1, 1, 3, 2, -4, -1, 2, 2, 0, 1, 1, 0, 2, 2, 3, 2, 2, 2, 4, 2, 2, 2, 2, 1, 1, 1, 1, 0, 1, 0, -2, 0, 1, 2, 1, 2, 0, 0, 2, 0, 1, 1, 1, 1, 2, 4, 3, 0, 1, 0, 0, 1, 0, 1, 0, 1, -3, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 2, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 1, 1, 1, 0, 0, 0, 0, 0, 2, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 1, 2, 1, -1, 0, -1, -2, -2, -2, -1, -1, 0, 0, 0, 0, -1, -1, 0, 2, 2, 2, 0, 1, 0, 1, 0, 1, 3, 0, 0, 1, 0, -1, -3, -1, -2, -3, 0, 0, 1, 0, 0, 0, 3, 4, 2, 2, 0, 0, 0, 0, 1, 1, 2, 1, 1, 0, 1, 0, 0, -2, -2, -2, -1, 0, 0, 0, 1, 2, 2, 4, 4, 3, 2, 2, 1, 0, 1, 0, 0, 0, 0, 1, 2, 2, -1, -2, -2, -2, 1, 1, 0, 0, 1, 2, 4, 5, 5, 4, 3, 2, 1, 2, 0, 1, 0, -1, 0, 1, 2, 0, 0, -1, -1, 0, 0, 1, 0, 0, 1, 2, 4, 4, 5, 2, 1, 1, 1, 1, 1, 0, -1, -1, 0, 0, 0, 1, 0, -2, -1, -1, 1, 1, 1, 2, 1, 2, 3, 5, 5, 4, 3, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 1, 1, 2, 3, 3, 2, 4, 5, 6, 4, 3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, -2, -1, 0, 3, 3, 4, 4, 3, 2, 4, 4, 4, 2, 2, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, -3, 1, 2, 2, 2, 3, 2, 1, 1, 3, 4, 2, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 1, 0, -4, 0, 1, 3, 4, 3, 2, 1, 1, 2, 2, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, -4, -1, 1, 2, 4, 4, 2, 2, 2, 0, 2, 2, 1, 2, 0, 1, 0, 1, 2, 2, 4, 3, 2, 2, 0, 0, -5, -3, 0, 2, 1, 2, 3, 1, 2, 1, 1, 2, 2, 0, 0, 1, 1, 1, 2, 2, 3, 2, 2, 1, -1, -1, -6, -4, -1, 0, 0, 1, 2, 3, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, -1, -2, 0, -7, -5, -3, -1, -2, 0, 0, 0, 2, 1, 1, 0, 0, 0, -1, -2, 0, 0, -1, 0, -1, 0, -2, -1, -2, -1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 1, 2, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 1, 0, 0, 1, 2, 2, 0, 1, 1, 0, -1, 1, 1, 1, 1, 1, 0, 0, -1, -1, -1, 0, -1, 1, 0, 0, 0, 0, 0, 1, 2, 2, 2, 1, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, -1, 0, 0, -1, 0, 0, 1, 2, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 1, 0, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, -12, -9, -6, -5, -5, -4, -2, -1, -2, 0, -2, 0, -1, -2, -3, -2, -2, -3, -5, -6, -6, -8, -5, -4, -5, -5, -9, -6, -5, -3, -2, -2, 0, -1, -2, -2, -1, -1, -1, 0, -2, -2, -1, 0, -2, -4, -5, -3, -3, -2, -3, -4, -9, -6, -3, 0, 1, 0, 0, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, -2, -1, -2, -1, -1, -1, -2, -7, -3, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 1, 2, 1, 2, -1, -7, -3, 0, 2, 1, 3, 2, 2, 2, 1, 1, 2, 0, 1, 2, 2, 1, 1, 1, 0, 0, 2, 3, 3, 4, 0, -6, -1, 0, 0, 3, 3, 3, 4, 3, 4, 4, 3, 2, 1, 2, 2, 2, 2, 3, 3, 1, 3, 3, 5, 4, 2, -5, 0, 1, 1, 3, 3, 2, 4, 4, 3, 4, 2, 3, 1, 1, 3, 3, 2, 2, 2, 3, 3, 4, 5, 5, 2, -3, 0, 2, 3, 2, 4, 4, 2, 3, 2, 4, 2, 1, 2, 4, 4, 2, 4, 1, 3, 1, 3, 3, 4, 4, 3, -4, 0, 4, 5, 3, 3, 4, 1, 2, 1, 1, 3, 2, 3, 4, 4, 2, 2, 1, 1, 3, 0, 2, 3, 2, 1, -2, 3, 4, 4, 5, 3, 2, 0, 1, 1, 0, 0, 2, 3, 4, 3, 4, 3, 1, 2, 1, 1, 2, 2, 1, 1, 0, 3, 5, 5, 4, 2, 3, 0, 0, 0, 1, 0, 0, 1, 3, 2, 2, 2, 1, 1, 0, 0, 0, 1, 1, 1, 1, 4, 5, 3, 4, 2, 2, 0, 0, 0, 0, 0, 0, 1, 1, 2, 3, 3, 0, 0, 0, 1, 0, 0, 0, -1, 0, 3, 3, 3, 3, 1, 2, 1, 1, 1, 1, 0, 0, 0, 2, 2, 4, 2, 1, 0, 0, 1, 0, -1, 0, -1, 0, 1, 4, 4, 4, 1, 2, 4, 3, 2, 3, 0, 0, 0, 1, 2, 1, 1, 1, 2, 3, 1, 0, -1, -2, -2, -2, 3, 4, 4, 5, 3, 5, 4, 4, 3, 2, 1, 0, 1, 2, 3, 1, 1, 1, 3, 4, 1, 2, 0, -2, -2, -2, 3, 4, 3, 3, 5, 4, 5, 4, 5, 2, 2, 2, 1, 1, 2, 1, 0, 0, 1, 3, 4, 2, 1, 0, -1, 0, 3, 2, 5, 4, 4, 5, 5, 5, 4, 2, 1, 2, 1, 1, 1, 2, 0, 0, 1, 1, 3, 3, 1, 1, 0, 0, 2, 4, 2, 3, 4, 5, 4, 5, 5, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 3, 1, 1, 0, 0, 1, 5, 4, 6, 4, 5, 5, 5, 5, 3, 2, 0, 0, 0, 1, 0, 0, 0, 2, 1, 1, 1, 0, 0, -1, -2, 0, 4, 3, 5, 5, 3, 5, 4, 5, 5, 2, 1, 0, 1, 1, 1, 0, 0, 0, 0, 2, 2, 1, 0, -1, -5, -1, 1, 3, 2, 4, 3, 3, 3, 2, 4, 2, 2, 2, 0, 2, 0, 0, 1, 0, 0, 0, 0, 2, 0, 0, -5, -2, 0, 1, 3, 3, 3, 1, 1, 2, 2, 2, 0, 1, 1, 1, 1, 1, 1, 1, 0, 2, 2, 1, 0, -1, -9, -4, -1, 1, 1, 2, 0, 0, 0, 0, 1, 2, 1, 0, 2, 1, 1, 0, 2, 2, 4, 4, 3, 1, 0, -2, -11, -6, -3, -1, 2, 1, 2, 0, 0, 0, 0, 2, 2, 0, 0, 1, 1, 2, 3, 2, 3, 3, 2, 1, -1, -3, -12, -8, -4, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 3, 2, 0, -1, -3, -13, -10, -7, -4, -3, -3, -1, 0, -1, -1, 0, 0, -1, -1, -3, -2, -1, -2, 0, 0, 0, 0, -2, -2, -5, -3, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 3, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 1, 1, 2, 1, 1, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 3, 1, 3, 1, 2, 0, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 3, 2, 2, 3, 2, 2, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 2, 1, 0, 0, 2, 2, 3, 3, 3, 3, 1, 2, 1, 1, 2, 0, 1, 0, 1, 1, 2, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 1, 1, 3, 4, 2, 1, 3, 3, 2, 2, 2, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 1, 3, 1, 3, 3, 3, 3, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 1, 1, 1, 2, 3, 2, 3, 1, 1, 1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 1, 1, 2, 2, 2, 2, 1, 0, 2, 1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 2, 0, 1, 1, 0, 0, 0, -1, 0, 1, 1, 0, -1, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 2, 2, 2, 0, 2, 1, 1, -1, -1, 0, -1, -1, 0, 0, -1, -2, 0, 0, 0, -2, -1, 0, 0, 0, 0, 2, 2, 2, 3, 1, 2, 2, 2, 0, 0, -1, -1, 0, 0, 0, 0, -2, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, 2, 3, 2, 2, 2, 1, 1, 1, 0, 0, 0, 1, 0, 0, -2, -2, 0, 0, -2, -1, -1, -1, 0, -2, 0, 1, 2, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, 0, -1, -1, 0, -1, 0, 2, 1, 1, 1, 3, 1, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -1, -2, -1, -1, 1, 1, 0, 1, 1, 0, 0, 2, 1, 2, 1, 1, 0, -1, -1, 0, 1, 0, 0, 0, 0, -2, -1, -1, -2, -1, 1, 1, 1, 1, 0, 1, 2, 3, 3, 3, 2, 1, 0, -1, 0, 0, -1, 0, 1, 1, -1, -1, -1, 0, -1, -1, 1, 0, 0, 0, 2, 2, 1, 1, 2, 2, 3, 1, 1, 1, -1, 0, 0, 0, 1, 1, 1, 0, -1, -1, 0, -1, 0, 1, 0, 0, 1, 1, 3, 2, 3, 3, 2, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -3, 0, -1, 1, 2, 2, 1, 0, 0, 2, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -3, -2, 0, 1, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -2, -2, -1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 3, 2, 0, 0, 0, 0, 2, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 2, 1, 2, 2, 1, 1, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -4, -4, -2, -1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -5, -3, -2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 1, 0, 1, 0, 0, -1, -5, -1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 2, 2, 1, 2, 2, 1, 0, -3, -3, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 2, 3, 2, 1, 2, 2, -3, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 2, 1, 0, 1, 0, 1, 2, 3, 3, -2, -2, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 1, 0, 1, 1, 2, 2, 2, -2, 0, 1, 2, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 2, 2, 1, -2, -1, 0, 3, 2, 0, 0, -1, -2, -1, 0, 0, 0, 0, 1, 0, 1, 0, 2, 1, 2, 2, 2, 2, 1, 2, 0, 1, 2, 3, 2, 2, -1, -2, -2, -1, 0, -1, -1, 0, 1, 0, 2, 0, 0, 0, 0, 2, 2, 0, 1, 2, 0, 1, 3, 3, 1, 0, -1, -2, -2, -3, -3, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 2, 1, 2, 2, 0, 2, 3, 3, 2, 0, 0, 0, -1, -1, -2, -2, 0, 0, 0, 2, 2, 0, 0, 2, 0, 1, 1, 1, 2, 0, 1, 1, 2, 1, 2, 1, 1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, 3, 2, 2, 2, 0, 1, 0, 0, 0, -1, -1, 0, -1, 1, 0, 0, 1, 0, 1, 0, 0, 2, 1, 1, 0, 1, 1, 3, 3, 3, 2, 1, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 3, 2, 1, 0, 0, 0, 2, 3, 4, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 1, 2, 2, 0, -1, -1, 2, 3, 3, 2, 2, 1, 1, 0, 0, -1, 0, 0, 0, 2, 1, 0, 1, 0, 0, 0, 2, 2, 2, 1, 0, -1, 1, 3, 1, 2, 2, 1, 0, 1, 0, -1, 0, 0, -1, 0, 1, 2, 1, 0, -1, 1, 0, 0, 1, 1, 1, -1, 1, 2, 3, 2, 3, 2, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, 0, 0, 2, 2, 3, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, -3, -2, 0, 2, 0, 1, 0, 1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, -4, -2, 0, 1, 2, 1, 2, 0, 0, 0, 0, 0, 2, 0, 0, 1, 1, 0, 2, 0, 2, 0, 1, 1, 0, 0, -4, -2, 0, 2, 2, 2, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 2, 1, 3, 3, 1, 0, 0, -5, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 1, 0, 3, 3, 3, 2, 1, -1, -5, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, -6, -4, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, -6, -4, -4, -1, -3, -1, 0, -1, 0, 0, -1, 0, -1, 0, -1, -1, 0, -1, -2, -1, 0, -1, -2, -1, -3, -2, -7, -4, -4, -1, -2, -1, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -3, -3, -3, -6, -3, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, -2, 0, -6, -2, -3, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -5, -3, -1, -1, -1, 0, 1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, 1, 1, 1, -3, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 2, 0, -4, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -3, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 2, 1, 2, -2, 0, 0, 1, 0, 1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 2, 0, 1, 1, 0, 0, 0, 2, 1, 2, -4, 0, 1, 1, 1, 0, 0, 0, -1, -1, -2, 0, -2, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 2, -2, 0, 2, 2, 1, 0, -1, 0, -1, -1, -3, -2, -1, 0, 0, 1, 1, 1, 1, 2, 0, 0, 1, 2, 1, 2, -1, 1, 3, 3, 2, 0, -2, -2, -1, -2, -1, -1, 0, 0, 0, 1, 0, 1, 3, 1, 0, 0, 0, 0, 1, 1, 0, 0, 2, 1, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 2, 1, 0, 1, 1, 1, 1, 2, 0, 1, 1, 3, 0, 1, 0, -1, -1, -2, -1, -3, -2, -2, 0, 0, 1, 0, 1, 2, 3, 2, 2, 1, 0, 0, 0, 1, 3, 3, 1, 0, 0, -1, -2, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 3, 2, 1, 0, 0, 1, 2, 3, 2, 1, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 3, 2, 1, 0, 1, 2, 3, 3, 2, 1, 0, -2, -1, 0, -1, -1, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 3, 0, 0, 0, 0, -1, 0, -2, -2, 0, 0, -1, 0, 0, -1, 0, -1, 1, 2, 1, 2, 0, 0, -1, 0, 3, 2, 0, 2, 1, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 1, 1, 2, 1, 0, -1, 1, 1, 3, 2, 1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, -2, 1, 0, 1, 2, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, -3, 0, 1, 2, 1, 3, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -3, -1, 0, 1, 2, 3, 2, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 0, -4, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 2, 2, 2, 2, 0, 1, 2, 3, 3, 2, 1, 1, -1, -3, -2, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 1, 0, 3, 3, 2, 2, 1, 0, 1, -3, -3, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 2, 1, 2, 0, 2, 3, 2, 2, 2, 0, -1, -1, -3, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 1, 0, 3, 3, 1, 2, 0, 0, -1, -4, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 1, 2, 1, 2, 3, 0, 1, 0, 0, 0, 3, 3, 2, -4, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 1, 1, 0, 1, 0, 2, 3, 2, 1, -5, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 2, 0, 0, 0, 1, 2, 2, 2, 2, 2, -3, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 2, 1, 1, 3, 3, 1, -6, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 0, 2, 1, 2, 2, 3, 1, -6, -3, -1, 0, -1, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 1, 2, 1, 1, 1, 3, -5, -3, -2, 0, 0, 1, 1, 1, 1, 1, 0, 1, 0, 1, 2, 2, 2, 2, 0, 0, 0, 1, 1, 3, 1, 2, -3, -2, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 1, -3, -3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, -1, -1, 0, 0, 0, 1, 0, -2, -1, 0, -1, 0, -1, -2, 0, -1, 0, -1, -1, -1, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 1, 0, 0, -4, -2, 0, -1, -1, -1, -3, -1, 0, -1, -3, -1, -1, -1, 0, 0, 2, 1, 0, -2, 0, 0, 0, 0, 0, 0, -4, -1, 0, -1, 0, -3, -1, -2, 0, -1, -2, -1, -2, -2, 0, 1, 0, 2, 0, 0, -1, 0, 0, -2, -1, -1, -3, -2, 0, 0, 0, -1, -2, 0, 0, 0, -2, 0, -1, -1, 0, 1, 0, 1, 0, 0, 1, 0, -1, -2, -1, -1, -2, 0, -1, -1, -1, 0, -1, 0, 1, 0, 0, -1, 0, -1, 0, -1, 1, 0, 0, 0, 2, 0, 0, -1, 0, 0, -2, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, -1, 0, -2, -2, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, -1, -2, -2, 0, -2, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, 1, 2, 1, 2, 0, -2, -1, -2, -3, -3, -1, -1, -1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 1, 1, 2, 0, 1, 2, 1, 1, 0, -1, -1, -3, -2, -2, -3, -1, -1, 0, 0, 1, 1, 0, 0, -1, -1, 0, 1, 1, 0, 0, 1, 0, 1, 2, 0, 0, -1, -2, -1, -2, -1, -2, -1, 0, 0, 0, 0, 1, 0, 0, -2, -1, 1, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, -1, -1, 0, -1, -2, -2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -2, -1, 0, 0, 0, 1, 1, 3, 3, 2, -2, 0, 1, 3, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 3, 2, 3, 1, 2, 2, -3, -1, 1, 1, 2, 1, 1, 2, 2, 1, 1, 1, 1, 0, 0, 0, 2, 0, 1, 2, 2, 3, 2, 2, 1, 2, -3, -2, 1, 0, 1, 2, 0, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 1, 2, 3, 1, 2, 1, 0, 1, 0, -2, 0, 0, 1, 0, 1, 2, 1, 1, 1, 1, 0, 1, 1, 0, -1, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 2, 2, 2, 0, 2, 0, -1, 0, -2, -1, -2, 0, 0, -1, -1, 0, 0, -1, 0, -9, -8, -7, -5, -5, -4, -5, -5, -4, -4, -4, -3, -4, -3, -2, -3, -4, -4, -3, -6, -4, -5, -5, -4, -6, -6, -9, -7, -3, -3, -3, -3, -2, -2, -3, -3, -3, -2, -2, -2, -1, -1, -2, -2, -1, -1, -2, -1, -2, -4, -3, -5, -6, -4, -2, -2, -2, -1, -2, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -3, -6, -3, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 2, 0, 0, 0, -5, -4, -2, -2, 0, 0, 0, 1, 0, 0, 1, 0, 2, 2, 1, 0, 2, 2, 2, 2, 2, 2, 1, 1, 1, 0, -4, -3, -1, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 1, 2, 2, 2, 1, 2, 0, 0, 1, 2, 3, 3, 1, -5, -2, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 2, 1, 2, 1, 1, 1, 1, 1, 1, 3, 2, 3, -2, 0, 2, 2, 2, 1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 2, 3, 2, 1, 1, 1, 1, 1, 4, 4, 2, 0, 1, 3, 3, 3, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 2, 2, 4, 4, 1, 1, 1, 2, 2, 3, 1, 0, 4, 5, 6, 4, 2, 0, -2, -3, 0, -1, -1, 0, 0, 0, 2, 2, 2, 3, 1, 2, 2, 2, 2, 2, 0, 1, 5, 6, 5, 3, 1, 1, 0, -2, -2, -2, 0, 0, 1, 2, 2, 0, 3, 2, 1, 2, 2, 2, 2, 1, 1, 1, 4, 5, 5, 4, 1, 1, 0, -1, 0, -2, -2, -1, 0, 0, 0, 2, 0, 2, 0, 1, 2, 2, 0, 2, 1, 1, 4, 5, 5, 4, 2, 1, 1, -1, -1, 0, -1, -2, -1, 0, 1, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 2, 4, 5, 6, 4, 4, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 2, 1, 0, 0, 1, 3, 4, 4, 3, 2, 2, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 2, 3, 3, 1, 0, -1, 1, 2, 4, 4, 3, 2, 1, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 2, 2, 3, 3, 1, 0, 0, 3, 3, 3, 4, 3, 3, 0, 0, 0, -2, -1, -2, -1, -1, 0, 0, 0, 1, 1, 2, 3, 1, 3, 2, 0, -1, 3, 2, 3, 4, 1, 2, 1, 0, 1, -1, -1, -2, -1, 0, 0, 1, 1, 1, 1, 0, 1, 2, 2, 1, 0, -3, 0, 2, 4, 4, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, -4, -1, 0, 2, 4, 2, 2, 0, 0, -1, 1, 1, 0, 0, 2, 0, 2, 1, 1, 0, 0, 1, 2, 1, 1, 1, -6, -2, 0, 2, 1, 2, 0, 0, -1, 1, 0, 1, 1, 0, 0, 0, 2, 2, 2, 1, 1, 2, 1, 1, 0, 0, -7, -3, -1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 3, 3, 3, 4, 5, 2, 1, 0, 0, -7, -5, -2, -1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 2, 2, 1, 2, 3, 3, 5, 4, 3, 0, 0, -2, -8, -5, -3, -3, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 3, 2, 2, 0, 0, -1, -2, -9, -7, -5, -3, -3, -3, -2, -1, 0, -1, -2, -1, -2, -1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, -2, -9, -9, -6, -4, -5, -4, -3, -1, -3, -1, -3, -2, -2, -3, -4, -2, -4, -2, -2, -3, -4, -4, -3, -5, -3, -5, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 2, 2, 2, 0, 1, 0, 0, 0, 0, 1, 3, 4, 3, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 1, 0, 0, 0, 2, 3, 3, 2, 3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 2, 2, 1, 3, 2, -1, -2, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 2, 1, 2, 1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 3, 2, -3, -1, -1, 0, 0, 1, 0, 0, 1, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, -1, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 3, 1, 1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, -1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, -1, 0, -1, -1, 0, -1, -2, -1, 0, -1, 1, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, -1, 1, 0, 0, 0, -1, 0, 0, -1, -1, -1, -2, -1, -1, -1, 0, 0, 1, 1, 0, -1, 0, -1, 0, 1, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, -1, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 2, 1, 0, 1, 0, 0, 0, -1, 0, -1, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 2, 1, 1, 0, 0, -1, -3, -2, -1, -1, -1, -1, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 2, 3, 2, 1, 1, 2, 0, 0, 0, -2, -3, -1, 0, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 2, 1, 1, 0, 0, 0, -2, -1, -2, -2, -3, -2, 0, 0, -2, 0, 0, -1, 0, 1, 0, 0, 0, 2, 2, 1, 2, 0, 1, 0, -1, 0, 0, 0, -2, -3, -1, 0, -1, 0, -1, -1, -1, 1, 1, 1, 1, 3, 0, 1, 2, 2, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 1, 1, 2, 3, 3, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 2, 2, 2, 1, 3, 3, 0, 1, 2, 0, 0, 1, 0, 1, 0, 0, 0, 0, 2, 0, 1, 0, 2, 0, 0, 1, 4, 1, 1, 1, 2, 1, 0, 0, 1, 0, 1, 0, 1, 0, 1, 1, 1, 2, 1, 2, 0, 2, 1, 2, 2, 4, 2, 2, 3, 1, 2, 1, 0, 1, 2, 1, 0, 0, 1, 0, 0, 3, 2, 2, 2, 2, 2, 3, 1, 2, 3, 2, 3, 3, 2, 1, 2, 2, 0, 0, 2, 0, 1, 3, 2, 1, 3, 3, 2, 2, 1, 2, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 1, -9, -7, -3, -4, -3, -1, -1, -1, -1, -1, -2, -2, -2, -2, -1, 0, -1, -1, 0, -2, -4, -3, -2, -4, -2, -4, -7, -4, -3, -3, -1, 0, -1, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, -2, 0, 0, -3, -7, -5, -1, -2, -2, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, -7, -3, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 2, 0, -6, -2, -1, -2, -1, -1, -1, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 1, 2, 2, 0, 1, -5, -3, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 2, 0, 2, 1, 1, -4, -1, 0, 0, 1, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 3, 1, 1, 0, 2, 2, 0, 1, 3, 1, -5, 0, 0, 1, 1, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 1, 1, 2, 1, 1, 2, 1, 2, 1, 3, 1, -3, 1, 2, 2, 2, 1, -1, -2, -2, -1, -1, -2, 0, 0, 1, 1, 1, 2, 2, 1, 2, 0, 0, 2, 1, 2, -1, 0, 1, 3, 2, 0, 0, 0, -2, -1, -1, 0, -1, 0, 0, 2, 0, 2, 1, 2, 0, 0, 0, 1, 0, 0, -2, 2, 3, 2, 1, 0, -1, 0, -1, -2, 0, -2, -1, 0, 1, 2, 3, 2, 1, 2, 1, 1, 1, 0, 1, 0, -2, 2, 3, 3, 1, 2, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, 2, 2, 1, 2, 2, 2, 2, 1, 0, -1, -1, 0, 3, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 2, 1, 0, 0, -1, -1, 0, 2, 2, 4, 1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 2, 0, 0, 1, 1, 1, 1, 1, 1, 0, -1, -1, 2, 3, 4, 3, 0, 1, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 2, 3, 2, 0, -1, 0, 2, 2, 2, 2, 1, 1, 0, 1, 0, 0, -2, 0, -1, 0, 1, 1, 1, 0, 0, 1, 2, 2, 1, 0, -1, 0, 1, 2, 4, 3, 1, 0, 0, 1, 0, 0, 0, -2, -1, -1, 0, 2, 2, 1, 1, 2, 0, 2, 2, 0, 0, -3, 0, 3, 3, 2, 3, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 2, 0, 0, -3, 0, 1, 1, 3, 2, 2, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -3, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6, -3, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 2, 1, 2, 2, 1, 1, 2, 1, 0, -2, -7, -4, -2, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 2, 1, 2, 2, 1, 0, 1, 1, 3, 2, 1, 0, 0, -6, -3, -4, -2, 0, 0, 1, 1, 0, 0, -1, 0, 1, 1, 2, 1, 2, 1, 1, 1, 1, 3, 1, 1, 0, -2, -8, -5, -4, -1, -2, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, -8, -7, -4, -3, -3, -1, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, -2, -2, 0, -2, -2, -3, -10, -7, -6, -6, -5, -3, -2, -3, -2, -2, -3, -2, -3, -2, -3, -1, -2, -3, -3, -4, -3, -4, -3, -5, -4, -5, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 1, 0, 0, -1, 0, 1, 0, -1, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, -1, 0, -1, -1, 1, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 1, 1, 0, 0, 0, -1, 1, 0, 0, 1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 1, 0, 0, 0, 1, 0, -1, 1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, -1, -2, -1, -2, -3, -3, -2, -2, -1, -2, -1, -1, -1, -1, -1, -2, -2, -1, -2, -2, -2, -4, -3, -1, -1, -2, 0, 0, -2, -2, 0, -2, -1, -1, -2, -1, -1, -2, -1, -2, -1, -1, -1, 0, -1, -1, -1, 0, -1, -2, -1, -1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, 0, 0, -1, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 2, 2, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 2, 2, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 1, 2, 1, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 0, 2, 2, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 2, 2, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 2, 2, 1, 3, 2, 2, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 3, 1, 3, 2, 1, 1, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, -2, -1, 0, -1, 0, 0, 0, 0, 2, 1, 2, 2, 1, 1, 1, 0, 0, 1, -1, -1, 0, 0, -2, -1, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 2, 1, 2, 1, 2, 1, 2, 1, 0, -1, 0, 0, -1, -1, -1, -3, -1, -1, -1, -2, -1, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 1, 1, 1, 0, 1, -1, 0, 0, 0, 0, -1, -1, -2, -1, 0, -1, 0, 1, 1, 0, 2, 2, 1, 0, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, 1, 1, 1, 2, 1, 1, 1, 0, 1, 2, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 2, 3, 2, 2, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 1, 0, 0, 0, 1, 0, 1, 1, 1, 2, 1, 0, 0, 0, 1, 1, 1, 1, 0, 1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 1, 0, 2, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 0, 1, 0, 0, 0, 0, 1, 0, 2, 2, 0, 0, 1, 0, 1, 0, 0, 1, 1, 1, 0, 0, 1, 1, 2, 0, 1, 1, 0, 0, 0, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 2, 1, 0, 0, 0, -1, -1, 1, 0, 0, 0, 1, 1, 0, 2, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 2, 1, 1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 2, 1, 1, 0, -1, 0, 0, 0, 0, 0, -2, 0, 0, -1, -3, -5, -3, -2, -3, -3, -2, -3, -3, -3, -2, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, -1, -1, 0, -2, 0, -2, -1, -2, -2, -1, -2, -1, 0, -2, 0, 0, 0, 0, 0, 1, 1, 2, 3, 2, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -2, -3, -2, -1, -1, 0, 0, -1, 0, 1, 2, 4, 3, 5, 4, 2, 2, 0, 1, 0, -1, 0, 0, -1, 0, 0, -2, -2, 0, 1, 1, 0, 0, 0, 0, 1, 2, 4, 5, 5, 5, 2, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 1, 0, 0, -1, 0, 0, 1, 3, 6, 7, 6, 5, 5, 2, 2, 1, 1, 0, 1, 1, 0, -1, 0, -2, -1, 0, 2, 2, 1, 0, 1, 2, 2, 4, 7, 8, 6, 7, 3, 4, 3, 3, 1, 0, 0, -1, -2, -2, -2, -3, 0, 1, 2, 2, 0, 1, 3, 5, 1, 4, 6, 8, 8, 6, 4, 5, 4, 3, 1, 1, 0, -2, -2, -2, -3, -2, -1, 0, 0, 2, 2, 1, 2, 3, 1, 4, 6, 8, 8, 6, 7, 6, 3, 2, 2, 0, 0, -1, -1, 0, 0, -2, -2, -1, 1, 0, 0, 2, 3, 4, 2, 3, 5, 8, 7, 7, 5, 3, 4, 1, 0, 0, 0, 1, -1, -1, -2, -1, -1, -1, -1, -1, 0, 0, 2, 4, 2, 3, 7, 7, 9, 7, 5, 4, 3, 2, 0, 1, 0, 0, 0, -1, -2, -1, -2, -3, 0, 0, 0, -1, 3, 4, 3, 3, 6, 9, 11, 8, 8, 5, 2, 3, 2, 0, -1, -1, -3, -2, -1, -3, -2, -2, -1, 0, 0, 0, 2, 5, 2, 4, 4, 6, 9, 7, 7, 4, 3, 2, 3, 0, -1, -2, -1, -2, -2, -3, -5, -4, -3, -1, -2, 0, 2, 6, 0, 2, 1, 3, 7, 6, 4, 5, 3, 4, 3, 0, -2, -2, -2, -2, -2, -3, -5, -4, -4, -2, -1, 0, 4, 6, 0, 0, 1, 3, 5, 3, 4, 2, 3, 3, 3, 0, -1, -3, -4, -3, -1, -2, -2, -2, -1, -2, -1, 0, 3, 5, 0, 1, 2, 3, 3, 3, 2, 2, 2, 4, 1, 0, -1, -2, -2, 0, 0, 1, 1, 0, 0, -1, 0, 0, 3, 3, 2, 4, 3, 4, 3, 3, 1, 2, 2, 2, 1, 0, 0, -2, -1, -1, 0, 3, 3, 0, 0, 0, 1, 2, 3, 6, 2, 2, 3, 2, 2, 1, 3, 4, 4, 2, 1, 0, -1, -1, -3, -1, 0, 2, 1, 1, 1, 1, 1, 2, 4, 6, 0, 2, 2, 3, 1, 1, 3, 2, 1, 0, 0, 0, -1, -2, -3, -2, -1, 1, 1, 1, 0, 1, 2, 2, 1, 2, 0, 0, 1, 2, 2, 3, 3, 1, 2, 0, 0, -1, -2, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 0, 0, 0, 0, 0, 3, 3, 2, 0, -1, -1, -1, -2, -1, 0, 1, 1, 2, 0, 0, -2, -2, 0, 1, 2, 4, -1, -1, 0, -1, -1, 1, 1, -1, -2, -2, -3, -3, -1, 0, 1, 1, 1, 3, 0, 0, -1, -1, 0, 1, 3, 4, 0, 0, 0, -1, -1, -1, 0, 0, -2, -2, 0, -1, -1, 0, -1, 1, 1, 1, 0, -2, -3, -2, 0, 2, 2, 3, 0, 1, 1, -1, 0, 0, 1, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, -1, 0, -2, -2, -1, 0, 1, 1, 2, -1, 1, 0, 1, 0, 1, 3, 2, 0, 0, 0, 0, 0, -2, 0, -1, -1, -1, -2, -3, -1, 0, 1, 2, 3, 3, 0, 1, 1, 1, 3, 4, 2, 4, 2, 0, 1, 0, 0, 1, 1, 0, -1, -1, -1, 0, 0, 1, 3, 4, 3, 5, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -4, -2, -1, 0, 0, 0, 1, 0, 0, 2, 1, 0, 2, 1, 3, 1, 2, 2, 1, 1, -1, 0, 0, -1, 0, -1, -5, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, -4, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 2, 2, -3, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 1, 1, 1, -1, -1, 0, -1, 0, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, -1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -2, 0, -1, -1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, -1, 0, 1, 0, 0, -1, -1, -3, -1, -3, -2, -2, -2, -1, 0, 0, 1, 0, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, -2, -3, -3, -5, -3, -3, -3, -2, -1, 0, 0, 1, 1, 1, 1, 1, 0, 1, 1, 2, 2, 0, 0, 2, 2, 0, -2, -4, -3, -3, -2, -2, -3, -1, 0, 0, 0, 1, 1, 2, 3, 2, 1, 0, 0, 0, 1, 2, 1, 2, 0, 0, -1, -3, -3, -3, -3, -4, -2, -2, -1, -1, 0, 0, 1, 2, 2, 1, 0, 2, 1, 1, 0, 1, 3, 3, 0, 0, 0, -2, -4, -2, -4, -3, -3, -1, 0, 0, 0, 1, 2, 0, 1, 1, 1, 2, 1, 0, 0, 0, 2, 1, 3, 0, 0, -2, -2, -3, -2, -3, -2, -2, -2, 0, 0, -1, -1, 0, 0, 2, 2, 0, 0, 0, 0, 0, 3, 3, 2, 2, 0, -2, -2, -2, -3, -3, -2, -2, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, -2, 0, 3, 2, 2, 1, 1, -2, -2, -1, -2, -2, -3, -1, -1, 0, -1, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 1, 1, 2, 0, 1, 0, 0, -2, -1, -3, -3, -3, -1, 0, 0, 0, 0, 0, -2, 0, 0, 1, 2, 2, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, -2, 0, -3, -4, -1, -1, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, -1, 0, -2, -3, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 0, 2, 2, 0, 0, 0, -1, 0, -1, -1, -2, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 3, 1, 1, 1, 0, 1, 0, 1, 1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, -2, 0, 2, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, -1, 0, 1, 1, 1, 1, 0, 0, 0, 1, 2, 0, 0, 0, 0, 1, 1, 1, 0, 2, 3, 1, 1, 1, 0, 1, -1, 0, 2, 2, 1, 1, 1, 0, 0, 0, 1, 2, 2, 1, 3, 3, 2, 2, 2, 2, 3, 3, 2, 2, 1, 0, -2, 0, 1, 1, 0, 1, 0, 2, 0, 0, 2, 1, 3, 1, 1, 2, 3, 1, 2, 4, 4, 4, 3, 2, 0, 0, -1, -1, 0, 0, 1, 0, 0, 1, 0, 2, 2, 1, 1, 2, 3, 3, 2, 2, 2, 3, 4, 3, 2, 2, 0, -1, 1, 1, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 2, 3, 3, 3, 1, 2, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 2, 4, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 2, 1, 1, 0, 1, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 2, 1, 1, 3, 3, 0, 0, 2, 0, 1, 2, 1, 0, 1, 1, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 1, 2, 2, 0, 1, 1, 0, 0, 1, 2, 2, 0, 1, 1, 1, 0, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 2, 0, 1, 3, 0, 2, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 3, 0, 1, 1, 2, 1, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 1, 0, 1, 1, 1, 1, 0, 1, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, 1, 1, 1, 1, 2, 2, 0, 1, 0, 1, 0, 1, 1, 0, -1, -1, -2, -2, -2, -3, 0, -1, -2, -2, -1, 0, 0, 0, 0, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -3, -2, -1, -1, -2, -1, 0, -1, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, -1, -2, -2, -3, -3, -3, -4, -2, 0, -1, -2, -1, -1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, -3, -4, -4, -2, -2, -2, -2, -1, -2, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -3, -2, -4, -4, -4, -3, 0, 0, 0, -2, -1, 0, 0, 0, 2, 3, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, -2, -1, -4, -3, -3, -2, 0, 0, -1, -1, 0, -1, 0, 1, 2, 3, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, -2, -2, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, -3, -3, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 2, 1, 0, -2, -3, -2, -1, 0, 1, 0, 0, 0, 0, 0, 0, 2, 1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, -1, -1, -1, 0, 1, 0, 0, 1, 2, 1, 1, 1, 1, 3, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 1, 2, 2, 0, 3, -1, 0, 0, 0, -1, 0, 1, 0, 2, 1, 0, 0, 0, -1, -1, 1, 1, 1, 2, 0, 2, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, -1, 0, 1, 1, 1, 1, 1, 0, 1, 0, 0, 2, 0, 0, 1, 0, 0, 0, 2, 0, 2, 2, 1, 1, -1, -1, -1, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 2, 0, 0, 0, 1, 0, 0, 2, 1, 0, 1, 0, 0, 0, 0, -2, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 4, 1, 1, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, 1, 1, 2, 3, 1, 0, 2, 2, 0, 1, 2, 2, 1, 1, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 3, 2, -6, -4, -2, -3, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -4, -5, -5, -8, -10, -5, -2, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 2, 2, 1, 1, 0, -1, 0, -3, -4, -5, -2, -3, 0, -1, 0, 0, 0, 2, 2, 0, 1, 1, 0, 2, 2, 2, 2, 3, 3, 1, 2, 2, 1, 0, 0, -2, -3, -1, 0, 0, 0, 0, 2, 1, 3, 1, 0, 0, 1, 1, 2, 1, 2, 2, 2, 3, 1, 1, 0, 0, 0, 0, -3, 0, -1, 0, 0, 0, 2, 2, 2, 1, 1, 0, 1, 0, 1, 2, 1, 1, 1, 1, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 1, 2, 0, 1, 0, 1, 0, 2, 1, 1, 2, 2, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 2, 2, 2, 2, 0, 1, 1, 2, 2, 0, 3, 3, 4, 4, 3, 0, 0, -1, -2, -1, -1, -1, 1, 0, 3, 4, 2, 2, 1, 1, 0, 2, 3, 1, 3, 1, 4, 5, 6, 4, 2, 1, -1, -2, -3, -1, 0, 0, 0, 1, 2, 2, 1, 2, 2, 2, 2, 2, 1, 3, 3, 5, 7, 8, 7, 5, 3, 0, -3, -3, -4, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 2, 1, 2, 2, 1, 2, 6, 8, 7, 7, 4, 3, -1, -2, -4, -2, -2, -1, 0, 0, 0, 0, 1, 1, 2, 3, 2, 2, 1, 2, 3, 1, 5, 8, 8, 5, 3, 3, 0, -2, -1, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 4, 4, 1, 1, 4, 6, 8, 6, 4, 3, -1, -2, -3, -1, -1, -2, 0, 0, 0, 0, -2, -1, 0, 0, 0, 3, 4, 3, 3, 1, 5, 9, 8, 8, 5, 2, 0, 0, -2, -2, -1, 0, -2, 0, 0, 0, 0, -1, 0, 1, 0, 3, 3, 4, 2, 0, 4, 7, 7, 7, 4, 2, 0, -2, -1, -3, -1, -1, -2, 0, 0, 1, 0, 0, 0, 0, 2, 2, 3, 4, 2, 0, 3, 5, 6, 3, 4, 2, 0, -2, -1, -1, -3, -2, -1, 0, 0, 2, 1, 0, 0, 0, 0, 3, 4, 4, 3, 0, 0, 2, 4, 2, 2, 1, 1, -2, -3, -1, -3, -1, -2, 0, 0, 1, 2, 1, 0, 0, 0, 1, 2, 3, 3, 0, -3, 1, 1, 1, 2, 2, 1, -2, -1, -2, -1, -1, 0, 1, 1, 2, 1, 2, 2, 0, 1, 1, 2, 3, 2, 0, -5, -1, 2, 3, 3, 2, 0, -1, 0, 0, 0, 0, 0, 3, 2, 1, 3, 2, 1, 0, -1, 0, 0, 1, 2, 0, -7, -3, 0, 1, 2, 2, 0, 0, -1, 0, 1, 0, 1, 2, 3, 1, 2, 1, 0, 0, 1, 0, 0, 2, 0, -1, -7, -3, 0, 1, 3, 1, 2, 0, 0, 0, 0, 0, 2, 2, 1, 2, 2, 3, 4, 2, 3, 3, 1, 2, 0, -1, -7, -3, -1, 0, 1, 3, 2, 0, 0, 1, 2, 1, 2, 2, 3, 2, 4, 2, 2, 3, 3, 4, 1, 1, 0, -2, -9, -5, -1, 0, 0, 1, 1, 1, 0, 1, 1, 1, 3, 3, 3, 2, 3, 1, 3, 2, 3, 3, 3, 0, -1, -2, -7, -4, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 3, 3, 0, 0, 0, 2, 1, 2, 3, 1, 1, -2, -3, -6, -3, -1, -1, 0, -1, 0, -1, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -4, -5, -6, -3, -2, -3, -3, -1, -2, -2, -2, 0, 0, 0, 0, -2, -1, 0, 0, -3, -2, -4, -4, -4, -4, -5, -6, -10, 1, -1, -1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 1, 0, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 6, 5, 4, 1, 3, 1, 3, 3, 4, 4, 2, 4, 2, 3, 3, 4, 2, 2, 3, 5, 7, 7, 7, 4, 3, 5, 7, 2, 1, 1, 1, 1, 1, 2, 0, 0, 2, 0, 1, 2, 3, 2, 2, 2, 4, 3, 3, 3, 5, 5, 2, 3, 5, 2, 1, 2, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 3, 1, 1, 2, 1, 2, 6, 2, 0, 2, 1, 1, 0, 1, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 5, 1, 1, 1, 0, 0, 1, -1, -1, -1, -2, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 2, 0, 0, 0, -1, 0, -1, 0, -2, -2, -2, 0, 0, 0, -1, -2, 0, -1, -1, -1, -3, -2, -2, -2, -2, -3, 2, 1, 0, -1, -1, -1, -1, -2, -2, 0, -1, -1, 0, 0, -1, -2, 0, -1, 0, -2, -3, -5, -4, -3, -4, -6, 0, 0, -1, -3, -2, -4, -2, -3, 0, -2, -1, -1, 0, 0, -2, -2, -1, -1, -2, -4, -5, -3, -3, -4, -5, -6, 0, 0, -1, -4, -4, -6, -5, -3, -1, -1, -1, -2, 0, -1, -1, -3, -1, -1, -1, -2, -2, -3, -3, -4, -4, -5, 0, -2, -3, -5, -6, -6, -6, -5, -1, -1, 0, -2, 0, -2, -2, -2, -1, -2, -1, -2, 0, -1, -2, -2, -4, -4, 0, -3, -2, -5, -7, -7, -7, -6, -3, -1, -1, 0, -2, 0, -2, -2, 0, -1, 0, 0, -1, -2, 0, -2, -2, -2, 0, -3, -3, -5, -4, -7, -6, -5, -3, -2, 0, -1, -1, 0, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, -1, -4, 1, -1, -3, -4, -5, -4, -4, -4, -4, -3, -1, 0, -1, -2, -2, 0, 0, 1, 0, 0, -2, -1, 0, 0, -1, -3, 1, -2, -2, -3, -4, -5, -4, -3, -4, -4, -1, 0, 0, -1, 0, 0, 0, -1, 0, -2, -3, -2, -2, -1, -3, -4, 0, -1, -3, -4, -4, -5, -4, -4, -4, -4, -3, 0, 0, 0, 0, 0, 0, 0, -1, -2, -4, -3, -3, -2, -4, -5, -1, -4, -3, -5, -5, -4, -5, -5, -6, -6, -2, 0, 0, 0, 0, 0, -1, -3, -4, -4, -4, -3, -2, -2, -5, -4, -2, -3, -4, -3, -5, -4, -4, -6, -5, -4, -5, -2, 0, 0, 0, 0, 0, -3, -2, -3, -3, -3, -3, -3, -4, -5, 0, -2, -1, -3, -4, -5, -5, -5, -6, -5, -4, -3, 0, 0, 0, -1, -3, -4, -3, -2, -3, -3, -4, -3, -4, -4, 0, 0, -1, -2, -3, -4, -5, -6, -5, -4, -3, -3, -2, -1, -1, -2, -4, -3, -3, -3, -4, -3, -3, -2, -2, -5, 3, 2, 0, 0, -1, -2, -3, -3, -4, -5, -4, -2, -1, -2, -1, -3, -3, -3, -3, -3, -3, -4, -2, -1, -2, -3, 5, 3, 1, 0, -1, -1, -2, -3, -1, -2, -2, -2, -2, -1, -2, -1, -3, -3, -4, -4, -4, -3, -3, -2, -2, -4, 6, 5, 1, 1, 0, -2, 0, -1, 0, -2, -1, -2, -2, -1, -3, -3, -2, -2, -3, -4, -3, -2, -2, -3, -1, -4, 7, 4, 3, 1, -1, -1, 0, -1, 0, 0, -1, 0, -2, -2, -1, -2, -1, -1, -2, -2, -1, 0, -2, -2, -2, -1, 7, 7, 4, 2, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 1, -1, -1, -1, -1, 9, 6, 4, 3, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 1, 2, 2, 4, 3, 4, 3, 0, 0, 1, 0, 8, 7, 5, 3, 2, 3, 0, 2, 0, 2, 2, 1, 3, 4, 4, 5, 5, 5, 7, 6, 6, 5, 4, 2, 3, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, -1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 2, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 2, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, -1, 0, 1, 0, 0, 1, 0, 1, 1, 1, 1, 1, 2, 0, 0, 1, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 1, 0, 1, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 2, 1, 1, 0, 0, 1, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 2, 2, 3, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 2, 2, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 1, 0, 2, 1, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 2, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, -1, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 1, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 4, 3, 2, 3, 2, 3, 3, 3, 3, 3, 4, 5, 5, 5, 5, 4, 5, 5, 5, 4, 5, 7, 5, 5, 5, 4, 2, 2, 1, 2, 2, 2, 4, 3, 3, 2, 1, 1, 2, 2, 3, 4, 3, 4, 3, 4, 5, 5, 4, 4, 4, 4, 3, 2, 0, 2, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 2, 3, 3, 4, 3, 2, 2, 2, 2, 1, 0, 2, 2, 1, 0, 0, -1, -2, -2, 0, 0, 0, 0, 1, 1, 2, 2, 1, 1, 1, 1, 1, 2, 2, 2, 1, 1, 1, 0, -1, 0, -1, -3, -2, -3, -1, -1, -1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 2, 0, 0, -1, -1, -1, -2, -1, -3, -2, -1, -2, -2, -1, -2, -1, 0, 0, 0, -2, -2, 0, 0, 0, -1, -1, 1, 0, 0, -1, -2, -3, -2, -1, -1, -3, -4, -2, -3, -1, -2, -1, -1, -1, -2, -2, -2, -2, -2, -1, -1, -1, 0, -1, -2, -2, -3, -3, -4, -2, -1, -3, -3, -4, -2, -3, -3, -2, -2, -2, 0, -2, -1, 0, -2, -2, -2, -1, 0, -1, -1, -4, -5, -4, -5, -3, -2, -4, -3, -4, -2, -3, -3, -1, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -2, -2, -4, -6, -5, -4, -3, -3, -4, -3, -3, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -5, -6, -5, -5, -5, -5, -5, -4, -3, -2, -3, 0, 0, 0, 0, 1, 0, 1, 0, 2, 2, 0, 0, -1, -1, -3, -4, -6, -6, -5, -5, -5, -5, -3, -4, -3, -2, -2, 0, 0, 0, 0, 1, 1, 0, 1, 2, 0, 0, 0, 0, -1, -3, -4, -6, -5, -5, -6, -5, -4, -2, -4, -4, -2, -1, 0, -1, -1, -1, 0, 1, 0, 0, 0, 2, 0, 0, -2, -3, -4, -4, -4, -6, -6, -5, -3, -4, -4, -2, -3, -1, 0, -2, -1, -1, -1, 0, 0, 0, 0, 0, 1, -1, -1, -3, -3, -4, -5, -6, -5, -4, -4, -4, -3, -2, -2, -1, -3, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, -3, -2, -4, -4, -5, -5, -4, -5, -3, -1, -1, -2, -2, -4, -2, -3, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, -1, -3, -4, -4, -6, -6, -5, -3, -1, 0, -2, -3, -2, -2, -1, -1, 0, 0, 0, 0, -1, 2, 1, 0, -1, 0, -1, -4, -3, -5, -5, -4, -3, -3, -1, -2, -3, -3, -3, -2, -2, 0, 0, -1, 0, 0, -1, 2, 1, 0, 0, 0, -1, -3, -3, -3, -3, -3, -3, -4, -2, -1, -2, -1, -2, -3, -2, -1, -1, 0, 0, 0, 0, 4, 4, 1, 0, 0, -1, -1, 0, -2, -1, -1, -2, -3, -3, -2, -1, -3, -3, -2, -1, -1, 0, 0, 0, 0, 0, 5, 3, 2, 1, 0, 1, 0, 0, -1, -1, 0, -1, 0, -2, -2, -1, -2, -3, -2, -2, 0, -1, 0, 0, 0, 1, 6, 4, 3, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 2, 2, 5, 5, 5, 2, 1, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 2, 1, 1, 7, 7, 4, 4, 3, 0, 2, 2, 2, 3, 2, 1, 1, 3, 2, 3, 3, 3, 4, 3, 4, 2, 2, 2, 3, 3, 6, 7, 7, 3, 3, 3, 2, 2, 3, 3, 2, 4, 4, 5, 4, 5, 4, 5, 5, 5, 7, 5, 4, 5, 5, 3, 6, 6, 5, 6, 5, 4, 4, 5, 3, 5, 5, 4, 5, 6, 6, 6, 7, 8, 8, 7, 7, 6, 7, 7, 4, 5, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 1, 0, -1, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -11, -8, -7, -7, -6, -5, -5, -6, -4, -5, -3, -3, -4, -4, -4, -3, -4, -5, -8, -9, -8, -9, -9, -8, -11, -12, -7, -6, -4, -3, -3, -4, -4, -4, -2, -3, -2, -3, -1, -2, -2, -2, -3, -3, -3, -5, -4, -4, -5, -7, -6, -10, -7, -3, -3, -1, -1, -3, -1, -2, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -1, -2, -4, -7, -5, -3, -1, -1, 0, -2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, -2, -4, -3, -3, -2, 0, 0, 1, 1, 0, 0, 2, 2, 1, 1, 0, 1, 1, 1, 1, 0, 0, 1, 1, 0, 0, -1, -2, -1, -1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 2, 1, 2, 1, 3, 2, 1, 1, 0, 1, 1, 2, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, -1, 0, 2, 1, 2, 2, 1, 0, 0, 1, 0, 2, 2, 2, 0, 0, 3, 1, 3, 2, 1, 0, -1, -2, -2, -2, 0, 0, 0, 1, 3, 2, 3, 2, 1, 2, 1, 1, 2, 2, 2, 1, 4, 6, 6, 4, 2, 0, -1, -4, -3, -3, -1, 0, 1, 2, 2, 3, 2, 3, 3, 1, 1, 1, 3, 4, 2, 3, 5, 8, 8, 5, 2, 0, -2, -4, -2, -1, -1, 1, 1, 2, 2, 2, 3, 3, 3, 2, 1, 3, 2, 2, 1, 6, 8, 7, 8, 6, 2, 0, -2, -3, -4, -3, -1, 1, 2, 2, 2, 2, 1, 1, 1, 1, 1, 3, 3, 2, 2, 5, 7, 7, 7, 4, 3, 1, -1, -3, -3, 0, -1, 1, 2, 1, 3, 1, 1, 1, 1, 2, 0, 3, 2, 2, 1, 6, 9, 6, 6, 5, 1, 1, 0, -1, -2, -2, 0, 0, 1, 2, 0, 1, 1, 2, 2, 0, 1, 2, 2, 1, -2, 5, 7, 7, 7, 6, 3, 0, 0, 0, 0, -1, 0, 2, 1, 1, 1, 0, 0, 1, 1, 0, 2, 1, 0, 0, -3, 5, 7, 6, 6, 4, 3, 2, 1, -1, 0, 0, -1, 0, 0, 1, 2, 0, 0, 1, 0, 2, 3, 2, 2, 1, -2, 5, 6, 5, 5, 3, 1, 1, 0, 0, -1, -1, -1, 0, 1, 1, 0, 1, 0, 1, 2, 3, 3, 3, 3, 2, 0, 3, 4, 5, 4, 4, 1, 1, 1, 1, -1, -1, -2, -1, 0, 2, 3, 2, 2, 1, 1, 1, 1, 3, 4, 2, 0, 1, 2, 4, 5, 3, 2, 1, 0, 0, 0, -2, -1, 0, 0, 1, 2, 3, 3, 0, 1, 0, 2, 1, 2, 2, -1, -2, 2, 1, 3, 4, 4, 1, 0, 0, 0, 0, 0, 0, 1, 3, 4, 2, 2, 1, 0, 2, 0, 2, 2, 1, 0, -3, 0, 0, 2, 4, 4, 2, 0, 0, 0, 1, 1, 0, 3, 1, 2, 2, 3, 1, 1, 2, 1, 0, 1, 1, -1, -5, -1, 0, 1, 3, 1, 1, 0, -1, 1, 1, 2, 2, 1, 2, 1, 1, 1, 3, 1, 3, 1, 2, 0, -1, -2, -7, -4, 0, 0, 1, 2, 0, 0, -1, 0, 0, 0, 1, 0, 1, 2, 2, 1, 2, 4, 3, 3, 2, 0, -1, -2, -9, -4, -2, 0, 1, 0, -1, -1, -1, -1, 0, 2, 1, 1, 2, 1, 2, 2, 3, 3, 5, 4, 0, 0, -2, -5, -10, -6, -4, 0, 0, 0, 0, -1, -1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 2, 1, 2, 1, 1, -1, -2, -5, -9, -7, -5, -3, 0, -1, 0, -1, -1, -2, -2, -1, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, -2, -1, -4, -6, -10, -9, -6, -4, -3, -3, -2, -2, -2, -1, -2, -3, -1, -4, -3, -3, -5, -5, -5, -4, -5, -5, -6, -6, -8, -10, 3, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 2, 1, 2, 2, 0, 2, 1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 2, 1, 1, 1, 3, 2, 2, 1, 0, 1, 1, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, -1, 1, 1, 1, 0, 2, 1, 1, 2, 1, 2, 1, 1, 0, 1, 1, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 2, 0, 2, 2, 1, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 2, 0, 2, 1, 2, 1, 2, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 3, 1, 0, 1, 1, 1, 2, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 2, 3, 0, 2, 1, 2, 0, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 2, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 1, 2, 1, 1, 2, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -2, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -2, -2, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, -1, 0, 0, 0, 0, 1, 0, 0, 1, 3, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, 0, -1, -2, 0, -1, 0, 0, 0, 1, 0, 0, 0, 2, 2, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, -1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 2, 1, 0, 0, 1, 0, 0, 0, 2, 1, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 2, 0, 0, 2, 2, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, -1, -1, 0, 0, 2, 1, 2, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, 2, 0, 2, 1, 1, 0, 0, 0, 2, 1, 1, 1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 1, 0, 1, 1, 0, 1, 1, 1, 1, 1, 1, 2, 0, 1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 2, 1, 1, 1, 0, 1, 1, 0, 1, 2, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, 0, 0, 1, 3, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 1, 4, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, -1, 0, 0, -1, -2, 0, 1, 1, 0, 0, 0, 0, 2, 0, 2, 1, 1, 1, 1, 0, 0, 0, -2, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 2, 0, 1, 2, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, 2, 2, 3, 3, 1, 2, 1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 3, 3, 2, 2, 2, 2, 1, 3, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 2, 3, 3, 2, 2, 3, 2, 3, 2, 2, 1, 1, 0, 0, -1, 0, 0, 0, 0, 2, 1, 2, 2, 2, 3, 1, 1, 2, 2, 2, 3, 3, 3, 3, 3, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 1, 1, 3, 2, 4, 4, 4, 1, 3, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 2, 1, 2, 2, 3, 4, 5, 3, 1, 2, 2, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 3, 3, 0, 3, 3, 3, 3, 4, 4, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, 2, 2, 3, 1, 1, 4, 3, 4, 4, 2, 2, 1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -2, 0, 0, 0, 1, 0, 4, 1, 1, 2, 3, 2, 3, 3, 2, 2, 2, 0, 0, 0, -1, 0, -1, 0, -1, -2, -2, -2, -1, 0, 0, 2, 4, 0, 0, 0, 0, 3, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 2, 3, 3, 0, 0, 0, 0, 1, 1, 1, 2, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 1, 1, 2, 0, 0, 0, 1, 3, 2, 2, 1, 2, 3, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 2, 1, 3, 0, 1, 1, 1, 1, 0, 0, 2, 2, 3, 2, 1, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 3, 3, 0, 0, 1, 2, 0, 2, 1, 2, 2, 2, 1, 2, 1, 0, 0, 0, 2, 1, 1, 0, 0, 1, 0, 1, 3, 2, 0, 1, 0, 1, 1, 3, 3, 2, 2, 2, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 2, 0, 0, 2, 0, 2, 0, 0, 0, 1, 1, 1, 3, 3, 1, 1, 2, 1, 2, 1, 1, 1, 2, 2, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 2, 1, 1, 2, 1, 0, 2, 0, 0, 1, 1, 1, 3, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 2, 2, 1, 2, 0, 1, 0, 1, 2, 2, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 2, 1, 1, 0, 1, 1, 0, 0, 1, 1, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, -2, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 2, 0, 0, 1, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, 0, 1, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 2, 0, 2, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 2, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 1, 2, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 2, 1, 0, 1, 0, 1, 1, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 2, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -2, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -2, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 1, 2, 0, 0, -1, 0, 1, 0, 0, 1, 1, 0, 0, 0, -2, -2, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 2, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 0, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 1, 0, 1, 2, 2, 2, 1, 2, 1, 1, 1, 2, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 3, 2, 2, 1, 2, 1, 2, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 2, 3, 4, 4, 2, 3, 3, 2, 3, 2, 1, 1, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 2, 3, 2, 3, 2, 3, 4, 2, 3, 1, 2, 3, 2, 2, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 3, 3, 4, 3, 4, 3, 3, 1, 2, 2, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 3, 1, 4, 4, 4, 3, 2, 1, 0, 1, 0, 0, 2, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 3, 3, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 2, 1, 3, 1, 2, 2, 2, 1, 0, 0, 1, 2, 0, 0, 0, 0, 1, -1, 1, 0, 0, 0, 0, 0, 1, 2, 2, 4, 2, 4, 3, 3, 3, 3, 2, 1, 0, 2, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 4, 4, 4, 4, 2, 2, 3, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 2, 3, 2, 2, 2, 3, 1, 3, 2, 2, 1, 0, 0, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 3, 2, 2, 2, 1, 1, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 2, 2, 3, 2, 3, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, -2, -1, 0, -2, -1, 0, 1, 2, 2, 1, 1, 2, 3, 2, 2, 1, 2, 0, 0, 1, 2, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 0, 1, 2, 1, 2, 1, 3, 2, 0, 2, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 2, 3, 2, 1, 1, 2, 2, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 1, -1, 0, 2, 3, 2, 3, 1, 2, 1, 2, 1, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 1, 0, 0, 1, 0, 2, 0, 2, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, 0, 0, -2, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, -2, -2, -1, -2, -2, -2, -1, 0, -2, -1, -1, 0, -1, -2, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -2, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, 0, -1, -2, 0, 0, -1, -1, 0, -1, 0, 2, 2, 2, 0, 1, 0, 1, 1, 2, 0, 0, 1, 0, 1, 1, 0, 0, -1, -1, 0, 0, -2, -1, 0, 0, 0, 0, 2, 3, 2, 2, 1, 1, 0, 1, 2, 0, 1, 2, 2, 0, 0, 1, 0, 1, 0, 0, -1, -1, -1, 0, 0, 2, 3, 3, 3, 4, 2, 2, 2, 2, 3, 1, 3, 1, 1, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 2, 3, 3, 2, 3, 2, 4, 3, 3, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, -2, 0, 0, 1, 1, 2, 3, 4, 3, 3, 2, 1, 1, 2, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 1, 2, 3, 4, 3, 2, 1, 1, 0, 0, 0, 2, 0, 0, 0, -1, 1, 0, 1, -1, 0, 0, 0, 0, 1, 0, 2, 4, 3, 3, 3, 2, 3, 2, 3, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 2, 2, 4, 3, 3, 4, 3, 2, 2, 2, 2, 2, 0, 1, 2, 1, 0, 1, 1, 1, 0, 0, -1, 1, 0, 3, 3, 2, 3, 3, 3, 4, 3, 2, 3, 1, 1, 1, 1, 0, 1, -1, -1, 0, 0, 1, 0, 0, -1, 0, 0, 1, 1, 3, 5, 3, 3, 3, 3, 4, 2, 2, 1, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 3, 3, 2, 3, 4, 4, 2, 3, 1, 1, 0, -1, 0, -1, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 1, 2, 2, 4, 2, 4, 3, 0, 0, 0, -2, 0, -3, -1, -1, -2, 0, -1, -2, -1, 1, 0, 0, 1, 1, 1, 1, 2, 1, 3, 3, 1, 1, 2, 0, 1, 1, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, 2, 0, 1, 0, 2, 2, 1, 1, 2, 3, 1, 3, 2, 2, 1, 2, 1, 1, 0, 0, 0, -1, -1, 0, 0, 2, 3, 1, 0, 1, 0, 2, 2, 1, 2, 2, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 2, 1, 2, 2, 1, 1, 1, 2, 2, 2, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 2, 1, 2, 2, 2, 1, 1, 0, 1, 2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 0, 0, 1, 0, 0, 2, 1, 0, 1, 1, 0, 1, 0, 1, 0, -1, -1, 0, 1, 1, 0, 0, 1, 1, 0, 1, 0, 0, -1, -1, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 3, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 2, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, -1, -1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, -4, -3, -1, -1, -2, -1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, -2, -2, -2, -2, -1, -1, -4, -4, -2, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -3, -3, -2, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, 0, 1, 0, 2, 0, 0, 1, 1, 0, 0, 0, 0, -3, -2, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 1, 1, 2, 1, -4, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 2, 1, 1, 1, 1, 1, 2, 2, 1, -3, -1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 2, -3, -1, 0, 2, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 2, 1, 1, 1, 0, 1, 1, 2, 1, -2, -1, 0, 2, 2, -1, -1, -2, -1, -1, -1, -1, 0, 0, 1, 1, 1, 2, 1, 1, 1, 1, 1, 3, 2, 2, 0, 0, 1, 0, 0, 0, -2, -1, -2, -3, -1, 0, -1, -1, 0, 0, 2, 1, 1, 2, 1, 2, 0, 1, 0, 2, 0, 2, 2, 1, 1, 0, -1, -2, -3, -2, -2, -2, -2, -1, 1, 1, 2, 2, 2, 1, 1, 1, 1, 1, 2, 0, 1, 1, 3, 0, 0, 0, -2, -4, -3, -3, -3, -3, 0, 0, 0, 0, 0, 3, 3, 3, 1, 2, 1, 1, 1, 2, 0, 3, 4, 3, 2, 0, -1, -2, -3, -1, -2, -3, -1, 0, 0, 0, 2, 0, 3, 1, 2, 1, 1, 1, 0, 0, 1, 3, 4, 3, 0, 1, -1, 0, -2, -2, -2, -1, 0, 0, 0, 0, 1, 1, 2, 1, 2, 2, 1, 1, 0, 0, 0, 3, 2, 2, 2, 1, 0, -1, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 3, 1, 0, 0, 0, 2, 3, 1, 1, 0, 0, 0, -2, -3, -2, -1, -2, -1, 0, 0, 0, -1, -1, 0, 1, 1, 1, 1, 0, -1, 1, 1, 3, 2, 1, 0, 1, 0, 0, -2, -2, -2, -2, -1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 2, 0, -1, 0, 2, 3, 2, 3, 0, 0, -1, -1, -2, -1, -1, -2, -2, 0, 1, 0, 0, -1, 0, 0, 1, 2, 1, 1, -1, 0, 1, 3, 2, 1, 1, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, -1, -1, 0, 0, 1, 1, 1, 1, -1, -2, 1, 1, 3, 3, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, -1, 0, 2, 2, 2, 1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 1, 0, 1, 1, 0, 1, 0, 0, -1, -3, 0, 1, 3, 2, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, -1, -3, -1, 0, 2, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 2, 1, 1, 0, 0, -2, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 1, 1, 2, 3, 1, 0, 0, -1, -5, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 3, 1, 2, 0, 0, 0, 0, -6, -2, -2, -1, 0, 0, 0, -1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, -1, -3, -6, -4, -3, -1, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -2, -2, -3, -2, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, -1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -2, -2, 0, -1, 0, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 2, 0, 1, 0, 1, 2, 0, 1, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 1, 2, 1, 1, 0, 1, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 1, 1, 1, 2, 2, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 1, 1, 2, 1, 2, 2, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 2, 2, 1, 2, 2, 3, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 2, 1, 1, 0, 0, 2, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 1, 2, 2, 2, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 2, 2, 1, 1, 0, 1, 2, 1, 0, 1, 1, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 2, 1, 3, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 2, 1, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 2, 0, 2, 0, 0, -1, 1, 1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 1, 1, 0, 1, 0, 2, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 2, 1, 0, 1, 0, 0, 1, 2, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 1, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 0, 0, 0, 0, 0, -7, -6, -4, -3, -2, -4, -2, -2, -1, -2, -1, -2, -2, -1, -1, -2, -2, -1, -3, -4, -3, -5, -4, -4, -5, -7, -5, -4, -3, -2, -2, 0, -1, -2, -2, 0, -2, -1, -1, -2, 0, 0, 0, 0, -1, -2, -1, -2, -3, -2, -2, -4, -5, -4, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, -6, -4, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, -3, -1, -2, -1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 2, 2, 2, -3, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, -3, 0, 2, 2, 2, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 2, 2, 0, 1, 1, 0, 0, 0, 2, 1, -2, 0, 2, 2, 2, 1, 1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 2, 3, 2, 1, 1, 1, 0, 0, 0, 3, 0, 2, 5, 5, 4, 3, 2, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, 1, 0, 2, 2, 0, 0, 1, 2, 3, 0, 5, 5, 5, 5, 3, 3, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 2, 0, 2, 2, 1, 1, 2, 2, 5, 7, 6, 7, 3, 2, 1, -1, -2, -1, -1, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 2, 1, 1, 5, 7, 7, 5, 3, 2, 1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 5, 7, 5, 6, 4, 2, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 2, 1, 0, 4, 7, 5, 5, 4, 1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 3, 1, 1, 2, 3, 5, 5, 5, 4, 2, 1, 1, 0, -1, -2, -2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 3, 0, 1, 3, 5, 5, 4, 3, 2, 1, 1, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, -1, 0, 1, 2, 3, 3, 3, -1, 2, 2, 5, 4, 4, 2, 0, 1, 0, -1, 0, -1, -2, 0, 2, 2, 0, 1, 0, 0, 1, 2, 3, 2, 2, -2, 1, 2, 3, 2, 4, 2, 1, 0, 0, 0, -1, 0, -1, 0, 1, 1, 0, 1, 0, -1, 1, 1, 2, 2, 1, -3, -1, 2, 3, 2, 4, 3, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 0, 0, -1, 1, 1, 2, 2, -5, -3, 0, 1, 1, 3, 3, 1, 0, -1, 0, 0, 1, 1, 2, 0, 1, 1, 0, 0, 0, 1, 0, 1, 1, 0, -6, -3, 0, 0, 2, 2, 1, 0, -1, -1, 0, 0, 1, 0, 0, 1, 2, 1, 2, 2, 1, 1, 2, 2, 0, 0, -8, -6, -3, 0, 1, 1, 1, 1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 1, 1, 1, 1, 0, 0, -8, -5, -3, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 0, 1, 1, 1, 2, 3, 3, 1, 0, 0, -8, -6, -3, -3, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 2, 2, 0, 0, -2, -8, -6, -5, -4, -2, -1, 0, -2, -1, -1, 0, -2, 0, 0, 0, 0, -1, -1, -2, 0, -1, 0, -1, 0, -1, -4, -8, -6, -6, -4, -4, -2, -2, -3, -2, -2, -2, -1, -2, -3, -2, -3, -1, -3, -4, -3, -4, -4, -3, -3, -5, -6, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, -1, 0, -1, 0, 1, 0, 0, 1, 0, 0, 2, 0, 1, 1, 1, 1, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 2, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 2, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 2, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 0, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 2, 1, 1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 2, 2, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 1, 1, 0, 0, 1, 0, 1, 0, 1, 1, 0, 1, 0, -1, -1, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 2, 1, 2, 2, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 1, 1, 2, 2, 2, 1, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 2, 2, 0, 0, 0, 1, 1, 1, 1, 0, 2, 1, 1, 1, 0, 0, 0, 1, 1, 0, -1, 1, 0, 1, 1, 1, 2, 0, 1, 1, 0, 0, 2, 2, 0, 0, 2, 1, 1, 2, 2, 1, 0, 0, 1, 1, 0, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 1, 0, 2, 1, 0, 1, 0, 2, 1, 2, 2, 2, 0, 0, 1, 0, 0, 0, 2, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 1, 0, 2, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 5, 3, 2, 2, 4, 4, 4, 6, 4, 3, 2, 2, 3, 4, 2, 4, 4, 6, 6, 5, 5, 2, 3, 3, 0, 2, 5, 4, 2, 2, 4, 3, 5, 4, 4, 3, 4, 2, 1, 1, 2, 5, 5, 5, 6, 4, 3, 4, 2, 1, 0, 0, 5, 4, 2, 2, 3, 5, 5, 4, 3, 2, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 0, 0, 0, 0, 1, 5, 4, 4, 3, 5, 4, 4, 4, 2, 2, 1, 1, 0, 0, 0, 1, 3, 2, 3, 0, 0, 0, 0, -1, 0, 0, 4, 3, 4, 5, 5, 3, 4, 2, 1, 2, 1, 1, 0, 0, 1, 0, 1, 1, 0, 0, -1, -1, 0, -3, -2, -2, 3, 2, 4, 4, 2, 4, 4, 2, 2, 2, 3, 1, 1, 1, 1, 0, 0, 1, 0, -1, -1, -3, -2, -4, -4, -3, 4, 4, 2, 3, 2, 4, 3, 4, 2, 3, 3, 2, 2, 3, 1, 0, 0, 0, -2, -2, -2, -1, -3, -3, -3, -5, 2, 3, 2, 2, 1, 3, 3, 3, 2, 4, 4, 4, 4, 3, 0, 0, 0, -1, -3, -4, -3, -3, -3, -4, -4, -5, 0, 0, 1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, -1, 0, -1, -2, -2, -1, -3, -3, -4, -3, -3, -4, 0, -1, 0, -1, 0, -1, 0, 1, 1, 1, 1, 1, 0, -1, 0, 0, 0, -2, -1, -1, -1, -1, -2, -4, -4, -3, -1, 0, 0, -2, 0, -1, -1, 0, 1, 0, 0, 0, 0, -1, -1, 0, -2, -2, -3, -2, 0, 0, 0, -1, -1, -2, -1, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -2, -2, 0, -1, -2, -2, -2, -1, 0, -1, 0, 0, -1, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, 1, -1, -1, -1, -3, -2, -1, -3, -2, -2, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 1, 1, 1, 2, 0, 0, 0, -1, -1, -1, -1, -2, -2, -5, -2, -2, 0, 0, 0, -1, -1, -1, -3, -1, 0, 0, 0, 0, 2, 0, 1, 1, 0, 0, 0, 0, -2, -3, -3, -4, -3, -4, -1, -1, 0, -1, 0, -3, -3, -2, 0, -1, 0, 0, 1, 0, 1, 0, 2, 1, 0, -1, 0, -2, -2, -4, -4, -2, -2, -3, -3, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 2, 2, 2, 1, 0, 0, -1, -2, -3, -1, -4, -4, -2, -3, -2, 0, 0, 1, -1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 1, -1, -1, 0, -1, 0, -1, -3, -3, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 2, 0, 0, 0, -1, -1, -1, -2, -1, -3, -2, -2, 0, -1, 0, 1, 2, 2, 2, 2, 3, 3, 3, 1, 1, 2, 0, 1, 0, -1, 0, -1, 0, 0, -2, -2, -2, -1, 0, 0, 1, 1, 1, 2, 2, 3, 3, 4, 3, 3, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -2, 0, -2, 1, 1, 2, 0, 1, 3, 3, 4, 5, 4, 3, 2, 3, 2, 1, 2, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 3, 2, 2, 2, 1, 3, 2, 4, 5, 3, 3, 1, 1, 1, 2, 1, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 4, 3, 2, 2, 0, 0, 2, 3, 2, 3, 2, 2, 3, 1, 2, 1, 3, 1, 2, 3, 2, 1, 0, 0, 0, 1, 6, 5, 6, 4, 1, 2, 1, 2, 4, 2, 3, 2, 1, 2, 2, 2, 1, 3, 1, 3, 1, 2, 1, 2, 1, 3, 7, 6, 5, 4, 3, 3, 2, 3, 5, 3, 3, 4, 2, 4, 4, 3, 2, 3, 2, 3, 3, 3, 5, 4, 5, 3, -2, -1, 0, -1, -1, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -2, -3, -4, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 2, 2, 1, 1, 0, 1, 1, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 2, 2, 0, 0, 1, 0, 1, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 2, 3, 2, 1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 2, 1, 1, 3, 4, 4, 3, 3, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 4, 2, 3, 4, 1, 0, 0, -1, 0, -2, 0, -1, 0, -1, -1, 0, -2, -1, 0, 0, 0, 1, 1, 0, 2, 3, 2, 3, 4, 2, 2, 0, -1, -1, 0, -1, -2, -1, 0, -2, 0, -1, -2, 0, 0, -1, 0, 1, 0, 2, 1, 2, 3, 4, 4, 2, 1, 1, 0, -1, -1, -2, -2, -1, -1, -1, -2, -2, -1, -2, 0, 0, 0, 0, 0, 2, 2, 2, 5, 4, 4, 3, 0, 0, -1, -1, 0, -1, -3, -3, -3, -2, -2, -1, -3, -1, -1, -2, 0, 1, 2, 1, 1, 4, 4, 4, 3, 2, 1, 0, 0, -1, -1, -2, -2, -4, -4, -2, -1, -2, -1, 0, -1, -1, 0, 0, 1, 1, 3, 2, 3, 4, 3, 3, 0, 0, -1, 0, -1, -1, -4, -2, -3, -1, 0, 0, 0, 0, 0, 0, 0, 2, 3, 4, 3, 0, 3, 2, 3, 1, 0, 0, 0, -2, -2, -3, -3, -2, -2, -2, 0, 1, 0, 0, 0, 0, 0, 0, 4, 4, 2, 0, 0, 1, 2, 1, 2, 0, -1, 0, -1, -1, -2, -2, -1, 0, 0, 1, 0, 1, -1, 0, 0, 0, 2, 2, 2, -1, -1, 0, 0, 0, 1, 0, 0, -1, -2, -2, -2, -1, 0, 1, 2, 1, 0, 0, 1, 0, 0, 0, 2, 2, 3, -2, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 1, 1, 1, 2, 2, 2, 1, 0, 0, 0, 1, 2, 1, -4, -3, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 1, 2, 2, 2, 3, 1, 0, 1, 0, 2, 0, 1, -4, -2, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 2, 1, 1, 3, 3, 1, 2, 2, 1, 1, 1, 3, 1, 0, -3, -1, -2, -1, -1, 1, 0, 1, 0, 1, 0, 1, 0, 1, 2, 1, 2, 2, 0, 2, 1, 3, 1, 0, 0, 0, -2, -3, -2, 0, 0, 0, 1, 1, 2, 0, 1, 2, 1, 1, 2, 1, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, -3, -2, -1, -1, 0, -1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -2, 0, -1, 0, 0, -1, 0, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -3, -4, -3, -3, -3, -1, -2, -1, -2, -3, -2, -3, -2, -1, -1, 0, -1, -2, -3, -3, -3, -1, -2, -3, -1, -2, -1, 0, 0, -1, -2, -2, -3, -1, 0, 0, -1, -1, -3, -1, 0, -1, -3, -3, -3, -3, -2, -2, -4, -2, -3, -3, -2, -3, -2, -2, -1, -1, -1, -1, 0, -1, -2, -2, -2, 0, -1, -1, -1, -3, -2, -3, -2, -2, -2, -1, -3, -3, -2, -3, -2, 0, -1, -2, -2, -1, -1, -1, -2, 0, 0, -1, -2, -1, -2, -2, -3, -4, -3, -1, -3, -2, -2, -2, -4, -5, -3, -2, -2, -1, 0, -2, -1, -2, -3, 0, -1, -1, -1, -3, -2, -2, -3, -2, -3, -1, -3, -2, -4, -1, -4, -4, -3, -4, -2, -2, -1, -1, -3, -3, -1, 0, 0, 0, -1, -1, -2, -2, -3, -2, -3, -1, -2, -2, -2, -2, -3, -4, -3, -2, -1, -3, -2, -3, -1, -1, -2, 1, 1, 0, 0, -2, -2, -3, -1, 0, -1, -3, -3, -4, -4, -3, -3, -3, -5, -2, -2, -2, -3, -2, -2, -1, -1, 0, 1, 0, 0, 0, -1, -3, -1, 0, 0, -2, -2, -2, -4, -4, -4, -4, -3, -3, -4, -4, -4, -4, -1, -2, 0, 0, 3, 2, 2, 1, 1, 0, 0, 0, 0, -2, -3, -3, -3, -3, -4, -4, -3, -3, -2, -5, -4, -3, -3, -2, 1, 3, 2, 4, 2, 2, 2, 0, 0, 0, -1, 0, -2, -1, -2, -2, -2, -3, -3, -2, -3, -3, -5, -4, -1, -2, 0, 2, 3, 4, 4, 1, 2, 0, 1, 0, 0, -1, 0, -3, -2, -2, -2, -2, -2, -3, -1, -5, -4, -4, -2, 0, 0, 2, 3, 3, 4, 3, 0, 0, 1, 2, 2, 0, -1, -2, -3, -2, -3, -3, -4, -3, -1, -3, -4, -3, -3, -1, 2, 1, 4, 4, 3, 3, 0, 0, 0, 0, 1, -1, -1, -1, -2, -2, -2, -3, -2, -3, -1, -4, -5, -2, -1, -2, 1, 3, 3, 5, 4, 3, 1, 1, 0, 1, 0, -1, -2, -1, -2, -2, -2, -3, -4, -4, -3, -4, -5, -4, -1, -1, 0, 3, 3, 4, 3, 1, 0, 0, 2, 0, 0, -2, -2, -2, 0, 0, -2, -2, -4, -3, -2, -4, -3, -2, -2, 0, 0, 3, 4, 6, 4, 1, 0, 1, 3, 1, 1, -1, 0, -1, -1, -1, -2, -1, -2, -3, -2, -2, -3, -2, -2, 0, 0, 2, 3, 3, 5, 2, 0, 1, 0, 2, 0, -1, -2, -2, -1, -1, 0, -1, -1, -2, -4, -3, -3, -4, -2, 0, 2, 1, 1, 3, 3, 2, 0, 0, 0, 0, 1, 0, 0, -1, -2, -1, -1, -1, -2, -2, -5, -3, -4, -4, -1, 0, 2, 0, 2, 1, 1, 0, 2, 0, 0, -1, -2, 0, 0, -3, -2, -2, 0, 0, 0, -1, -2, -3, -3, -2, 0, 0, 1, 0, 2, 2, 1, 0, 2, 1, 0, -2, -2, -1, -2, -4, -2, -3, 0, -2, 0, -1, -1, -2, -3, -2, -1, 0, 0, 1, 2, 2, 0, 0, 0, 1, -1, -3, -3, -3, -3, -2, -3, -2, -1, -1, 0, -2, -1, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, -3, -4, -4, -4, -1, -3, -3, -3, -2, -1, -2, -1, -1, -3, 0, 0, -1, 0, -1, 1, 2, 0, 0, 0, 1, 0, -2, -4, -4, -2, -2, -3, -2, -3, -3, -2, -2, -3, -4, -1, -2, 1, 1, -2, -3, 0, 1, 0, -1, 0, 0, 0, -3, -4, -4, -2, -2, -2, -2, -1, -3, -3, -4, -4, -3, -4, -2, -1, 0, -2, -3, 0, 0, -1, -2, -1, 0, -1, -3, -3, -3, -3, -3, -1, -2, -2, -2, -3, -2, -3, -2, -3, -3, -1, -2, -2, -3, -2, -1, -2, -3, -2, -1, -2, -4, -4, -3, -3, -1, -2, -2, -2, -1, -4, -3, -3, -2, -2, -1, -2, -1, -3, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 3, 2, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 2, 1, 1, 2, 2, 1, 0, 0, 0, 1, 1, 2, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 2, 1, 4, 3, 3, 1, 1, 1, 0, 1, 2, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 2, 1, 3, 3, 1, 2, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 1, 2, 1, 2, 2, 3, 1, 3, 1, 1, 2, 1, 0, 0, 0, 0, 1, 0, 1, 0, 2, 2, 0, 1, 2, 0, 1, 1, 1, 2, 3, 2, 3, 3, 4, 2, 2, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 2, 2, 2, 0, 0, 1, 3, 2, 3, 2, 3, 1, 2, 1, 2, 0, 1, 2, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 3, 3, 2, 3, 1, 2, 2, 2, 1, 3, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 4, 4, 2, 2, 1, 3, 1, 3, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 2, 3, 4, 3, 5, 4, 3, 2, 3, 2, 3, 1, 1, 0, 1, 0, 0, 0, -1, 0, 1, 0, 1, 1, 0, 1, 0, 0, 1, 2, 3, 3, 2, 3, 1, 2, 3, 1, 1, 1, 1, 0, 0, -1, -1, -2, 0, 0, 1, 2, 1, -1, 0, 0, 0, 1, 1, 1, 2, 2, 1, 1, 1, 1, 0, 2, 1, 0, 0, -2, -2, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 2, 3, 2, 2, 2, 2, 2, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 2, 1, 0, 3, 2, 1, 2, 1, 2, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 2, 0, 0, 1, 1, 0, 1, 1, 0, 2, 0, 0, 0, 0, 2, 0, 0, 1, 1, 0, 2, 1, 1, 0, 0, 1, 0, 1, 2, 0, 0, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 1, 0, 2, 0, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, 0, 0, 2, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 1, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -2, -1, -1, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 2, 0, 1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 1, 0, 1, 1, 0, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 2, 0, 1, 1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 2, 2, 2, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 3, 1, 2, 1, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, 1, 2, 2, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 1, 1, 0, 0, 1, 0, 0, 1, 2, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, -2, 0, -2, -1, -1, -1, -1, 1, 1, 1, 1, 2, 2, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, -1, -1, -3, -3, -1, -2, -1, -1, -2, -2, -1, 0, 0, 0, 2, 3, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -4, -2, -4, -2, -2, -2, -2, -1, -2, -2, 0, 0, 0, 0, 2, 1, 2, 2, 1, 0, 0, -1, 0, -1, -1, -2, -3, -3, -4, -4, -2, -2, -2, -1, -2, -2, -1, 0, 0, 0, 2, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, -2, -4, -4, -5, -3, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 1, 1, 0, -1, -1, -4, -3, -3, -2, -2, -2, -2, 0, -1, -1, 0, 0, 1, 2, 2, -1, 1, 1, 1, 1, 2, 1, 1, 1, 0, 0, -2, -4, -4, -3, -3, -2, -1, 0, -1, -1, 0, 0, 1, 1, 3, 0, -1, 0, 1, 2, 2, 1, 0, 0, 0, 0, -2, -2, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 1, 0, 2, 1, 2, 1, 2, 0, 0, -1, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 1, -1, 0, 0, 0, 0, 2, 1, 2, 1, 0, -1, 0, -1, 0, 0, 2, 2, 1, 1, 0, 0, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, 1, 0, 0, 2, 1, 1, 1, 1, 0, 0, 2, 2, 0, 0, 0, 0, 0, 1, 2, 2, 2, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 3, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 2, 0, 1, 1, 3, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 2, 0, 1, 1, 0, 0, 1, 0, 2, 3, 2, 0, 0, 0, 0, -1, 0, 1, 0, 0, 2, 1, 0, 0, 1, 1, 2, 1, 1, 0, 1, 0, 0, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 2, 1, 0, 0, 1, 2, 1, 1, 0, 0, -1, 0, 0, -2, -1, 0, 0, 0, 0, -1, 0, 2, 2, 4, 1, 0, 2, 2, 1, 0, 0, 0, 2, 0, 0, -1, -1, -2, 0, -2, -1, 0, -1, 0, -1, 0, 0, 2, 1, 2, -11, -9, -8, -7, -7, -7, -7, -5, -4, -6, -4, -4, -4, -4, -5, -5, -8, -9, -9, -10, -11, -8, -8, -8, -10, -12, -9, -8, -5, -6, -3, -5, -4, -4, -5, -4, -3, -4, -3, -2, -2, -4, -5, -6, -7, -6, -5, -5, -4, -6, -6, -9, -6, -5, -3, -2, -3, -1, -1, -2, -3, -3, -3, -3, -3, -1, 0, 0, -2, -3, -1, -2, -2, -3, -2, -3, -5, -8, -5, -2, -2, -1, -2, -1, 0, 0, 0, 0, -2, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -2, -5, -3, -3, -3, -1, 0, 0, 0, 1, 2, 1, 1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, -2, -3, -2, -2, 0, 0, 1, 2, 2, 2, 1, 0, 0, 1, 1, 1, 2, 2, 0, 1, 0, 0, 0, 1, 3, 0, -2, -2, 0, 0, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 2, 1, 2, 1, 1, 1, 0, 1, 0, 1, 2, 1, 0, 0, 0, 3, 2, 2, 1, 1, 0, -1, -1, 0, 0, 1, 2, 4, 3, 2, 2, 2, 2, 0, 0, 3, 2, 1, 0, 1, 3, 6, 6, 5, 2, 0, -2, -2, -1, -2, 0, 0, 1, 3, 3, 3, 3, 2, 2, 1, 2, 3, 3, 3, 0, 2, 7, 8, 8, 4, 2, 0, 0, -2, 0, -2, 0, 0, 1, 2, 2, 3, 2, 3, 1, 1, 2, 0, 2, 2, 0, 5, 7, 7, 7, 5, 1, 0, -1, -2, -2, -1, 0, 1, 2, 3, 1, 1, 2, 2, 1, 1, 1, 0, 1, 0, 0, 4, 6, 6, 7, 5, 2, 1, 0, 0, -3, -1, 0, 0, 1, 1, 2, 1, 1, 2, 0, 1, 2, 2, 2, 0, -1, 4, 5, 6, 5, 4, 3, 3, 1, 0, 0, 0, -1, 0, 2, 2, 0, 1, 0, 2, 1, 2, 1, 0, 0, 0, -3, 5, 6, 6, 7, 5, 4, 3, 2, 0, -1, -1, 0, 0, 1, 0, 1, 1, 0, 1, 2, 2, 2, 0, 0, -2, -3, 6, 6, 6, 7, 6, 4, 3, 2, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 3, 3, 1, 1, 0, -1, -6, 5, 6, 5, 5, 4, 3, 4, 3, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 2, 1, 3, 0, -1, -4, 4, 6, 4, 5, 3, 3, 3, 1, 2, 0, -1, -1, 0, 0, 1, 1, 0, 0, 1, 2, 2, 3, 3, 1, 0, -4, 1, 4, 4, 6, 5, 4, 2, 1, 1, 0, -1, -1, -1, 0, 1, 0, 1, 0, 0, 1, 1, 0, 2, 1, 0, -2, 2, 2, 4, 5, 4, 2, 1, 0, 0, 0, -1, 0, -1, 1, 1, 1, 1, -1, 0, 0, 1, 0, 1, 1, 0, -1, -1, 0, 3, 5, 5, 3, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -3, -3, 0, 0, 3, 3, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -2, -3, -5, -3, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 2, 1, 0, -1, -3, -5, -7, -3, -1, 0, 0, -1, -2, -1, -2, -1, -1, 0, 0, 0, 1, 0, 0, 1, 2, 4, 3, 1, 0, -1, -2, -5, -8, -6, -3, -2, 0, -1, -2, -1, -3, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 3, 2, 1, -1, -2, -4, -6, -11, -7, -4, -3, -2, -4, -4, -2, -3, -2, -1, -2, -3, -2, -3, -3, -3, -2, -1, 0, 0, -1, -2, -4, -5, -8, -12, -9, -6, -4, -5, -6, -4, -3, -4, -5, -5, -5, -5, -4, -4, -5, -5, -5, -5, -4, -5, -6, -6, -8, -9, -11, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, -1, 0, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, -3, -1, -2, 0, -1, -1, -2, -2, -1, 0, 0, -2, -1, -1, -2, 0, -1, -3, -2, -2, -2, -1, -3, -2, -4, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -2, 0, -1, -1, 0, -1, -4, 0, 0, 1, 1, 1, 0, 0, 1, 1, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, -3, 0, 0, 1, 2, 0, 0, 1, 0, 1, 1, 0, 0, 2, 2, 1, 1, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 2, 0, 1, 1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 1, 2, 1, 1, 3, 2, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, -1, 0, 2, 1, 2, 2, 0, 2, 2, 0, 0, 0, 1, 0, 1, 2, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 2, 1, 3, 1, 1, 2, 0, 0, -1, 0, -1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 3, 2, 3, 1, 3, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 3, 5, 5, 4, 3, 3, 2, 1, 0, -1, -1, -1, 0, 2, 2, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 2, 2, 3, 2, 1, 0, 1, 0, 0, 0, -1, 0, 0, 1, 2, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 3, 3, 2, 1, 2, 0, 1, 0, 0, -1, 0, 0, 1, 2, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 2, 2, 2, 1, 2, 1, 1, 1, 0, 0, 0, 0, 2, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 3, 2, 3, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 4, 2, 1, 2, 3, 0, 0, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 1, 1, 1, 0, 0, -1, 2, 2, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 1, 0, 0, 1, 2, 0, -2, 2, 2, 0, 2, 1, 1, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, -2, 0, 2, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 2, 1, 1, 0, -1, 0, 0, 0, 1, 1, 2, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 2, 1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 1, 0, -1, -2, -2, -1, 0, 0, 2, 0, 0, 0, -1, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, -2, 0, -2, -2, -2, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, -1, -1, -2, -2, -2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, -1, 0, -2, -1, -2, -2, -2, -1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, -1, -2, -2, -4, -4, -3, -2, -2, -1, -1, -1, -1, -1, 0, 0, -1, -2, -2, -2, -2, -3, -2, -2, -2, -2, -2, -2, -3, -4, 5, 3, 1, 2, 2, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 1, 3, 3, 3, 3, 2, 1, 2, 3, 2, 3, 3, 3, 2, 2, 1, 2, 2, 3, 2, 2, 2, 0, 0, 0, 0, 2, 2, 3, 3, 2, 1, 2, 0, 0, 1, 2, 4, 3, 4, 2, 3, 3, 4, 4, 3, 3, 1, 1, 0, 0, 0, 0, 1, 3, 3, 2, 0, 0, 1, 0, 2, 1, 3, 5, 4, 3, 6, 5, 3, 4, 4, 4, 2, 1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 2, 5, 5, 5, 5, 6, 4, 3, 3, 2, 2, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, -1, -1, 4, 5, 6, 4, 6, 5, 4, 5, 3, 4, 4, 3, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, -3, -2, 2, 6, 5, 5, 5, 5, 4, 5, 4, 4, 4, 3, 3, 3, 1, 0, 0, 0, -1, -1, 0, 0, -1, -2, -3, -1, 2, 5, 4, 6, 5, 4, 6, 5, 3, 4, 5, 4, 2, 2, 1, 0, -1, -1, -3, -2, -1, -2, 0, -2, -3, -1, 0, 1, 3, 2, 4, 3, 4, 4, 4, 2, 2, 2, 1, 0, -1, -1, -1, -2, -3, -3, -1, 0, 0, -2, -3, -2, 0, 0, 1, 0, 0, 1, 3, 3, 1, 3, 2, -1, -2, -2, -2, -4, -3, -2, -3, -4, -3, -2, 0, -3, -2, -2, 1, -1, -2, 0, 0, 1, 0, 0, 0, 0, 0, -1, -3, -4, -4, -2, -3, -3, -4, -5, -4, -2, -3, -2, -1, -1, 0, -2, -2, -1, -1, 0, 0, 0, 0, 0, -1, -1, -4, -4, -5, -4, -1, -3, -2, -3, -3, -3, -3, -2, -2, 0, -3, -2, -1, 0, 0, 0, 1, 1, 0, 0, 0, -2, -4, -5, -4, -3, -1, -3, -3, -4, -3, -2, -3, -2, 0, 0, -2, -1, 0, 0, 2, 3, 2, 1, 3, 3, 1, -1, -3, -5, -4, -4, -2, -2, -2, -3, -2, -1, -2, -2, 0, 0, -4, -4, -3, -1, 1, 3, 2, 4, 3, 3, 2, 0, -2, -2, -2, -3, -2, -3, -4, -2, -2, -2, -1, -2, 0, 0, -5, -4, -3, -2, 0, 1, 3, 3, 3, 4, 3, 1, 0, -1, -2, -2, -2, -2, -2, -3, -3, -3, -3, -2, -1, 0, -3, -4, -2, 0, 1, 0, 1, 3, 3, 3, 2, 2, 0, -1, -2, -2, -1, 0, 0, -2, -2, -2, -4, -2, -1, 0, -1, -1, -2, -1, 0, 2, 1, 4, 4, 2, 3, 2, 0, -1, -2, 0, -1, 0, 0, 0, 0, -2, -4, -1, -2, -1, 0, -1, 0, 0, 0, 2, 3, 3, 4, 5, 3, 4, 2, -1, -1, -2, 0, 0, 0, 0, 0, -2, -3, -3, -1, -1, 0, 0, 0, 0, 0, 2, 2, 3, 5, 5, 4, 5, 3, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 3, 5, 6, 5, 5, 4, 3, 1, 1, 0, 0, 0, 0, -1, -1, -2, -2, -2, -2, -2, 1, 1, 0, 2, 1, 1, 4, 5, 4, 6, 5, 3, 3, 2, 0, 0, 0, 1, 0, 0, 0, 0, -3, -2, -3, -1, 2, 1, 0, 1, 1, 2, 3, 4, 4, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -2, -1, -3, -2, 0, 3, 1, 1, 1, 0, 1, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, -1, -1, 0, 2, 4, 3, 2, 0, -1, 0, 1, 2, 2, 1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 2, 3, 3, 2, 1, 1, 1, 0, 2, 3, 3, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 2, 3, 5, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 2, 1, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, 2, 0, 1, 0, -1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 2, 1, 0, 0, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, 1, 2, 0, 0, -1, 0, -3, -2, -2, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -2, 0, -1, 0, -1, 1, 1, 0, 1, 0, -1, -3, -2, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 3, 2, 1, 0, -1, 0, -2, -4, -3, -1, -1, -1, 0, 0, -1, -1, -1, -1, 1, 0, 0, 0, 0, -1, 0, 0, 3, 2, 1, 1, 0, -2, -2, -2, -2, -1, -2, -1, -1, -1, -1, -1, -2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 4, 3, 0, 1, 0, 0, -2, -3, -1, -2, -1, -1, -2, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 2, 0, 0, 0, -1, -1, -2, -1, -2, -4, -3, -1, -2, -1, 0, -2, -1, 0, 0, -1, -1, 1, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, -2, -1, -2, -3, -1, -2, -2, -2, 0, 0, 0, 0, -1, 0, -1, 0, 1, 1, 1, -1, 1, 0, 1, 0, 0, -2, -2, -2, -2, -1, -3, -2, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -2, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -2, -3, -1, 0, 0, 1, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, -1, 0, -3, -1, -1, -2, -2, 0, 1, 0, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -2, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 2, 0, 1, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 2, 2, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, -1, 0, 2, 1, 1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 2, 1, 2, 0, 2, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -2, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -2, -2, 0, -1, -1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 0, 0, -1, 0, -1, 1, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, -1, 0, 1, 0, 0, 0, 1, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 1, 1, 0, 2, 1, 2, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 2, 0, 2, 2, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, -1, 1, 1, 0, 1, 0, 1, 0, 1, 0, 1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 0, 2, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, -1, -1, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -7, -5, -6, -3, -3, -3, -3, -2, -3, -2, -3, -1, 0, -2, -2, 0, -1, -2, -1, -3, -4, -3, -5, -4, -5, -6, -6, -5, -3, -3, -3, -1, 0, 0, -2, -1, 0, -1, 0, -2, 0, -1, 0, -1, -1, -3, -1, -2, -4, -2, -4, -2, -6, -5, -1, -1, 0, 0, 0, -1, 0, -2, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -2, -2, -5, -3, -2, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -5, -2, -2, 0, 0, 0, 0, 0, 1, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, -4, -3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 2, 2, -3, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 1, 1, 0, 1, 0, 1, 3, -3, -1, 0, 2, 1, 2, 1, 1, -1, 0, 0, 0, -1, -1, 0, 0, 1, 2, 0, 0, 2, 1, 2, 0, 1, 1, -3, 0, 3, 2, 4, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 1, 2, 1, 0, 1, 1, 0, 1, 4, 3, 3, 3, 2, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 3, 2, 2, 1, 1, 2, 0, 3, 3, 3, 3, 3, 1, 1, 1, 0, -1, -1, -1, 0, 1, 0, 2, 1, 0, 2, 1, 1, 0, 1, 1, 2, -1, 1, 3, 3, 3, 3, 2, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 0, 3, 3, 3, 4, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 2, 1, 0, 3, 4, 4, 4, 2, 1, 0, 0, 1, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 2, 1, 2, -1, 1, 4, 3, 3, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 2, 1, 0, 2, 3, 3, 3, 3, 2, 1, 1, 0, 1, -1, -1, 0, 0, 0, 0, 1, 0, -1, 0, 1, 2, 3, 3, 1, -3, 1, 2, 1, 2, 1, 1, 1, 1, 0, 0, 0, -2, 0, 0, 1, 0, 1, 1, 0, 0, 1, 2, 3, 3, 1, -2, -1, 1, 2, 1, 3, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 2, -3, 0, 1, 0, 0, 2, 3, 1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, -6, -3, -1, 0, 0, 1, 2, 0, -1, -1, 0, 0, 0, 1, 2, 2, 2, 2, 1, 0, 0, 0, 1, 0, 0, 0, -6, -5, -1, -1, 0, 1, 1, 2, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 1, 0, 1, 2, 0, -7, -4, -2, -1, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 2, 1, 1, 1, 1, 1, 2, 0, 1, 1, -6, -4, -4, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 2, 2, 0, 0, -7, -5, -4, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 0, 2, 0, 0, -5, -5, -3, -2, -1, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, -1, -1, -2, -1, -1, -1, 1, 0, 1, 0, 1, 1, 2, 1, 3, 3, 2, 2, 1, 2, 1, 1, 0, 0, 1, 0, 2, 0, 0, 0, -1, -1, 0, 0, 1, 1, 1, 0, 2, 0, 2, 1, 2, 2, 2, 1, 2, 1, 1, 1, 1, 0, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -1, 0, -1, 0, 1, 0, 0, 0, 1, 0, 1, 2, 1, 1, 1, -1, -1, 0, 0, 0, 0, -1, -1, 0, -2, -2, 0, -2, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -2, 0, 0, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 1, 0, 0, 0, -1, -1, 0, -2, -1, 0, 0, -1, -3, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -2, 0, -2, -1, -2, -3, -1, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, -1, -1, -2, -2, -1, -2, -3, -3, -2, -2, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, -1, -3, -3, -5, -3, -3, -3, -1, -2, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 0, -2, -4, -4, -5, -3, -4, -1, -2, -2, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 1, 2, 0, 0, 1, 0, -1, -2, -4, -3, -4, -4, -4, -3, -2, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 2, 1, 1, 0, 1, 0, 0, -2, -2, -3, -4, -3, -3, -2, -2, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 2, 0, 0, 1, 0, -1, -1, -1, -4, -2, -3, -1, -2, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 2, 0, 0, 0, -1, -2, -2, -2, -3, -3, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -3, -2, -3, -2, -1, -2, -1, 0, 0, -1, -1, 0, 0, -1, 0, 1, 0, 0, 0, -2, 1, 0, 0, 1, 0, -2, -2, -2, -4, -3, -3, -3, -1, 0, -1, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, -2, 0, 0, 1, 0, 0, 0, 0, -1, -1, -4, -3, -2, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 2, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -2, -3, -3, -3, -1, 0, -1, 0, -1, -2, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, -1, -1, -1, -1, -3, -1, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 3, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 3, 3, 1, 1, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 2, 2, 1, 0, 0, 1, 1, 2, 3, 0, 0, 0, 0, 0, 2, 2, 2, 2, 2, 1, 0, 1, 0, 1, 3, 2, 2, 2, 0, 1, 0, 1, 0, 1, 2, 0, 0, 0, 0, 2, 3, 1, 2, 1, 3, 1, 3, 1, 3, 3, 3, 5, 3, 2, 0, 1, 0, 0, 1, 3, 2, 2, 0, 1, 2, 0, 3, 3, 3, 3, 3, 2, 2, 3, 3, 3, 4, 4, 3, 3, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, 2, 2, 2, 1, 1, 2, 0, 0, 2, 2, 4, 4, 4, -2, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 2, 1, 0, 0, 1, 1, 2, 1, 4, 3, 3, -3, 0, -1, 0, -1, 0, 0, -2, 0, -2, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 2, 3, 3, 2, 2, -3, -2, 0, -1, 0, -1, 0, 0, 0, 0, -2, -2, -1, -1, -2, -1, -1, -1, 0, 1, 0, 0, 1, 3, 2, 2, -4, -3, -2, -2, 0, -1, -1, 0, -1, -1, -1, -2, -1, -1, -2, 0, -2, -1, 0, 0, 0, 0, 1, 2, 2, 2, -4, -2, -1, -1, 0, -2, -2, -1, -2, 0, -1, -1, -2, -1, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -5, -3, -2, -1, 0, 0, -1, -1, 0, -2, -1, -1, -3, 0, 0, -2, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, -5, -3, -2, -2, 0, -1, 0, 0, -2, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, -4, -4, -2, 0, 0, 0, 0, -1, -1, 0, -2, 0, -2, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -3, -3, -2, -1, 0, -1, 0, -1, -1, -2, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -4, -2, 0, 0, -1, 0, 0, -3, -1, -1, -2, -3, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, -4, -1, 1, 0, 0, -1, 0, -1, -1, -1, -3, -1, -2, -2, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 1, -2, -2, 1, 0, 0, -2, -2, -2, 0, -2, -1, -3, -2, 0, 0, 1, 0, 0, -1, 0, -1, 0, -2, -2, 0, 0, -3, -2, 0, 0, 0, -1, -1, -1, -1, -1, -3, -2, -2, -1, 0, 0, 0, 0, -1, 0, -1, -2, -1, -2, 0, 0, -2, -2, 0, 0, 0, -2, -1, -1, -3, -2, -3, -2, -2, -2, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, -2, 0, -1, 0, 0, 0, -2, -2, -1, -2, -3, -2, -2, -2, 0, 0, -1, -1, 0, -1, -2, -1, 0, 0, 1, 1, -1, 0, 1, 0, 0, -1, -1, -1, -2, -3, -2, -2, -1, -1, -1, -1, -2, -2, -1, -3, -2, -2, 0, 0, 0, 2, 0, 0, 1, -1, 0, -1, -1, -2, -1, 0, -1, -2, -2, -1, -1, -3, -1, -1, -1, -1, -1, -1, 0, 0, 1, 0, -1, 1, 0, 0, -1, -1, 0, -1, -1, 0, 0, -3, -2, -2, -2, -2, -3, -3, -1, -1, -2, 0, 1, 0, 0, 2, -1, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, -3, -4, -3, -4, -3, -3, -1, -1, 0, 1, 1, 0, 2, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, -3, -1, -3, -2, -1, 0, 0, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, 1, 1, 2, 3, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 2, 2, 2, 3, 4, 4, 4, 0, 0, 1, 0, 0, 0, 0, 0, 2, 1, 2, 1, 2, 3, 2, 2, 1, 1, 2, 2, 3, 4, 2, 3, 2, 3, 0, 0, 0, 1, 1, 0, 2, 2, 1, 2, 3, 4, 4, 2, 3, 1, 3, 2, 1, 1, 1, 1, 3, 3, 2, 2, 1, 2, 1, 2, 3, 3, 3, 1, 4, 2, 3, 3, 3, 4, 2, 1, 0, 0, 1, 1, 2, 1, 1, 1, 1, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, -1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, -1, 0, -1, -1, 0, -1, 0, 0, -1, -1, -1, 0, 1, 0, 1, 2, -1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 2, 0, 0, -1, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -2, 0, -1, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 2, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -2, -1, -2, -1, -1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 2, 0, 0, 0, 1, 1, 0, -1, -1, -1, 0, -1, -2, -1, -2, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 0, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, -1, -1, -2, -1, -1, -1, -1, 0, 1, 0, 0, 1, 0, 0, 2, 1, 2, 0, 1, 1, 2, 0, 0, 0, 0, -1, -2, -1, -1, -2, -1, -1, -1, 0, 0, 0, 1, 1, 0, 1, 2, 1, 2, 0, 0, 2, 2, 1, 1, 0, 0, -1, -2, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 2, 1, 0, 2, 0, 0, -1, -2, -2, -2, -2, -2, -2, -1, 0, 0, -1, 0, -1, 0, 1, 0, 2, 3, 1, 1, 2, 1, 0, 2, 0, 0, -2, -1, -1, -3, -2, -1, -2, -1, -2, 0, -2, 0, 0, -1, 0, 1, 1, 2, 0, 1, 1, 1, 0, 1, 0, -1, 0, 0, -3, -2, -4, -2, -2, -2, -1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 1, 0, 2, 0, 1, 1, 0, -1, 0, -1, -4, -2, -3, -2, -3, 0, 0, -1, 0, 0, 0, 2, 0, 3, 2, 1, 1, 1, 0, 2, 1, 0, 0, 0, -1, -3, -3, -3, -4, -3, -2, -1, 0, 0, 0, 0, 0, 1, 2, 2, 3, 0, 1, 0, 1, 1, 0, 0, -1, -1, 0, -2, -1, -3, -2, -3, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 3, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -3, -2, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 3, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, -2, -1, -3, -1, 0, 0, 0, 2, 1, 1, 1, 0, 2, 1, 2, 2, -2, -1, -1, 0, 0, 0, 0, 0, -1, -2, -1, -2, -2, 0, 0, 1, 1, 2, 0, 2, 0, 0, 0, 0, 1, 2, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -2, 0, 0, 0, 1, 2, 1, 1, 1, 1, 0, 2, 1, 2, 2, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 1, 2, 2, 3, 1, 1, 2, -1, 0, -1, 0, -1, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 2, 2, 3, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 2, 2, 1, 4, 4, 6, 7, 7, 6, 7, 5, -1, -2, 0, 0, 0, -2, 0, -2, -1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 3, 3, 5, 5, 5, 4, 3, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 3, 3, 2, 3, 4, -2, -2, -2, 0, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 2, 3, 2, 3, -1, -3, 0, -1, 0, -1, 0, -2, -2, -3, 0, -1, -2, 0, -2, 0, -1, -1, 0, 0, 0, 1, 0, 1, 1, 1, -3, -2, -1, -2, -1, -1, -1, 0, -3, -2, -3, -1, -1, -1, -1, -2, -1, 0, 0, -1, -1, -1, -2, -1, -1, -1, -1, -4, -4, -3, -2, -2, 0, -2, -1, -4, -3, -4, -2, -1, -1, -2, 0, -1, -2, -2, -1, -1, -3, -3, -2, -1, -2, -4, -4, -4, -3, -3, -1, -2, -2, -3, -4, -2, -3, -3, -1, -1, 0, 0, 0, -2, -1, -3, -1, -3, -3, -1, -4, -2, -3, -2, -2, -3, -1, -1, -3, -2, -3, -4, -4, -2, -1, 0, -2, -1, -1, -1, -2, -3, -1, -4, -1, -2, -2, -3, -1, -1, -1, -2, -2, -3, -2, -1, -3, -3, -2, -2, -2, -1, -1, -2, -1, -1, -2, -1, -3, -2, -1, -1, -2, -3, -2, -2, 0, 0, 0, -2, -2, -2, -1, -3, -2, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -2, 0, 0, -1, 0, -1, -1, -2, 0, -2, 0, -1, -1, 0, 0, 1, 0, 0, 1, 1, 0, -1, -1, 0, -2, -2, -1, 0, -1, 0, -1, -2, -2, -3, -1, -3, -2, 0, -1, 0, 1, 0, 0, 1, 0, 1, 0, -1, 0, 0, -3, -2, -1, -1, -2, 0, -2, -2, -3, -3, -3, -2, -2, 0, 0, -1, 0, 0, -1, -1, -2, 0, -1, -1, -1, 0, -2, -1, -1, -1, 0, -1, -2, -2, -2, -3, -3, -1, 0, -1, 0, 0, -1, -2, -1, -1, -1, -1, -1, 0, -2, 0, -2, -2, 0, -3, -2, -2, -2, -2, -3, -3, -2, -2, -1, 0, -1, 0, -3, -1, -3, -3, -3, -1, -1, -2, 0, -1, -2, -2, 0, -1, -3, -1, -4, -3, -5, -3, -4, -1, -2, -1, -1, -2, -2, -2, -2, -2, -2, -2, -1, 0, -1, 0, 0, -1, 0, -1, -3, -2, -4, -4, -6, -3, -4, -3, 0, -2, -2, -2, -3, -2, -3, -3, -3, -2, -1, 0, 0, -1, 0, 0, 0, -1, -2, -2, -3, -4, -3, -4, -2, -3, 0, -2, -1, -2, -4, -4, -2, -3, -3, -3, -1, -1, -1, -1, 1, 1, 0, -2, -3, -2, -3, -3, -3, -3, -1, 0, -2, -1, -2, -4, -3, -4, -4, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -4, -3, -2, -3, -1, -1, -1, -3, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, -3, -2, -1, -2, -1, -1, -1, -2, -3, -2, -3, -1, -3, -1, 0, -1, -1, 0, 1, 2, 3, 1, 0, 0, -2, -2, -2, -1, -1, -3, 0, -1, -2, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 1, 2, 2, 3, 1, 0, 0, 0, -1, -2, -1, -1, -2, -1, 0, 0, -1, 0, 0, 1, 1, 2, 2, 2, 1, 0, 0, 1, 2, 1, 3, 1, 0, 1, -1, -2, -2, -2, -1, 0, 0, 0, 0, 2, 0, 2, 2, 3, 3, 3, 1, 1, 1, 1, 2, 3, 4, 2, 3, 1, 2, 0, 0, 0, 0, 0, 0, 0, 2, 3, 4, 3, 4, 4, 4, 5, 4, 2, 1, 2, 4, 3, -8, -7, -4, -4, -4, -2, -3, -2, -3, -1, -3, -3, -4, -4, -4, -3, -3, -3, -5, -4, -5, -4, -5, -4, -4, -5, -7, -5, -3, 0, 0, -1, 0, -2, -1, 0, -3, -2, -2, -2, -1, -3, -3, -1, -2, -2, -2, -2, -2, 0, -1, -3, -4, -2, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -4, -2, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 2, 0, -3, 0, -1, -1, 1, 0, 0, 1, 1, 1, 1, 1, 2, 2, 0, 1, 1, 1, 0, 2, 0, 0, 2, 2, 2, 1, -4, -1, 0, 0, 0, 0, 1, 1, 2, 2, 2, 0, 0, 0, 2, 1, 1, 1, 1, 0, 0, 2, 3, 2, 3, 3, -1, -1, 1, 1, 1, 1, 1, 2, 1, 0, 0, 0, 0, 1, 1, 3, 2, 2, 0, 0, 1, 2, 2, 2, 3, 2, 0, 0, 3, 3, 2, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 3, 3, 2, 1, 2, 1, 1, 2, 2, 0, 1, 2, 5, 2, 2, 0, -1, -1, 0, 0, -1, -1, 0, 1, 1, 1, 1, 1, 2, 3, 2, 2, 3, 2, 2, 0, 3, 5, 4, 3, 2, 0, 0, 0, 0, -1, -2, 0, 0, 1, 2, 1, 2, 2, 0, 1, 1, 1, 2, 2, 2, 2, 5, 5, 4, 4, 4, 1, 1, -1, -1, -2, -1, 0, 1, 2, 2, 1, 0, 1, 0, 0, 0, 2, 2, 2, 2, 1, 4, 5, 4, 4, 2, 2, 1, 1, 0, 0, -1, 0, 0, 1, 1, 1, 1, 0, 1, 0, 2, 2, 1, 0, 0, 1, 3, 6, 5, 4, 2, 2, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 5, 4, 5, 4, 3, 2, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 0, 0, 3, 4, 4, 2, 4, 1, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 3, 1, 1, 1, 0, 3, 3, 3, 4, 3, 2, 2, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 2, 3, 3, 3, 2, 0, 0, 1, 3, 3, 2, 2, 2, 3, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 2, 2, 2, 2, 0, 0, 1, 3, 2, 2, 3, 2, 1, 0, 1, 0, -1, 0, 0, 0, 2, 1, 2, 1, 0, 1, 1, 3, 1, 1, 0, -2, 1, 0, 3, 4, 2, 1, 1, 2, 0, 1, 0, 1, 0, 1, 1, 0, 0, 1, 0, 1, 1, 1, 1, 2, 1, -2, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, -4, -3, -2, 1, 1, 0, 0, 0, 0, 0, 1, 1, 2, 0, 2, 1, 0, 2, 1, 0, 2, 2, 1, 2, 0, 0, -6, -4, -2, 0, 0, 2, 0, 0, 0, 0, 1, 0, 0, 0, 2, 1, 1, 2, 2, 2, 2, 3, 2, 1, 0, 0, -8, -5, -4, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 2, 2, 1, 2, 3, 3, 2, 1, 0, 0, -1, -9, -5, -4, -2, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, -1, -1, -10, -8, -4, -3, -3, -1, -1, -2, -1, -1, 0, 0, -2, 0, -1, 0, 0, -2, 0, -1, 0, -1, -1, -3, -3, -2, -9, -8, -8, -5, -4, -4, -4, -2, -2, -1, -1, -1, -3, -2, -4, -4, -4, -4, -3, -5, -3, -6, -5, -6, -4, -4, 2, 2, 3, 2, 2, 3, 1, 2, 1, 2, 1, 1, 2, 3, 1, 0, 2, 1, 0, 0, 1, 1, 2, 0, -2, -3, 3, 2, 1, 1, 2, 0, 1, 2, 2, 1, 0, 1, 2, 1, 2, 1, 0, 0, 1, 2, 2, 0, 0, 0, 0, -2, 4, 2, 1, 1, 2, 1, 1, 1, 0, 1, 0, 1, 1, 0, 0, 2, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 1, 0, 0, 2, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, -1, 0, -2, 0, 3, 1, 1, 0, 0, 1, 1, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -2, -2, -1, 4, 1, 2, 1, 1, 1, 1, -1, 0, 0, -2, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, -2, 0, -2, -2, 2, 1, 0, 0, 0, 1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -3, -3, 2, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, -3, -1, -1, -2, -1, -1, 2, 2, 2, 0, 0, -1, -2, -2, -2, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, 3, 2, 0, 1, 0, -2, -2, -4, -1, 0, -1, 1, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -2, -1, 1, 1, 1, 0, -1, -1, -3, -4, -2, -3, -1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, -1, 2, 1, 1, 0, -1, -1, -2, -4, -4, -3, -1, -1, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 3, 1, 0, 0, 0, -2, -1, -1, -3, -2, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -2, 4, 1, 1, 0, 0, -1, -3, -3, -3, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -2, 4, 0, 0, 0, -1, 0, -1, -3, -4, -2, -2, -1, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, 0, 0, -2, -3, 0, 1, 0, 0, -1, -1, -1, -2, -2, -2, -2, -2, -1, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -3, 0, 0, -1, -1, 0, -1, -2, -2, -3, -3, -3, -2, -1, 1, 2, 1, 1, -1, -1, 0, -1, -2, -1, 0, -1, -2, 0, 0, 0, 0, 0, -1, -2, -2, -4, -3, -3, -2, 0, 2, 2, 0, 1, 0, 0, -1, -2, -1, -2, -2, -2, -2, 0, 0, 0, 0, 1, 0, -1, -1, -3, -1, -1, 0, 0, 2, 1, 1, -1, 0, 0, -1, -2, 0, -1, -1, -2, -2, 1, 0, 1, 1, 0, 0, 0, -2, -2, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -2, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -2, -4, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, -1, -1, -2, -3, 1, 2, 3, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, -1, -2, -4, 2, 3, 3, 2, 0, 0, -1, 0, 0, 0, 0, 2, 0, 2, 0, 1, 0, 1, 1, 1, 2, 0, 0, 0, 0, -2, 3, 2, 2, 1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 2, 0, 0, 1, 0, 2, 2, 1, 1, 0, -1, -1, 4, 2, 4, 2, 1, 1, 0, 0, 1, 0, 0, 2, 1, 2, 1, 2, 1, 0, 1, 0, 2, 1, 0, 0, 0, -3, -4, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 1, 1, 0, 0, 0, 1, 2, 3, 4, 3, -4, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 2, 3, 3, 3, -4, -3, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 2, 1, 2, 3, 4, 4, 3, -3, -2, -2, -1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 2, 1, 3, 4, 2, -5, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 2, 3, 3, 3, 2, -5, -3, -3, -1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 1, 1, 1, 0, 1, 1, 1, 4, -6, -3, -2, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 2, 1, -4, -3, -2, 0, 0, 0, 1, 0, 2, 1, 1, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 3, -5, -2, -1, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, -4, -2, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, -4, -1, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 3, 1, 1, -1, -1, -1, -1, 0, 0, 0, -3, 0, 1, 0, 1, 0, 0, -1, -1, -1, -1, -1, -2, -1, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -3, 0, 2, 1, 2, 0, 1, 0, 0, 0, -1, -1, 0, -2, 0, 1, 1, 1, 0, -1, -1, 0, 0, -2, 0, 0, -1, 0, 2, 1, 0, 1, 0, 1, 0, -1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 1, -2, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, -1, -1, -2, -1, 0, -1, 0, 0, 1, -1, 0, 0, 1, 0, 1, 2, 0, 1, 1, -1, -1, -2, -2, -2, 0, -1, -1, -2, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 1, 1, 2, 1, 1, 1, 1, 0, -2, -2, -1, -2, -1, -1, -2, 0, -1, 0, -1, 0, 0, 0, 0, -2, 1, 2, 1, 2, 0, 3, 2, 1, 0, 0, 0, -1, -1, -3, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 2, 2, 3, 0, 1, 2, 1, 1, 0, -1, -2, -2, -1, -3, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, -2, 0, 1, 1, 3, 2, 2, 2, 0, 1, 1, 0, -1, -1, 0, -3, -1, -1, 0, 0, 0, 1, 0, 2, 2, 2, -1, 0, 0, 2, 1, 1, 1, 0, 0, 1, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 4, 2, -2, 0, 0, 1, 1, 2, 1, 1, 1, 2, 0, 2, 0, 0, 1, 0, 0, 0, 0, 1, 3, 3, 2, 4, 3, 3, -1, -1, 0, 1, 0, 1, 2, 2, 3, 2, 3, 1, 1, 2, 2, 1, 1, 1, 2, 2, 2, 4, 4, 2, 3, 3, -1, 0, 0, 1, 0, 2, 1, 2, 2, 2, 2, 2, 1, 2, 2, 0, 1, 2, 2, 4, 4, 5, 5, 4, 2, 2, -1, 0, 0, 0, 1, 2, 2, 3, 4, 3, 2, 3, 1, 3, 2, 1, 2, 2, 3, 2, 3, 4, 1, 3, 1, 1, -1, 0, 0, 0, 1, 0, 2, 3, 2, 3, 2, 3, 1, 1, 2, 2, 0, 1, 0, 1, 0, 2, 2, 1, 1, 1,
    -- filter=0 channel=6
    -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 2, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 2, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, 1, -1, -1, 0, 0, 0, -1, 0, 0, 2, 1, 0, 1, 1, 2, 0, 2, 2, 1, 1, 1, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -2, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -1, -1, 0, -1, -1, -1, 0, 0, -1, 1, 0, 0, 0, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, -2, -1, -2, -2, 0, -1, 0, -2, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -2, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, -1, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -2, -1, -2, 0, 0, 0, -1, -1, -1, 0, -1, -2, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, -2, 0, 0, 0, -1, 0, -1, 0, 0, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 1, 0, -1, -1, -2, 0, -2, -1, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, 0, -1, 0, 0, 0, -1, -3, -1, -2, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, -2, -2, -1, -1, -1, -2, -2, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -2, 0, 0, -1, 0, -1, 0, -1, -1, -2, -1, -2, -1, 0, -2, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, -2, 0, -2, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, -2, -1, -1, 0, -1, 0, -1, 0, -1, 0, -2, -2, -1, -2, -2, 0, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, 0, -1, 0, -3, 0, 0, 0, 0, -1, -3, -3, -1, -2, 0, -2, -2, -1, -1, -2, 0, -1, 0, 0, -1, 0, -2, 0, -1, -1, -2, 0, 0, 0, -2, 0, 0, 0, -1, -1, -2, -1, -3, -2, -2, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -2, 0, 0, 0, 0, -2, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -2, -2, -1, -1, 0, 0, 0, -1, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 2, 2, -1, 0, -1, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 3, 1, 0, 0, -1, 0, 1, 1, 0, -1, -1, -3, -2, -2, -2, 0, 2, 0, 0, 1, 0, 0, -1, 0, 1, -1, 0, 2, 1, 0, 0, 0, 1, 0, 0, -1, -1, 0, -2, -2, 0, 1, 1, 1, 1, 1, 1, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 3, 2, 1, 0, 0, 0, 1, 2, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 1, 2, 2, 0, -1, 1, 1, 2, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 1, 2, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 3, 2, 2, 3, 1, 2, 0, 1, 0, 1, 0, 1, 3, 3, 2, 0, -1, -2, 0, 0, 1, 1, 0, 1, 3, 2, 2, 4, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 1, 2, 1, 0, 0, -1, -1, -1, -1, 0, 0, 2, 3, 3, 4, 4, 3, 2, 1, 2, 0, 0, 0, 0, 0, 2, 2, 2, 1, 1, -1, -1, 0, 0, 0, 0, 1, 4, 2, 3, 2, 2, 3, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, 3, 3, 4, 5, 2, 3, 2, 0, 2, 0, 1, 2, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, -1, -1, 0, 1, 2, 3, 3, 3, 2, 3, 1, 1, 2, 0, 2, 2, 1, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 2, 4, 3, 4, 4, 2, 2, 0, 3, 2, 2, 2, 1, 0, 0, 1, 1, 1, 2, 0, -1, 1, 0, 0, 2, 2, 3, 5, 4, 3, 4, 1, 1, 1, 2, 2, 2, 0, 1, 1, 0, 3, 2, 3, 1, 0, -1, 1, 1, 1, 1, 2, 4, 4, 5, 4, 2, 3, 1, 2, 3, 3, 2, 0, 0, 0, 0, 1, 3, 2, 2, 0, 0, 0, 1, 2, 2, 3, 5, 5, 4, 3, 2, 2, 3, 4, 2, 2, 2, 1, 0, 0, 1, 2, 3, 2, 2, 1, 1, 1, 1, 2, 1, 2, 5, 3, 4, 4, 1, 3, 2, 2, 2, 2, 2, 0, 0, 0, 0, 3, 3, 4, 4, 1, 0, 0, 0, 2, 0, 1, 2, 4, 2, 2, 1, 2, 2, 0, 0, 1, 0, 1, 0, 1, 3, 2, 5, 2, 2, 1, 0, 0, 1, 1, 0, 2, 2, 5, 2, 3, 2, 1, 0, 0, 0, 0, 0, 0, 1, 2, 3, 3, 4, 1, 0, 0, 0, 1, 0, 0, -1, 2, 2, 4, 3, 2, 1, 0, 1, 0, 0, 0, 1, 1, 1, 3, 3, 1, 1, 1, 0, 0, -1, 1, 0, -1, 0, 2, 3, 3, 3, 0, 1, 2, 0, 0, 0, 0, 0, 3, 2, 3, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 1, 0, -1, 0, 1, 3, 1, 2, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 3, 1, 2, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 2, 1, -1, -1, -1, 0, 0, -2, 0, 0, 0, 0, 2, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 1, 2, 0, 0, 0, 0, 0, -1, 0, -2, 0, 1, 1, 2, 2, 1, 1, 1, 2, 3, 1, 1, 0, 0, -1, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, -2, -1, 0, 2, 1, 2, 1, 1, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -2, -2, -3, 0, 0, 0, 1, 1, 1, 2, 3, 1, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, -1, -1, 0, 0, -1, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -2, -2, 0, -1, -1, -1, 0, -1, -2, -2, -1, -1, 0, 0, -2, -1, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, 0, -2, -2, -1, -2, -1, -1, -1, -2, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -2, -1, 0, -1, -1, 0, -1, 1, 0, 1, 1, 1, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 1, 1, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, 0, -1, 0, -1, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 2, 1, 0, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 0, 1, 1, 0, 2, 2, 2, 3, 2, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 2, 2, 1, 1, 1, 1, 1, 2, 1, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 2, 0, 0, 1, 0, 0, 0, 1, 0, -1, 1, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 1, 0, 2, 1, 2, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -2, 0, 0, -2, -1, -2, -1, -2, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -2, 0, -2, -2, 0, -2, -1, -1, -3, -2, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -2, -2, -1, -3, -1, -2, -2, 0, -2, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, 0, -1, -2, -2, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 1, 0, 2, 2, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -2, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -2, -2, -1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -2, -1, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, -1, -1, -2, -2, -3, 0, -2, -1, -2, -2, 0, 0, 1, 1, 0, 1, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -3, -2, -2, -1, -1, -1, 0, 0, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -2, -1, -1, 0, 0, 0, 1, 2, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, -1, -2, -1, -2, -2, -1, -1, -1, -1, 0, 0, 1, 2, 1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, -2, -1, -2, -2, -2, -2, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -2, 0, -2, -2, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 1, 1, 2, 1, 1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 2, 0, 0, 1, 0, -1, 0, 0, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 1, 0, 0, 2, 1, 2, 0, 0, 1, 0, 2, -1, 0, -1, -1, 0, -1, 0, 0, 2, 1, 1, 1, 0, 0, 1, 0, 1, 1, 0, 1, 1, 1, 1, 2, 2, 1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 3, 2, 1, 1, 0, 0, 0, 0, -1, -1, -2, -3, -2, -2, -4, -2, -1, 0, -1, 0, 0, -1, -2, 0, -1, -3, 2, 1, 0, 0, -1, -1, 0, -1, -1, -1, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, -1, -2, -2, -1, 4, 1, 0, 0, 0, 0, -1, 0, -2, -2, 0, -2, 0, -1, 0, 0, 0, 2, 0, 0, 0, -1, 0, -1, 0, -1, 4, 1, 2, 1, 0, 0, -1, -1, -2, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 2, 2, 1, 1, 0, 0, -1, -2, -1, -2, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 3, 1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, -2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, -2, 1, 1, 1, -1, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, -1, 0, -1, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 3, 2, 1, 1, 0, 0, 0, -1, -2, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 4, 4, 2, 3, 3, 2, 1, 0, 0, 0, -2, -3, -3, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, 1, 3, 4, 4, 5, 3, 1, 1, 1, 0, 0, 0, -1, -1, -3, -2, -1, 0, 0, 0, -1, 1, -1, 0, 1, 1, 2, 4, 5, 5, 5, 4, 2, 1, 1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 3, 4, 6, 6, 4, 4, 1, 0, 1, 1, -1, 0, 0, -1, -3, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 4, 4, 6, 4, 5, 4, 3, 0, 1, 0, 0, 0, -1, -1, -2, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 2, 4, 5, 6, 4, 4, 2, 2, 0, 0, 1, 0, -1, -1, -2, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 3, 3, 4, 4, 4, 5, 1, 1, 1, -1, 0, 0, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 2, 1, 2, 2, 3, 3, 5, 5, 3, 4, 3, 0, 0, 0, -1, -1, -1, -1, 0, -1, 1, 2, 0, 0, 0, -1, 2, 1, 1, 2, 2, 3, 3, 3, 4, 3, 1, 0, -1, -1, -2, -2, -2, -3, 0, -1, 0, 1, 0, 0, 0, 0, 3, 3, 1, 2, 0, 2, 3, 2, 2, 2, 0, 0, -2, -2, -1, -2, -3, -2, -1, 0, 0, 2, 1, 0, 0, -1, 3, 1, 2, 0, 0, 0, 0, 3, 0, 1, 0, 0, -1, -3, -2, -3, -3, -2, 0, 0, 1, 1, 0, 0, -1, -3, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -2, -4, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 3, 0, 0, 0, -1, -1, 0, 0, -2, -2, -1, -3, -3, -2, -3, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 2, 1, 0, 0, 0, 0, -1, -2, -1, -2, -2, -3, -3, -1, 0, -1, -1, 1, 1, 0, 0, 0, 1, 0, 0, -1, 3, 1, 1, 0, 0, -1, 0, 0, -1, -3, -4, -1, -2, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, -2, -2, -2, -3, -2, -1, -1, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 3, 2, 1, 0, 1, 0, 0, 0, -3, -4, -3, -4, -2, -1, 0, 0, 2, 0, 0, 0, 0, 0, 1, 0, 1, 2, 8, 5, 4, 2, 3, 1, 1, 1, -2, -2, -3, -6, -6, -6, -4, -3, -2, 0, 0, 0, 0, 2, 3, 2, 3, 1, 5, 3, 2, 2, 1, 1, 0, 0, -1, -3, -5, -5, -5, -6, -3, -2, -1, 0, 0, 1, 0, 0, 3, 4, 4, 1, 4, 1, 2, 1, 0, 0, 1, 0, -1, -4, -5, -4, -3, -4, -2, -1, -1, 0, 0, 1, 0, 0, 0, 2, 2, 1, 1, 2, 0, 1, 0, 0, 0, -1, 0, -3, -4, -2, -3, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 2, 0, 0, 1, -1, -1, -1, 0, -2, -2, -4, -2, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, -2, -2, -2, -1, -2, -1, -1, -1, -1, 0, 0, -1, 0, -1, -1, 0, 1, 0, 0, -3, -3, 1, 0, -1, -1, -1, -3, -3, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -1, 0, 0, 0, -1, -3, -5, 1, 0, -1, 0, -1, 0, -1, 1, 0, 1, 3, 2, 0, 1, 0, 0, -1, -2, -3, -3, -2, 0, -1, -1, -3, -7, 2, -1, 0, 0, 0, 0, 3, 1, 2, 3, 4, 3, 3, 3, 2, 1, 0, -2, -3, -4, -2, -2, -2, -1, -2, -5, 0, -1, -2, 0, 1, 2, 5, 6, 6, 7, 6, 5, 4, 5, 5, 3, 0, -2, -3, -3, -4, -3, -3, -1, -2, -5, -1, -1, -2, 0, 2, 3, 5, 8, 8, 8, 9, 9, 8, 8, 6, 5, 2, -1, -3, -4, -4, -4, -2, -2, -3, -5, -1, 0, 0, 0, 3, 5, 6, 7, 8, 9, 10, 9, 9, 7, 9, 8, 5, 0, -2, -3, -3, -3, -2, -3, -4, -5, -1, -1, -1, 1, 3, 3, 6, 7, 6, 9, 9, 7, 9, 7, 7, 7, 4, 0, -2, -4, -3, -2, -2, -2, -2, -4, -2, -2, 0, 0, 2, 6, 6, 6, 8, 9, 8, 9, 7, 7, 6, 7, 3, 0, -2, -6, -3, -1, 0, 0, -1, -2, -2, -1, 0, 1, 3, 4, 8, 7, 7, 7, 6, 7, 7, 6, 8, 6, 4, 0, -2, -5, -4, -2, 1, 0, 0, -1, -3, 0, 1, 1, 1, 4, 6, 8, 6, 5, 5, 4, 5, 7, 6, 5, 2, 0, -1, -2, -3, -1, 0, 0, 0, 1, -1, 0, 0, 0, 2, 4, 7, 6, 4, 4, 5, 5, 3, 3, 3, 4, 1, 1, -1, -1, -1, 0, -1, 0, 2, 0, -1, 0, 2, 1, 0, 5, 7, 7, 4, 4, 3, 4, 3, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 3, 4, 5, 4, 1, 1, 0, 0, -1, -2, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, -2, 0, -1, 0, 0, 1, 2, 0, 0, 0, 0, -1, -2, -5, -5, -3, -1, 0, 0, 0, -1, -1, -1, 0, -3, 0, -3, -2, -1, -1, 0, 0, -1, -1, -1, -2, -3, -4, -4, -6, -6, -1, 0, 0, 0, -1, 0, -1, -2, -2, -1, -1, -3, -4, 0, -1, 0, -2, -3, -3, -3, -5, -5, -7, -5, -6, -3, -1, 0, 1, 1, 1, 1, 0, 0, 0, -2, 0, 0, -3, -2, 0, -1, -2, -3, -5, -5, -4, -7, -7, -8, -6, -5, -2, 0, 1, 0, 1, 1, 1, 2, 1, 0, 1, 0, -1, 0, 0, -1, -1, -4, -4, -6, -6, -7, -7, -6, -5, -2, 0, 0, 0, 1, 1, 2, 3, 2, 2, 1, 3, 0, 0, 0, 0, 0, 0, -4, -4, -6, -6, -6, -7, -5, -6, -2, 0, 0, 0, 2, 2, 2, 3, 4, 3, 1, 3, 2, 0, 1, 1, 2, 1, 0, -4, -6, -5, -6, -7, -5, -5, -5, -1, 0, 1, 0, 1, 2, 3, 2, 1, 2, -4, -2, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 2, 0, 0, 1, 0, 2, 3, 3, 5, 5, 5, 8, -4, -1, -1, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 3, 4, 5, -3, -2, 0, 0, 0, 0, -1, -1, -2, -2, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 2, 1, 3, 4, -3, -2, -1, 0, 0, 0, 0, 0, -1, -2, -2, -2, -2, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 2, 3, 2, -2, -2, 0, 0, -1, 0, 0, -1, -1, -3, -2, -3, -2, -1, -2, -3, 0, 0, -2, 0, 0, 0, 0, 0, 1, 2, -2, 0, 0, 0, -1, 0, -2, -1, -1, -2, -2, -2, -2, -3, -2, -3, -1, -3, -1, -1, 0, 0, 0, -1, 0, 1, -1, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, -2, -3, -4, -1, -3, -1, -1, 0, -1, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -2, -2, -2, -3, -2, -3, -3, -2, -1, 0, -1, 0, 0, 0, -3, -1, -1, -1, 0, -1, 0, -2, -1, 0, -1, 0, 0, 0, -1, -2, -1, -3, -2, -2, -2, -1, 0, 1, 0, 1, -1, 0, 0, -1, 0, 0, 0, -2, -1, -1, -1, -1, 0, -1, -2, -2, -3, -3, -3, -3, -3, -1, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, -1, -1, -1, -2, -1, 0, -1, -1, -2, -3, -1, -3, -3, -4, -2, -1, 0, 0, 0, 1, 0, 2, 1, 0, -1, -1, -1, -1, -2, -2, 0, -1, 0, 0, -1, -1, -1, -3, -1, -3, -2, -2, -1, 0, 0, 1, 0, 2, 2, 1, 0, -2, -1, -3, -2, -1, 0, -1, -1, -1, -1, -2, -1, -1, -2, -2, -4, -2, -1, 0, 0, 0, 1, 2, 3, 1, 0, 0, -2, -3, -2, -3, -1, -1, 0, 0, -1, -2, -1, 0, 0, -3, -2, -3, -2, 0, 0, 0, 0, 0, 2, 0, 0, -2, -3, -2, -2, -2, -3, -3, -1, -2, -2, -1, -1, 0, -1, -2, -3, -4, -1, -1, 0, 0, 0, 0, 1, 1, 0, -2, -3, -3, -3, -3, -3, -1, -2, -3, -3, -1, -1, 0, 0, -2, -4, -2, -1, 0, 0, 0, -1, 0, 1, 0, 0, -2, -2, -3, -2, -1, -3, -2, -2, -1, -3, -1, 0, 0, 0, -3, -2, -2, 0, 0, 0, 1, -2, 0, 2, 1, 0, -1, -1, -2, -2, -2, -1, -2, -1, -3, -2, -2, 0, 0, 0, -1, -2, -1, 0, 0, 1, 1, -3, 0, 0, 0, -2, -2, -2, -3, -3, -3, -2, -3, -4, -2, -3, -1, -1, 0, 0, 0, -1, -2, -1, -1, 1, 1, -4, -1, 0, 0, 0, -2, -3, -2, -3, -3, -3, -2, -3, -3, -4, -3, -1, 0, 0, 0, -1, -1, 0, 0, 0, 2, -3, 0, 0, 0, 0, 0, -3, -2, -1, -2, -3, -2, -3, -2, -3, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -3, -2, -4, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 2, 3, -3, -1, 0, 0, -1, 0, 0, 0, -1, -2, -1, -3, -2, -3, -2, -1, -1, 0, 0, 0, 0, 0, 1, 1, 2, 3, -2, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 5, 4, -3, -1, 0, 0, 0, 0, 0, -2, -1, -2, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, -1, 1, 1, 2, 3, 5, -4, -2, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 3, 4, 5, 5, 0, 1, 1, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -1, -2, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, -1, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -2, 0, 0, 0, -1, 0, -2, -2, -1, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, -1, -1, 0, 0, 0, 1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, 2, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 1, 1, 0, 1, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 1, 1, 1, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 2, 0, 1, 2, -3, 0, 1, 3, 0, 0, 0, 0, 1, 1, 0, 1, 1, 2, 1, 1, 2, 3, 4, 4, 6, 7, 8, 8, 9, 9, -2, 0, 1, 0, 1, 2, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 2, 2, 2, 4, 3, 5, 6, 7, 6, -1, -1, 0, 1, 1, 1, 0, 1, 0, -2, -1, -3, -1, -2, -2, 0, 0, 0, 0, 1, 1, 1, 1, 4, 4, 5, -3, -2, 0, 0, 0, 0, -1, 0, -2, -3, -4, -2, -2, -2, -2, -2, -2, 0, 0, 0, 0, 0, 1, 1, 2, 4, -4, -1, 0, 0, 0, -1, -1, -2, -4, -3, -5, -3, -3, -4, -2, -4, -3, -2, -1, -1, -1, 0, 0, 0, 2, 3, -4, -2, -1, 0, 0, -2, -2, -1, -2, -4, -4, -4, -3, -3, -5, -3, -3, -3, -1, -1, 0, 0, 0, 0, 0, 0, -4, 0, -1, 0, -1, -2, -2, -4, -4, -2, -1, -3, -3, -4, -5, -3, -5, -4, -2, 0, 0, 0, 0, 0, -1, 1, -2, 0, 0, 0, 0, -2, -2, -3, -2, -1, 0, -2, -3, -2, -4, -3, -3, -2, -2, -3, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, -2, -2, -3, -2, -1, 0, 0, -1, -1, -2, -4, -4, -3, -3, -2, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 1, 1, 0, -1, -1, -2, -3, -4, -4, -2, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, 0, -2, -4, -5, -3, -3, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -3, 0, 0, 0, 0, 0, -1, -1, 0, -1, -2, -2, -4, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, -2, -2, -3, -1, -1, -2, 0, 0, 0, 0, -1, -1, 0, 0, -1, -2, -3, -2, -1, 0, -1, 1, 2, 1, 0, -1, -3, -2, -4, -4, -2, -3, 0, 0, 0, -1, 0, 0, 0, -1, -2, -4, -4, -3, -2, -1, -2, 0, 1, 2, 1, -1, -3, -4, -3, -3, -4, -2, -2, -1, 0, -1, 0, 0, 1, 0, -2, -2, -2, -3, -2, -2, -2, 0, 0, 1, -1, -1, -3, -4, -4, -4, -2, -2, -1, 0, 0, 0, 1, 2, 1, -1, -3, -5, -4, -4, -3, 0, -1, -1, 0, 0, 0, -1, -1, -4, -2, -4, -2, 0, 0, -1, -1, -2, 0, 0, 1, -1, -2, -3, -2, -2, -2, 0, 0, -1, 0, 0, 0, -1, -2, -3, -4, -2, -2, -2, 0, -2, 0, -2, -2, -1, -1, -1, -1, -2, -2, -2, 0, 1, 1, -3, -1, 1, 0, -2, -1, -3, -2, -4, -3, -2, -3, -2, -2, -2, -2, -2, -1, -1, -2, -1, -2, 0, 0, 0, 1, -2, -1, -1, 0, -1, -3, -4, -4, -3, -4, -3, -4, -5, -4, -3, -2, -2, -1, -2, -1, -1, -1, 0, 0, 1, 2, -3, 0, 0, 0, -1, -2, -4, -3, -2, -1, -2, -5, -5, -5, -4, -4, -1, -1, -1, -1, 0, -1, -1, 0, 0, 1, -2, 0, 1, 0, 0, -1, 0, -2, -3, -1, -2, -3, -5, -4, -4, -3, -2, 0, 0, 0, 0, 0, 0, 2, 3, 2, -2, 0, 0, 1, 0, 1, 0, 0, -1, 0, -3, -3, -3, -4, -3, -1, 0, 0, 0, 1, 0, 0, 0, 3, 4, 5, -2, 0, 0, 0, 0, 0, 0, 1, 0, -1, -2, -2, -3, -1, -2, -1, 0, 1, 1, 0, 1, 1, 3, 3, 5, 8, -3, 0, 1, 0, 0, 0, 1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 3, 3, 5, 7, 9, -3, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 1, 0, 1, 0, 1, 0, 2, 3, 4, 5, 5, 7, 9, 1, 0, 0, 0, 0, 0, -1, -2, 0, -2, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -2, -1, -1, -1, 0, -1, 0, -1, 0, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -3, -2, -2, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, -2, -1, -2, -3, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, -2, -1, -3, -2, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -3, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -3, -3, -3, 0, -1, 0, 0, 0, 2, 0, 0, -1, 0, 2, 1, 0, 0, 0, 0, -1, 0, 0, -2, -1, -2, -2, -4, -3, -4, -1, -2, 0, 1, 1, 2, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -3, -3, -4, -4, -2, -2, -3, -1, 0, 2, 1, 1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 1, -1, 0, -1, -2, -4, -3, -5, -4, -4, -3, -2, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -3, -2, -4, -4, -4, -4, -2, -1, -1, 0, 1, 1, 0, 2, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -2, -2, -3, -3, -2, -2, -2, -2, 0, 0, 1, 0, 2, 2, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, -2, -2, -2, -3, -2, -2, -2, 0, 0, 1, 2, 0, 1, 0, 1, -1, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, -1, -1, -3, -2, -3, -2, 0, 0, 0, 2, 1, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 1, 2, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 2, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 2, 1, 3, 3, 4, 3, 3, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, -1, 0, 1, 1, 0, 2, 2, 3, 3, 3, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 1, -1, -1, 0, 0, 0, 0, 1, 1, 2, 3, 1, 3, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 2, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 1, 1, 0, 0, 0, 0, 2, 3, 2, 2, 0, 1, 1, 2, 2, 1, 0, 0, 0, -1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 2, 2, 1, 0, 1, 1, 1, 2, 1, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, -1, -2, -3, -4, -3, -3, -2, -1, -1, 0, 1, 0, 1, 1, 1, 3, 3, 5, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -4, -3, -3, -2, -1, -1, 0, 0, 1, 0, 0, 1, 1, 1, 4, 2, -1, 0, 0, 1, 0, -1, 0, 0, -2, -1, -2, -4, -4, -3, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 2, -1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -3, -4, -4, -4, -3, -2, -3, 0, -2, -2, 0, 0, 1, 0, 1, 0, -2, -1, -1, 0, 0, -1, 0, 0, -2, -2, -3, -4, -2, -3, -3, -2, -1, -2, -3, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, -2, -2, -3, -2, -3, -2, -3, -2, -2, -2, -2, -1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -2, 0, 0, -2, -1, -2, -2, -2, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 2, 1, 0, 0, -1, 0, -3, -3, -2, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 2, 4, 3, 0, 0, 0, 0, -3, -2, -1, -1, -1, -1, -1, -2, 0, -1, -2, 0, 0, 1, 1, 2, 1, 2, 2, 4, 4, 3, 4, 3, 1, 0, -1, -1, -3, -3, -1, -1, -2, -1, 0, -1, 0, -1, 0, 0, 2, 2, 1, 2, 3, 3, 5, 3, 2, 3, 2, 0, -1, -1, -1, -2, -1, -1, -2, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 4, 4, 4, 3, 3, 1, 0, 0, -3, -2, -2, -3, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 2, 3, 4, 4, 2, 4, 2, 2, 1, 0, -2, -3, -2, -2, 0, -1, -2, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 2, 4, 3, 3, 4, 3, 2, 2, 0, -2, -2, -1, -1, 0, -1, -3, -1, -1, -2, -2, -2, 0, 1, 1, 0, 2, 3, 2, 2, 3, 2, 3, 2, 0, 0, -2, -2, -3, -1, -1, 0, -2, -1, 0, -2, -2, 0, -1, 1, 0, 0, 2, 1, 3, 2, 4, 3, 3, 1, 0, 0, -2, -4, -2, -1, -1, -1, -1, -2, 0, 0, -2, -1, -2, -1, 0, 0, 0, 2, 2, 0, 0, 0, 1, 0, 0, -2, -2, -2, -3, -1, 0, 0, -2, -1, -1, -2, -2, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, -1, -1, -2, -1, -2, -1, -1, -2, -2, 0, 0, -3, -2, 0, -2, 0, -2, -1, -2, 0, 0, 0, 0, -1, -1, -2, -1, -2, -3, -2, -2, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -2, -1, -2, -3, -2, -3, -1, -1, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -3, -3, -4, -2, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, -4, -3, -1, -1, -1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, -2, -2, -2, 0, -1, 0, 0, 0, 1, 1, 2, 3, 4, 3, 1, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, -3, -3, 0, 0, 1, 0, 1, 2, 0, 3, 1, 4, 4, 5, 0, 0, 1, 1, 2, 0, 0, 0, 1, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 3, 4, 4, 0, 0, 2, 0, 2, 2, 2, 1, 2, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 3, 3, 4, 6, 5, 4, 0, 1, 2, 0, 3, 0, 0, 1, -1, -2, -1, -1, -3, -3, -1, 0, 0, 0, 0, 1, 1, 1, 3, 3, 3, 4, 1, 1, 0, 0, 1, 1, 0, -1, -1, -1, -1, -4, -4, -2, -2, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 4, -1, 1, 0, 0, 0, 0, 0, -1, 0, -2, -2, -4, -4, -3, -2, -2, -2, 0, -1, 0, 0, 0, 1, 2, 2, 3, -1, -1, -1, 0, -1, 0, 0, 0, 0, -3, -1, -4, -4, -3, 0, -2, 0, 0, -1, -1, 0, 0, 0, 0, 2, 2, -2, -1, 0, 0, 0, 0, 0, 0, 0, -2, -3, -2, -3, -1, -2, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -2, -3, -3, -1, 0, 0, -1, -1, 0, -2, 0, 0, 0, 0, 1, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, -2, -2, 0, -1, -1, 0, 0, 0, -1, -1, 0, -2, -1, 0, 0, 0, 0, -2, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 1, 1, 0, 0, 0, 0, -2, -1, -1, -1, -1, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 2, 1, 3, 3, 0, 0, 0, 0, -1, -3, -2, -2, 0, -1, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 2, 3, 3, 3, 2, -1, -2, -3, -2, -1, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 3, 4, 2, 1, 0, -1, -1, -2, -2, -2, -2, -2, -1, -2, 0, 0, 0, 0, 0, 1, 3, 1, 2, 2, 3, 4, 4, 3, 3, 2, 0, -1, -2, -1, -3, -1, -2, -1, -1, -2, 0, 0, 0, 0, 1, 1, 1, 0, 2, 2, 3, 4, 2, 3, 1, 1, 0, -1, -1, -2, -3, -3, -1, -1, -2, -2, 0, 0, 0, 0, 0, 0, 2, 0, 2, 1, 4, 4, 3, 4, 1, 2, 1, 1, -1, -1, -2, -2, -2, -2, -1, -2, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 3, 3, 2, 1, 1, 3, 0, 0, -2, -2, -3, -2, -2, -3, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 1, 4, 2, 4, 1, 0, 1, 0, -1, -2, -3, -1, -1, -2, -1, -3, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 3, 1, 3, 2, 2, 0, 0, -2, -1, -3, -2, -1, -1, -1, -3, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 2, 0, 0, 1, 0, -1, 0, -1, -1, -2, -3, -2, -1, -2, 0, -2, -2, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -2, 0, -1, 0, -1, -2, -1, -2, -2, -1, -4, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, -1, -2, -2, 0, -1, 0, 0, 0, 0, -1, -1, 0, -3, -1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -2, -2, -2, -3, -1, -1, -1, 0, -1, -1, 0, -1, -1, -1, -1, -1, -2, 0, 0, 0, 1, 0, 0, -1, -1, -2, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, -1, -1, -1, -3, -3, -3, -2, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 2, 0, 0, 0, -1, -1, -2, -2, -2, -2, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 2, 2, 1, -1, 0, 0, 0, 2, 1, 0, 0, -1, -2, 0, 0, -1, -2, -1, 0, -1, -1, 0, 0, 1, 1, 1, 3, 3, 2, 0, 0, 0, 2, 3, 0, 0, 0, -1, -1, -1, -2, -1, -1, 0, -1, 0, -1, 0, 0, 0, 1, 3, 3, 3, 4, -2, -2, 0, 0, 0, 0, -2, -1, -2, -1, -2, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, -2, -2, 0, 0, -1, 0, 0, 0, -2, -2, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 1, 1, 2, -3, -2, -1, 0, -1, 0, -1, 0, -3, -2, -3, -1, -2, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, -3, -1, -1, -1, 0, 0, -1, -1, -2, -3, -2, -1, -1, -1, -2, -1, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, -3, -1, 0, -1, 0, -1, -1, -1, -3, -3, -1, -3, -3, -2, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, -2, -2, -1, -2, -2, -2, -2, -3, -3, -2, -2, 0, 0, -2, -1, -2, -2, 0, -1, 0, 0, -1, -1, -1, -1, -2, -1, -2, 0, -2, 0, -1, -3, -3, -4, -1, -1, -2, -1, -1, -1, 0, -1, 0, -2, 0, 0, -1, 0, -1, -1, -2, -3, 0, 0, -1, 0, -2, -1, -3, -3, -3, -3, -2, -2, -1, 0, -1, 0, 0, -3, -1, 0, -1, -1, 0, -1, -1, -3, 0, 0, 0, 0, 0, 0, -3, -2, -2, -4, -2, -2, -2, 0, 0, 0, 0, -3, -2, 0, 0, 0, 0, -2, 0, 0, -1, -2, 0, -1, 0, 0, -2, -2, -1, -2, -3, -1, -2, 0, 0, -1, 0, -2, -1, 0, 1, 0, -2, -2, 0, -1, 0, 0, -1, 0, -1, 0, -2, -1, -2, -3, -2, -3, -1, 0, 0, 0, 0, 0, 1, 1, 0, -1, -1, -1, -3, -3, -1, 0, -1, 0, -1, -1, -1, -3, -1, -2, -3, -4, -1, -2, -1, -1, -1, 0, 0, 0, 0, -2, -1, -1, -3, -3, -1, -1, -1, -2, -1, 0, -1, -1, -2, -3, -4, -4, -3, -3, 0, -1, -1, 0, 0, 0, 0, -1, -3, -2, -1, -2, -1, -1, -1, -1, -1, -1, -1, 0, -1, -1, -3, -3, -4, -2, -2, -2, -3, 0, 0, 0, 0, 0, -1, -2, -2, -2, -2, -1, -2, -1, -2, 0, -1, 0, -1, -1, -2, -3, -3, -3, -3, -2, -1, -2, 0, 0, 0, -2, -1, -1, -3, -2, -1, -1, -1, 0, 0, -1, 0, 0, 0, -2, -3, -4, -3, -1, -2, -1, -2, -2, 0, 0, 0, -1, 0, -1, -3, -2, -3, -2, -2, -2, -1, -1, -1, -1, -1, 0, -1, -2, -2, -2, -1, 0, -1, -2, 0, 0, 0, -1, -2, -3, -3, -3, -1, -3, -3, -1, -1, -2, -2, -2, -2, -1, -2, -1, -2, -1, -2, -1, -1, -2, 0, 0, 0, 0, -2, -3, -3, -1, -1, -1, -3, -3, -3, -3, -1, -2, -2, -1, 0, -2, -1, -1, -1, 0, 0, -2, 0, 0, 0, -2, -2, -2, -2, -3, -2, -3, -3, -2, -3, -3, -1, -1, -1, -1, 0, 0, -1, 0, -1, -1, -1, -3, 0, 1, 0, 0, 0, -1, 0, -2, -2, -2, -2, -3, -4, -2, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, -1, -2, -2, -1, -3, -3, -4, -4, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, -3, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -3, -2, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 2, -3, 0, 0, 0, 0, -1, -1, -1, -2, -1, -2, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 2, 2, 3, -4, -1, -1, -1, 0, -2, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 5, 4, -5, -3, -1, 0, -2, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 4, 5, 5, 2, 1, 2, 3, 3, 1, 2, 1, 1, 0, 0, -1, -1, 0, 0, 1, 1, 0, 2, 4, 2, 2, 3, 5, 5, 4, 0, 1, 0, 0, 2, 2, 2, 0, 0, 0, -1, -1, -2, -2, 0, 1, 0, 1, 2, 2, 2, 1, 2, 3, 3, 2, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -3, -3, -1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 2, 0, 0, 0, 1, 0, 0, 0, -1, -2, -3, -4, -3, -3, -3, -1, -1, 0, 0, -1, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, -1, -1, -2, -4, -4, -4, -5, -4, -2, -1, -1, -1, -1, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, -3, -2, -4, -4, -3, -2, -3, -4, -1, -1, -1, -1, 0, 0, 0, 2, 2, 0, 0, 0, 0, -1, 0, -1, 0, -2, -2, -1, -1, -1, -1, -1, -2, -1, -1, -3, -1, -1, -1, 0, 1, 1, 1, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -2, -2, -2, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 1, 2, 2, 0, 1, -1, 0, -2, -1, -1, 0, 0, 0, 0, 0, -2, -1, -2, 0, 0, 0, 0, 0, 1, 1, 2, 4, 2, 2, 2, 2, 1, -1, -1, -2, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 2, 2, 3, 3, 3, 3, 1, 0, 0, -1, -1, -1, -2, -2, -1, 0, -2, -2, -2, -1, 0, 0, 0, 1, 0, 1, 1, 2, 3, 3, 4, 3, 1, 0, 0, 0, -2, -3, -2, -1, -1, -2, -1, -1, -2, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 2, 3, 1, 2, 2, 0, 0, -2, -3, -2, -3, -2, -1, -1, -2, -1, 0, -2, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 3, 2, 0, -2, -2, -2, -1, -1, 0, 0, -2, -1, -1, -2, -1, 0, 0, 1, 1, 1, 0, 0, 1, 1, 2, 1, 3, 1, 1, -1, -2, -2, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 2, 2, 1, 2, 2, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 0, 1, 1, 0, 0, -2, -2, -2, -2, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, -2, 0, 0, -1, -1, 0, -2, -2, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -2, 0, 0, 0, 0, 0, -1, -1, -2, -4, -3, -1, -2, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, -1, 0, -2, -1, -1, -4, -3, -4, -4, -2, -2, 0, 0, 0, -2, -1, -1, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -3, -3, -5, -5, -4, -3, -2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -4, -4, -5, -3, -2, -3, 0, 0, 0, -1, -1, 0, 1, 0, 2, 1, 1, 0, 1, 0, 1, 0, -1, 0, -3, -4, -3, -3, -3, -4, -1, -2, -1, 0, 0, -1, 0, 1, 2, 2, 5, 0, 1, 2, 0, 1, 1, 0, -1, -2, -1, -3, -1, -3, -3, -1, -1, 0, 0, 0, 0, 0, 0, 2, 3, 5, 5, 1, 1, 2, 2, 0, 1, 0, 0, -1, 0, 0, -1, -2, -2, -2, 0, 0, 0, 0, 0, 1, 2, 3, 5, 6, 5, 0, 0, 1, 1, 2, 3, 3, 2, 2, 1, 1, 0, 0, 1, 1, 1, 0, 0, 1, 1, 1, 3, 5, 5, 5, 6, -2, -2, -1, -2, -1, -1, 0, 0, -1, 0, -1, -1, -2, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, -2, 0, -2, 0, -1, 0, 0, -1, -2, -1, 0, 0, 0, -2, 0, 0, 0, 0, -1, -2, -2, 0, -1, -1, 0, 0, -1, -1, -1, -1, -2, -1, -2, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -2, -2, -2, 0, 0, -1, 0, 0, 0, 0, -2, 0, 0, -2, -1, -1, -1, -1, -2, 0, -1, 0, -2, 0, -1, -1, -1, -3, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -2, -1, -2, 0, 0, 0, 0, 0, 0, -2, 0, -2, -1, 0, 0, -1, -2, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -2, 0, -2, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, -2, -2, -1, -1, 0, -1, -1, -1, -1, -1, -2, 0, -1, 0, 0, 0, -1, -1, 0, -3, -2, -1, -1, -1, -2, -1, 0, -2, -1, -1, -1, 0, 0, 0, -2, -1, -2, -2, 0, 0, 0, -1, -1, 0, -2, -3, -1, -2, 0, -2, -2, -2, -2, -1, -1, -1, 0, 0, 0, 0, -1, -1, -2, -1, -2, 0, -1, -2, 0, -1, -1, -2, -3, -1, 0, -1, -2, -2, -2, -1, -2, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -2, 0, -2, -2, -1, 0, 0, -1, 0, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -1, 0, -2, -1, -2, 0, -1, -2, 0, -1, -1, -2, -1, -2, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -3, -1, -1, -2, -2, -2, 0, -2, -1, 0, -1, -2, -1, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -2, -1, -2, -1, -1, -1, -2, -2, -2, -1, -1, -2, -1, -3, -1, -2, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, -2, -1, -1, -1, -2, -1, 0, 0, -1, -1, -2, -2, -1, -2, -1, -2, -1, 0, -1, -1, 0, 0, -1, -1, 0, -1, -2, -2, -2, -3, -2, -1, -1, -1, -2, 0, -2, -1, -2, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, -2, -2, -2, -1, -1, -1, -1, -2, -1, -2, -1, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, -2, -3, -3, -3, 0, 0, -1, 0, 0, -3, -2, -1, -1, -2, 0, -1, 0, -1, -2, -2, -2, 0, -1, -1, -1, -1, -1, -2, -1, -3, -1, -1, -1, -2, -2, -2, -1, -1, -1, -2, -1, -2, 0, 0, -1, -1, -1, 0, -2, 0, -1, -2, 0, -1, -1, -2, 0, 0, 0, -1, -2, 0, -1, -1, -1, -2, -1, -2, -2, -1, -1, -2, 0, -1, 0, -1, -1, -2, -1, -1, -1, -2, 0, -1, 0, -1, -1, -2, -2, -2, -1, -3, -2, -2, -3, -2, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, -1, -2, 0, 0, -1, -1, -1, -1, 0, -2, -1, 0, -2, -2, -1, -2, -1, 0, -1, -2, -1, 0, 0, 0, -1, -2, -2, -1, -1, -1, -1, 0, -1, -2, -1, 0, -2, -2, -1, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 1, -2, -2, -1, 0, -1, -1, 0, 0, -1, 0, 0, -2, -1, -1, 0, -2, -1, -1, -2, -1, 0, 0, 0, 0, 1, 1, -3, -2, -2, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, -2, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 3, 1, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 1, 2, 2, 4, 3, 5, -1, 0, 1, 1, 1, 2, 0, 0, 0, 0, -2, 0, -2, -1, -1, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 3, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -3, -2, -2, -2, -1, 0, 0, 0, -1, -1, 1, 0, 0, 1, 1, 0, -1, -1, 0, 0, 0, 0, -2, 0, 0, -3, -2, -3, -2, -2, -2, -2, -1, -1, 0, 0, 0, 1, 0, 1, 0, 1, -2, 0, -1, 0, 1, 0, 0, -2, -2, -3, -1, -2, -2, -2, -1, -3, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 1, 1, 0, -1, 0, -3, -2, 0, -2, -1, -1, -3, -1, -3, -1, -3, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, -2, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, -2, -1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 3, 3, 2, 1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, -2, -1, 0, 0, 1, 0, 0, 2, 1, 0, 2, 2, 3, 3, 2, 1, 1, 0, 0, -1, 0, -3, -2, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 3, 3, 2, 2, 1, 2, 0, 0, -1, -1, -2, -2, -2, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 3, 2, 0, 0, -1, -1, -2, -2, -3, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 2, 2, 1, 0, 0, 3, 1, 2, 0, -1, -3, -2, -2, -1, -1, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 1, 2, 2, 3, 3, 3, 1, -3, -2, -4, -2, 0, 0, -1, -1, 0, 0, 0, -1, 1, 1, 1, 0, 1, 2, 2, 1, 2, 2, 3, 1, 1, 0, -3, -3, -3, -2, -2, -1, -2, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 2, 2, 1, 2, 1, 2, 0, 1, 0, -3, -2, -3, -2, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 2, 1, 1, 1, 0, 0, 0, -1, -2, -1, -1, -1, -1, 0, -2, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, -1, -1, -1, 0, 0, 1, -1, 0, 0, 0, 0, -2, -1, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, -1, -1, -1, -1, -2, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, -1, -2, -2, -1, -2, -1, -2, 0, -2, -1, -1, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, -2, -1, -1, -1, -2, -3, -1, -2, -2, -2, -2, -1, -1, -1, -1, 0, 1, 1, 1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, -3, -3, -2, -2, -2, -1, -1, 0, -1, -1, 0, 0, 1, 2, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -2, -2, -2, 0, 0, -1, -1, 0, -1, 0, 1, 0, 1, 2, 3, 0, 0, 2, 2, 0, 1, 0, 1, 0, 0, 1, 0, -1, -2, 0, -1, 0, -1, 0, 0, 2, 2, 1, 3, 2, 4, 0, 0, 2, 1, 1, 0, 2, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 2, 3, 0, 1, 2, 2, 0, 2, 3, 2, 1, 2, 2, 2, 3, 1, 1, 0, 2, 0, 0, 1, 3, 4, 4, 4, 5, 4, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, -1, 0, -1, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 1, 1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 1, 0, -1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, -1, 1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 2, 2, 2, 2, 1, 3, 2, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 2, 2, 1, 1, 2, 2, 0, 1, 3, 2, 1, 1, 2, 2, 2, 2, 2, 2, 0, 1, 0, 1, 0, 0, 0, 1, 2, 1, 0, 2, 2, 1, 0, 1, 2, 2, 2, 0, 2, 0, 2, 0, 1, 0, 0, 0, 1, 0, 1, 1, 2, 1, 1, 0, 1, 0, 2, 1, 0, 0, 3, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, -1, -1, -2, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 2, 0, 1, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, -2, -2, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -2, 0, -2, -2, -1, 0, -1, -1, 0, 0, 1, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -2, -2, -2, -1, 0, -2, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, -1, -1, -1, -1, -3, -2, -3, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, -3, -2, -3, -2, -1, -1, 0, 0, 2, 1, 0, 0, 0, -1, 0, 1, 1, 2, 2, 1, 2, 0, 0, 0, -1, 0, -1, -3, -2, -3, -2, -1, 0, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 1, 2, 1, 2, 1, -1, 0, -2, -2, -1, -2, -3, -2, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 2, 2, 1, 0, 0, 0, -2, -1, -2, -1, -2, -1, -2, -3, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, -2, -1, 0, -1, -2, -1, -2, 0, 0, 2, 2, 1, 0, 1, 1, 1, 0, 1, 0, 1, 1, 0, -1, -1, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 1, 2, 1, 2, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 2, 1, 2, 3, 1, 1, 2, 1, 0, 0, 0, 0, 1, 2, 1, 1, 1, -1, -1, -1, -2, 0, -1, 0, 0, 0, 2, 2, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -2, -1, -2, -1, 0, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -2, -1, -2, -1, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -1, -1, -1, 1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, -1, -1, 0, -2, 0, 0, 0, 0, 1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -2, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, -1, -2, -1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 1, 1, 1, 2, 0, 1, 1, 1, 1, -1, 0, 0, 0, -1, -1, 0, 0, 1, 1, 1, 2, 1, 0, 1, 0, 2, 2, 1, 2, 2, -1, 1, 0, 1, 0, 0, -1, -1, -1, 1, 1, 3, 1, 2, 1, 1, 0, 0, 0, 0, -1, -2, -2, 0, -1, -2, 1, 2, 3, 0, 1, 0, 0, 0, 0, 3, 3, 2, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, -2, -2, -3, 3, 3, 1, 1, 2, 1, 2, 1, 3, 3, 2, 1, 0, -2, -1, -1, 0, 0, 1, 0, 0, 0, -3, -3, -2, 0, 2, 1, 0, 1, 1, 2, 2, 2, 1, 2, 1, 0, 0, -2, -1, -1, 0, 1, 1, 2, -1, -2, -4, -3, -2, -1, 1, 2, 0, 1, 0, 1, 1, 2, 1, 0, 0, 0, -1, -1, -2, -1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 2, 0, 0, -1, -2, -2, -2, -3, 0, 0, 0, -1, -2, -1, 0, -1, 0, 1, 0, -1, -2, 0, -1, 0, 1, 0, 1, 0, -2, -4, -2, -3, -4, -3, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -2, 0, -1, 0, 0, 1, 0, -1, -3, -4, -3, -4, -3, -3, -1, 0, 1, 1, 2, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 1, 0, -3, -3, -5, -7, -7, -6, -4, -2, 0, 1, 3, 1, 2, 0, -1, 0, 0, 0, 0, 0, -2, -1, -2, -2, -1, -1, -3, -4, -5, -5, -6, -5, -4, -3, -2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -2, 0, -2, -3, -4, -6, -6, -6, -5, -4, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, -2, -2, -2, -2, 0, 0, -2, -1, -4, -5, -4, -4, -4, -3, -3, -1, -2, -1, 0, 1, 2, 0, 2, 0, -1, -1, -1, -1, -2, -1, -2, 0, 0, -1, -3, -5, -4, -4, -2, -2, -3, -1, -2, 0, 2, 1, 1, 0, 0, -1, -1, -2, -1, -2, -1, -2, 0, -2, -2, -2, -4, -4, -4, -3, -5, -3, -2, -2, 0, 2, 3, 1, 0, 0, 0, -1, -1, -1, 0, -1, -2, -4, -1, -1, 0, -1, -3, -4, -5, -6, -4, -4, -3, -1, 0, 3, 4, 1, 1, 0, -1, -1, -1, -2, -1, -1, -3, -5, -2, -1, -1, -2, -2, -5, -3, -2, -2, -2, 0, 1, 2, 3, 3, 1, 1, 0, 0, -2, 0, -2, -2, -1, -3, -4, -3, 0, -1, 0, -2, -3, -1, 0, 0, 1, 0, 1, 2, 1, 1, 1, 1, 1, -1, 0, -1, -1, -2, -1, -3, -4, -2, -2, 0, 0, 0, 0, 2, 2, 2, 2, 1, 3, 1, 1, 1, 1, 1, 1, -1, -1, 0, -1, -2, -1, -3, -3, -1, -1, 0, 2, 2, 2, 3, 3, 3, 2, 0, 0, 1, 0, 2, 1, 2, 0, -1, 0, -1, -1, -1, -3, -3, -2, -1, -1, 0, 1, 3, 2, 2, 4, 1, 0, 0, 0, 0, 0, 2, 2, 1, 1, -1, -2, -1, -2, -2, -3, -1, -1, -1, 0, 1, 0, 1, 2, 3, 3, 1, 0, -3, -1, 0, 1, 1, 3, 1, 1, -1, -2, -3, -2, -2, -2, -1, -1, 0, 2, 1, 1, 1, 2, 2, 2, -1, -1, -1, 0, 1, 1, 1, 1, 2, 0, -1, -1, 0, 0, -2, -2, -2, 0, 0, 1, 1, 1, 1, 1, 2, 1, 0, -1, 0, 1, 2, 2, 2, 3, 2, 0, 0, -1, -1, -1, -1, -1, -2, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 3, 3, 3, 4, 3, 0, 0, 0, 0, 0, 0, -2, -2, -2, -1, -2, -1, 0, -1, -1, 0, 1, 1, 0, 0, 2, 3, 2, 1, 2, 2, 0, 1, 0, 1, 0, -1, -2, -2, -3, -2, -2, -2, -1, 0, -1, 0, 0, 0, 1, 4, 3, 3, 1, 0, 0, 2, 0, 2, 2, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 1, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 0, 1, 0, 0, 0, -2, -2, -3, -4, -4, -4, -3, -2, 0, 0, 0, 1, 2, 3, 3, 5, 5, 1, 2, 2, 1, 1, 0, -1, 0, 0, -2, -3, -3, -5, -4, -2, -1, -2, 0, 0, 0, 1, 0, 3, 2, 4, 3, 1, 2, 0, 1, 0, 0, -1, -2, -1, -3, -4, -3, -5, -3, -2, -2, 0, -1, -1, 0, 0, -1, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -2, -4, -3, -2, -2, -2, 0, -1, -1, 0, -2, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, -1, -2, -2, -1, -4, -3, -2, -3, -2, -1, -1, -2, -3, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, -2, -1, -3, -2, -2, -1, 0, -1, -1, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, -2, -2, -1, 0, -1, 0, -1, -2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, -4, -2, -1, 0, -1, -2, -3, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 1, 2, 1, 4, 3, 1, 0, -1, -3, -2, -1, -2, -1, -2, -2, -2, 0, 0, 0, 0, 0, 0, 2, 2, 3, 2, 4, 5, 4, 5, 3, 4, 2, -1, -1, -3, -2, -3, -2, -1, -3, -2, 0, 0, 0, 0, 1, 0, 2, 3, 2, 3, 3, 5, 5, 6, 5, 3, 3, 0, -1, -2, -2, -1, -2, -1, -3, -2, -1, 0, 0, 1, 0, 3, 3, 4, 4, 4, 4, 6, 7, 5, 5, 5, 4, 0, -1, -3, -3, -2, -2, -2, -3, -3, -2, 0, 1, 1, 0, 1, 1, 3, 1, 3, 4, 7, 6, 5, 4, 4, 2, 2, 0, -1, -3, -4, -3, -4, -3, -1, -1, 0, 0, -1, 0, 1, 2, 2, 2, 2, 3, 5, 5, 5, 5, 5, 4, 1, -1, -1, -2, -3, -2, -3, -2, -1, -1, -1, 0, 0, -1, 1, 2, 2, 3, 3, 5, 5, 5, 4, 5, 5, 4, 2, 1, -1, -4, -4, -4, -2, -1, -1, -2, -1, 0, 0, 0, 0, 0, 2, 1, 3, 3, 3, 5, 5, 5, 4, 3, 1, 0, -2, -3, -2, -4, -4, -2, -2, -1, 0, -1, 0, 0, 0, 0, 2, 2, 1, 2, 4, 5, 4, 2, 3, 2, 1, 0, -1, -3, -3, -3, -2, -2, -2, -2, -1, -1, 0, -1, 1, 1, 0, 1, 2, 1, 3, 3, 2, 0, 0, 1, -1, 0, -1, -3, -3, -3, -4, -1, 0, -2, -2, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, -2, -2, -1, -2, -3, -3, -3, -2, 0, -2, -1, -2, -1, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, -3, -1, -1, -2, -1, -2, -2, -2, -1, -2, -1, -1, 0, 0, -1, 0, -1, 0, 0, -2, -2, -1, -1, -2, -2, -1, -1, -2, -1, -1, -1, -1, -1, -1, -1, 0, -2, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -2, -2, -3, -4, -3, -1, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, -2, -2, -3, -2, -2, -4, -3, -3, -2, -1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 1, 2, 1, 1, 0, -2, -1, -2, -2, -4, -3, -2, 0, 0, -1, 0, 0, 0, 1, 1, 0, 3, 3, 3, 2, 1, 1, 1, 1, 0, 0, 0, -3, -3, -2, -3, -4, -1, -1, -1, -1, 0, 0, 1, 1, 3, 3, 4, 3, 4, 1, 2, 2, 2, 1, 2, 1, -1, -1, -1, -2, -2, -3, -1, 0, 0, -1, 0, -1, 1, 2, 3, 2, 3, 4, 4, 0, 0, 0, 0, -1, -1, -2, -1, -2, -2, -2, -2, -2, -2, -1, -1, 0, -1, -2, -1, -2, -1, -1, 0, 0, -2, 2, 2, 0, 0, 0, 0, 0, -1, -1, -3, -1, -1, -2, -1, -1, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, -2, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 1, 1, 1, 0, 0, -2, 0, -1, -1, -1, -1, -2, 0, -2, 0, -1, 0, 0, -1, 0, 0, -2, -1, 0, -1, 0, 2, 0, 1, -1, -1, 0, -1, -1, -1, -1, 0, -1, 0, 0, -1, -2, 0, 0, -2, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, -1, -1, 0, -1, -1, 0, -1, -1, 0, 0, -2, -1, -1, -2, -1, -2, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -2, -2, -1, -1, -1, -1, -2, -1, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -1, -2, -2, -1, -1, -1, -2, -1, -2, -1, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 2, 2, 0, 0, 0, -1, -1, -2, -1, -1, -2, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 2, 1, 0, -1, -1, 0, -2, -3, -2, -2, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 2, 3, 2, 2, 2, 0, 0, -2, -1, -3, -3, -1, -2, -2, -1, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 1, 2, 2, 2, 3, 1, -1, -2, -2, -3, -3, -2, -3, -3, -1, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 1, 2, 0, 0, -2, -3, -2, -3, -3, -2, -3, -2, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 1, 2, 3, 1, 2, 0, -2, -2, -3, -2, -2, -1, -2, -2, -1, 0, 0, 1, 0, 0, -1, 2, 1, 0, 1, 1, 0, 2, 3, 1, 0, 0, -2, -3, -3, -2, -2, -2, -2, -2, 0, 0, 1, 1, 0, 0, 0, 1, 2, 2, 2, 2, 2, 2, 1, 2, 0, 0, -2, -3, -2, -3, -3, -3, -2, -1, 0, 0, 1, 0, 0, 0, -1, 2, 2, 1, 3, 1, 2, 2, 0, 0, 0, 0, -2, -1, -2, -3, -2, -2, -1, -1, 0, 0, 0, 1, 0, 0, -1, 1, 1, 2, 3, 1, 0, 0, 2, 1, 0, 0, -1, -1, -2, -1, -3, -3, -1, -1, 0, 0, 1, 0, 1, 0, -1, 3, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, 3, 2, 2, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, -2, -2, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 1, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 1, -1, 0, -1, 0, 1, 0, 0, 0, 2, 0, 1, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -2, 1, 2, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 0, 0, 1, 0, 0, 0, 0, -1, -1, 1, 1, 2, 3, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 1, 1, 1, 1, 0, 0, 1, 0, 1, 1, 7, 4, 4, 3, 3, 3, 3, 0, -1, -2, -5, -7, -8, -8, -5, -2, -2, 0, 0, 1, 2, 2, 2, 3, 4, 2, 6, 4, 2, 1, 1, 1, 0, 0, -1, -2, -4, -8, -6, -6, -5, -2, -1, 0, 1, 0, 0, 0, 1, 2, 2, 2, 3, 3, 2, 1, 0, 0, 0, -2, -4, -3, -7, -7, -6, -5, -3, -2, 0, -1, 0, 0, 0, 0, 1, 2, 1, 1, 2, 1, 0, 0, -1, -1, -1, -4, -5, -6, -7, -6, -6, -6, -3, -2, -1, 0, -2, -1, 0, 0, 0, 2, 0, 0, 3, 0, 1, 0, -1, 0, -2, -3, -5, -6, -5, -6, -4, -4, -3, -2, -3, -1, -2, -1, 0, 0, 1, 1, 0, -2, 2, 0, -1, 0, 0, 0, -1, -3, -4, -3, -4, -3, -2, -3, -1, -3, -2, -3, -2, 0, 0, 0, 1, 0, 0, -3, 3, 1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, -1, -3, -3, -2, -1, 0, 0, 0, 0, -2, -4, 1, 1, 0, 0, 0, 1, 2, 2, 3, 4, 5, 4, 2, 3, 1, 0, -1, -1, -2, -3, -3, -1, -1, 0, -3, -5, 2, 0, 0, -1, 0, 1, 2, 4, 6, 7, 6, 6, 6, 5, 4, 2, 1, -1, -2, -3, -3, -2, -2, -1, -4, -7, 1, 0, -1, 0, 1, 2, 7, 7, 9, 8, 9, 9, 8, 9, 8, 7, 3, 0, -2, -2, -5, -3, -4, -4, -5, -6, 0, -2, 0, 0, 1, 4, 6, 7, 9, 8, 10, 11, 10, 9, 11, 8, 6, 2, 0, -1, -2, -4, -3, -5, -5, -6, -3, -2, 0, 0, 2, 4, 5, 7, 8, 9, 10, 10, 9, 10, 10, 7, 5, 4, 2, 0, -2, -3, -4, -3, -3, -5, -3, -2, 0, 0, 2, 5, 5, 7, 8, 9, 8, 9, 9, 8, 9, 7, 6, 4, 2, -1, -1, -3, -3, -3, -3, -3, -4, -1, 0, 1, 1, 5, 7, 8, 7, 8, 7, 7, 8, 9, 9, 9, 8, 6, 1, 0, -2, -2, -2, 0, -1, -1, -3, -1, 0, 0, 2, 4, 6, 6, 6, 6, 7, 6, 8, 8, 10, 9, 5, 5, 2, 0, -1, -2, -2, -1, 0, 0, -3, -1, 0, 1, 4, 5, 7, 8, 7, 8, 7, 7, 8, 8, 7, 5, 5, 2, 0, 0, -2, -1, -1, 0, 0, 1, -2, 0, 0, 1, 3, 5, 5, 6, 7, 5, 6, 6, 5, 4, 3, 1, 0, 0, -2, -2, -1, -2, -1, 0, -1, 1, -2, -1, 0, 0, 1, 1, 4, 5, 3, 3, 2, 2, 2, 0, -1, -2, -3, -2, -3, -1, 0, 0, -1, -1, -1, -1, -1, -1, -1, -2, 0, 0, 0, 2, 1, 1, 0, -1, 0, -2, -4, -3, -5, -4, -2, 0, 0, 0, 0, -2, -2, -1, 0, -1, -2, -1, -1, 0, 0, 0, -1, 0, -2, -3, -2, -4, -3, -4, -3, -3, -1, 0, 0, 0, 0, -1, -2, -2, 0, 0, -1, -1, 0, 0, -1, -2, -3, -4, -3, -3, -4, -5, -6, -5, -3, -2, -1, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, -1, 0, 0, -2, -3, -4, -5, -5, -7, -6, -4, -4, -2, -2, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, 0, -1, -1, -1, -4, -5, -5, -5, -4, -6, -7, -5, -2, -2, 0, 0, 0, 1, 1, 3, 1, 3, 1, 3, 3, 0, 0, 0, 0, -2, -1, -3, -3, -2, -5, -4, -4, -5, -4, -2, -1, 0, 1, 2, 1, 1, 4, 3, 2, 5, 4, 2, 0, 0, 0, 0, 0, -2, -3, -3, -3, -4, -4, -2, -1, 0, 0, 0, 2, 2, 2, 3, 4, 4, 4, 5, 4, 3, 1, 3, 2, 2, 0, 1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 2, 2, 2, 4, 5, 4, 4, 4, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, -1, 4, 5, 2, 1, 0, 0, 0, 0, -1, -3, -5, -6, -6, -4, -4, -1, -2, 0, -2, -1, 0, 0, 1, 1, 1, 2, 5, 2, 2, 2, 0, 0, 0, -1, -2, -3, -5, -5, -3, -1, -2, -1, -1, 0, -1, -2, -1, 1, 1, 3, 3, 2, 3, 2, 3, 2, 0, 0, 0, 0, -2, -3, -2, -3, -2, 0, -1, 0, -1, -1, -2, -2, -1, 0, 1, 3, 1, 1, 3, 4, 2, 2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 1, 2, 1, 0, 1, 4, 4, 3, 0, 0, 1, 3, 2, 1, 0, 0, 1, 3, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 3, 4, 4, 1, 0, 0, 0, 2, 3, 1, 1, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 1, 1, 1, -1, 0, 2, 2, 3, 0, 0, 0, 2, 1, 2, 3, 2, 2, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 2, 3, 1, 0, 1, 2, 3, 1, 2, 2, 3, 2, 1, 2, 2, 2, 1, 0, 0, 0, 0, 0, -3, -1, 0, -2, 2, 1, 0, 0, 0, 1, 3, 2, 0, 1, 3, 2, 2, 2, 4, 4, 1, 0, 0, -2, -1, -1, -2, -2, -2, -1, 3, 1, 1, 2, 1, 2, 1, 1, 1, 1, 2, 1, 3, 4, 4, 2, 2, 1, -1, 0, -2, -2, -1, -1, 0, -2, 3, 3, 3, 1, 1, 1, 3, 2, 0, 3, 1, 3, 1, 4, 4, 3, 2, 0, 0, -2, -2, 0, -1, 0, 0, 0, 5, 3, 2, 1, 3, 3, 2, 0, 2, 4, 4, 2, 4, 3, 5, 2, 2, 0, -2, -1, 0, 0, 0, 1, 0, 0, 6, 4, 1, 2, 2, 2, 2, 0, 3, 3, 3, 3, 4, 4, 5, 3, 1, -1, -3, -1, 0, 2, 2, 0, 1, 2, 5, 3, 2, 1, 3, 3, 0, 1, 1, 3, 5, 4, 6, 7, 7, 5, 1, -3, -3, -1, 0, 1, 1, 2, 2, 2, 5, 3, 0, 0, 0, 2, 2, 1, 1, 2, 3, 4, 6, 7, 6, 2, 0, -2, -2, 0, 0, 1, 1, 2, 2, 1, 5, 3, 1, 0, 1, 2, 2, 0, 0, 2, 3, 3, 4, 4, 3, 1, 1, 0, -1, 0, 0, 2, 1, 0, 2, 1, 4, 2, 1, 0, 0, 1, 2, 0, 0, 1, 1, 3, 2, 4, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 4, 2, 1, 0, 0, 1, 2, 2, 1, 1, 2, 3, 2, 3, 2, 2, 1, 0, 0, 0, 2, 0, 0, -2, 0, -1, 4, 2, 1, 0, 0, 3, 4, 2, 0, 0, 1, 1, 1, 1, 1, 3, 3, 1, 1, 0, 1, 0, 0, -1, -1, 0, 3, 2, 0, 1, 2, 2, 3, 0, 0, 0, 1, 0, 0, 0, 0, 2, 4, 3, 1, 0, 0, -1, -2, -2, -1, 0, 4, 1, 2, 2, 3, 1, 0, -1, 0, 0, 0, 1, 2, 0, 2, 2, 3, 2, 1, 0, 0, -2, -2, 0, 1, 2, 3, 1, 2, 2, 2, 1, -1, -1, 0, 0, 0, 0, 0, 0, 2, 3, 3, 1, 0, 0, -1, 0, 0, 0, 0, 0, 3, 3, 5, 5, 2, 0, -2, -2, -1, 0, 0, 0, 0, 0, 1, 1, 3, 1, 0, 0, 0, 1, 1, 0, 0, 0, 2, 4, 4, 4, 2, 1, -1, -1, -1, -1, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 2, 1, 2, 1, 0, 3, 4, 4, 5, 4, 3, 0, -1, -2, -2, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 1, 1, 1, 1, 0, 0, 3, 3, 4, 5, 4, 3, 0, -1, -2, -1, -2, -2, -1, -1, 0, -1, -1, -2, -1, 0, 1, 3, 2, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, -1, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, -2, -1, -2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, -2, -2, -1, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, -1, -1, -2, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -2, -2, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, -1, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 7, 6, 4, 2, 1, 0, 0, -2, -1, -2, -4, -4, -4, -4, -4, -4, -3, -2, -1, 0, 0, 2, 4, 4, 5, 6, 6, 6, 4, 3, 2, 0, -1, 0, -3, -3, -5, -6, -5, -3, -4, -3, -3, -2, 0, -2, 0, 0, 1, 4, 3, 5, 4, 4, 3, 2, 1, 0, 0, 0, -1, -2, -4, -3, -2, -3, -3, -3, -2, -2, 0, -1, 0, 0, 0, 1, 3, 4, 3, 2, 3, 0, 0, 0, 0, 0, -1, -2, -3, -2, -1, -2, -1, 0, -2, -2, 0, -1, 0, 0, 0, 1, 2, 2, 3, 2, 2, 0, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, -2, -3, 0, 0, -1, 0, 0, 0, 0, 2, 1, 2, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -2, 0, -2, -2, -1, -2, -1, -1, 0, 1, 1, 2, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -2, -2, 0, -2, 0, -1, 1, 0, 0, -1, 0, 1, 0, 0, 0, 1, 2, 0, 0, 2, 1, 2, 0, -1, -1, -2, -2, -3, -2, -1, -2, -1, 3, 0, 0, 0, 0, 1, 0, 0, 1, 0, 2, 3, 2, 3, 3, 2, 0, -1, -1, -3, -2, -3, -1, 0, -2, -2, 2, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 3, 3, 4, 4, 2, 1, 0, 0, -1, -1, -2, -1, 0, -1, -1, 1, 0, 1, 0, 0, 2, 0, 3, 2, 3, 5, 5, 5, 5, 6, 4, 2, -1, 0, -3, -1, 0, 0, -1, -1, 0, 2, 1, 0, -1, 0, 1, 1, 1, 4, 3, 6, 5, 6, 6, 6, 3, 3, 0, -2, -1, 0, -2, -1, 0, 0, 0, 2, 1, -1, 0, 0, 1, 0, 2, 4, 4, 5, 7, 8, 7, 7, 5, 1, -1, -1, -2, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 2, 4, 6, 6, 7, 7, 6, 5, 2, 0, -3, -2, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, 0, 2, 3, 3, 3, 6, 7, 7, 6, 4, 1, -1, -2, -1, -2, 0, 0, -1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 2, 1, 2, 3, 4, 5, 6, 4, 2, 0, 0, -1, -1, 0, 0, -2, -1, -1, 0, 0, 0, -1, -2, -2, 0, 1, 0, 1, 0, 1, 3, 3, 5, 3, 1, 0, 0, -1, 0, -2, -3, -1, -1, -1, -1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 2, 0, 0, -1, 0, -2, -2, -2, -3, -2, -2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 1, -1, -1, 0, 0, -3, -3, -1, -3, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -3, -2, -2, 0, 1, 0, 2, 0, 0, 0, -1, 0, -1, 0, 0, -1, -2, -2, 0, 0, 0, 0, -1, 0, -1, -2, -2, 0, 0, 1, 2, 2, 1, 2, 1, -1, -1, -2, -2, -2, -2, -1, -2, -1, 0, 1, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, 4, 2, 2, 2, 1, -1, -2, -3, -3, -2, -1, -2, -2, 0, -1, 0, 0, -1, 0, 0, 0, 0, 2, 0, 1, 0, 3, 4, 3, 3, 3, 1, 0, -1, -2, -3, 0, -2, 0, -1, 0, 0, 0, -1, 0, 0, 0, 2, 2, 3, 1, 1, 5, 5, 4, 4, 4, 3, 0, -2, -2, -3, -3, -2, -1, 0, 0, 0, 0, 0, -1, 1, 3, 3, 2, 3, 1, 2, 5, 6, 3, 5, 4, 3, 0, -1, -3, -4, -4, -3, -3, -1, 0, -2, -2, -1, -1, -1, 1, 3, 2, 4, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 1, -1, 0, -1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 7, 5, 5, 5, 5, 5, 4, 2, 0, 0, -1, -2, 0, -2, -1, -1, 1, 3, 4, 3, 3, 6, 4, 7, 6, 7, 4, 3, 3, 1, 1, 1, 2, 1, 1, -1, -3, -3, -3, -4, -2, 0, 0, 2, 1, 1, 2, 2, 3, 4, 6, 6, 3, 1, 2, 1, 0, 0, -1, 0, -2, -2, -4, -4, -5, -3, -2, 0, 1, 0, 0, 0, 1, 1, 2, 2, 4, 3, 1, 0, 1, 0, 0, -1, 0, -2, -2, -4, -5, -7, -5, -4, -2, 0, 0, -1, 0, 0, 0, 0, 0, 2, 2, 1, 2, 1, 1, 0, 0, 0, -4, -4, -5, -6, -6, -5, -5, -4, -2, -2, -1, -2, 0, -1, 0, 0, 2, 0, 1, 0, 3, 0, 0, 0, 0, -2, -2, -4, -4, -3, -3, -5, -4, -3, -2, -1, -3, -3, -1, -2, 0, 0, 2, 0, 0, -2, 3, 1, 0, 1, 0, 0, -3, -3, -1, -1, -1, -1, -2, 0, -1, -1, -1, -3, -2, -2, 0, 1, 2, 0, -1, -2, 2, 1, 1, 0, 0, 0, 0, -1, 1, 2, 3, 2, 0, 0, 0, 0, -1, -4, -3, -3, 0, 0, -1, -1, -1, -4, 3, 1, 0, 0, 0, 1, 1, 2, 2, 4, 5, 4, 4, 2, 3, 1, 0, -3, -3, -2, -3, 0, 0, -1, -2, -3, 0, 0, 0, 0, 0, 1, 3, 4, 7, 7, 7, 7, 7, 6, 5, 2, 0, -1, -2, -3, -3, -2, -2, -1, -1, -3, 1, 0, 0, 0, 2, 1, 3, 5, 5, 8, 7, 8, 8, 8, 7, 4, 1, 0, -2, -3, -3, -3, -4, -3, -3, -4, -1, 0, -1, 0, 0, 2, 4, 4, 4, 4, 8, 7, 8, 6, 7, 5, 4, 1, -1, -2, -4, -3, -4, -2, -4, -4, -1, -1, -2, 0, 0, 2, 2, 2, 3, 4, 5, 5, 5, 6, 5, 7, 6, 4, 0, -1, -3, -4, -2, -2, -2, -3, -2, 0, 0, -1, 0, 1, 4, 3, 3, 4, 4, 5, 4, 6, 6, 7, 6, 5, 2, -2, -3, -2, -1, -2, -2, -2, 0, -2, 0, 0, 1, 2, 4, 3, 2, 4, 4, 3, 4, 5, 5, 7, 6, 3, 1, -2, -2, -2, 0, 0, 0, 0, -2, -1, 0, 1, 0, 1, 3, 4, 2, 5, 4, 4, 3, 4, 6, 6, 5, 3, 1, -2, -3, -2, -1, 0, 1, 1, 0, -2, 0, 0, 0, 1, 1, 3, 3, 3, 4, 3, 3, 3, 2, 2, 2, 2, -1, -2, -1, -2, 0, 0, 0, 3, -1, -2, -1, 0, 0, 0, 1, 1, 3, 3, 2, 1, 1, 1, 0, -1, -1, -1, 0, -3, -1, -1, 0, -1, 2, 1, 0, 0, 0, -1, -3, -1, 0, 0, 0, -1, 0, 0, 0, -2, -3, -2, -2, -2, -1, -1, -1, -2, -1, -1, 0, 0, 0, -1, -1, -2, -2, -2, -2, 0, -2, -3, -3, -3, -3, -3, -4, -4, -3, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -2, -3, -2, -4, -4, -5, -5, -5, -5, -3, -3, -2, 0, 0, 0, 0, 0, 0, 1, 0, 3, 1, 0, -2, 0, 0, -1, -1, -4, -5, -6, -4, -5, -5, -5, -4, -3, 0, 1, 1, 0, 0, 0, 2, 1, 2, 4, 2, 0, 0, 1, 0, 0, -2, -3, -4, -4, -4, -5, -5, -3, -4, -2, 0, 1, 0, 0, 1, 1, 2, 3, 6, 6, 2, 1, 1, 1, 0, 0, -1, -3, -3, -3, -3, -5, -4, -3, -3, 0, 0, 0, 1, 1, 2, 2, 3, 5, 6, 5, 4, 2, 1, 2, 0, 1, 0, 0, 0, 0, -2, -2, -3, -1, -1, 0, 1, 0, 3, 2, 1, 2, 4, 5, 6, 5, 5, 3, 1, 1, 2, 2, 3, 1, 2, 1, 1, 0, 0, 0, 0, 0, 1, 2, 3, 2, 3, 4, 6, 8, 7, 0, 0, 1, 0, -1, -1, -2, -2, -2, -1, -1, -1, 0, 0, -1, -3, -3, -1, -2, -2, -2, 0, -1, -2, 0, -2, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, 0, -1, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, -2, 0, -1, 0, 0, 1, 1, 0, 0, 0, -1, 0, -2, 0, -2, 0, -2, -2, -2, -1, -1, -1, -1, -1, -2, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, 2, 1, 0, 0, -1, 0, 0, -1, 0, -1, -1, -2, 0, 0, -1, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, -1, -2, 0, -1, -1, -2, -1, -1, 0, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -2, -2, -2, -2, -1, -1, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, -1, -2, -1, -2, 0, -1, 0, -1, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -2, -2, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 2, 1, 0, 0, 0, -1, -2, -3, -1, -2, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 1, 0, 0, 0, -2, -1, -2, -1, -3, -3, -2, -1, 0, 0, -1, 0, 0, 0, -1, 1, 1, 1, 1, 1, 1, 0, 1, 2, 0, -1, -1, -1, -3, -2, -2, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 2, 0, 2, 2, 1, -1, -1, -2, -2, -2, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 2, 1, 0, 0, -1, 0, -2, -1, -3, -2, 0, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, -1, 0, -2, -3, -1, -1, -1, -2, 0, 0, 0, 0, 0, -1, 0, -1, 1, 1, 0, 1, 1, 0, 1, 1, 2, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 2, 2, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 2, 1, 1, 0, 1, 1, 1, 0, 2, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, 1, 0, 1, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, -2, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 2, 1, 2, 1, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 1, 2, 1, 2, 2, 0, 1, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 2, 1, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, -1, 1, 1, 0, 2, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, 0, -1, 0, 0, -1, -1, -1, -3, -2, -2, -1, -1, 0, 0, 1, 2, 1, 0, 1, 1, 0, 0, 0, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, -3, -3, -2, 0, -2, 0, 0, 1, 1, 2, 2, 1, 0, 0, 0, 1, -1, 0, -1, -1, 0, 1, 0, 0, 0, -1, -2, -3, -1, -1, -1, -2, 0, 1, 2, 0, 2, 1, 1, 0, 0, 1, 0, -2, -1, -2, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -3, 0, -1, 0, 0, 0, 2, 2, 1, 1, 0, 1, -1, -1, -1, -1, 0, 0, 0, -1, 0, -1, -2, -2, 0, -2, -1, -1, 0, -1, 0, 1, 2, 3, 1, 0, 2, 1, 0, -2, 0, 0, 0, 0, 0, 0, -1, 0, -3, -2, -2, -3, -3, -1, -3, -2, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -3, -2, -2, -2, -2, -1, 0, 2, 3, 3, 3, 0, -1, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, -2, 0, -1, -2, -4, -2, -2, -2, 0, 0, 2, 3, 3, 3, 1, 0, 0, 0, 0, 0, -1, -1, -2, 0, -1, 0, -1, -1, -3, -1, -2, -1, -1, 0, 0, 1, 1, 2, 1, 2, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 3, 1, 2, 1, 1, 0, 0, 0, -1, -1, -2, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 2, 1, 3, 2, 1, 2, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, -1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 0, 2, 0, 0, 0, -1, -1, 0, -2, -1, -1, 0, 0, 0, 1, 0, 0, 0, 2, 1, 0, 1, 1, 1, 2, 2, 1, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 1, 1, 3, 2, 2, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, 2, 2, 2, 3, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 3, 1, 1, 3, 0, 0, 2, 1, 0, 2, 0, 1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 1, 0, 0, 2, 1, 3, 2, 1, 1, 2, 2, 1, 0, 2, 1, 2, 1, 1, 0, 1, 0, 0, 0, -1, -1, -1, 0, -2, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -2, 0, -1, -1, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, -1, -2, -1, -2, 0, -1, 0, -2, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, -2, 0, 0, -1, -2, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, -1, -2, -2, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, -2, -1, -1, -1, -2, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, -2, -1, -2, -1, -1, 0, -2, -1, -1, -1, -1, -2, -2, 0, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -2, -1, 0, 0, 0, -2, 0, 0, -2, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, -2, -1, -2, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -2, 0, -2, -2, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, 0, -2, 0, -2, 0, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -2, -2, -2, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, -1, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, -1, 0, -3, -1, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -2, -3, -2, -2, 0, 0, -2, -1, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, -2, -1, -1, -2, -1, 0, -2, -2, -1, 0, 0, -1, -1, -1, -1, -1, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, -2, -2, -2, 0, -2, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, -1, -2, -1, -1, -2, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, -2, -2, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 1, 0, 1, 0, 1, 2, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, -2, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, 1, 1, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, 0, 1, 2, -1, -1, -1, 0, -1, -1, -1, -2, -1, -1, -1, -3, -1, -1, -1, -1, 0, 0, 2, 2, 1, 2, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, -3, -3, -2, -3, -1, -2, -1, 0, 1, 2, 3, 2, 2, 0, 0, 1, 0, 0, 0, 0, -2, -2, -2, -2, -2, -3, -3, -3, -4, -2, -1, -1, 0, 0, 0, 0, 1, 3, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, -1, -2, -1, -3, -3, -3, -3, -1, -1, -1, 0, 1, 1, 2, 2, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -2, -2, -1, -1, -3, -3, -1, -2, -1, 0, 1, 1, 0, 0, 1, 1, 0, 2, 0, 1, 0, 0, 0, -1, -1, -1, 0, -1, -2, -1, -3, -3, -1, -1, -2, 0, 1, 1, 1, 3, 1, 2, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, -2, -2, 0, -2, -1, -2, 0, -2, -2, 0, 1, 2, 2, 2, 2, 2, 0, 2, 1, 0, -1, 0, 0, -2, -1, -2, -2, 0, -1, -2, -2, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 2, 0, 1, 1, 1, -1, -1, 0, -2, -2, -2, -2, -2, -1, -1, -1, 0, 0, 1, 1, 3, 2, 1, 1, 1, 1, 0, 0, 0, 1, 0, -1, -1, -1, -2, -1, -3, -2, -1, 0, 0, 0, 0, 2, 1, 1, 2, 3, 2, 1, 1, 1, 0, 1, 1, 2, 1, 0, 0, 0, -1, -2, -2, -1, 0, -1, 0, 0, 1, 3, 2, 1, 3, 3, 2, 1, 2, 1, 0, 0, 0, 2, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 1, 1, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, -1, -1, 0, -2, 0, 0, 0, 1, 2, 0, 2, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 1, 1, 2, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 1, 0, 1, 0, 0, 0, 1, 2, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 2, 2, 0, -1, 0, 0, 0, 1, 1, 2, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 1, 1, 0, 3, 1, 1, 2, 1, 2, 1, 0, 1, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 0, 0, 0, 2, 1, 1, 0, 0, 0, -2, 0, -1, -1, -1, 0, -1, 0, 0, 1, 2, 2, 1, 2, 1, 1, 0, 1, 2, 2, 2, 2, 2, 0, 0, -1, -2, -1, -1, 0, -1, -1, -2, -2, 0, 0, 0, 0, 2, 0, 1, 0, 0, 2, 2, 2, 3, 2, 1, 0, -1, 0, 0, -2, -1, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, 1, 1, 0, 1, 2, 2, 3, 1, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 0, 2, 2, 1, 2, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 2, 0, 1, 0, 2, -1, -1, -3, 0, -2, -1, -2, -2, -2, -2, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 2, 1, 0, -1, -1, -1, -2, -2, -2, -2, -2, -2, 0, -1, -2, -2, 0, 0, 0, 0, 1, 2, 0, 1, 0, 1, 0, 0, 1, 0, 0, -1, -2, -1, -2, -3, -3, -2, -2, -1, -2, -3, -1, -1, -1, 0, 0, 0, 3, 3, 2, 1, 0, 0, 0, 0, -1, 0, -2, -1, -3, -3, -4, -3, -3, -4, -2, -3, -2, -2, -1, 0, 0, 2, 2, 3, 0, 0, 1, 1, 0, 0, 0, -2, -2, -3, -2, -2, -4, -3, -5, -4, -3, -4, -2, -1, -2, 0, 0, 2, 2, 3, 1, 2, 0, 0, 0, 0, 0, -1, -2, -1, -3, -3, -3, -4, -3, -3, -4, -3, -2, -3, -1, 0, 0, 0, 2, 2, 3, 1, 0, 0, 0, 2, 0, -2, -1, -1, -3, -3, -3, -3, -3, -5, -3, -3, -2, -1, -1, -1, 1, 1, 1, 2, 2, 2, 0, 1, 0, 0, -1, -1, 0, 0, -2, -4, -4, -3, -2, -3, -4, -3, -3, -2, 0, 0, 0, 1, 3, 3, 3, 1, 1, 0, 0, 1, 0, 0, 0, -2, -3, -4, -2, -3, -4, -3, -2, -2, -3, -3, 0, -1, 0, 2, 1, 3, 3, 2, 0, 0, 0, 0, -1, 0, -2, -1, -3, -2, -2, -2, -3, -3, -2, -1, -2, 0, -1, 0, 1, 0, 2, 3, 1, 2, 1, 1, 0, 0, -1, -1, -3, -4, -3, -2, -3, -2, -3, -1, -2, -2, 0, 0, 2, 0, 2, 1, 1, 0, 1, 1, 1, 0, 1, -1, -2, -1, -3, -3, -3, -3, -3, -3, -1, -2, 0, 0, 1, 2, 1, 2, 1, 1, 1, 0, 2, 1, 1, 0, 0, 0, -1, 0, -3, -1, -3, -2, -1, -1, 0, -1, -1, 1, 0, 1, 3, 3, 2, 1, 1, 1, 0, 0, 1, 0, 2, 0, 0, -1, 0, -1, -2, -1, -2, 0, -1, 0, 0, 1, 1, 2, 1, 2, 3, 2, 1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, -2, 0, -1, 0, -1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 2, 2, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, -1, -1, -1, -2, -2, -2, 0, 0, 0, 0, 0, 1, 1, 3, 3, 3, 5, 4, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -3, -4, -2, -3, -1, 0, 0, 0, 0, 0, 1, 0, 2, 3, 3, 2, -1, 1, 1, 0, 0, -1, -1, -1, -2, -3, -3, -4, -2, -2, -2, 0, -2, -1, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, -1, -1, -1, -3, -2, -4, -4, -3, -3, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 2, 0, -2, 0, 1, 0, 0, 0, -1, -2, -3, -1, -3, -4, -3, -2, -1, -1, -2, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -2, -2, -2, -2, -1, -1, -1, -3, -2, -3, -2, -1, 0, 0, 1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, -1, 0, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, -2, -3, -3, -1, -2, -1, 0, -2, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 2, 2, 2, 3, 1, 0, -2, -2, -3, -1, -1, 0, -1, -2, -1, 0, -1, 0, 1, 0, 0, 0, 1, 1, 1, 2, 3, 4, 4, 3, 3, 0, -1, -1, -2, -1, -1, -2, -2, -3, -3, -1, -1, 0, 0, 1, 0, 2, 0, 1, 2, 3, 3, 4, 4, 4, 3, 3, 0, -2, -3, -3, -3, -3, -2, -2, -2, -1, 0, 0, 0, 0, 1, 0, 0, 2, 1, 3, 2, 4, 3, 3, 3, 2, 0, 0, -1, -2, -2, -3, -1, -1, -2, -1, 0, 1, 0, 0, 0, 1, 1, 1, 2, 2, 4, 4, 3, 5, 3, 4, 3, 0, -2, -2, -2, -3, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 2, 2, 2, 3, 4, 4, 5, 4, 1, 0, -2, -2, -4, -4, -1, -1, -2, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 2, 2, 4, 3, 3, 3, 2, 0, -2, -4, -4, -3, -2, -2, -1, -1, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 2, 4, 2, 3, 4, 1, 1, 0, 0, -2, -1, -2, -1, -1, 0, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 2, 0, -1, -2, -2, -4, -3, -2, -2, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, -2, -2, -3, -4, -2, -3, -2, 0, -2, -1, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, -2, -1, -1, -2, -3, -1, -2, -1, -2, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, -2, -1, -1, -1, -3, -2, -2, 0, 0, -1, 0, -1, 0, -1, -1, -2, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, -3, -2, -2, -3, -2, -1, -1, -1, -1, -1, -1, -1, -1, -1, 0, 1, -1, 0, 1, 0, 0, 0, -1, -1, -2, -1, -1, -3, -4, -3, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 2, 2, 0, 2, 1, 1, 2, 1, 0, 0, -2, -1, -1, -1, -2, -3, -2, -2, 0, 0, 0, 0, 0, 0, 1, 3, 3, 3, 0, 1, 0, 2, 1, 1, 0, -1, -2, -1, -1, -2, -3, -2, -1, 0, 0, 0, 1, 1, 2, 1, 2, 3, 3, 4, 0, 2, 2, 2, 1, 2, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 3, 3, 4, 4, 5, 0, 2, 3, 1, 2, 2, 1, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 2, 3, 3, 5, 5, 5, 6, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, -1, 1, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, -1, 0, 1, 0, 0, 0, 0, -1, 0, 1, -1, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, -1, -1, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 1, 2, 2, 1, 2, 2, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 2, 1, 0, 1, 0, 1, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -2, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 1, 0, -1, -2, -2, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 2, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 4, 3, 3, 4, 4, 3, 3, 1, 0, 0, 0, -1, -3, -1, -3, -2, 0, 0, 0, 1, 1, 1, 2, 2, 3, 4, 2, 2, 0, 1, 2, 1, 0, 0, 0, -1, -1, -3, -2, -2, -1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 4, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, -3, -4, -4, -4, -3, -1, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 1, 1, 0, 0, 1, 1, -2, -2, -1, -1, -2, -4, -5, -5, -2, -2, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, -1, -3, -1, -2, -4, -3, -4, -1, -2, -2, 0, 0, -1, 0, 0, 1, 0, 0, 0, 2, 1, 0, 0, 1, 0, 0, -2, -2, -2, -1, -3, -2, -2, -2, -1, -1, -2, -1, 0, 0, 0, 1, 0, 1, -1, 2, 0, 1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, -2, 0, 0, 0, 0, 2, 0, -2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 1, -1, -2, 0, 0, -1, -1, 0, 0, 0, 1, 1, 2, 1, 2, 2, 1, 2, 0, 0, 0, -1, -2, -2, -2, 0, -1, -2, -1, 0, 0, -1, 0, -1, 0, 1, 2, 2, 2, 2, 2, 4, 4, 3, 2, 1, 1, 0, 0, -2, -3, -1, -1, -2, -2, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 3, 2, 5, 4, 2, 3, 2, 2, 0, -1, -2, -2, -3, -1, -1, -2, 0, 0, 0, 0, -1, 0, 0, 2, 1, 2, 2, 3, 3, 2, 2, 4, 4, 3, 2, 0, 0, -2, -2, -2, -2, -3, -1, -1, -1, 0, 0, 0, 2, 2, 2, 0, 1, 2, 2, 3, 3, 4, 3, 3, 3, 1, 0, -1, -1, -2, -2, -2, -1, -1, 0, -1, 0, 0, 0, 2, 2, 0, 1, 0, 3, 3, 3, 3, 2, 3, 3, 1, -1, -2, -1, -1, 0, -1, -1, -1, -1, -1, -1, 0, 2, 2, 0, 0, 0, 3, 2, 2, 4, 2, 3, 4, 3, 1, 0, -1, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 1, 1, 1, 3, 2, 2, 1, 0, -1, -3, -1, 0, -1, 0, -2, -1, -1, 0, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -2, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -2, 0, -2, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, -2, -2, 0, -1, -2, -2, -3, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -2, -2, -1, -3, -3, -4, -2, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, -1, -1, -1, -2, -2, -1, -1, -3, -4, -2, -2, -3, -4, -2, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -2, -1, -3, -3, -3, -4, -4, -4, -1, -2, 0, 1, 1, 1, 0, 0, 0, 2, 3, 3, 0, 0, 0, 0, 0, -1, -3, -2, -1, -1, -3, -4, -4, -2, -3, 0, 0, 0, 0, 0, 0, 1, 1, 2, 3, 1, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, -2, -1, -3, -2, -1, 0, 0, 0, 1, 1, 2, 2, 1, 1, 3, 3, 0, 2, 1, 1, 0, 1, 0, -1, 0, -1, -1, -2, 0, 0, 0, -1, 1, 1, 1, 2, 2, 3, 3, 3, 2, 3, 1, 1, 1, 2, 2, 3, 1, 1, 1, 0, 0, 0, 1, 1, 1, 1, 2, 2, 3, 1, 2, 4, 5, 5, 0, -1, -1, 0, -1, 0, -2, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 1, 0, -1, -2, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, -2, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, -2, -1, -2, -2, -1, -1, -1, -1, -1, -1, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -2, -2, -1, -2, -1, -2, 0, -1, -1, 0, 1, 0, 0, 0, 1, 0, 0, 1, -2, -1, 0, 0, -1, 0, -1, 0, -1, 0, -2, -1, 0, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -2, -2, 0, 0, 0, 0, -1, 1, 0, 2, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, 0, 0, -2, -1, 0, -1, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -2, -1, 0, -1, -1, -1, -1, -2, 0, -1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, -1, -1, -1, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -2, -1, -1, 0, 0, -1, 0, 0, -2, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 2, 2, 2, 2, 1, 1, 1, 0, 1, 0, 1, 1, 0, 7, 5, 3, 0, 0, 0, 0, -2, -1, -4, -3, -4, -6, -5, -3, -3, 0, 0, -1, 0, 0, 0, 1, 3, 2, 3, 5, 4, 3, 1, 1, -1, 0, -1, -3, -2, -3, -3, -3, -2, -2, -2, -1, 1, 0, 1, 1, 2, 2, 2, 2, 4, 4, 3, 4, 1, 0, 0, 0, 0, -1, 0, -2, 0, -2, -1, -1, -1, 0, 2, 1, 3, 2, 1, 2, 3, 3, 3, 4, 4, 3, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 3, 1, 2, 1, 1, 3, 5, 3, 2, 1, 0, 0, 2, 1, 3, 1, 2, 2, 1, 0, 0, 0, 1, 1, 1, 3, 1, 0, 1, 1, 3, 3, 4, 3, 1, 1, 0, 0, 1, 3, 2, 2, 2, 1, 2, 0, 0, 0, 1, 1, 1, 1, 2, 0, 1, 1, 2, 2, 1, 2, 1, 0, 0, 0, 1, 2, 2, 3, 2, 3, 2, 0, 2, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, -1, 0, 0, 0, 1, 1, 3, 2, 3, 3, 1, 3, 2, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, -1, 1, 2, 3, 2, 2, 2, 2, 3, 2, 2, 3, 3, 1, 0, 0, -2, -2, -1, -1, 0, 0, 0, 2, 0, 0, 0, 0, 2, 4, 4, 4, 3, 1, 0, 1, 4, 2, 3, 2, 1, 0, -1, 0, -1, 0, 0, 1, 0, 2, 0, 0, 0, 1, 2, 3, 5, 3, 5, 3, 2, 4, 2, 2, 2, 2, 1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 2, 1, 3, 4, 6, 5, 6, 4, 4, 5, 4, 3, 3, 3, 0, 2, 1, 0, 2, 3, 2, 0, 0, 3, 2, 1, 2, 2, 5, 4, 4, 7, 5, 4, 6, 6, 5, 4, 3, 2, 2, 0, 0, 1, 4, 2, 2, 1, 0, 2, 1, 2, 3, 4, 4, 5, 6, 6, 6, 6, 7, 7, 7, 4, 4, 3, 2, 0, 2, 4, 3, 2, 2, 2, 0, 2, 2, 3, 4, 5, 5, 7, 6, 5, 6, 6, 6, 5, 5, 4, 2, 0, 2, 2, 2, 2, 3, 3, 2, 2, 1, 2, 2, 2, 2, 3, 3, 4, 5, 4, 4, 4, 3, 4, 4, 4, 3, 2, 2, 1, 2, 2, 4, 4, 4, 3, 0, 1, 2, 3, 2, 3, 4, 6, 5, 6, 2, 2, 3, 4, 4, 3, 3, 3, 3, 2, 3, 3, 5, 5, 2, 1, 0, 0, 1, 0, 0, 3, 3, 6, 4, 4, 4, 2, 3, 2, 4, 1, 3, 3, 3, 2, 3, 4, 4, 3, 2, 0, 0, 0, 0, 1, 0, 2, 3, 4, 5, 4, 3, 2, 3, 3, 3, 1, 1, 2, 3, 3, 3, 2, 1, 3, 1, 0, 0, 1, 1, 0, 0, 2, 2, 3, 2, 3, 3, 3, 2, 2, 1, 1, 0, 2, 1, 3, 2, 2, 3, 2, 2, 0, 1, 2, 0, 0, 0, 1, 2, 2, 2, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 1, 2, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 2, 1, 1, -1, 2, 0, 0, 0, 0, -1, -1, -2, -4, -4, -3, -2, -1, -2, -1, 0, 0, 0, 0, 0, 2, 2, 3, 2, 0, 0, 3, 3, 1, 2, 2, 0, 0, -2, -4, -4, -5, -3, -4, -4, -1, -1, 0, 1, 2, 1, 4, 4, 3, 1, 0, 0, 3, 3, 4, 2, 3, 0, -1, -3, -4, -5, -6, -6, -6, -4, -2, -2, 0, 1, 1, 2, 4, 3, 3, 3, 1, 1, 4, 3, 3, 2, 2, 1, -1, -3, -5, -8, -7, -8, -7, -3, -3, -1, 0, 0, 1, 1, 2, 3, 2, 1, 1, 4, 5, 2, 1, 1, 0, 0, 0, 2, 0, 0, 0, -1, -3, -4, -2, -1, 0, -1, 1, 0, 0, -1, -1, -1, 0, -2, 4, 3, 1, 1, 2, 1, 1, 0, 0, -1, -1, -1, -3, -2, -1, 1, 1, 1, 2, 0, 0, 0, 0, 0, -1, -1, 3, 2, 0, 0, 2, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 2, 1, 0, 0, 0, 1, 1, 0, 0, 4, 2, 1, 2, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 2, 0, 1, -1, 1, 1, 1, 1, 0, 0, -1, -1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, -1, 0, 3, 2, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 0, -2, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -2, 1, 1, 0, 0, 1, 0, 1, 1, 2, 3, 2, 2, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -3, 1, 0, -1, 0, 1, 1, 3, 4, 5, 3, 4, 4, 3, 3, 1, 1, 0, -1, 0, -1, -2, 0, 0, 0, -2, -2, 0, 0, -1, 0, 0, 3, 4, 5, 5, 4, 5, 5, 4, 2, 2, 2, 0, 0, 0, -1, -2, -1, -2, -2, -2, -3, 0, -1, 0, 0, 2, 3, 5, 6, 5, 5, 4, 5, 3, 2, 2, 1, 2, 0, 0, -1, 0, -1, 0, 0, -2, -1, 0, 0, -1, 0, 3, 4, 5, 6, 6, 6, 4, 4, 5, 2, 3, 1, 1, 1, 0, 0, -1, 0, -1, 0, 0, -2, -2, 0, 0, 0, 3, 3, 5, 7, 5, 4, 3, 3, 2, 3, 3, 2, 2, 2, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 4, 4, 6, 6, 6, 4, 5, 2, 3, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, -1, 1, 3, 2, 5, 6, 6, 6, 3, 4, 3, 3, 3, 2, 3, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 2, 2, 4, 4, 5, 6, 5, 3, 4, 3, 4, 3, 2, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 5, 4, 4, 5, 4, 4, 3, 2, 1, 1, 0, -1, -1, -1, 0, 0, 2, 1, 1, 0, -1, 1, 1, 0, 2, 1, 2, 3, 3, 4, 2, 1, 1, 0, 0, -1, -2, -2, -1, -1, 0, 1, 2, 0, 0, 0, -2, 1, 0, 1, 0, 2, 2, 2, 2, 3, 2, 1, 1, -1, 0, -2, -2, -1, 0, 0, 0, 1, 0, 1, 1, 0, -3, 1, 0, 0, 0, 0, 2, 1, 2, 1, 0, 0, -1, -1, -2, -3, -3, -1, 0, 0, 1, 1, 1, 1, 0, -2, -2, 0, 1, 0, 0, -1, 1, 0, 0, 0, 0, -1, -2, -1, -2, -2, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, -1, -2, -2, -1, -2, -1, -2, -3, -2, -2, 0, 0, 1, 1, 2, 1, 1, 1, 0, 0, 2, 1, 0, -1, 0, 0, 0, -3, -3, -4, -2, -2, -2, -1, -2, -1, 0, 0, 0, 1, 1, 2, 1, 0, 1, 0, 4, 1, 0, 1, 0, 0, -1, -2, -4, -4, -4, -2, -3, -1, 0, -1, 0, 0, 1, 0, 1, 2, 2, 0, 1, 0, 4, 0, 1, 0, 2, 0, 0, 0, -1, -3, -3, -3, -2, 0, 0, 0, 1, 2, 1, 1, 1, 1, 1, 1, 1, 0, 4, 2, 1, 1, 1, 1, 0, 0, -2, 0, -1, -1, 0, 0, 1, 1, 2, 3, 2, 3, 1, 2, 1, 2, 2, 0, -2, -2, -2, -1, 0, -1, 0, -1, -1, 1, 0, 1, 0, 0, 0, -2, 0, -1, -3, -1, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 1, 2, 0, 0, 0, 0, -1, 0, -2, 0, -1, -1, 0, 0, -2, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, 1, 0, 2, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, -1, 1, 1, 0, 0, 2, 2, 1, 2, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 0, 2, 1, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 1, 2, 1, 2, 1, 0, 0, 2, 0, 1, 0, 1, -1, 0, 0, -1, 0, 1, 0, 0, -2, -1, 0, 0, 1, 1, 3, 2, 3, 0, 1, 1, 0, 0, 1, 2, 0, 0, 0, -1, -1, 0, -1, 0, 0, -2, -2, 0, 0, -1, -1, 0, 0, 3, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, -1, 0, -1, 0, 0, -1, -3, -2, -2, -1, 0, 0, 1, 1, 2, 1, 0, 1, 0, 0, 0, 2, -1, 0, 1, 0, 0, 0, 0, -2, -1, -1, -3, -2, -2, -3, 0, 0, 0, 1, 0, 1, 2, 1, 0, 0, 2, 1, -2, 0, 0, 1, -1, 0, 0, 0, -2, -2, -2, -3, -2, -3, -1, -1, -2, 0, 0, 1, 1, 1, 0, 2, 0, 1, -3, 0, 0, 0, 0, 0, -1, -2, -2, -3, -4, -2, -2, -4, -2, -2, -1, -2, 0, 1, 2, 1, 0, 0, 1, 1, -2, 0, 0, 0, 0, -1, -3, -2, -2, -1, -2, -3, -2, -3, -2, -1, -2, 0, 0, 1, 2, 0, 1, 1, 1, 0, 0, -1, 0, 0, -1, -2, 0, -1, 0, -2, -4, -2, -1, -3, -1, -1, -2, 0, 0, 2, 2, 0, 1, 0, 0, 0, -1, 0, 0, -2, 0, 0, 0, 0, -1, 0, -3, -2, -3, -1, 0, -2, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 2, 1, 0, -1, -2, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -2, -2, -1, 0, 0, 0, 1, 0, 0, 1, 2, 2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, 0, -1, 0, 0, 1, 0, 1, 0, 3, 1, 2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -3, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -2, -3, -2, -1, -1, -1, -1, -1, 0, 0, 1, 0, 2, 0, 2, 0, 1, 0, 0, 0, 0, -1, -2, -2, -2, -1, -2, -1, -1, -1, 0, 0, -2, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, -3, -2, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -2, 0, 0, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 1, 0, -2, -1, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, -1, 0, -1, 0, -2, -2, -2, -2, -1, -1, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, -1, -1, -1, -1, 0, 0, 0, 0, -2, -1, -1, 0, -1, -2, -2, -3, -1, -2, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, -2, -2, -1, 0, 0, -1, 0, -2, -3, -1, -1, -2, -2, -2, -1, -1, -1, 0, -1, 0, 2, 0, 1, 0, 0, -1, -1, 0, 0, -1, 0, -2, -1, -2, -1, -1, -3, -2, -3, -1, -3, -2, -1, -2, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -2, -1, -3, -2, -2, -2, -1, -2, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -2, -2, -1, -3, -3, -2, -3, -1, -2, -1, 0, -1, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, -2, 0, 0, -1, -1, -1, -1, -3, -2, -2, -1, -2, -1, -1, 0, -1, 0, 0, 0, 2, 1, 0, 0, 0, -2, 0, 0, 0, 0, -2, -1, -3, -1, -1, -2, -2, 0, -1, -2, -1, -1, 0, 0, 0, 3, 1, 0, 0, -1, -1, -1, -1, 0, -2, -1, -2, -1, -3, -3, -2, -1, -2, -1, 0, -2, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, -2, -2, -1, -1, -1, -1, -2, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, 2, 0, 0, 0, 0, -1, 0, -1, -2, -2, -3, -2, -2, -2, -2, -3, -1, -1, -1, 0, 0, 0, 1, 2, 1, 2, 0, 0, -1, -1, 0, -1, -1, 0, 0, -2, -2, -2, -3, -1, -1, -1, -1, 0, 0, 0, 0, 2, 2, 1, 2, 0, 1, 0, 0, -1, 0, 0, 0, 0, -2, -1, -1, -1, -3, -3, -1, -1, 0, 0, 0, 1, 2, 2, 2, 2, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, -2, -3, -3, -2, 0, 0, -1, 0, 2, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, -2, -2, -1, -1, -1, 0, -1, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -2, -2, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 2, 1, 1, 1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, -2, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 2, 0, 1, 0, 0, -1, -2, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 1, 2, 1, 0, 0, 0, -2, -1, -1, -1, 0, 0, -1, -1, 0, 0, 1, 0, 1, 1, -1, -1, 0, 1, 0, -1, 2, 0, 0, 0, 0, -1, -1, -2, -2, -1, 0, 0, 0, 0, -1, 1, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 2, 1, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, -1, 1, 2, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, -1, 0, 0, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, -1, 1, 1, 1, 0, 1, 0, 0, -1, 0, -1, -1, -1, -1, -2, -1, 0, -1, 0, 0, 1, 1, 2, 0, 0, 0, 1, 0, 0, 3, 2, 1, 0, 0, -1, -2, -2, -1, -2, -1, 0, 0, -1, 0, 0, 0, 1, 2, 2, 0, 0, 0, 1, 0, 2, 3, 4, 3, 2, 0, -1, 0, -2, -2, -3, -2, -1, -1, 0, 0, 0, 2, 1, 2, 1, 0, 1, 0, 1, 1, 3, 4, 2, 4, 1, 0, 0, -1, -2, -2, -2, -3, -1, -1, 0, 0, 1, 1, 2, 2, 2, 2, 1, 0, 1, 1, 3, 5, 3, 4, 1, 0, -2, -2, -3, -2, -4, -3, -1, 0, 0, 1, 0, 2, 1, 2, 2, 0, 0, 0, 1, 1, 3, 4, 4, 3, 3, 0, 0, -2, -2, -2, -3, -2, -2, -1, 0, 0, 1, 2, 1, 2, 0, 1, 1, 0, 1, 2, 2, 4, 4, 3, 3, 0, -2, -2, -2, -1, -2, -3, -1, -2, 0, 0, 2, 2, 2, 2, 0, 1, 0, 0, 2, 3, 4, 3, 4, 4, 3, 0, -2, -2, -3, -2, -2, -3, -3, -2, 0, 2, 1, 2, 1, 0, 0, 1, 2, 1, 1, 3, 3, 3, 3, 2, 1, 1, -2, -1, -2, -3, -2, -3, -3, 0, 1, 1, 3, 3, 2, 0, 0, 2, 1, 1, 1, 1, 3, 2, 2, 3, 0, 0, -1, -1, -4, -2, -2, -1, -2, 0, 1, 1, 2, 2, 1, 2, 0, 1, 2, 0, 1, 2, 2, 1, 3, 1, 2, 0, 0, -3, -2, -2, -1, -2, -1, 0, 0, 2, 1, 2, 0, 1, 1, 1, 2, 1, 1, 1, 2, 1, 1, 2, 2, 1, 0, -2, 0, -1, -2, 0, -1, -1, 0, 1, 2, 2, 0, 0, -1, 2, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 2, 0, 0, 2, 3, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 1, 1, 1, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -2, -1, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 2, 0, 1, 0, 0, -1, -1, -2, -1, -1, 0, 0, 1, 2, 1, 0, 1, 0, 1, 0, 0, 2, 0, 1, 2, 3, 3, 2, 0, 0, 0, 0, -2, -1, -1, 0, 0, 2, 1, 2, 2, 2, 1, 0, 1, 1, 0, 1, 2, 1, 1, 4, 3, 5, 3, 4, 3, 2, 0, 1, 1, 1, 1, 0, 0, 2, 2, 3, 3, 3, 4, 7, 7, 7, 9, 6, 0, 0, 0, 1, 1, 1, 1, 1, 0, -1, -1, -2, -1, -1, 0, 1, 2, 2, 2, 1, 1, 3, 4, 5, 6, 5, 0, 0, 1, 1, 0, 0, 0, 0, -1, -2, -4, -3, -1, -1, 0, -1, 0, 0, 1, 0, 1, 0, 2, 4, 6, 6, 0, 0, -1, 0, -1, 0, -1, -1, -2, -6, -5, -4, -4, -1, -3, -3, -2, 0, -1, 0, 1, 0, 1, 3, 4, 4, 0, -1, 0, 0, 0, 0, -3, -3, -4, -4, -5, -5, -5, -4, -3, -4, -4, -1, 0, 0, 1, 0, 0, 0, 2, 0, 0, 0, 0, 0, -2, -3, -3, -5, -4, -4, -5, -3, -5, -4, -4, -4, -2, -1, -1, 0, 0, 0, 2, 0, 1, -1, -1, 0, 0, 0, 0, -3, -5, -4, -3, -3, -3, -4, -4, -4, -2, -2, -3, -1, -1, 0, 0, 1, 2, 1, 0, -2, 0, 0, -1, 0, -1, 0, -2, -3, -3, -1, -2, -1, 0, -2, -3, -1, -3, -2, 0, -1, 0, 1, 1, 1, 0, -2, 0, -1, 0, 0, 0, -2, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, -1, -3, -2, -1, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 1, 1, 2, 2, 1, 0, -2, -2, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 2, 2, 1, 0, -2, -2, -1, -2, -2, -3, -2, -2, -2, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 2, 2, 2, 1, 3, 2, 1, 0, -1, -1, -3, -1, -1, -2, -3, -2, 0, -1, -1, -2, -1, -1, -2, -2, -2, 0, 0, 1, 0, 2, 1, 3, 4, 1, 0, -2, -3, -2, -2, -3, -2, -1, 0, -1, -1, -2, -2, -2, -3, -3, -3, -2, 0, 0, 1, 2, 1, 4, 4, 3, 0, -2, -3, -3, -2, -1, -2, -1, 0, 0, -2, -1, -1, -1, -1, -3, -1, -1, 0, 1, 1, 2, 4, 4, 4, 3, 0, -2, -4, -1, -1, 0, 0, 0, -2, -1, -2, -1, -2, -2, -1, 0, -1, 0, 0, 1, 2, 1, 4, 4, 3, 0, -2, -3, -3, -2, -2, 0, 1, 2, -1, -1, -1, -1, -1, 0, 0, -2, -1, 0, 0, 1, 0, 0, 2, 3, 2, 1, -1, -3, -3, -3, -2, 1, 2, 3, -1, 0, -1, -1, -3, -2, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -3, -2, -2, -2, 0, 1, 2, -2, 0, -1, -4, -3, -2, -1, 0, -1, -1, -3, -2, -2, -3, -2, -2, -1, 0, -2, -2, -1, -2, 0, 0, 2, 3, -2, -1, -1, -3, -3, -4, -1, -1, -2, -2, -4, -3, -4, -2, -3, -2, -1, 0, -2, -2, -1, -1, -1, 0, 2, 3, -1, 0, 0, -3, -3, -1, -2, -1, -3, -2, -5, -5, -4, -5, -3, -2, -2, -1, 0, -1, 0, -1, 1, 2, 3, 3, 0, 0, 0, 0, 0, 0, -2, -3, -3, -3, -4, -4, -5, -5, -4, -2, 0, 0, 0, 0, 0, 0, 1, 2, 4, 5, 1, 0, 0, 0, 0, 0, 0, -3, -3, -3, -2, -3, -3, -2, -3, -3, -1, 0, 0, 0, 0, 1, 1, 4, 7, 7, 1, 2, 0, 0, 1, 0, 0, -2, 0, -2, -2, -2, -2, -3, -2, -1, 0, 0, 1, 0, 1, 2, 3, 8, 9, 8, 2, 0, 2, 0, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 1, 2, 2, 3, 5, 7, 10, 8, 0, 2, 1, 3, 2, 3, 1, 3, 4, 2, 3, 2, 1, 0, 0, 0, 0, 3, 2, 3, 3, 5, 7, 9, 10, 10, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 3, 2, 4, 3, 4, 2, 2, 2, 0, 2, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 3, 1, 3, 2, 3, 2, 3, 3, 1, 0, 2, 0, 1, 0, 0, -1, 0, -1, -2, -1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 3, 3, 3, 2, 2, 1, 1, 0, 0, 0, 0, -1, -1, -2, -3, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 1, 2, 0, 0, 0, 0, 0, -2, -3, -1, -4, -3, -1, -2, 0, -2, 0, -1, 0, -1, -1, -1, 0, 1, 2, 1, 1, 0, 1, 1, 0, 0, -2, -3, -3, -2, -4, -2, -2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 1, 2, 1, 0, 0, -1, -2, -1, -3, -3, -2, -1, -1, -2, -2, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 2, 0, 0, 1, 0, -1, -1, -1, -2, 0, -1, -1, -2, -3, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -2, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 1, 1, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, -1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, 0, -2, -1, -1, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, -1, -1, 1, 0, 1, 0, 1, 0, 1, 1, 0, -2, -2, -1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, -1, -2, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, -1, -2, -2, 0, 0, 0, 1, 1, 3, 1, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, -1, -2, -1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 0, 1, 0, 0, -1, -1, -1, 0, 0, -2, -1, -1, 0, 0, -2, -1, -1, 0, 1, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, -2, -1, 0, -2, -2, 0, 0, -1, -1, 0, 0, 0, 2, 0, 2, 0, 1, 1, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 1, 1, 0, -1, 0, 0, 0, 0, -2, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 3, 4, 5, 2, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 4, 5, 2, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 3, 4, 3, 4, 2, 0, 1, 0, 0, 0, 0, 2, 3, 3, 2, 2, 1, 3, 1, 1, 2, 3, 2, 1, 2, 2, 3, 4, 3, 4, 4, 3, 1, 0, 1, 0, -2, -4, -5, -5, -3, -2, -3, -5, -2, -4, -2, -3, -3, -3, -1, 0, -1, 0, -1, 0, 4, 2, 2, 0, -1, -1, -2, -3, -4, -3, -3, -1, -2, -1, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 4, 4, 1, 0, 0, 0, -1, -3, -1, -2, -1, -1, -1, 0, 0, 0, 0, 1, 2, 2, 2, 0, 0, 0, -1, 0, 4, 4, 3, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 2, 4, 1, 0, 0, 1, 1, 4, 3, 4, 1, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 1, 0, 1, 1, 2, 2, 2, 0, 0, 0, 1, 4, 5, 3, 3, 0, 1, 2, 1, 1, 2, 3, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 3, 5, 2, 0, 0, 0, 2, 2, 1, 3, 3, 2, 1, 1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 1, 2, 4, 2, 3, 2, 1, 4, 2, 4, 2, 1, 2, 2, 1, 1, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, 0, 2, 3, 3, 2, 1, 3, 3, 6, 5, 3, 3, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 1, 2, 2, 4, 6, 5, 6, 3, 3, 1, 0, 0, 0, -1, -1, 0, 1, 1, 0, 0, 1, 0, 2, 2, 2, 5, 4, 4, 4, 5, 5, 8, 8, 4, 3, 0, 1, 0, 0, -1, -1, 0, 0, 2, 0, 3, 3, 2, 2, 1, 2, 5, 4, 2, 5, 4, 6, 8, 8, 8, 4, 2, 0, -1, 0, 0, 0, 0, 1, 2, 2, 3, 4, 3, 3, 0, 0, 5, 5, 3, 4, 6, 7, 8, 8, 7, 6, 4, 2, 1, 0, -1, -1, -1, 0, 0, 2, 2, 4, 4, 2, 1, -1, 5, 5, 6, 6, 8, 7, 9, 9, 8, 6, 4, 3, 2, 0, 0, -1, -1, 0, 0, 1, 5, 4, 5, 2, 2, 0, 4, 4, 7, 5, 8, 9, 8, 8, 8, 4, 3, 2, 1, -1, 0, -1, -1, 0, 0, 3, 3, 5, 5, 4, 0, 0, 5, 5, 6, 7, 9, 8, 8, 9, 7, 4, 4, 0, 0, 0, -1, 0, 0, 0, 2, 1, 5, 6, 5, 4, 2, -1, 4, 5, 4, 5, 5, 6, 6, 7, 7, 5, 3, 2, 0, 0, 0, 0, 0, 0, 1, 3, 6, 6, 7, 5, 1, 0, 2, 3, 3, 5, 5, 6, 6, 6, 6, 6, 3, 1, 1, 1, 1, 2, 2, 2, 3, 4, 5, 5, 5, 3, 0, -1, 4, 3, 3, 3, 3, 4, 6, 5, 4, 5, 4, 1, 0, 0, 1, 2, 4, 4, 4, 2, 4, 3, 3, 3, 1, 0, 4, 3, 4, 3, 3, 5, 6, 6, 6, 4, 4, 2, 2, 0, 1, 3, 3, 2, 2, 2, 2, 4, 3, 2, 2, 0, 6, 5, 1, 2, 3, 3, 5, 3, 4, 4, 3, 3, 0, 0, 0, 2, 2, 1, 2, 1, 1, 3, 3, 3, 1, -2, 3, 3, 1, 3, 1, 2, 4, 3, 1, 3, 2, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 2, 1, 0, -2, 2, 3, 1, 0, 0, 2, 3, 1, 0, 1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, -2, 2, 3, 3, 1, 0, 1, 0, 0, -2, -1, 0, -1, -1, 0, 0, 0, 2, 2, 0, 1, 1, 2, 0, 0, 0, 0, 4, 1, 3, 3, 0, 0, -1, 0, -2, -3, -2, -2, -2, -1, 0, 1, 2, 1, 0, 1, 2, 1, 1, 2, 0, 1, 2, 2, 3, 1, 2, 0, -1, -2, -4, -4, -6, -4, -2, -3, -1, -1, 0, 1, 2, 1, 2, 2, 2, 1, 1, 0, 2, 2, 2, 1, 0, 0, 0, -1, 0, -1, -1, -2, -3, -1, -3, -1, -2, 0, -1, 0, -1, -1, 0, -1, 0, -2, 1, 1, 0, 0, -1, -1, 0, -1, -1, -2, -3, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, -1, -2, -2, -1, -2, -2, -1, -1, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 2, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, -2, -3, 0, 0, -1, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -2, -3, 0, 0, 0, 0, 1, 0, 1, 1, 2, 3, 3, 1, 1, 2, 0, 0, 0, 0, -3, -1, -2, -1, 0, -1, -3, -4, 0, 0, 0, 0, 1, 3, 2, 5, 4, 4, 4, 3, 2, 3, 0, 1, -1, -2, -1, -3, -2, -1, -3, -2, -2, -2, 0, 0, 0, 2, 1, 4, 5, 4, 5, 4, 4, 4, 4, 3, 3, 1, 0, -2, -1, -2, -3, 0, -1, -1, -1, -4, 0, 0, 0, 1, 2, 5, 4, 4, 4, 5, 5, 5, 3, 3, 2, 0, 0, -2, -3, -2, -3, -1, -1, -2, -2, -3, 0, 0, 0, 2, 1, 3, 5, 5, 3, 5, 5, 3, 4, 2, 2, 2, 0, -2, -2, -2, -2, 0, 0, -1, -1, -2, 0, 0, 0, 0, 4, 4, 5, 4, 4, 4, 3, 4, 4, 4, 2, 2, 0, -1, -2, -2, -1, 0, 0, 0, 0, -2, -1, 0, 0, 1, 4, 4, 4, 3, 5, 4, 3, 3, 2, 1, 1, 2, 0, -1, -2, -1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 2, 2, 4, 4, 4, 5, 2, 3, 2, 3, 2, 0, 1, 0, -1, -2, -1, -2, 0, 1, 1, 0, 0, 0, 1, 1, 2, 2, 4, 5, 5, 3, 2, 3, 1, 2, 1, 0, 0, 0, -2, -2, -2, 0, 0, 1, 1, 0, -1, 0, 0, 0, 2, 1, 3, 4, 3, 2, 1, 1, 0, 0, -1, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 1, 1, 1, 0, 0, -2, -1, -2, -2, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 0, 2, 0, 0, 0, 0, -1, -1, -3, -1, -2, 0, -1, 0, 0, -1, 0, -1, 0, -1, 1, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, -1, 0, -1, 0, 0, -3, -2, -2, -1, -2, -1, -1, -2, -2, -1, 1, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, -2, -3, -3, -2, -2, -3, -4, -3, -2, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -2, -2, -4, -3, -2, -2, -3, -2, -2, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, -1, -3, -3, -3, -3, -2, -3, -3, -1, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -3, -4, -2, -3, -3, -3, -1, -1, 0, 0, 0, 0, 1, 1, 2, 1, 1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, -1, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -2, 0, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -2, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, 0, -1, -2, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, 2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 0, 1, 0, 1, 1, 2, 4, 2, 2, 2, 2, 0, 0, 0, 0, 1, 0, 2, 0, 2, 2, 2, 2, 2, 1, 3, 2, 2, 1, 2, 2, 1, 2, 2, 2, 0, 2, 0, 1, -1, 0, -1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 2, 1, 1, 1, 0, 1, 0, -2, -1, -1, -1, 1, 1, 0, 1, 1, 1, 1, 1, 1, 2, 0, 0, 1, 0, 0, 1, 0, 2, 0, 0, 0, -1, -3, -2, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, -1, -1, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 2, 0, 0, 0, 0, -1, -1, 0, -2, -2, -1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 0, 1, 0, 2, 1, 0, 1, 1, 0, 0, -1, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 1, 1, 2, 2, 2, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 2, 1, 3, 1, 2, 1, 2, 3, 4, 2, 3, 0, 0, 0, -1, -1, 0, -1, -1, 0, -2, 0, -1, 0, -1, 1, 2, 2, 3, 0, 2, 2, 4, 4, 3, 2, 2, 1, 0, 0, 0, 0, -1, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 3, 3, 2, 2, 1, 2, 1, 1, 1, 0, 0, -2, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 2, 2, 1, 2, 2, 3, 1, 3, 1, 1, 2, 3, 2, 0, -1, -2, -1, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 2, 2, 2, 3, 2, 1, 3, 2, 1, -1, -1, -1, 0, -2, -2, 0, 0, 1, 0, 1, 0, 0, 0, 1, 2, 1, 3, 3, 2, 4, 2, 3, 4, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 1, 3, 1, 3, 1, 2, 1, 1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 2, 0, 1, 0, 1, 0, 1, -1, 0, -1, 0, -1, 0, -1, -2, 0, -2, 0, 0, 1, -1, 0, 0, 0, 1, 0, 0, 1, 0, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, -3, -2, -1, -2, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, -1, -1, -2, -1, -2, 0, -2, -3, 0, -1, 0, 1, 0, 1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, -1, -1, 0, 2, 2, 2, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 2, 3, 4, 2, 1, 0, 0, 0, -1, -2, -3, -2, -4, -3, -4, -4, -4, -3, -1, 0, 0, 0, 0, 1, 3, 2, 4, 3, 2, 2, 2, 1, 0, -1, -2, 0, -1, -4, -3, -3, -4, -3, -3, -3, -2, 0, 0, 0, 0, 0, 3, 3, 3, 2, 1, 2, 2, 0, 0, 0, -1, 0, -1, -4, -5, -4, -3, -3, -3, -2, -2, -1, -1, 0, -1, 0, 1, 2, 2, 1, 1, 2, 1, 1, 0, -1, -1, 0, -1, -2, -4, -2, -2, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -3, -1, -3, -2, -1, -1, 0, -1, 0, -2, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, -1, -1, -1, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -2, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, -2, -3, -3, -1, -1, -1, -1, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 3, 2, 3, 3, 2, 0, -1, -2, -2, -2, -1, -1, -1, -2, -2, 0, 0, 0, -1, 0, 2, 0, 0, 3, 3, 2, 3, 2, 3, 5, 2, 0, -1, -1, -1, -1, -1, -1, -2, -2, -2, 1, 0, 0, 0, 0, 1, 2, 1, 2, 4, 4, 4, 5, 6, 3, 3, 0, 0, -1, -1, -3, -2, -1, 0, -1, -2, 0, 0, 0, 0, 1, 1, 2, 2, 4, 4, 6, 5, 7, 5, 5, 4, 2, 0, -2, -2, -2, -1, -1, -1, -1, -2, 0, 0, 0, 0, 1, 1, 1, 2, 4, 5, 5, 5, 6, 6, 5, 3, 3, 0, 0, -3, -2, -2, -2, -1, -2, -2, 0, -1, 0, 0, 0, 1, 2, 1, 2, 4, 6, 5, 6, 5, 6, 5, 3, 0, -2, -2, -4, -1, -2, 0, 0, 0, 0, 0, -2, -1, 0, 1, 1, 0, 2, 3, 4, 5, 6, 6, 5, 5, 3, 1, -2, -3, -1, -1, 0, -1, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 1, 4, 5, 3, 5, 4, 4, 3, 1, 0, -1, -2, -3, -3, -2, -2, 0, -2, -2, -1, 0, 0, 0, 0, 1, 0, 1, 2, 4, 2, 4, 4, 3, 3, 2, 0, 0, -2, -2, -3, -3, -3, -2, -1, -1, 0, -1, 0, -2, 0, 1, 0, 0, 2, 1, 1, 3, 1, 1, 0, 0, 0, -1, -3, -1, -3, -1, -3, -1, -2, -2, 0, 0, -2, -1, -1, 0, 1, 1, 0, 2, 0, 0, 0, 0, -1, -1, -1, -1, -1, -2, -2, -3, -3, -1, -2, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, -1, -1, -1, -1, -1, -2, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, -1, -2, -1, -1, -2, 0, -2, 0, -1, -2, -1, -1, -1, 0, -2, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -2, 0, -1, -1, 0, -3, -1, -2, -3, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 1, 1, -1, -1, -2, -2, -1, -2, -3, -3, -3, -2, 0, -1, 0, 0, -1, 0, 0, 0, 1, 2, 1, 0, 0, 0, 2, 2, 1, -1, -3, -2, -1, -2, -2, -4, -2, -2, 0, -1, -1, 0, 0, 1, 1, 1, 2, 2, 2, 1, 0, 2, 2, 1, 1, 0, -2, -2, -1, -1, -2, -3, -3, -1, 0, 0, 0, 0, 0, 1, 2, 3, 4, 4, 2, 2, 1, 2, 4, 3, 3, 2, 0, -2, -3, -3, -2, -4, -3, -2, 0, -2, 0, 0, 0, 1, 1, 3, 4, 4, 4, -3, -4, -1, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, -1, -2, -2, -1, -1, 0, 0, 0, -1, -1, -3, -1, -1, -1, -1, 0, -1, -2, -2, -1, -2, -2, -1, -2, -1, -1, 0, -1, -2, -2, -1, 0, 0, -1, 0, 0, -3, 0, -1, -1, -1, -1, 0, -1, -2, -1, -2, 0, -1, -1, -1, -1, 0, -1, 0, -1, -2, 0, 0, -1, 0, -1, -1, -2, -1, -1, 0, -1, -2, -1, -2, -2, -1, -2, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -2, -2, 0, 0, 0, 0, -2, -1, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -2, 0, -2, -2, -1, -1, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -2, -2, -2, -1, -1, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, -2, -2, -1, 0, -1, -2, -2, -2, 0, -1, -1, -1, -1, 0, -1, 0, 0, -2, -1, 0, -1, 0, -2, 0, -2, -1, 0, -4, -2, -1, -1, -1, -2, -2, -2, -3, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -2, 0, -1, 0, -2, -2, -1, 0, -1, -2, -3, -2, -1, -1, -1, 0, 0, 0, -1, 0, -1, -1, -2, 0, -1, -2, -2, -1, -2, 0, -2, -4, -2, -1, -2, -2, -1, -2, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -2, -3, -1, -2, -2, -1, -2, -2, -1, -2, -1, -1, -3, -3, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, -2, 0, -1, -2, -2, -1, -2, -1, -2, -1, -2, -2, -2, -1, -3, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -2, -2, -3, -1, 0, -2, -2, -2, 0, -2, 0, -2, -3, -2, -1, -2, -1, -1, -1, 0, 0, -1, 0, -1, -1, -1, -1, -2, -3, -3, -3, -3, -3, -2, -1, 0, -2, -2, -3, -1, -2, -2, -2, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, -2, -3, -1, -2, -2, -1, -2, -1, 0, -1, -3, -2, -2, -1, 0, 0, -2, -1, -1, -1, 0, 0, -1, 0, -1, 0, -3, -2, -2, -2, -2, -3, -2, -2, 0, -2, -1, -3, -2, -2, -2, 0, 0, -2, 0, 0, -1, -1, -1, 0, -2, 0, -2, -2, -1, -4, -2, -2, -2, 0, 0, -1, -1, -2, -3, -2, -1, -1, -2, -1, -2, 0, -1, -1, 0, -1, -1, -1, -1, -3, -2, -2, -2, -2, 0, -1, 0, 0, -2, -2, -2, -2, -1, -1, -2, 0, -1, -1, -2, 0, -1, 0, 0, -1, -2, -1, -2, -2, -2, -2, -1, 0, -1, 0, 0, -2, -2, -1, -2, -1, -2, -2, -1, 0, -1, -1, -1, -1, -3, -2, -2, -1, -1, -1, -1, -3, 0, 0, 0, 0, 0, -1, -2, -2, -2, -2, -1, -1, -1, -1, -2, -2, -2, -2, -1, -2, 0, -1, -2, 0, -2, -2, 0, -1, 0, 0, 0, 0, -1, -1, -2, -1, -2, -1, -3, -3, -2, -1, -2, -1, -1, -2, -1, -2, 0, -1, -2, -1, -1, -1, -1, 0, 0, -2, -1, -2, -1, -1, -2, -1, -2, -1, -3, -2, -1, -2, 0, 0, -2, -2, -1, -2, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -2, -3, -3, -2, -2, -2, -2, -2, -1, 0, 0, -1, 0, 0, -3, -1, 0, 0, 0, 0, -1, 0, -1, -2, 0, -2, -2, -2, -1, -2, -3, -2, 0, -2, -1, -2, -1, 0, -1, -1, -4, -2, -1, 0, -1, 0, -1, -1, -1, -1, -2, -1, -2, -2, -2, -1, 0, -2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, -1, 0, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 3, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -2, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, -1, -2, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, -2, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, -1, -2, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -2, -1, -1, -2, -1, 1, 1, 0, 0, -1, 0, 0, -1, -1, -1, -2, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -2, -2, 0, -1, 1, 0, 0, 0, -1, 0, -2, -1, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, -1, 0, -1, 0, -1, 0, 0, 1, 0, 1, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, -1, -1, -1, 0, 1, 0, 0, 0, 0, 2, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, -3, -3, -2, -2, -1, 0, 1, 0, 0, 0, 1, 2, 1, 1, -1, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, -3, -2, -3, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, 0, -2, -3, -1, 0, 0, 0, -1, 0, 0, 0, 2, 0, 1, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, -2, -1, 2, 0, 1, 1, 0, 0, -1, -2, -2, -1, 0, -1, 0, -1, 0, -2, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 1, 1, 1, 0, 1, -1, -1, -1, -1, -2, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, -2, -1, 2, 0, 0, 1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 1, 2, 1, 0, 0, 1, 1, 0, -1, -1, 0, 0, 0, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 1, 2, 0, 1, 1, 0, 1, 0, 0, 1, 1, 0, 2, 1, 2, 1, 2, 0, 0, 1, 0, -1, 0, 1, 0, 3, 3, 4, 3, 3, 2, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 2, 1, 2, 5, 3, 3, 3, 1, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, -2, -2, -1, -1, -1, 0, 0, 0, 2, 1, 3, 3, 5, 3, 3, 2, 1, 0, 0, 0, -2, -2, -2, -2, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 2, 1, 2, 2, 5, 3, 2, 2, 0, 1, 0, 0, -3, -3, -2, -1, -2, -1, 0, 1, 0, -1, -1, 0, 0, 1, 0, 1, 2, 2, 4, 1, 1, 2, 1, 1, 0, -1, -1, -1, -2, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 4, 3, 0, 1, 0, 0, 0, -2, -3, -1, -3, -1, -2, -1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 1, 2, 3, 2, 0, 0, 0, 0, 0, -2, -2, -2, -3, -4, -2, -1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 3, 1, 1, 1, 0, 0, -2, -2, -2, -2, -3, -2, -2, -2, 0, 0, 0, 1, 0, 1, 0, -1, -1, 1, 1, 3, 2, 1, 0, 0, -1, -2, -3, -2, -3, -2, -3, -3, -1, -2, -1, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 2, 2, 0, 0, 0, -1, -4, -5, -3, -3, -4, -3, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 0, -1, -3, -5, -4, -3, -4, -4, -1, -2, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 3, 1, 0, -1, -3, -4, -4, -4, -3, -4, -2, -2, -2, 0, 0, 0, 1, -1, -1, -1, -1, -1, 0, 1, 2, 2, 4, 1, 0, 0, -3, -4, -3, -5, -4, -4, -3, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, -1, 1, 1, 3, 1, 3, 0, 0, -2, -3, -4, -5, -5, -5, -4, -2, -3, -3, -2, -1, -1, 0, 0, 0, -1, 0, 0, 1, 2, 1, 3, 3, 0, 0, -2, -1, -4, -3, -3, -4, -5, -3, -3, -1, 0, -2, -1, 0, 0, 0, -1, -1, 0, 1, 1, 2, 2, 4, 1, 0, -1, -2, -3, -3, -3, -4, -3, -4, -3, -3, -2, -2, 0, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 0, 0, 0, -2, -4, -3, -2, -4, -4, -1, -2, -2, -3, -1, -2, -1, 0, -1, 0, 0, 0, 0, -1, -1, 4, 1, 0, 0, -2, -1, -3, -2, -2, -3, -3, -3, -3, -3, -1, -1, -1, -1, -1, 0, -1, -1, 0, 0, -1, 0, 4, 2, 1, 0, -1, -1, -2, -2, -1, -1, -2, -3, -3, -2, 0, 0, 0, -2, -2, -1, -3, -3, -1, -1, 0, 1, 3, 4, 2, 0, 0, -2, -1, -1, -2, -3, -4, -3, -2, -1, 0, -1, 0, -1, -2, -2, -3, -3, -2, -2, 0, 2, 4, 4, 2, 2, -1, 0, -2, -2, -1, -2, -2, -3, 0, 0, 0, 0, -1, -1, -3, -3, -3, -4, -3, -1, 0, 1, 6, 5, 4, 1, 1, 0, -2, 0, 0, -2, -2, 0, 0, -1, 0, 0, -1, -2, -3, -4, -3, -4, -2, -2, -1, 2, 6, 5, 4, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, -2, -3, -3, -3, -3, -2, -3, 0, 2, 6, 6, 5, 3, 2, 1, 1, 1, 0, 0, 1, 1, -1, -1, -1, 0, -3, -3, -2, -2, -4, -2, -3, -1, 0, 0, 7, 7, 5, 4, 3, 2, 3, 1, 1, 1, 0, 0, 0, 0, -2, -1, -3, -1, -1, -1, 0, -3, -2, 0, 0, 1, 5, 5, 6, 6, 4, 2, 4, 3, 1, 3, 1, 1, 0, 0, 0, 0, -2, -1, -2, 0, -1, -1, -1, 0, 0, 1, 2, 3, 3, 3, 4, 3, 4, 3, 1, 2, 2, 1, 1, 0, 0, 0, 0, 2, 2, 2, 3, 3, 4, 5, 5, 5, 1, 1, 3, 3, 2, 3, 2, 2, 2, 0, -1, -1, -1, 0, 1, 1, 1, 2, 1, 0, 2, 3, 3, 3, 3, 3, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -2, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 3, 1, 3, 1, 0, 1, 0, 1, 0, 0, 0, -1, -3, -4, -2, -2, -2, -2, 0, 0, -2, -2, 0, 0, 0, 0, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, -3, -2, -4, -3, -4, -3, -3, -1, -2, -1, -1, 0, -1, -1, 0, 2, 0, 0, 2, 1, 1, 1, 0, 0, 0, -1, -3, -3, -3, -2, -2, -2, -3, -2, -2, -2, -1, -2, 0, 0, 0, 0, 0, 2, 2, 2, 0, 1, 0, 0, 0, -1, -1, -2, -1, -2, 0, 0, 0, -2, -1, -2, -1, 0, -2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -2, -1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 1, 0, 0, 0, -2, 0, 0, -2, 0, 1, 0, 0, 1, 0, 0, 1, -1, -1, 0, -1, 0, 1, 2, 3, 2, 1, 0, 1, 0, 0, 0, -1, -2, -1, -2, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 2, 2, 2, 2, 0, 1, 0, 0, -1, -1, -1, 0, -2, 0, -1, 0, 1, 0, 0, -2, -1, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, -1, -2, -2, -2, 0, -1, 0, 0, 0, 0, -1, 0, -2, -1, -2, 0, -2, -1, -1, 0, 0, 1, 0, 0, 0, 2, 1, -1, -2, -1, -1, 0, 0, 0, 0, 0, -1, -1, -3, -1, -1, -2, -2, 0, -1, 0, 0, 0, 0, 2, 2, 1, 0, 0, -1, -1, -2, 0, 0, 2, 0, 0, -1, -1, -1, -3, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 2, 0, -1, -1, -1, -1, 0, 1, 2, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, -1, -2, 0, 0, 2, 1, 0, 0, -1, 0, -2, -1, -1, -2, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 3, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, -1, -1, -2, -1, -2, -2, -1, -1, 0, 1, 2, 2, 0, 0, 0, 0, -1, -3, -2, -2, -2, -2, -2, 0, -2, -1, -3, -3, -2, -3, -2, 0, -2, 0, 0, 1, 0, 2, 0, 0, 1, -1, -1, -3, -2, -1, -1, -3, -1, -2, -2, -3, -4, -3, -2, -1, -2, -1, 0, -1, 0, 0, 1, 3, 0, 0, 1, 0, -2, 0, -1, -1, 0, -1, -3, -2, -2, -4, -3, -3, -2, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 1, 0, 0, 0, -1, 0, 0, -2, -2, -2, -1, -2, -2, -1, -1, 0, -1, 0, 0, 0, 0, 1, 3, 3, 2, 1, 1, 0, 0, 0, 0, -1, 0, 0, -2, -3, -1, -2, -2, -1, -2, 0, 1, 0, 0, 0, 1, 1, 3, 6, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 1, 0, 0, 1, 0, 2, 4, 5, 1, 2, 0, 0, 1, 0, 1, 1, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 4, 4, 7, 2, 1, 1, 2, 2, 2, 2, 3, 3, 3, 4, 5, 4, 2, 1, 0, 2, 0, 1, 2, 4, 4, 4, 6, 6, 7, 6, 3, 2, 1, 1, 0, 0, -1, -2, -2, -5, -7, -6, -6, -5, -3, -1, 0, 0, -1, -1, 0, 1, 1, 1, 0, 3, 3, 1, 1, 0, 1, 0, 0, -1, -2, -4, -4, -5, -3, -2, -2, -1, 0, 0, 0, 0, 1, 1, 0, 2, 1, 3, 2, 1, 1, 1, 0, -1, -1, -1, -3, -3, -2, -3, -2, -2, -2, 0, 1, 1, 0, 0, 1, 0, 1, 1, 1, 1, 2, 0, 0, 0, 0, 0, -1, 0, -2, -2, -3, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, -1, -2, 1, 1, 2, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -4, 1, 0, 1, 0, 0, 0, 1, 2, 2, 4, 2, 2, 1, 3, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -3, 1, 0, 0, 0, 0, 1, 0, 2, 3, 5, 2, 3, 1, 2, 3, 0, 0, -1, -1, 0, -1, 0, -1, -2, -3, -5, 0, 0, 0, 0, 1, 1, 3, 4, 4, 4, 5, 3, 2, 4, 3, 2, 0, -1, 0, -1, -1, -2, -1, -3, -3, -5, 0, 0, 0, 0, 1, 3, 5, 4, 4, 5, 4, 5, 5, 6, 5, 4, 2, 1, -1, 0, -2, -1, -1, -2, -3, -3, 0, 0, 0, 2, 1, 3, 5, 3, 4, 4, 6, 5, 5, 5, 7, 6, 3, 2, 0, 0, -1, -3, -2, -1, -2, -4, 0, 0, 0, 2, 2, 3, 5, 4, 5, 5, 5, 5, 7, 7, 5, 5, 4, 1, 0, 0, 0, -2, -1, 0, -2, -1, 0, 0, 0, 0, 2, 4, 3, 6, 6, 7, 6, 5, 5, 6, 6, 5, 4, 1, 0, -2, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 2, 4, 6, 4, 4, 5, 7, 7, 7, 7, 7, 6, 3, 0, -2, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 2, 2, 4, 4, 5, 5, 7, 6, 6, 7, 8, 7, 5, 3, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 1, 1, 3, 3, 5, 3, 6, 5, 5, 7, 7, 7, 6, 4, 3, 1, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 1, 0, 2, 4, 5, 4, 4, 4, 4, 4, 5, 4, 4, 2, 2, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 1, 0, 0, 1, 2, 4, 5, 2, 3, 4, 3, 2, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, -1, 0, -2, 0, 0, -1, 0, 0, 0, 3, 3, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, 0, 0, -1, -2, 0, 2, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -2, 1, 0, -2, 0, 1, 1, 1, 1, 0, 0, -1, 0, -1, -1, -1, -1, 1, 1, 1, 0, 1, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -3, 0, -1, -3, -2, -2, -2, 0, 1, 1, 0, 0, 0, 1, 0, 2, 0, 0, 2, 0, 0, 0, 0, 0, -1, -2, -3, -1, -2, -3, -3, -2, -1, 0, 0, 0, 0, 1, 2, 1, 2, 3, 0, 0, 1, 1, 0, 1, 1, 0, -2, -2, -3, -1, -3, -4, -3, -2, -1, 0, 1, 0, 0, 0, 0, 3, 3, 1, 1, 1, 1, 1, 1, 0, 3, 2, 0, 0, -3, -2, -2, -5, -4, -4, -1, 0, -1, 0, 0, 1, 2, 1, 2, 2, 2, 0, 3, 1, 1, 2, 3, 3, 0, 0, -2, -2, -4, -5, -4, -3, -3, -2, -1, 0, 0, 2, 2, 3, 2, 2, 1, 1, -5, -5, -4, -2, -1, -2, -3, -3, -2, -1, -3, -1, -2, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -5, -3, -3, -2, -1, -1, -1, -2, -2, -2, -1, -2, -1, -2, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -5, -4, -2, -1, 0, -1, 0, -2, -1, -2, -1, -2, 0, -2, -2, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -4, -4, -3, -1, -1, -1, 0, 0, -2, -1, -1, -2, -2, -2, -2, -2, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, -4, -2, -2, 0, -1, 0, 0, 0, -1, -1, -1, -2, -1, -2, -2, -1, 0, 0, -1, -2, 0, 0, 0, 0, 0, -2, -5, -2, -1, -2, 0, -1, -2, 0, -1, -1, -1, 0, -1, -1, -1, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, -4, -2, -2, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -1, 0, 0, 0, 0, -1, -2, -5, -4, -2, -1, -2, -2, -2, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -2, -2, -1, -1, 0, 0, 0, 0, -2, -5, -2, -2, -1, -1, -2, -2, -1, -1, 0, 0, 1, 1, 0, 0, 0, -1, 0, -2, -2, 0, -1, -1, 0, 0, 0, -4, -3, -2, -1, 0, -1, -1, -2, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, -1, 0, -3, -3, -1, -2, 0, -1, -2, 0, -1, -1, 0, 0, 0, 1, 0, 0, -1, 0, -1, -3, -2, -2, -1, 0, 0, -2, -3, -3, -1, -1, -2, -2, -1, -2, -2, 0, 0, 0, 1, 0, 1, 0, 1, 0, -1, -1, -3, -2, -1, -2, -2, -2, -4, -1, -1, -1, -1, -3, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -2, -1, -2, -1, -2, -3, -2, -3, -1, -1, -1, -1, -3, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -3, -2, -1, 0, -2, -2, -2, 0, -1, -2, -1, -1, -1, -2, -1, 0, 0, 0, 0, 1, 0, 1, 0, -1, -1, -1, -1, -3, -2, -1, -2, -4, -1, -1, -1, -2, -3, -2, -2, -1, -2, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, -2, -2, -1, -4, -2, 0, -2, -1, -3, -2, -1, -2, -2, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -2, -1, -1, -1, -1, -2, -4, -1, -2, -1, -2, -1, -1, -3, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -2, 0, -1, -1, -4, -1, -1, -1, -2, -2, -2, -1, -2, -2, 0, -1, -2, -1, -2, 0, -1, 0, 0, 0, -2, -3, -2, 0, 0, -2, -4, -3, 0, -2, -2, -3, -2, -2, -1, -1, -1, -1, 0, -2, -1, -1, -1, -1, 0, -1, 0, -2, 0, -2, -1, -1, -4, -1, -2, -2, 0, -2, -2, -1, 0, -2, -2, -1, -3, -1, -1, -1, 0, 0, 0, -1, 0, 0, -2, 0, -1, -1, -4, -3, -2, 0, -1, 0, -2, -2, -3, -1, -2, -2, -2, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, -3, -1, 0, -1, 0, 0, -2, -2, -2, -1, -1, -3, -3, -1, -3, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, -5, -3, -2, 0, -2, 0, 0, 0, -2, -1, -2, -2, -2, -1, -2, -1, -2, 0, -1, 0, 0, -1, 0, 1, 1, 1, -6, -2, -1, -1, -2, -1, -1, 0, -2, -1, -2, -1, -2, -2, -1, -3, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, -6, -3, -1, -2, -1, -2, -2, -2, 0, -1, -2, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 1, 0, 0, 2,
    -- filter=0 channel=7
    3, 2, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 2, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 2, 2, 0, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, -2, 0, -1, -1, 0, 0, -1, 0, 0, 3, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -2, -1, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, 1, 2, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, 0, -1, 0, 0, 0, 0, -1, 0, -1, 2, 2, 0, 0, 0, 1, 0, 1, 0, 0, -1, -1, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 3, 3, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -2, 0, 2, 2, 1, 1, 1, 1, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, -1, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, -1, -1, -1, 3, 0, 0, 0, 0, 2, 1, 1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -2, 0, 3, 0, 0, 0, 1, 1, 0, 1, 0, -2, -3, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, -1, 0, -2, -1, 0, 0, -1, 0, 1, 0, 0, 0, 1, 1, 1, 1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, 2, 0, 0, 0, 0, 1, 1, 0, -1, -2, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 2, 2, 1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, 0, 2, 1, 1, 0, 1, 1, 0, 0, -1, -1, -2, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 1, 0, 0, 2, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 2, 0, 2, 1, 1, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, -1, -1, 2, 1, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -2, -1, 0, -1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 3, 1, 0, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, 3, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, -1, 2, 2, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 2, 2, 1, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 3, 2, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 4, 2, 1, 0, -2, 0, -1, -1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, -1, -3, -1, -3, -2, 2, 0, 0, 0, -1, -2, -2, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, -1, 0, -2, -3, 2, 0, 0, -1, -1, -2, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 2, 1, 0, -1, -1, -1, 0, 0, 0, 2, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 3, 0, -1, -2, -1, -1, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, -1, 2, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, -1, 3, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 3, 3, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, -1, 4, 2, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 2, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 1, 1, 2, 0, 0, 1, -1, -1, -1, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 0, 0, -1, 0, 0, 0, 0, 0, 2, 2, 0, 1, -1, -1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 3, 1, 0, 0, 0, 0, 2, -1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 1, 0, 0, 1, 2, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, 0, -1, -1, -1, -1, 1, 0, 2, 0, 1, 0, 0, 0, 3, 0, 1, 1, 2, 0, 0, 0, 0, 2, 2, 1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 3, 1, 1, 2, 1, 0, 1, 1, 2, 1, 0, 2, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, -1, 0, 3, 1, 1, 0, 0, 0, 0, 0, 0, 2, 1, 2, 0, 1, 0, 1, 0, 1, 1, 1, 2, 1, 0, 1, -1, 0, 4, 2, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 1, 0, 2, 2, 0, 1, 1, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 1, 1, 0, 0, 1, 1, 2, 2, 1, 0, 1, 0, 1, 0, 3, 0, 1, 0, 0, -1, 0, -1, 1, 0, 2, 1, 0, 0, 1, 1, 1, 2, 2, 2, 2, 1, 1, 1, 0, 0, 3, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 0, 1, 2, 1, 0, 0, 0, -1, 2, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 2, 1, 0, -1, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -2, -2, -3, 3, 2, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, -2, -1, -2, -3, -4, 0, 1, 2, 2, 1, 1, 2, 1, 2, 3, 2, 4, 3, 4, 2, 2, 2, 4, 2, 2, 2, 3, 2, 3, 4, 6, 0, 1, 3, 2, 1, 1, 2, 2, 0, 1, 0, 0, 3, 2, 1, 1, 1, 1, 1, 1, 1, 2, 2, 1, 3, 4, 0, 1, 3, 2, 1, 1, 1, 0, 0, -1, 0, 0, 0, 2, 1, 3, 2, 2, 0, 0, 0, 1, 1, 0, 0, 2, 0, 1, 3, 3, 1, 1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 1, 3, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 3, 2, 0, 2, 1, 0, 0, -1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 2, 1, 1, 0, 1, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 2, 2, 1, 0, 0, 0, -1, -2, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 2, 1, 1, 0, -1, -2, -3, -4, -3, -1, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 2, 2, 0, 1, 1, 0, -1, -1, -4, -3, -3, -3, -2, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, -1, 2, 3, 2, 2, 1, 0, -1, 0, -1, -4, -3, -3, -2, -2, 0, 0, 2, 2, 2, 0, 0, 0, 0, 0, 2, 0, 2, 2, 2, 1, 0, 0, 0, 0, -1, -3, -5, -3, -2, 0, 0, 1, 2, 3, 0, 0, 0, 0, -1, 0, 2, 0, 2, 2, 3, 0, 0, 0, 0, -2, -2, -2, -4, -4, -1, -1, 0, 1, 4, 1, 0, 0, 0, 0, 1, 0, 3, 0, 3, 2, 1, 0, 0, -1, -1, -2, -3, -3, -5, -3, -3, -1, 0, 2, 3, 3, 2, 0, 0, 1, 0, 2, 2, 0, 1, 2, 0, 0, 0, 0, -2, -3, -3, -3, -5, -4, -3, -3, 0, 2, 3, 4, 2, 1, 0, 0, 1, 1, 3, 0, 2, 2, 2, 0, 0, -2, -2, -1, -3, -5, -6, -6, -3, -3, 0, 2, 4, 3, 3, 0, 1, 1, 1, 0, 3, 0, 1, 0, 0, 1, 0, 0, -2, -2, -3, -3, -3, -4, -3, -3, -1, 2, 2, 2, 2, 1, 0, 1, 2, 1, 3, -1, 1, 2, 0, 1, 0, 0, 0, -2, -3, -4, -4, -2, -3, -2, 0, 1, 2, 2, 1, 2, 1, 1, 0, 1, 3, 0, 1, 0, 0, 0, 1, 0, -1, -2, -2, -3, -2, -4, -3, -2, -1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 3, 0, 0, 1, 1, 1, 0, 0, 0, -2, -1, -3, -3, -2, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 2, 1, 0, 0, 0, -2, 0, -1, -2, -2, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 1, 2, 0, 0, 1, 2, 1, 0, 0, 0, -2, 0, -1, 0, -1, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 2, 2, 2, 1, 0, -1, 0, 0, 0, -2, -1, 0, 0, 0, 0, -2, 0, -1, 0, 0, 1, 0, 1, 2, 0, 1, 2, 1, 1, 1, 0, 0, 0, -1, 0, -2, 0, 0, 0, -1, 0, -1, 0, 1, 1, 0, 2, 2, 1, 3, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 2, 1, 1, 3, 1, 4, -1, 1, 2, 2, 3, 2, 1, 1, 1, 0, 2, 1, 1, 1, 1, 0, 1, 0, 1, 1, 1, 3, 4, 3, 4, 4, -1, 2, 2, 4, 3, 3, 1, 1, 3, 4, 4, 4, 4, 2, 2, 3, 0, 1, 2, 2, 2, 5, 3, 4, 4, 6, 0, -1, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, -2, 0, 0, 1, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 2, 2, 2, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 1, 2, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 1, 1, 1, 1, 2, 1, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 2, 2, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 3, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 2, 1, 2, 2, 3, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 1, 2, 1, 2, 2, 3, 3, 2, 2, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 1, 1, 3, 1, 3, 3, 1, 1, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 1, 0, 2, 3, 2, 2, 3, 2, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 2, 2, 2, 2, 2, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, -1, -1, 0, 1, 0, 2, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 1, -1, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 2, 1, 1, 0, 1, 0, 2, 1, 1, 2, 0, 1, 1, 0, 0, 0, -2, 0, -1, 0, -1, 0, 0, 2, 1, 1, 1, 1, 1, 1, 2, 1, 2, 1, 0, 0, 1, 0, 0, 0, -1, -1, -2, 0, 0, 0, 1, 2, 1, 1, 2, 2, 2, 2, 2, 2, 2, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 1, 2, 1, 2, 2, 2, 3, 3, 3, 3, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 2, 1, 2, 2, 1, 2, 2, 2, 1, 1, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 3, 1, 2, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 3, 2, 1, 2, 1, 2, 1, 1, 0, 1, 2, 0, 0, 1, 1, 0, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 1, 2, 0, 0, 3, 0, 1, 1, 0, 2, 0, 1, 0, 0, 0, 1, 1, 0, 0, 2, 1, 1, 2, 2, 1, 1, 2, 2, 1, 0, 1, 2, 0, 0, 2, 1, 2, 0, 0, -1, -1, 0, -1, -1, 0, 1, 1, 3, 2, 2, 1, 3, 0, 2, 1, 0, 2, 0, 1, 2, 2, 1, 2, 0, -1, -1, 0, -2, -1, -2, 0, 1, 2, 2, 1, 3, 3, 3, 2, 1, 2, 0, 0, 0, 0, 2, 2, 3, 0, 2, 0, 0, 0, -2, -1, -2, 0, 0, 0, 0, 0, 2, 1, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 3, 3, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 2, 2, 0, 1, 0, 1, 0, 1, 1, 2, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 1, 0, 0, 2, 1, 2, 2, 1, 1, 3, 2, 1, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 1, 1, 1, 1, 2, 2, 1, 4, 3, 1, 2, 3, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 2, 0, 2, 1, 1, 1, 2, 3, 3, 3, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 3, 0, 1, 2, 2, 0, 1, 0, 1, 2, 1, 2, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 2, 1, 1, 0, 0, 0, 2, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 2, 0, 1, 2, 1, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -2, -2, -2, -4, -3, -1, 0, -1, 0, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 2, 2, 1, 3, -3, -2, -2, 0, 0, -1, 0, -2, -1, -2, -1, -1, -1, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 2, 2, 4, -5, -3, -1, 0, 0, 0, -1, -1, -2, -2, -2, -2, -2, -1, -1, 0, -2, 0, 0, 0, 0, 0, 0, 1, 3, 2, -3, -1, 0, 0, 0, -1, 0, -1, -2, -3, -4, -3, -2, -2, -3, -2, -2, 0, 0, -1, -1, -1, 0, 1, 1, 2, -3, -2, 0, 0, 0, 0, 1, 0, -2, -3, -3, -2, -3, -3, -1, -1, -1, 0, 0, 0, 0, -2, -1, 1, 1, 2, -2, -1, 0, 0, 0, 0, 1, 0, -1, 0, -3, -1, -3, -2, -2, -2, -2, -1, 0, -2, 0, 0, -1, 1, 0, 2, -3, -2, -1, 1, 0, 0, 2, 2, 0, 0, 0, -2, -2, -1, -1, -3, -2, -2, -2, -2, -1, 0, -2, 0, 0, 2, -5, -3, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, -1, -1, -2, -3, -3, -2, -3, -2, 0, 0, -1, 0, 0, 0, -4, -3, -1, 0, 0, 1, 0, 2, 2, 0, 1, -1, -2, -1, -3, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, -2, -3, -2, 0, 0, 0, 0, 2, 0, 2, 0, 0, -1, 0, -1, -1, -1, -2, -1, -1, 0, 0, 0, -1, 0, 1, -3, -3, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 0, 1, 0, 0, -1, -2, 0, 0, 1, -1, 0, 0, 0, 1, -2, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, -3, 0, 0, 0, 0, -1, 1, 0, 0, 1, 2, 1, 1, 2, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -2, 0, -1, -1, 0, 0, 0, 0, 0, 1, 2, 2, 2, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 2, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 2, -1, -2, 0, 0, -1, 0, 0, 1, 0, 2, 2, 1, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, -2, -3, -2, 0, 0, 0, 0, 1, 0, 2, 1, 1, 1, 2, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 2, -3, -3, -2, -1, -1, 0, 0, 2, 1, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, -3, -3, -1, -1, 0, 0, 2, 3, 1, 3, 2, 1, 2, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -3, -2, -2, 0, 1, 0, 2, 2, 1, 3, 2, 2, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, -4, -3, 0, -1, 0, 2, 0, 2, 3, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 1, 0, 1, 2, -3, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 1, 1, 0, 3, -3, -3, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, -1, -1, -2, -2, 0, -1, 0, -1, 0, 2, 1, 3, -3, -2, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, -2, -2, -1, 0, -1, -1, 0, 0, 0, 0, 2, 1, 2, 3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 3, 2, 4, 4, -4, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 1, 1, 3, 3, 4, 5, 5, -5, -2, -2, 0, 0, 0, 0, 1, 2, 4, 6, 8, 10, 11, 10, 10, 9, 8, 5, 6, 4, 4, 6, 6, 7, 10, -6, -2, -2, -1, -1, -1, -1, 0, 0, 1, 2, 3, 6, 6, 7, 6, 4, 4, 2, 3, 3, 3, 4, 3, 4, 7, -6, -3, -3, -1, -2, -1, -1, 0, 0, 1, 0, 1, 1, 4, 3, 3, 3, 3, 1, 0, 0, 3, 3, 2, 3, 6, -6, -3, -3, -2, -1, -1, 0, 0, 0, -1, -1, 0, 1, 1, 1, 2, 2, 1, 1, 1, -1, 0, 1, 2, 1, 3, -5, -2, -1, -1, -2, -1, 0, -1, -2, -4, -1, -1, -1, 0, 0, 2, 2, 3, 2, 0, 0, -1, 0, 2, 3, 4, -5, -1, 0, -1, 0, -2, 0, -1, -3, -5, -3, -4, -1, 0, 0, 1, 3, 3, 3, 2, 0, 1, 2, 2, 3, 3, -4, -1, 0, 2, 1, 0, 0, -3, -3, -4, -4, -3, -2, -2, -1, 1, 1, 3, 3, 2, 1, 0, 2, 2, 3, 4, -5, -2, 1, 1, 2, 0, 0, 0, -2, -3, -6, -4, -6, -5, -2, 0, 0, 0, 2, 1, 0, 0, 1, 0, 0, 2, -5, -1, 0, 2, 1, 0, 2, 1, 0, -2, -3, -5, -6, -8, -4, -3, 0, 1, 4, 2, 1, 0, 0, 1, 1, 2, -5, -2, 1, 2, 1, 1, 1, 0, 0, 0, -2, -5, -7, -8, -7, -4, 0, 3, 3, 4, 1, 1, 1, 1, 0, 3, -5, -3, 0, 1, 2, 0, 0, 0, 1, 0, -3, -6, -8, -8, -4, -2, 1, 4, 8, 5, 3, 2, 1, 1, 1, 2, -4, -2, 0, 1, 0, 0, -1, -3, -2, -2, -2, -4, -6, -5, -3, -2, 4, 7, 10, 9, 5, 3, 2, 1, 0, 2, -6, -3, 0, 1, 0, -1, -2, -3, -3, -1, -2, -5, -5, -4, -3, -1, 5, 10, 12, 11, 8, 5, 3, 2, 2, 2, -4, -3, 0, 0, -1, -2, -3, -4, -4, -3, -5, -4, -7, -5, -4, 0, 4, 9, 13, 13, 9, 6, 3, 1, 0, 2, -4, -1, 0, 0, -1, -2, -3, -3, -2, -2, -5, -6, -6, -8, -5, -2, 1, 6, 10, 9, 7, 5, 3, 1, 1, 1, -5, -1, 0, -1, 0, -1, -3, -3, -3, -3, -3, -5, -6, -7, -8, -3, 0, 3, 6, 7, 6, 3, 2, 1, 1, 1, -3, -2, -1, -1, -2, -2, -2, -3, -1, -3, -4, -4, -4, -7, -7, -4, -1, 1, 4, 3, 2, 0, 0, 0, 2, 2, -3, -1, 0, 0, -1, 0, -1, -3, -3, -2, -2, -2, -3, -3, -4, -3, -1, 2, 4, 3, 1, 0, 0, 0, 0, 3, -4, -2, 0, -1, -1, 0, -1, -3, -2, -1, -1, 0, -2, -1, -1, 0, 0, 3, 4, 3, 3, 0, -1, 0, 1, 3, -6, -4, -2, 0, 0, 0, 0, -2, -2, -4, -2, 0, -1, 0, 0, 3, 1, 2, 3, 5, 3, 2, 0, 0, 0, 2, -5, -4, -2, -1, 0, 1, 1, 0, 0, -3, -1, -1, 0, 0, 2, 1, 1, 2, 4, 4, 3, 3, 3, 1, 1, 2, -4, -4, -1, -1, 0, 0, 0, 1, 2, 0, 0, 1, 0, 2, 2, 0, 0, 1, 0, 2, 2, 2, 2, 2, 1, 3, -4, -4, -2, -2, 0, 0, 0, 2, 1, 1, 0, 1, 0, 0, 2, 1, 0, -1, -2, -1, -1, 0, 0, 1, 1, 4, -3, -2, -1, -1, 0, 0, 0, 2, 1, 0, 2, 1, 2, 1, 0, 0, -1, -1, -1, -1, -2, 0, 0, 2, 2, 5, -5, -2, -1, -1, -2, -1, 0, 1, 0, 2, 3, 2, 3, 3, 2, 1, 1, 0, 0, -1, -1, -1, 0, 1, 3, 5, -2, 0, 0, 0, 1, 0, 0, 0, 1, 4, 5, 5, 6, 7, 6, 5, 4, 3, 1, 0, 0, 1, 3, 5, 4, 7, 5, 4, 1, 0, -1, -4, -4, -4, -3, -1, 0, 1, 2, 2, 2, 0, -1, -1, -2, -3, -3, -2, -3, -4, -4, -5, 5, 0, 1, -1, 0, -2, -2, -1, 0, 0, 0, 1, 1, 1, 1, 0, -1, -2, -2, -2, -2, -3, -3, -2, -4, -3, 4, 2, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 2, 3, 2, 0, 0, 0, -1, -1, -1, -2, -1, -1, -2, -3, 3, 1, 0, 0, 0, -2, -2, 0, 0, 2, 1, 3, 2, 1, 2, 1, 0, 0, 0, -1, 0, -1, 0, -1, -1, -2, 4, 2, 0, 0, 0, -1, -1, 0, 0, 0, 1, 2, 1, 3, 1, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, -1, 4, 2, 1, 0, 0, 0, 0, 0, 0, -1, 1, 1, 1, 2, 1, 2, 0, 0, -1, -1, 0, 0, 0, 0, 0, -2, 4, 2, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 5, 1, 2, 0, 0, 0, 0, 1, 2, 1, 3, 2, 2, 2, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 5, 2, 1, 1, 3, 2, 2, 1, 3, 4, 4, 4, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 1, 0, 2, 1, 0, 1, 3, 4, 6, 6, 5, 2, 0, -1, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 2, -1, 0, 0, 0, 0, 1, 1, 0, 2, 6, 5, 6, 4, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -2, -3, 0, 0, 0, -1, 0, -1, 2, 5, 6, 4, 4, 1, -1, -3, -2, 0, 1, 0, 0, -1, -1, 0, -1, -1, -5, -4, 0, 0, 0, 0, 0, 0, 3, 5, 4, 6, 2, 0, -1, -2, 0, 0, 0, 0, 0, 0, 1, 0, -2, 0, -5, -3, -1, 0, 0, -1, -1, 0, 2, 4, 4, 5, 2, 0, -1, -1, -1, -1, 1, 1, 1, 1, 1, 0, 0, 0, -3, -1, 0, 1, 0, 0, 0, 2, 4, 5, 5, 5, 2, 2, -1, -1, -3, -1, 0, 0, 0, 0, 0, -1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 2, 6, 5, 4, 1, 1, -1, -3, 0, 0, 1, 0, 0, 0, 0, 0, -2, 3, 1, 1, 0, 0, 0, 0, 0, 1, 3, 3, 4, 4, 1, 0, 0, -1, -1, 0, 2, 0, 0, 0, -1, 0, -1, 5, 1, 0, 1, 0, 0, 0, 1, 1, 3, 3, 4, 2, 1, 2, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 6, 1, 0, 1, 0, 0, 0, 2, 4, 4, 4, 3, 2, 1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 4, 1, 2, 1, 1, 1, 0, 2, 4, 2, 2, 2, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, -1, 5, 1, 1, 2, 1, 0, 1, 1, 1, 1, 2, 1, 0, 0, 1, 0, 0, 1, 1, 2, 0, 0, 0, 1, 0, -2, 4, 1, 0, 0, 1, 2, 1, 1, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, -3, 4, 0, 0, 1, 1, 0, 0, 1, 0, 2, 1, 3, 3, 2, 2, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -3, 4, 0, -1, 0, 1, 1, 0, 0, 0, 2, 3, 3, 4, 4, 1, 2, 1, 0, 0, 0, -1, -2, -2, -1, -1, -3, 4, 0, 0, 0, 1, 0, 0, -2, 0, 1, 2, 3, 4, 3, 2, 2, 2, 0, 0, -1, 0, -3, -2, -1, -3, -3, 7, 1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 2, 4, 2, 3, 2, 0, 1, -1, 0, -2, -2, -3, -4, -4, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, -2, -1, -1, -1, -1, 0, -1, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 2, 0, 0, 0, 1, 0, 0, 0, 1, -2, -1, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, -2, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, -1, 1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 2, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 2, 2, 1, 2, 2, 1, 0, 0, 1, 0, 0, -1, -1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 2, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 2, 2, 0, 1, 2, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 9, 4, 0, -2, -4, -4, -4, -5, -2, -2, 2, 4, 3, 4, 5, 3, 1, 0, 0, -2, -3, -2, -3, -4, -3, -4, 6, 1, 0, -3, -3, -4, -3, -4, -2, 0, 1, 4, 4, 3, 3, 1, 0, 0, 0, -1, -2, -2, -1, -2, -2, -4, 4, 0, -1, -3, -2, -3, -3, -1, 0, 0, 1, 2, 3, 4, 3, 2, 1, 0, -1, 0, 0, -1, -2, 0, 0, -3, 5, 1, -1, -2, -3, -2, -1, 0, 0, 0, 1, 2, 3, 4, 3, 3, 0, 0, 1, 0, 0, -1, -1, -1, -1, -1, 5, 0, 0, 0, -3, -2, -3, 0, 0, 1, 2, 2, 3, 3, 2, 3, 2, 1, 2, 2, 0, 0, 0, 0, 0, -1, 5, 2, 0, 0, -2, -1, -2, -2, -1, -1, 1, 1, 1, 3, 1, 2, 3, 2, 1, 2, 1, 0, 0, 0, 1, 0, 7, 1, 1, 0, 0, -2, -3, -1, -2, 0, 0, 0, 1, 1, 2, 1, 3, 2, 1, 1, 2, 2, 2, 1, 2, 1, 8, 4, 2, 0, 1, -1, 0, 0, 0, 2, 1, 3, 1, 0, 0, 0, 0, 1, 2, 2, 2, 2, 1, 1, 0, 0, 5, 2, 0, 1, 0, 0, 0, 2, 3, 3, 4, 2, 2, 0, -1, -2, -1, 0, 3, 3, 1, 2, 1, 1, 0, 0, 6, 2, 0, 1, 0, 1, 2, 2, 2, 4, 5, 4, 2, 0, -2, -2, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 4, 0, 0, 1, 0, 1, 0, 0, 1, 5, 6, 6, 5, 0, -2, -2, -3, 0, 0, 3, 1, 0, 0, -1, -1, 0, 0, -1, -1, 0, 1, 2, 1, 0, 0, 3, 5, 5, 3, 1, -2, -3, -2, 0, 3, 3, 3, 1, 0, 0, -1, -1, 0, -3, -4, -1, 1, 0, -1, 0, 0, 2, 3, 3, 2, 0, -2, -3, -2, 0, 4, 5, 4, 4, 2, 0, 0, -2, 0, -5, -4, -1, 1, 1, 0, 0, 1, 3, 3, 4, 1, 0, -2, -2, -3, 0, 2, 5, 5, 2, 2, 1, 0, -1, 1, -3, -2, 0, 0, 2, 0, 1, 2, 3, 5, 5, 2, 0, -1, -4, -2, -1, 1, 3, 3, 1, 1, 0, 0, 0, 1, -2, 0, 0, 3, 1, 3, 1, 2, 5, 5, 3, 3, 0, -1, -3, -3, 0, 0, 2, 2, 2, 1, 0, -1, -1, 2, 1, 0, 0, 1, 1, 0, 0, 3, 4, 3, 4, 3, 0, -2, -1, -2, 1, 3, 2, 2, 1, 1, 0, 0, -2, 6, 1, 0, 0, 1, 1, 0, 0, 1, 3, 3, 1, 2, 0, 0, 0, 0, 0, 3, 3, 1, 2, 0, 0, -1, -1, 6, 1, 0, 0, 0, 0, 0, 0, 1, 2, 3, 1, 1, 0, 1, 0, 1, 1, 2, 2, 2, 3, 1, 0, 0, -1, 5, 1, 0, 0, 0, 1, 1, 2, 2, 1, 1, 0, 0, 0, 0, 1, 2, 2, 4, 4, 4, 3, 4, 3, 0, 0, 6, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 3, 4, 4, 4, 3, 1, 1, 0, 4, 1, 0, -1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 1, 0, 0, 1, 1, 2, 2, 1, 3, 2, 2, 0, -1, 5, 0, 0, 0, -1, 0, -2, -1, 0, 1, 2, 3, 3, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, -2, -1, 5, 0, 0, 0, -1, -2, -2, -1, 0, 1, 3, 3, 4, 2, 3, 2, 2, 1, 0, 0, 0, -1, -2, 0, -3, -4, 7, 1, 0, 0, 0, -1, -2, 0, 0, 1, 3, 4, 5, 4, 4, 4, 2, 1, 0, 0, -1, -3, -4, -2, -2, -4, 8, 4, 1, 1, 0, 0, 0, -2, 0, 0, 2, 4, 4, 5, 6, 3, 4, 3, 0, 0, 0, -3, -2, -3, -3, -6, -1, -2, 0, -1, 0, 0, 0, -1, -1, -1, 1, 1, 1, 2, 2, 1, 2, 2, 0, 0, 1, 0, 0, 0, 1, 0, -2, -1, -1, 0, 0, -1, -1, -1, 0, -1, 1, 2, 1, 2, 2, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 2, 2, 2, 1, 0, -1, -1, -1, 0, -1, -1, -2, -1, 0, 0, -2, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, -1, -1, -2, -1, 0, -3, -2, -1, 0, 0, -2, 0, 0, 1, 0, 1, 0, 0, 0, 0, 2, 0, 1, 1, 0, 0, -1, -2, -2, -3, -2, -2, -2, -1, 0, 0, -3, 0, 0, 0, 1, 2, 2, 0, 3, 2, 2, 1, 1, 0, 1, -1, 0, -3, -3, -3, -3, -3, -1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 2, 1, 1, 2, 2, 0, 1, 0, 1, 0, 0, -1, 0, -1, -1, -3, -1, 0, 0, 0, -2, -1, 0, 0, 0, 1, 2, 3, 3, 3, 3, 1, 0, 2, 0, 1, 1, -1, -1, -2, -2, -1, 0, -2, -1, -1, -2, -1, 0, 0, 0, 0, 1, 1, 2, 4, 3, 2, 2, 1, 2, 0, 0, -1, -2, -1, -1, -3, -2, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 2, 2, 3, 2, 2, 3, 2, 1, 0, 0, -1, -3, -1, -3, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 3, 2, 2, 2, 2, 0, 0, 0, -2, -3, -2, -3, -2, -2, -2, -1, -1, -2, -1, 0, 0, 0, 0, 1, 1, 4, 3, 4, 3, 3, 3, 0, 0, 0, -2, -3, -4, -4, -2, 0, 0, -2, -2, -2, 0, -1, 1, 1, 0, 1, 3, 4, 3, 4, 3, 2, 3, 2, 2, 0, -1, -2, -2, -3, -3, -2, -2, 0, -1, -1, 0, 0, 0, 0, 2, 1, 3, 1, 2, 3, 3, 2, 1, 0, 0, 0, 0, -2, -4, -4, -1, -2, -1, -1, 0, -1, -2, -1, 0, 0, 0, 0, 3, 3, 2, 3, 1, 0, 0, 1, 1, 0, 0, -2, -2, -3, -1, 0, 0, 0, -1, -3, 0, 0, 0, 0, 1, 2, 2, 2, 1, 2, 0, 2, 1, 0, 0, 0, 0, -3, -4, -2, -1, 0, 0, 0, 0, -3, -3, -1, 1, 0, 0, 2, 3, 2, 2, 0, 0, 0, 1, 0, 0, 0, -2, -1, -3, -3, -2, 0, -2, 0, 0, -2, -1, 0, 0, 0, 1, 2, 3, 2, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, -3, -2, -2, -1, 0, 0, -3, -3, -1, 0, 1, 1, 3, 3, 1, 2, 0, 0, 0, -1, -2, -1, -2, -1, -2, -3, -3, -1, -1, 0, -1, -1, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -2, -2, -3, -1, -2, -3, -1, -2, -2, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -1, 0, -2, -2, -1, -1, 0, -1, -1, -3, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -2, 0, 0, 0, -1, -1, -2, -1, -1, 0, -1, -2, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, -2, -2, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -2, -3, -1, -1, -2, -1, -2, -2, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 1, 1, 0, 0, 0, -1, -1, -1, -2, -2, -2, -1, -2, -1, -1, -1, -2, -2, -2, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 3, 2, 0, 0, -2, -2, -3, -1, 0, 1, 1, 0, 3, 2, 3, 4, 2, 2, 0, 0, 0, -2, -1, -3, -2, -2, 3, 0, 0, -1, -2, -2, -1, 0, 0, 1, 2, 0, 2, 2, 1, 2, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 2, 0, -1, -2, -2, -2, 0, -1, 0, 0, 1, 2, 1, 0, 2, 0, 2, 1, 1, 0, 0, -1, 0, -2, -1, 0, 3, 0, -2, -2, -2, -2, -3, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, 3, 0, -1, -1, -1, -1, -3, -3, -1, -1, -1, 0, 0, 0, 1, 2, 3, 2, 1, 3, 1, 1, 1, 1, 0, -1, 3, 2, 0, -1, 0, -1, -1, -3, -2, -2, -1, 0, -1, -1, 1, 0, 1, 2, 2, 2, 3, 2, 2, 1, 0, 0, 6, 1, 1, -1, -1, -2, -2, -3, -3, -2, -3, 0, -1, 0, 0, 1, 0, 1, 2, 2, 2, 3, 1, 2, 0, 0, 5, 2, 1, 0, 0, 0, 0, -2, -1, 0, 0, -1, -1, -2, -3, -2, -1, 0, 1, 2, 1, 2, 1, 0, 1, 0, 4, 2, 0, 0, 1, 0, -1, -1, 0, 0, -1, 0, -3, -3, -3, -2, -1, 0, 0, 1, 2, 1, 1, 0, 0, -1, 4, 1, 1, 0, 1, 1, -1, -1, -1, 0, -1, 0, -4, -3, -5, -4, -2, -1, 2, 2, 3, 2, 1, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -1, -3, -5, -5, -4, -1, 1, 4, 5, 5, 4, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, -1, -3, -1, -2, -3, -4, -3, -2, 0, 2, 5, 6, 6, 6, 3, 1, 1, 0, 0, -2, -2, -2, -1, -1, 0, -1, -2, -3, -1, -2, -2, -2, -2, -1, 0, 2, 5, 7, 7, 5, 3, 2, 0, 0, 0, -1, -1, -1, 0, 0, 0, -2, -1, -1, -2, -2, -2, -3, -5, -3, 0, 1, 4, 5, 6, 4, 4, 1, 1, -1, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -4, -5, -3, 0, 1, 4, 5, 5, 4, 1, 1, 0, 0, 3, 2, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, -3, -5, -3, -3, 0, 1, 3, 3, 3, 2, 2, 2, 0, -1, 3, 2, 0, -1, -1, 0, 0, 0, -2, -1, 0, 0, -3, -4, -2, -2, -1, 0, 1, 4, 4, 2, 1, 2, 0, 0, 3, 1, 0, -1, 0, 0, -2, -2, -3, -2, -2, -1, -1, -2, -3, -2, -1, 0, 1, 3, 3, 3, 2, 1, 1, 0, 2, 0, 0, -2, -1, -2, 0, -1, -2, -4, -2, -3, -1, -3, -1, 0, 2, 1, 4, 5, 4, 4, 3, 1, 2, 0, 3, 1, 0, -1, 0, 0, -1, -1, -3, -2, -3, -2, -3, -1, -1, 0, 2, 2, 5, 5, 4, 3, 3, 2, 1, 0, 2, -1, 0, -2, -3, -3, -1, -3, -2, -1, -2, -1, -1, -2, -1, 0, 1, 3, 2, 2, 4, 2, 2, 1, 1, 1, 1, 0, -1, -2, -2, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 2, 1, 1, 2, 0, 0, 0, 4, 0, -1, -2, -1, -2, -2, -2, -1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 5, 1, 0, 0, -2, -1, -2, 0, 0, 1, 1, 2, 1, 3, 1, 1, 1, 2, 0, 0, 1, -1, 0, -1, -1, 0, 6, 2, 0, 0, 0, 0, -1, -1, 0, 1, 2, 2, 4, 2, 3, 3, 2, 3, 3, 1, 0, -1, 0, -1, -1, -2, 7, 3, 3, 1, 2, 1, 0, 0, 0, 1, 4, 4, 5, 5, 4, 4, 4, 4, 3, 2, 1, 0, 0, 0, 0, 0, 4, 4, 2, 0, 0, -1, -1, 0, 1, 0, 3, 2, 3, 4, 5, 4, 4, 3, 2, 1, 0, 0, 0, -1, 0, 0, 5, 3, 0, 0, -1, -1, -2, -2, 0, 0, 0, 3, 1, 2, 2, 1, 0, 1, 0, 0, 0, 0, 0, -2, 0, -1, 4, 1, 0, -2, -2, -3, 0, -1, -1, 1, 0, 0, 2, 1, 2, 2, 1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 5, 1, -1, -2, -1, -2, -2, -2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 0, 0, -2, -3, -3, -2, -2, -1, -2, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 4, 2, 1, 0, 0, 0, -2, -2, -3, -2, -3, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 1, 4, 3, 0, 1, 0, -1, -1, -2, -3, -4, -4, -3, -3, -1, 0, 0, 0, 1, 1, 1, 0, 2, 2, 1, 1, 2, 7, 3, 2, 0, 0, 0, -1, -1, -3, -2, -3, -2, -2, -2, -2, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 7, 4, 0, 0, 0, 0, 0, -2, -1, -3, -3, -3, -2, -2, -3, -4, -1, 0, 0, 0, 2, 1, 0, 1, 0, 1, 4, 2, 1, 0, 0, 0, 0, 0, 0, -2, -3, -1, -3, -4, -4, -4, -1, 0, 0, 0, 1, 2, 0, 0, 0, 0, 4, 0, 0, 0, 1, 1, 0, 0, -2, -3, 0, -1, -1, -3, -3, -3, -2, 0, 1, 2, 3, 1, 1, 1, 0, 0, 1, 0, -1, 0, -1, 0, -1, -2, -2, -1, -1, -2, -2, -2, -2, -3, -3, 0, 3, 4, 4, 3, 1, 1, 1, 1, 1, -1, -2, -2, 0, -1, -1, -3, -2, -2, -2, -1, -1, -3, -2, -3, -1, 2, 4, 4, 4, 4, 2, 0, 0, 0, 2, -1, -3, -2, -1, 0, 0, -1, -3, -1, -1, 0, 0, -3, -2, -3, 0, 1, 3, 5, 4, 3, 2, 0, 0, 1, 3, 0, -1, -2, -2, 0, -1, -3, -2, -1, -1, 0, -2, -2, -4, -2, -1, 2, 3, 5, 5, 4, 3, 1, 0, 1, 4, 2, 0, 0, 0, 0, -1, -2, -3, -1, -1, -1, -2, -2, -4, -3, 0, 0, 3, 2, 3, 3, 2, 1, 0, 0, 4, 2, 1, 0, -1, 0, 0, -1, -1, -1, -1, -2, -2, -4, -4, -4, 0, 0, 2, 1, 1, 3, 1, 1, 0, 0, 4, 2, 0, 0, -1, 0, 0, -1, -2, -1, -2, -3, -3, -3, -3, -3, -2, 0, 1, 1, 2, 2, 0, 0, 0, 1, 4, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -3, -2, -3, -3, -2, 0, 0, 2, 2, 3, 1, 1, 1, 2, 0, 4, 0, -1, 0, 0, -1, -1, 0, -1, -3, -2, -2, -3, -3, -1, -2, 0, 0, 1, 2, 1, 3, 1, 2, 2, 0, 4, 1, 0, 0, -1, 0, -1, -1, -1, -2, -1, -1, -3, -1, -1, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, 0, 5, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, 0, -1, -1, 0, 0, 0, 0, 1, 2, 0, 1, 0, 1, 0, 4, 2, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 5, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, -2, -1, 5, 3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 0, 0, 0, -1, 0, 0, -2, -3, -1, 0, 0, 8, 4, 2, 1, 1, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 1, 0, 0, 0, 0, -2, -3, -1, -2, 0, 5, 1, 0, -2, -2, -2, -1, -2, -2, 0, 0, 1, 1, 1, 0, 0, -1, 0, -1, -1, -3, -3, -5, -5, -5, -7, 2, 1, -1, -2, -2, -2, -1, 0, -1, -1, 0, 1, 1, 0, 0, -1, -1, -2, -2, -2, -2, -3, -3, -3, -3, -5, 3, 0, 0, -2, -2, -1, -1, 0, 1, 0, 0, 0, 1, 0, 0, -1, -1, -2, 0, 0, 0, -1, -1, -3, -3, -4, 2, 0, -1, -2, -2, -2, -1, 0, -1, -1, 0, -1, 0, 0, 1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -2, -3, 3, 1, -1, -1, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -2, -3, 4, 1, 0, -2, -1, -2, -1, 0, -1, -2, -1, -1, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, -1, 4, 1, 1, 0, 0, -2, -1, -1, 0, -1, -1, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 5, 2, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -2, 0, 1, 0, 0, 1, 0, -1, -1, -1, 4, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, -2, -2, 0, 2, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 3, 1, 0, -1, -1, -1, 0, 0, -1, 0, 0, -2, 0, 0, -2, 0, -1, -2, 0, 0, -1, 0, -1, 0, 0, 1, 1, 1, 0, -2, -3, -1, 0, 0, 1, 0, 0, 0, -1, -2, -2, 0, -3, -2, -1, -1, 0, -2, 0, 0, 0, 2, 2, 1, 0, 0, -1, -1, 0, 0, 0, 2, 0, 0, 0, -1, -1, -1, -3, -3, -1, 0, -1, -2, -2, 0, 2, 2, 2, 3, 0, 0, -2, -1, -1, 0, 1, 1, 1, 0, 0, 0, -3, 0, -4, -2, -2, 0, 0, 0, 0, 1, 3, 3, 3, 2, 0, -1, -1, -1, -2, 0, 1, 1, 2, 0, 0, 0, -2, 0, 0, -2, -1, 0, -1, -2, 0, 1, 3, 5, 4, 2, 0, -1, -1, -1, -1, 0, 0, 1, 1, 0, 0, 0, -3, 1, 0, 0, 0, -2, 0, -1, -1, 1, 4, 4, 2, 2, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, -1, 4, 1, -1, 0, 0, -3, -2, -1, 1, 1, 3, 2, 2, 1, -1, -1, -2, 0, 1, 1, 1, 0, 0, 0, -1, -2, 4, 0, 0, -1, -2, -1, 0, 0, 2, 1, 2, 0, 0, 0, 0, -2, 0, 0, 0, 1, 1, 2, 0, 0, 0, -2, 4, 0, 0, 0, -1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 2, 0, 1, 0, 0, -2, 4, 2, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, -2, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 5, 2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -3, 3, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, -1, -2, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -3, -3, -4, 3, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, -1, -2, -3, -2, -2, -3, -6, 6, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 1, 1, 1, 1, 0, 0, 0, -1, -3, -4, -3, -4, -5, 7, 2, 0, 0, 0, -1, 0, -2, -1, -1, 0, 0, 2, 1, 1, 2, 1, 2, 0, 0, -1, -3, -4, -4, -6, -7, 3, 1, 0, 0, -2, -1, -3, -2, -1, 0, 1, 2, 3, 4, 5, 3, 3, 2, 2, 2, 1, 1, 1, 1, 0, 2, 1, 0, -1, 0, -3, -2, -1, -1, 0, -1, 1, 1, 2, 2, 4, 3, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -2, -2, -3, -2, -1, 0, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, -2, -2, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -2, -2, -2, -2, -2, -1, -2, -2, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 3, 1, 0, -1, 0, -2, -1, -2, -3, -3, -1, -2, -1, -2, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 3, 2, 0, 0, 1, 1, -1, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 4, 0, 1, 0, 1, 2, 1, 1, 2, 1, 0, 0, -1, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 1, 1, 3, 2, 3, 2, 1, 0, -2, -4, -3, -3, -2, -2, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 2, 1, 3, 2, 0, 3, 2, 0, -1, -3, -6, -6, -5, -2, -1, 0, 0, -1, -2, -1, -2, -1, -1, -1, 0, 2, 2, 2, 1, 1, 2, 0, 2, 1, -1, -3, -5, -5, -4, -3, 0, 0, 0, 0, 0, -2, -2, -2, 0, -3, -1, 0, 0, 2, 1, 0, 0, 0, 2, 0, -1, -4, -4, -4, -4, 0, 1, 1, 1, 1, 0, -1, -2, -1, -1, -2, -1, 0, 0, 1, 0, 0, 2, 1, 0, 0, -2, -2, -4, -3, -3, -1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 1, 1, 1, 1, 2, 1, 0, -2, -5, -4, -2, 0, 1, 2, 2, 2, 1, 0, -1, 0, 1, -1, 0, 0, 0, 0, 3, 2, 2, 2, 1, 0, 0, -3, -4, -4, -4, -1, 0, 2, 2, 2, 0, 0, -1, -2, 2, 1, 0, 0, 0, 0, 2, 2, 2, 2, 2, 1, -1, -3, -4, -5, -3, -1, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, 2, 1, 2, 1, 0, 0, 0, 0, -2, -4, -4, -2, 0, 0, 0, 0, 0, -1, -2, -2, -2, 2, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 1, -2, -2, -2, -2, -2, -1, 1, 0, 1, 0, 0, 0, -2, -2, 1, 0, 0, 0, 0, 1, 2, 0, 0, -1, -1, -1, -3, -2, -3, -2, 0, 0, 1, 1, 3, 1, 0, 1, -1, -1, 1, 0, 0, 0, 0, 2, 2, 0, 0, -1, -1, -1, -2, -1, -1, -1, 0, 2, 3, 2, 1, 2, 1, 0, 0, -1, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, -2, -1, -3, 0, -2, 0, 0, 1, 0, 1, 0, 1, 1, 1, 1, 0, 1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, -1, -2, -1, -3, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, -1, 0, 0, -1, 3, 1, -1, -1, -1, -2, 0, -1, -2, 0, 0, 0, 0, 2, 0, 0, 0, -1, -1, -2, -2, -1, -1, 0, 0, 0, 2, 2, 0, -1, -1, -2, -2, -3, -2, 0, 0, 1, 2, 1, 2, 2, 2, 1, 1, 0, -1, -1, -1, -1, -1, 0, 6, 3, 2, 1, 0, 0, -2, -2, -2, -1, 0, 2, 2, 4, 3, 5, 4, 5, 4, 1, 0, 1, 1, 1, 2, 1, 2, 0, 1, 0, -1, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, -2, -1, -2, -2, -2, -4, 0, 1, 1, -1, 0, -2, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, -1, -1, -1, -2, -4, -4, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -2, -1, -4, 0, 0, 0, -1, -1, -1, -3, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, -2, -2, -3, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -3, 1, 0, 0, -1, -2, -1, -2, -2, -2, -2, -2, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -2, 1, 1, 0, 0, -1, 0, -2, -2, 0, -2, -2, 0, -1, -2, -1, 0, 0, 0, 0, 2, 1, 0, 0, -1, 0, 0, 2, 0, 1, 0, 0, 0, -1, -2, -2, 0, -1, -1, 0, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -1, 2, 2, 2, 0, 0, 0, 0, 0, -1, 0, -2, -2, 0, 0, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -1, 1, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, -1, -2, -3, -1, -2, 0, 1, 1, 1, 0, -1, 0, -1, 0, -2, 1, 2, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, -2, -2, -1, -1, -2, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 2, 1, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -2, -2, -2, -1, 0, 1, 2, 1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -2, -3, -1, 0, 0, 0, 2, 2, 1, 0, -1, -1, 0, -1, 0, 0, 0, 1, -1, -1, -1, 0, 0, 0, 0, -1, 0, -3, -1, 0, 0, 2, 1, 0, 1, 1, -1, -1, -2, 1, 1, 0, 0, 0, -1, -1, -2, 0, 0, -1, 0, -2, -3, -2, -1, -1, 1, 1, 1, 0, 0, 0, 0, -1, -1, 3, 1, 0, 0, 0, -2, -3, -2, 0, 0, 0, -2, -3, -3, -3, -2, -1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 2, 2, 1, -1, 0, -3, -2, -1, -3, 0, 0, -1, -2, -1, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 3, 1, 1, -1, -1, -3, -2, -1, -2, -1, 0, -1, 0, -3, -2, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 2, 1, 0, 0, -1, -3, -3, -3, -1, -1, -2, -3, -2, -1, 0, -2, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, -1, -1, -2, -1, -1, -3, -2, -1, -3, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -2, 2, 1, -1, -1, -2, -2, -2, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 2, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -2, -2, -1, -2, 2, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, -1, -2, 3, 2, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -2, -2, -3, -3, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, -1, -2, -1, -3, -4, -2, -3, 5, 3, 0, -1, -2, -2, -2, -2, 0, -1, 0, 0, 1, 3, 1, 2, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, 3, 1, -1, -1, -1, -2, -2, -1, -1, 0, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, 3, 0, -2, -2, -1, -2, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 4, 0, -1, -2, -2, -1, -2, -1, -2, -1, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 4, 1, 0, -2, -1, -2, -2, -3, -1, -1, -2, -1, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 3, 1, 0, -1, -1, -2, -2, -1, -2, -3, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 6, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 1, 1, 0, 2, 1, 0, 0, 0, 4, 2, -1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 0, -2, 0, -2, 0, 1, 1, 0, 0, 1, 1, 0, 0, 4, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -4, -3, -4, -2, 0, 0, 1, 0, -1, -1, -1, -1, 0, -1, -2, 0, -1, 0, 0, 0, -2, 0, 0, 0, -1, -1, -2, -3, -2, -1, 0, 0, 2, 1, 0, -1, 0, -1, 0, -2, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -2, 0, 1, 3, 1, 1, 0, -2, -2, 0, -3, -4, -1, -1, 1, 0, 0, -1, 0, 0, 0, 0, -1, -2, -2, -2, 0, 1, 3, 3, 2, 0, 0, 0, 0, 1, 0, -3, -3, -1, 0, 0, 0, -1, 0, 1, 1, -1, -3, -2, -4, -2, 0, 1, 2, 3, 1, 0, 0, 0, -2, 1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 1, 0, -1, -2, -2, -4, -1, 0, 0, 2, 1, 0, 0, 0, 0, -1, 3, 0, 0, -2, 0, 0, 0, 0, -1, 1, 0, 0, -1, -2, -2, -2, -2, 0, 0, 0, 0, 0, 0, -2, 0, -2, 2, -1, 0, -1, -2, -1, 0, -1, -1, 0, 0, 0, -2, -1, -3, -4, -1, 0, 0, 2, 1, 1, 1, -1, -2, 0, 4, 0, -2, 0, -1, -1, 0, 0, -2, -1, 0, -1, -1, -2, -2, -2, -1, 0, 0, 1, 0, 2, 0, 0, 0, 0, 2, 0, 0, -1, 0, -1, 0, -1, -2, -2, -1, -3, -2, -2, -2, -1, -2, 0, 0, 1, 1, 1, 0, 1, 1, 0, 4, 0, -1, 0, 0, -1, -1, -2, 0, -2, -2, -3, -2, -1, -1, -2, -1, 1, 1, 1, 2, 2, 3, 2, 0, 0, 3, 0, -1, -1, -2, -1, -1, 0, -2, -3, 0, -1, 0, 0, -2, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 3, 0, -1, -2, -3, -3, -2, -3, 0, -2, 0, -1, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 3, 0, -1, -3, -2, -3, -3, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, 4, 0, 0, -1, -2, -1, -3, -2, -1, -2, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 6, 1, 0, -1, 0, -1, -3, -3, -2, 0, -1, 0, 0, 1, 1, 3, 3, 1, 1, 0, 0, 0, -1, 0, 0, 0, 9, 3, 3, 2, 1, 0, -1, 0, 0, 0, 0, 2, 2, 4, 3, 3, 3, 2, 3, 3, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, -1, -2, -2, -1, 0, -1, 1, 0, 1, 1, 2, 1, 2, 2, 2, 1, 2, 3, 2, 2, 2, 0, -2, -1, 0, -1, -1, -1, -2, -2, 0, 0, -1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 1, 1, 2, 1, 2, -1, 0, -2, 0, 0, 0, 0, -1, 0, -2, -2, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 1, 2, 0, 0, -1, 0, 1, -1, 0, 0, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 1, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -2, 0, -1, 0, 0, 0, 0, 0, 1, 0, 2, 3, 3, 2, 1, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 3, 3, 3, 2, 1, 0, -1, 0, -2, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 2, 2, 2, 1, 3, 3, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 1, 3, 2, 1, 3, 2, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -2, 0, 0, 1, 2, 2, 2, 2, 3, 3, 2, 2, 0, 0, 0, 1, 1, 0, 0, 0, -2, -3, -1, -2, 0, 0, -1, 0, 0, 1, 3, 1, 1, 3, 1, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, -2, 0, 0, 2, 3, 3, 2, 1, 1, 0, 2, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, 1, 3, 4, 4, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -2, 0, 0, 1, 3, 3, 2, 2, 2, 1, 2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, -2, 0, 1, 2, 3, 2, 2, 1, 2, 1, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -2, 0, 0, 0, 2, 3, 3, 1, 2, 3, 3, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, -1, 0, -2, 0, -1, 1, 1, 2, 1, 1, 1, 3, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 2, 2, 3, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 2, 2, 3, 2, 1, 0, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, 1, 3, 2, 4, 3, 1, 0, 1, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, -2, -1, 0, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, -2, 0, -1, 0, 0, 1, 1, -1, -1, 0, 0, -1, 0, -1, -2, -2, -2, -1, 0, -2, 0, 0, 0, 0, 0, 1, -2, 0, -1, -1, 0, 0, 0, 0, 0, -2, 0, -1, -1, -1, -2, -2, -2, -2, 0, -1, 0, -1, 1, 0, 1, 0, -1, -2, -1, 0, 0, -1, -1, -1, -1, -2, -1, -1, -1, -1, -1, -1, -1, -2, -2, 0, 0, 0, 1, 0, 0, 1, 0, 2, 3, 2, 2, 4, 3, 1, 0, 0, 2, 3, 2, 3, 2, 3, 2, 3, 3, 3, 3, 0, 1, 1, 1, 3, 2, 1, 2, 2, 2, 2, 1, 0, 0, 0, 1, 1, 1, 1, 1, 2, 1, 1, 1, 1, 2, 0, 0, 0, 0, 3, 2, 2, 2, 1, 1, 1, 0, -2, 0, -1, 1, 1, 0, 1, 2, 1, 1, 0, 3, 2, 2, 1, 1, 2, 2, 3, 1, 0, 0, 1, 1, 2, 0, 0, 0, 2, 2, 0, 0, 0, 2, 3, 0, 0, 1, 2, 2, 0, 0, 3, 2, 2, 0, 0, -1, 1, 1, 2, 1, 1, 2, 4, 2, 1, 0, 2, 2, 4, 1, 1, 3, 1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 2, 2, 3, 4, 2, 5, 4, 1, 0, 1, 2, 2, 4, 2, 1, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 3, 2, 4, 2, 2, 2, 2, 2, 0, 1, 2, 2, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 1, 1, 2, 2, 2, 2, 1, 2, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, -2, -1, 0, 2, 0, 1, 1, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 3, 0, -1, -4, -2, 1, 3, 3, 3, 2, 1, 1, -1, -2, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, -1, -1, 3, 0, -1, -2, 0, 3, 4, 5, 3, 1, 0, 2, 1, 1, 0, 1, 1, 1, -1, 0, -1, 0, -1, 0, -1, -1, 2, 2, 0, 0, 3, 6, 8, 6, 5, 3, 1, 2, 1, 0, 2, 2, 0, -1, -2, -2, -1, -1, 0, 0, -1, 0, 3, 3, 0, 3, 5, 6, 8, 5, 4, 2, 0, 0, 1, 0, 2, 1, 1, -2, -2, -3, -4, -2, 0, 1, 0, 0, 4, 2, 2, 3, 6, 9, 9, 7, 2, -1, -3, -1, -2, 0, 0, 2, 2, 0, 0, -2, -1, -1, 0, 0, 0, 1, 2, 1, 3, 5, 6, 9, 11, 6, 4, 0, -2, -4, -1, -1, 0, 1, 1, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 2, 4, 5, 9, 11, 10, 8, 4, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, 0, 1, 1, 3, 5, 6, 9, 10, 7, 4, 2, 2, 0, -1, -1, -1, -3, -3, -3, -2, 0, -2, 0, 0, 0, 0, 0, 0, 1, 3, 5, 5, 7, 7, 5, 4, 2, 1, 0, -1, -1, -1, -3, -1, -2, -2, -3, -3, 0, -1, 0, 0, 0, 3, 1, 2, 3, 2, 2, 3, 3, 4, 3, 1, 0, -1, 0, 0, -1, 0, 0, 0, -2, -1, -1, -1, -1, -1, 0, 2, 1, 0, 0, 2, 1, 1, 3, 3, 4, 2, 2, 0, 1, 2, 1, 1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 3, 0, 0, 1, 1, 1, 1, 4, 4, 5, 4, 1, 1, 1, 1, 0, 1, 2, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 1, 3, 4, 4, 5, 2, 1, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 2, 2, 3, 3, 4, 3, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 1, 2, 2, 1, 2, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, -1, -2, -1, 1, 0, 0, 0, 0, -2, -1, -2, -1, -2, -2, 0, -2, 0, 0, 2, 2, 2, 2, 1, 1, 0, -1, -1, -3, 0, 0, -2, 0, 0, -2, -1, -2, -3, -3, -3, -4, -3, -2, -2, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 4, 1, 1, 1, -1, -2, -2, -1, 0, 0, 3, 3, 4, 4, 5, 3, 3, 3, 1, 1, 0, 0, -3, -2, -1, -2, 3, 2, -1, -1, -3, -1, -2, -2, 0, 0, 2, 2, 2, 4, 2, 2, 1, 0, 0, -1, -2, 0, -1, -2, -2, -1, 2, 1, -1, -1, -2, -2, -2, 0, 0, 0, 2, 3, 2, 3, 1, 2, 2, 1, 0, 0, -2, -2, -2, -2, -1, 0, 3, 1, 0, -3, -2, -2, -3, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 2, 0, -1, -2, -2, -3, -3, -1, -1, -1, -1, -2, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 3, 1, 1, -1, -2, -4, -4, -4, -3, -4, -3, -3, 0, -1, -1, 1, 1, 0, 2, 2, 1, 1, 2, 2, 1, 0, 4, 1, 0, 1, 0, -3, -3, -4, -6, -4, -4, -3, -3, -2, -1, -1, 0, 1, 1, 2, 2, 2, 1, 1, 0, 1, 5, 2, 0, 0, 0, -2, -2, -3, -5, -6, -4, -5, -3, -4, -3, 0, 0, 2, 0, 2, 2, 2, 0, 0, 0, 0, 6, 1, 2, 1, -1, -2, -1, -3, -3, -4, -3, -4, -3, -3, -4, -3, -2, 0, 1, 2, 2, 1, 0, 2, 0, 2, 5, 2, 0, 0, 1, 0, -2, -1, -2, -2, -3, -2, -3, -3, -5, -5, -1, 0, 1, 2, 2, 2, 3, 0, 0, 1, 2, 0, 0, 0, 0, 0, -1, -2, -2, -2, -3, -3, -4, -4, -5, -4, -2, 0, 2, 3, 4, 4, 3, 1, 1, 0, 0, -1, -1, -1, -2, -2, -1, -3, -4, -3, -1, -2, -4, -5, -6, -3, -1, 1, 3, 5, 7, 6, 2, 2, 1, 0, -1, -3, -3, -2, -3, -3, -2, -2, -4, -3, -1, -3, -4, -5, -5, -2, 0, 3, 6, 8, 8, 7, 3, 2, 1, 0, -1, -3, -2, -3, -3, -3, -2, -3, -3, -2, -2, -1, -3, -2, -5, -2, 0, 4, 6, 8, 7, 6, 4, 1, 1, 1, 0, -1, -1, -3, -2, -3, -3, -3, -2, -1, -1, -2, -4, -4, -5, -3, 0, 1, 5, 7, 5, 6, 3, 1, 0, 1, 1, 0, -1, -1, -2, 0, -3, -2, -3, -2, -2, -1, -4, -6, -4, -4, -3, 0, 4, 4, 4, 3, 3, 0, 0, 1, 3, 1, 1, 0, 0, -1, -2, -1, -2, -2, -3, -3, -5, -5, -5, -4, -1, 1, 1, 3, 2, 2, 1, 0, 0, 1, 3, 0, 0, 0, 0, 0, -2, -3, -3, -2, -2, -2, -4, -4, -3, -4, -1, 0, 0, 2, 1, 3, 2, 0, 0, 0, 3, 1, -1, -1, -1, -1, -1, 0, -1, -2, -3, -3, -4, -3, -3, -1, 0, 1, 1, 2, 3, 3, 3, 0, 1, 0, 2, 1, -1, 0, 0, 0, -2, -1, -3, -2, -2, -4, -3, -3, -1, 0, 0, 2, 4, 4, 3, 4, 2, 1, 2, 1, 3, 0, 0, 0, -2, -2, 0, -3, -3, -4, -4, -2, -2, -1, -1, 1, 0, 2, 4, 3, 2, 3, 3, 1, 0, 0, 3, 0, -1, -2, 0, 0, -1, 0, -2, -2, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 0, 0, 1, 0, -1, -2, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 2, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 2, 2, 0, 1, 0, 0, -1, -2, -1, -1, -2, -1, -2, 3, 2, 0, 0, 0, 0, -1, 0, 0, 2, 1, 0, 1, 1, 3, 1, 0, 1, -1, 0, 0, -2, -1, -2, 0, -2, 5, 2, 0, 1, 0, 0, -1, 0, 0, 1, 3, 2, 2, 3, 3, 2, 3, 1, 0, 0, -1, -1, -2, -1, 0, -2, -3, -2, -1, 0, 0, 0, -1, -2, -1, -1, -2, -1, -1, -1, -1, -2, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 1, 0, 1, 1, 0, 0, -2, -2, -1, -1, -2, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, -2, -2, -1, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 1, 0, -1, 1, 1, 1, 0, 1, 0, 0, 0, 0, -2, -1, -1, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -2, -1, 1, 1, 1, 2, 1, 2, 2, 1, 0, -1, 0, 0, -1, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 0, 2, 1, 0, 0, -1, -1, 0, -1, 0, -2, -1, -2, -1, -1, 0, -2, -1, -1, -2, 0, -1, 0, 2, 1, 1, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 1, 1, 1, 2, 1, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, -2, 0, 0, 0, 1, 2, 1, 3, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -2, 0, 0, 0, 1, 2, 0, 3, 2, 2, 2, 2, 2, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 1, 1, 1, 1, 1, 2, 2, 2, 2, 2, 0, -1, 0, -1, 0, -1, 0, -1, -1, 0, -2, -1, -1, 0, 0, 2, 2, 2, 2, 3, 3, 2, 2, 1, 1, 0, 1, 0, -2, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, 2, 2, 3, 1, 1, 3, 2, 2, 0, 1, 0, -2, -1, -2, -1, -1, 0, 0, 1, -1, -2, 0, 0, 0, 1, 0, 2, 1, 2, 1, 2, 1, 2, 1, 0, 1, -1, -1, -2, -2, 0, 0, 0, 0, 1, -3, 0, -1, 0, 0, 0, 1, 1, 2, 3, 1, 0, 1, 2, 0, 1, 0, 0, 0, -2, 0, 0, -1, 1, 1, 0, -1, -2, -1, 0, 0, 1, 2, 2, 2, 2, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, -2, -3, 0, -1, 0, 2, 2, 2, 3, 2, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -3, -2, 0, 0, 1, 2, 3, 2, 4, 3, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, -1, -1, 0, 0, 2, 2, 2, 2, 3, 2, 1, 1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 2, 1, 3, 1, 2, 1, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, -2, 0, -1, 0, -2, 0, -1, 0, 0, 0, 1, 0, 1, -2, -1, 0, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, -2, 0, -2, -1, -2, -1, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 1, 1, 0, -1, 0, -2, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, -2, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -2, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 1, 1, 1, 2, 1, 1, 0, -1, -1, -3, -1, -2, -3, -1, 0, 1, 3, 3, 7, 8, 10, 10, 9, 7, 7, 5, 4, 3, 3, 3, 6, 6, 9, -1, -2, -4, -2, -3, -2, -2, -1, 1, 2, 2, 4, 5, 7, 6, 4, 4, 4, 1, 3, 3, 3, 3, 4, 4, 7, -4, -5, -2, -4, -2, -3, -2, -1, 0, 0, 0, 0, 2, 2, 2, 2, 3, 1, 1, 0, 0, 1, 1, 1, 3, 5, -3, -4, -4, -3, -2, -2, -3, -1, 0, 0, 0, 0, 0, 1, 2, 0, 1, 1, 1, 0, 0, -1, 0, 1, 2, 4, -4, -1, -1, -1, -2, -1, -2, -3, -3, -3, -2, -1, 0, 1, 0, 2, 3, 1, 3, 2, 1, 0, 1, 1, 2, 4, -2, -1, 0, 0, 0, -1, -3, -3, -3, -3, -1, -2, -2, 0, 0, 1, 1, 1, 3, 3, 1, 1, 0, 2, 3, 4, -1, -1, -2, 0, -1, -1, -2, -2, -2, -1, -2, -2, 0, -1, 0, 0, 0, 2, 2, 3, 3, 1, 1, 0, 1, 3, -1, -1, 0, 0, 0, -1, -1, 0, 0, -2, -1, -1, -2, -2, -3, -2, -1, 0, 0, 1, 1, 3, 1, 2, 0, 2, -1, -3, -1, -1, 0, 0, 0, 0, 0, -1, -1, -2, -2, -4, -5, -5, -3, -1, 0, 1, 1, 2, 0, 1, 0, 2, -3, -3, 0, 1, 0, 1, -1, -1, 0, -1, 0, -1, -3, -5, -6, -5, -3, -2, 2, 3, 5, 2, 2, 0, 0, 2, -3, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, -2, -4, -5, -6, -6, -2, 2, 6, 7, 7, 4, 2, 2, 0, 2, -4, -3, -1, -1, -1, 0, 0, -2, -2, 0, 0, -1, -3, -3, -4, -4, -1, 4, 8, 10, 8, 6, 4, 2, 0, 1, -2, -2, -1, -2, -1, -1, -1, -1, -1, -1, 0, -1, -2, -3, -4, -3, 0, 3, 7, 9, 9, 6, 3, 2, 1, 2, -4, -2, -1, -2, -2, -2, -2, -1, 0, -2, 0, 0, -3, -6, -6, -5, -2, 2, 6, 9, 8, 7, 5, 2, 1, 1, -1, -1, -1, -3, -1, -1, -1, -1, -1, -1, 0, -2, -2, -6, -6, -5, 0, 2, 4, 7, 6, 4, 3, 1, -1, 0, 0, -3, -1, -1, -2, 0, 0, 0, 0, -1, 0, -1, -3, -5, -7, -6, -1, 1, 4, 5, 2, 1, 0, -1, 0, 1, -1, -2, -1, -1, 0, -1, 0, 0, 0, -1, 0, -1, -2, -5, -6, -5, -2, 0, 2, 4, 2, 2, 1, -1, 0, 2, -3, -2, -3, -1, -2, 0, 0, 0, -1, -2, -3, -3, -3, -3, -3, -3, -2, 0, 3, 3, 3, 3, 0, 0, 0, 2, -3, -2, -2, -1, -1, 0, 1, 0, -3, -4, -4, -3, -1, -1, -1, 0, 0, 2, 4, 4, 5, 3, 1, 2, 2, 2, -3, -3, -3, -2, -2, -1, 0, -1, -1, -3, -4, -2, 0, -1, 0, 0, 2, 1, 2, 4, 4, 3, 2, 1, 2, 3, -2, -3, -3, -4, -3, -1, -1, -2, -2, -2, -2, -1, -1, 0, 0, 1, 1, 1, 2, 2, 0, 0, 2, 2, 1, 3, -1, -4, -5, -3, -4, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 5, -1, -2, -3, -3, -4, -4, -3, -2, -1, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, 0, 0, 2, 2, 4, 0, -1, -3, -3, -4, -2, -4, -3, -3, -1, -1, 0, 1, 1, 1, 2, 2, 0, 0, -1, 0, 0, 0, 1, 4, 6, 0, 0, 0, 0, -1, -2, -3, -2, -1, -1, 1, 3, 4, 6, 6, 4, 5, 4, 3, 1, 0, 0, 3, 3, 4, 8, 2, 1, 2, 2, 1, 0, -1, 0, 0, 2, 5, 6, 8, 11, 9, 9, 9, 8, 7, 5, 6, 7, 6, 7, 10, 12, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 1, 1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, -1, 0, 1, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 4, 3, 2, 2, 2, 2, 4, 4, 3, 4, 3, 2, 3, 1, 0, 1, 0, -2, -4, -2, -4, -2, -3, -5, -2, 1, 2, 4, 3, 3, 1, 1, 2, 3, 3, 2, 2, 3, 4, 2, 1, 0, 1, -3, -4, -2, -3, -2, -5, -3, -4, 1, 4, 3, 4, 2, 1, 1, 1, 2, 4, 2, 3, 3, 3, 3, 4, 2, 1, -1, -4, -3, -3, -2, -5, -4, -1, 1, 5, 3, 3, 0, 0, 0, 1, 3, 2, 2, 2, 3, 3, 3, 3, 2, 2, 0, -3, -2, -2, -2, -3, -3, -1, 4, 6, 5, 1, 2, 0, 0, 1, 1, 1, 0, 1, 0, 3, 3, 3, 1, 0, 0, -2, -1, -1, 0, -1, -3, -2, 5, 5, 3, 3, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 1, 2, 1, 1, 0, -1, -2, 0, 0, 0, -1, -1, 3, 5, 4, 1, 0, 0, 0, -1, -3, -4, -3, -3, -2, -2, 0, 0, 1, 0, 0, -2, 0, 0, 0, -2, -1, -2, 3, 5, 4, 3, 1, 1, 0, -2, -3, -6, -5, -5, -6, -3, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, 3, 4, 5, 5, 3, 1, 0, -2, -3, -6, -8, -8, -6, -4, -1, 1, 3, 2, 1, 0, 0, -1, 0, -2, 0, 0, 2, 3, 6, 6, 2, 1, -1, -2, -6, -8, -10, -9, -8, -3, 0, 2, 5, 4, 2, 1, 0, -1, -1, 0, 0, 0, 3, 2, 5, 4, 3, 0, -1, -4, -7, -7, -10, -9, -7, -3, 0, 2, 4, 4, 4, 1, 1, 0, 0, 1, 1, 1, 1, 3, 4, 2, 1, -2, -4, -6, -6, -9, -9, -8, -7, -2, 1, 3, 5, 6, 5, 3, 0, 0, 0, 0, 0, 2, 0, 1, 1, 1, 0, -3, -3, -5, -8, -9, -9, -8, -7, -1, 0, 4, 6, 7, 7, 3, 0, 0, 0, -1, 1, 2, 1, 2, 2, 0, 0, -2, -6, -6, -8, -6, -8, -7, -6, -1, 0, 3, 6, 7, 5, 3, 2, 0, 0, 0, 0, 3, 0, 2, 2, 1, 0, -2, -4, -5, -6, -7, -8, -8, -7, -3, 0, 3, 3, 5, 4, 2, 0, 0, 0, 1, 1, 3, 2, 3, 1, 0, 0, -2, -3, -5, -5, -8, -9, -8, -5, -3, -1, 2, 4, 2, 3, 2, 0, 0, 0, 0, 2, 2, 3, 4, 4, 3, 0, 0, -3, -5, -4, -4, -7, -7, -6, -3, 0, 0, 3, 0, 1, 0, 0, 0, 0, 2, 0, 2, 3, 5, 4, 4, 1, 0, -1, -2, -2, -4, -6, -6, -5, -4, -1, 1, 1, 1, 0, -2, -2, 0, 0, 0, 0, 0, 3, 5, 5, 4, 2, 0, -1, 0, -3, -5, -6, -4, -3, -2, 0, 1, 1, 0, -1, -1, -2, -2, -1, 0, -2, 1, 3, 3, 4, 2, 1, 2, 0, -1, -3, -3, -5, -5, -2, -1, 0, 1, 0, -1, 0, -2, 0, -1, -2, -2, 0, -1, 1, 3, 4, 2, 4, 2, 1, 0, -1, -3, -3, -1, 0, 0, 2, 0, 0, -2, -2, -1, -2, 0, -1, -2, -2, -2, 2, 2, 3, 4, 4, 3, 1, 1, 0, 0, -1, -1, 0, 0, 2, 0, -1, -2, -1, -1, 0, -1, 0, 0, -2, 0, 1, 3, 2, 5, 4, 2, 3, 2, 0, 0, 0, 0, 2, 3, 1, 0, -1, -2, -2, 0, -1, -1, -1, -1, -1, -1, 0, 1, 1, 4, 5, 4, 2, 2, 1, 2, 2, 0, 3, 3, 2, 0, -1, -2, -2, -4, -3, -2, -2, -3, -1, -1, 0, 1, 2, 3, 3, 2, 2, 3, 4, 3, 2, 4, 2, 4, 2, -1, -2, -2, -2, -3, -3, -3, -3, -3, -3, -1, 0, 1, 4, 4, 4, 2, 3, 3, 4, 6, 4, 5, 3, 3, 0, 0, 0, -2, -2, -4, -4, -3, -3, -4, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -2, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 1, -1, 0, 0, -1, 1, 1, 0, 1, 1, 1, 0, 1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 2, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 2, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, -1, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 2, 3, 1, 3, 2, 2, 1, 2, 0, -1, -3, -2, -3, -4, -4, -5, -4, 1, 1, 0, 0, -1, 0, 0, 0, 0, 2, 1, 3, 3, 3, 2, 1, 1, 1, -1, -1, -3, -3, -4, -5, -3, -4, 0, 1, 0, -1, 0, -1, -2, 0, 0, 2, 1, 1, 3, 2, 3, 1, 2, 2, 0, -1, -1, -2, -3, -3, -2, -4, 1, 0, 1, 0, 0, -2, 0, -1, 1, 0, 1, 0, 1, 0, 1, 3, 1, 0, 0, -2, -1, -1, 0, -1, -2, -1, 3, 1, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 4, 2, 1, 0, -1, -2, -1, -2, -2, -2, -3, -3, -2, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 3, 4, 3, 0, 0, 0, -3, -3, -5, -6, -6, -6, -5, -2, 0, 1, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 5, 4, 2, 3, 0, -1, -3, -2, -3, -5, -8, -8, -6, -4, -3, -1, 0, 1, 1, 1, 2, 2, 2, 1, 0, 0, 3, 4, 5, 2, 0, 0, -1, -3, -5, -5, -7, -8, -7, -4, -1, 0, 0, 1, 3, 2, 3, 1, 2, 2, 0, 0, 4, 3, 4, 3, 2, 1, -1, -2, -6, -5, -7, -9, -6, -4, -1, 0, 0, 4, 2, 2, 2, 3, 2, 0, 1, 1, 3, 3, 3, 3, 2, 0, -2, -4, -4, -7, -6, -6, -7, -4, -2, 0, 1, 4, 3, 4, 5, 4, 2, 1, 2, 1, 1, 1, 2, 1, 0, -2, -2, -3, -6, -7, -6, -6, -5, -3, -1, 0, 1, 4, 5, 6, 5, 3, 3, 2, 2, 1, 0, 0, 0, 0, 0, -2, -3, -4, -6, -6, -6, -5, -4, -3, 0, 0, 2, 6, 6, 8, 6, 4, 3, 1, 2, 1, 0, 0, 0, 0, -1, -1, -5, -4, -6, -7, -7, -6, -5, -3, -2, 1, 2, 5, 7, 9, 5, 4, 3, 2, 1, 3, 0, 1, 1, 0, 0, -1, -4, -4, -6, -7, -7, -7, -5, -3, -2, 0, 2, 4, 5, 7, 6, 4, 4, 3, 2, 1, 1, 1, 1, 0, -1, -3, -3, -4, -5, -7, -6, -5, -4, -4, -3, 0, 0, 3, 5, 4, 4, 3, 2, 1, 1, 1, 2, 1, 1, 0, 0, -1, -4, -5, -5, -6, -6, -6, -5, -5, -3, -2, 0, 0, 2, 1, 3, 2, 1, 1, 2, 3, 3, 3, 1, 0, 0, 0, -2, -3, -5, -6, -7, -5, -4, -3, -1, 0, 0, 0, 1, 2, 2, 1, 3, 2, 1, 2, 2, 1, 1, 2, 0, 0, 0, -1, -3, -4, -7, -5, -4, -1, -1, 0, 0, 0, 1, 1, 3, 3, 3, 1, 1, 2, 1, 2, 1, 0, 0, 0, -2, -1, -4, -3, -5, -5, -2, -1, 0, 1, 0, 2, 2, 3, 2, 2, 1, 1, 1, 0, 1, 2, 1, 0, 1, 0, 0, -2, -1, -3, -4, -1, 0, -1, 0, 0, 1, 1, 2, 3, 2, 3, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 1, 0, 0, 1, 1, 1, 1, 1, 1, 0, -1, 0, -1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 1, 0, 0, 1, 0, -1, -1, -1, -1, -2, -2, -2, -3, -1, -2, 1, 0, 0, 1, 0, 1, 1, 1, 2, 1, 2, 3, 2, 3, 0, 0, -1, 0, -2, -2, -3, -3, -3, -5, -2, -2, 1, 0, 1, 1, 1, 0, 0, 2, 3, 2, 3, 1, 2, 2, 2, 0, 0, 0, -3, -2, -3, -4, -4, -3, -4, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, -1, 1, 0, 0, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 1, 1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, -1, 1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, -1, 1, -1, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, -1, 1, 0, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -2, -3, -4, -4, -3, 0, 2, 3, 5, 8, 9, 8, 8, 7, 6, 3, 5, 2, 2, 3, 5, 5, 6, -3, -2, -3, -1, -3, -4, -2, -2, 0, 0, 2, 2, 5, 4, 5, 4, 2, 2, 1, 0, 1, 2, 2, 3, 3, 2, -4, -3, -2, -1, -3, -2, -2, 0, 1, 0, 1, 1, 1, 1, 2, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 2, -3, -2, -3, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, -4, -2, -2, 0, -2, -2, -2, 0, -1, -2, -1, -2, 0, -2, -1, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 1, -2, -2, 0, 0, 0, -1, 0, -2, -2, -1, -1, -1, -2, -1, -2, 0, 1, 1, 0, 2, 0, 0, 1, 2, 2, 3, -3, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, -2, -3, 0, 1, 1, 1, 2, 1, 1, 1, 1, 0, 2, -4, -3, -2, -1, 1, 0, 1, 1, 2, 1, 2, 0, 0, -1, -3, -2, -1, 1, 0, 0, 0, 0, 1, 0, 2, 1, -3, -4, -3, -1, 0, 0, 0, 2, 4, 3, 3, 2, 0, -4, -4, -3, -2, -1, 1, 1, 0, 1, 1, 0, 0, 1, -3, -3, -3, 0, 1, 0, 0, 1, 3, 4, 4, 1, -1, -4, -7, -5, -2, 0, 0, 1, 1, 0, 0, 0, 0, 0, -5, -4, -1, 0, 0, -1, 0, 1, 1, 4, 4, 1, -2, -4, -7, -7, -3, 0, 2, 5, 3, 2, 0, 0, 0, -1, -5, -5, -2, -1, 0, 0, 0, 0, 1, 4, 4, 0, -3, -6, -8, -7, -2, 0, 5, 6, 3, 2, 0, -1, -2, -2, -6, -5, -2, -1, 0, -1, 0, -1, 2, 1, 2, 2, -1, -5, -7, -4, -3, 1, 5, 8, 4, 2, 0, -2, -2, 0, -4, -5, -2, -1, -1, 0, -1, 0, 2, 2, 2, 1, -1, -5, -6, -7, -3, 1, 5, 6, 4, 3, 0, 0, -2, -3, -4, -4, -4, -2, -2, 0, 1, 0, 1, 3, 2, 1, -2, -4, -7, -6, -4, -1, 2, 4, 4, 1, -1, -2, -2, -2, -4, -4, -3, -1, 0, 0, 1, 3, 3, 3, 1, 1, -1, -6, -6, -7, -3, -2, 1, 2, 0, -1, -2, -2, -2, -3, -5, -3, -4, 0, 0, 0, 1, 2, 3, 1, 1, 1, -2, -4, -7, -5, -3, -1, 1, 0, -1, 0, -2, -1, -2, -1, -4, -5, -2, -2, 0, 2, 4, 2, 1, 0, 0, 1, 0, -3, -4, -5, -2, 0, 0, 2, 0, 0, -3, -1, -2, -2, -4, -4, -3, 0, 1, 3, 3, 2, 0, 0, 0, 0, -1, -3, -1, -3, -2, 0, 1, 3, 3, 0, 0, 0, -2, -1, -4, -4, -2, -1, 0, 1, 3, 1, -1, -2, 0, 0, 0, -1, -2, -1, 0, 1, 3, 2, 2, 2, 0, 0, 0, 0, -2, -4, -2, 0, 0, 0, 0, 1, 0, 0, -2, 0, -1, -1, -1, 0, 0, 1, 1, 0, 2, 0, 0, 0, 0, 1, -4, -2, -3, -1, -1, -1, -1, 0, -1, -1, -2, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, 1, 1, 0, 2, -4, -2, -3, -4, -3, -4, -1, -2, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, -2, -3, -3, -2, 0, 0, 1, 2, -1, -3, -3, -4, -3, -4, -3, -1, -1, 0, -1, 0, 1, 0, 0, 2, 1, 0, 0, -2, -1, -2, -1, 0, 0, 2, -1, -1, -2, -1, -2, -3, -3, -1, -2, 0, 0, 0, 3, 3, 3, 5, 4, 2, 3, 0, 0, 0, 1, 3, 2, 3, 1, 0, 1, 1, 0, -1, -3, -2, -1, 1, 2, 4, 6, 8, 9, 10, 9, 6, 7, 5, 3, 4, 6, 6, 5, 8, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 1, -1, -1, 0, 0, 1, 0, 0, -1, 0, -2, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, -1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 1, -1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 1, 0, 0, -1, 0, -1, 1, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -2, 0, 0, 0, 2, 0, 2, 1, 2, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 1, 1, 0, 1, 0, 1, 1, 2, 1, 1, 2, 1, 0, -1, -1, -1, 0, -1, 0, 0, 1, -2, 0, 0, 0, 0, 1, 1, 0, 1, 1, 2, 0, 1, 0, 1, 1, 0, -1, 0, -2, -1, -1, -1, 0, 0, 1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 1, 0, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 0, 1, 2, 1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, -2, -1, -1, 0, 0, 0, 2, 2, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 2, 3, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -3, -1, -1, 0, 0, 2, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, 0, 0, 0, 0, 1, 0, 1, 3, 1, 1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -2, -1, 0, 0, 0, 1, 2, 0, 2, 2, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 1, 1, 1, 0, 0, 0, -2, -1, -1, 0, 0, 1, 1, 0, 1, 1, 1, 0, -2, -1, 0, 0, 0, -1, -1, 0, 0, 1, 1, 1, 1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, 1, 1, 0, -2, 0, 0, 0, 0, -1, -1, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -2, -2, -2, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -2, -1, 0, -1, -1, -1, -1, -2, -2, -2, -1, -1, -2, 0, 0, -1, 0, 0, 0, 2, 2, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -2, -3, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, 1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 1, 1, 0, 2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 1, 1, 0, 0, 1, 0, 1, 1, -1, -2, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 2, 1, 0, 0, 0, 1, -1, -1, 0, 1, 1, -1, -1, 0, 0, 1, 1, 1, 2, 0, 0, 1, 0, 0, 0, 2, 0, 0, 1, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 2, 2, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, -1, 1, 1, 1, 1, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 2, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 1, 1, 1, 2, 3, 2, 3, 1, 2, 1, 1, 0, 0, 0, 2, 1, 0, -1, -1, -1, -1, 0, 0, 0, 1, 1, 1, 3, 1, 4, 3, 3, 2, 1, 0, 0, 1, -1, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 1, 3, 2, 3, 4, 4, 4, 2, -1, 0, -2, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, -1, -1, 0, 1, 1, 0, 1, 2, 3, 5, 4, 4, 2, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, -1, -1, 0, 2, 4, 6, 5, 3, 2, 2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 3, 5, 4, 4, 1, 1, 1, 1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 2, 1, 2, 2, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 2, 1, 1, 0, 2, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 2, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, -2, 0, -1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 2, 2, 1, 2, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 1, 1, 1, 2, 2, 2, 3, 2, 1, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 2, 1, 1, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 1, 0, 1, -1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, -1, -1, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 1, 1, 0, 0, 2, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, -1, 0, 0, 0, 2, 0, 0, 2, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 2, 2, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -2, -1, 0, 0, -1, 0, 0, 1, 1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 3, 1, 2, 1, 2, 2, 1, 3, 3, 3, 2, 2, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, -1, 0, 2, 1, 1, 0, 1, 1, 1, 0, 2, 2, 1, 1, 2, 2, 1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 2, 0, 1, 1, 0, 0, 0, 0, 1, 2, 3, 1, 2, 3, 2, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 3, 3, 1, 2, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 1, 0, 0, 2, 2, 1, 2, 2, 2, 3, 2, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, -2, -2, -1, 0, 0, 1, 0, 0, 2, 1, 2, 1, 3, 3, 1, 2, 0, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 2, 2, 3, 1, 2, 3, 1, 2, 2, 1, 1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 2, 3, 2, 2, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, -1, 0, 0, -1, 0, 0, 0, 1, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 2, 1, 1, 2, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, -1, 0, 0, 2, 2, 1, 1, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 2, 1, 2, 2, 1, 1, 0, 1, 1, 0, -2, 0, -1, 0, -1, -2, -2, 0, 0, 1, 1, 0, 2, 2, 2, 2, 1, 2, 1, 0, 2, 1, 1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 2, 2, 0, 0, 0, 2, 0, 2, 1, 0, 0, 0, 0, -1, 0, -2, -1, -1, -1, 0, 0, 0, 0, 2, 0, 0, 2, 2, 1, 1, 0, 0, 2, 0, 2, 0, -1, -1, -1, 0, 0, -2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 1, 2, 0, 0, 1, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 1, 2, 3, 3, 3, 4, 2, 4, 3, 4, 2, 2, 1, 2, 0, 1, 0, 0, -1, -1, -2, -2, 0, 0, 1, 1, 2, 1, 2, 3, 2, 2, 1, 2, 3, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 1, 3, 3, 2, 2, 1, 0, 1, 1, 2, 3, 3, 1, 1, 1, 1, 0, 1, 0, 0, -1, 0, -1, -2, -2, 0, 0, 2, 1, 0, 0, 1, 1, 0, 2, 2, 3, 1, 2, 2, 2, 2, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 2, 1, 2, 3, 4, 1, 0, 2, 2, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 1, 2, 2, 1, 2, 2, 3, 3, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -2, -3, 0, 0, 1, 1, 0, 1, 2, 2, 3, 2, 3, 3, 2, 3, 1, 2, 1, 1, 0, 1, -1, -1, 0, -2, -2, -1, 1, 2, 2, 2, 1, 0, 0, 1, 2, 1, 2, 3, 3, 3, 2, 3, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 1, 4, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 3, 0, 2, 0, 0, 0, -1, -2, 0, -1, 0, 0, 1, 2, 1, 1, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 2, 2, 1, 1, 1, 0, -1, -1, -2, -1, -2, 0, 1, 1, 2, 0, 0, 0, 1, 0, 2, 2, 0, 1, 1, 2, 0, 1, 0, 0, -1, -2, -2, -2, -1, -1, -1, 1, 2, 1, 1, 3, 0, 2, 0, 0, 2, 0, 2, 0, 1, 0, 0, 2, 0, 0, 0, 0, -2, 0, -1, -1, -1, 2, 3, 2, 3, 3, 0, 2, 2, 3, 2, 2, 0, 0, 2, 1, 1, 2, 1, 1, 0, -1, 0, -2, 0, -1, 0, 0, 2, 2, 3, 3, 0, 0, 1, 0, 1, 0, 0, 1, 0, 2, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 2, 2, 2, 0, 1, 1, -1, 0, 0, -1, 0, 0, 0, 1, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 1, 0, 0, 2, 0, 2, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, 0, 2, 0, 1, -1, -1, 0, 0, -1, 0, 1, 0, 0, 1, 0, 2, 3, 2, 1, 0, 0, 0, -1, -1, -2, -2, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 1, 2, 2, 0, 1, 3, 3, 2, 3, 3, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 3, 3, 2, 2, 2, 2, 3, 2, 1, 0, 1, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, 1, 1, 0, 2, 2, 3, 2, 1, 3, 1, 3, 2, 3, 3, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 2, 1, 1, 2, 1, 2, 2, 1, 1, 0, 1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 2, 0, 2, 2, 3, 2, 2, 2, 2, 1, 1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, 4, 2, 1, 0, 0, -3, -1, -1, 0, 0, 1, 2, 3, 4, 2, 2, 0, 0, 1, 0, -1, -2, -3, -2, -3, -2, 3, 0, 0, 0, -2, -1, -2, -1, -1, 0, 1, 2, 3, 1, 1, 0, 1, 1, 0, 0, -2, -1, -3, -2, -4, -4, 3, 0, 0, 0, -3, -3, -1, -2, 0, 0, 1, 0, 0, 0, 0, 2, 0, 0, 0, 0, -1, 0, -1, -1, -2, -1, 4, 1, 0, -1, -2, -3, -3, -3, -2, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 4, 0, 0, 0, -2, -3, -3, -2, -4, -2, -2, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 4, 1, 0, -1, -2, -2, -3, -3, -3, -3, -3, -1, -2, -1, 0, 0, 2, 1, 0, 0, 2, 1, 2, 0, 0, 0, 5, 1, 1, 0, 0, -1, -3, -2, -2, -3, -2, -2, -2, -1, -3, 0, 0, 0, 2, 2, 0, 1, 1, 0, 0, 0, 6, 1, 0, 0, -1, -1, -2, -1, -2, -2, -1, -1, -3, -2, -3, -2, -1, 0, 1, 2, 2, 1, 1, 0, 0, 0, 5, 1, 1, 1, 1, 0, 0, -2, -2, 0, -2, -2, -4, -3, -3, -4, -3, 0, 2, 2, 2, 1, 1, 0, 0, 0, 3, 0, 0, 1, 0, 0, -2, -1, -2, 0, 0, -3, -4, -5, -4, -4, -2, -1, 1, 2, 2, 2, 1, 0, -1, -1, 2, 0, 0, 0, 0, 0, -2, -2, -1, -2, -1, -3, -4, -5, -6, -3, -2, 0, 2, 3, 4, 2, 0, -1, -1, -1, 1, -2, 0, -1, -1, -2, -1, -1, -3, -1, -1, -1, -4, -4, -5, -3, -1, 1, 3, 6, 4, 3, 2, 0, 0, -1, 0, -1, -1, -1, 0, 0, -3, -3, -3, -2, 0, -2, -2, -3, -5, -3, 0, 2, 5, 6, 5, 4, 0, 0, -1, -1, 1, 0, -2, -1, -2, -2, -1, -2, -2, -2, 0, -1, -3, -3, -4, -3, 0, 1, 5, 5, 4, 2, 3, 0, 0, -2, 1, 0, -2, -2, 0, -2, 0, -1, 0, 0, -1, -2, -3, -4, -4, -4, -1, 2, 2, 3, 4, 2, 0, 0, -1, -2, 2, 1, -1, 0, -1, -1, -2, -2, -2, 0, 0, -2, -4, -6, -5, -4, -2, 0, 2, 3, 3, 3, 1, 0, -1, 0, 2, 1, 0, 0, 0, -1, 0, 0, -2, -1, -3, -3, -4, -5, -6, -4, -2, 0, 1, 2, 3, 2, 1, 1, 0, 0, 3, 1, 0, 0, -1, 0, -1, 0, -2, -1, -3, -2, -4, -4, -3, -2, 0, 1, 2, 3, 3, 1, 1, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, -2, -2, -2, -3, -4, -3, -5, -3, -2, 0, 0, 2, 3, 2, 3, 2, 0, 0, -1, 3, 0, 0, -1, 0, -1, -1, -2, -3, -2, -4, -5, -4, -4, -2, -1, 1, 1, 3, 3, 3, 3, 2, 2, 0, 0, 2, 0, 0, 0, -1, -1, -1, -1, -1, -3, -3, -4, -2, -2, -2, 0, 0, 2, 3, 3, 3, 3, 2, 1, 1, 0, 2, 0, -1, -1, -1, -2, -2, -1, -1, -2, -1, -2, 0, 0, 0, 0, 1, 1, 2, 2, 1, 0, 0, 1, 0, -1, 2, 0, -1, -2, -1, -2, -2, -2, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, -1, -1, -1, -1, -1, 3, 1, -1, 0, 0, -1, -1, -2, 0, 0, 0, 0, 2, 0, 3, 2, 0, 1, 1, 0, -1, -2, -2, 0, -2, -2, 6, 1, 0, 0, 0, 0, -2, -1, 1, 1, 2, 2, 3, 4, 2, 3, 3, 2, 0, 0, -1, 0, 0, -2, 0, -3, 8, 4, 3, 1, 0, 0, -1, 0, 0, 2, 4, 5, 6, 5, 5, 5, 5, 4, 3, 2, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 1, 1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, 1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, -1, -1, -1, -2, -1, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 3, 1, 0, 0, 0, -1, -2, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, -2, -2, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 2, 2, 0, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, -1, -1, 0, 0, 1, 0, -1, 0, -1, -1, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, -2, -1, -2, 0, -3, -1, 0, 0, 2, 2, 4, 6, 6, 7, 5, 4, 5, 2, 3, 2, 2, 4, 4, 3, 0, 0, -2, -2, -2, -2, -2, -1, 0, -1, 0, 0, 2, 1, 3, 4, 2, 1, 1, 1, 2, 2, 0, 3, 2, 3, 0, -1, -2, -2, -1, -3, -2, 0, 0, 1, 0, 0, 0, 0, 2, 1, 2, 0, 1, 1, 0, 0, 0, 0, 1, 2, 0, -1, -3, 0, -1, -2, -2, -3, 0, -1, 0, 0, 0, -1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, -1, -2, -1, -1, -1, -2, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 1, 1, 2, 0, 2, 1, 0, 0, 0, 1, 0, -1, 0, -1, 0, -1, -1, -2, -2, -1, 0, -1, -1, -1, 0, 0, 0, 2, 1, 1, 2, 1, 0, 0, 2, 2, 0, 0, -2, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -2, -2, 0, 1, 1, 1, 1, 0, 0, 1, 1, 0, -2, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, -1, -2, -2, -1, 0, 0, 2, 0, 1, 1, 1, 1, 0, 0, 0, -1, -1, 1, 1, 1, 1, 0, 1, 1, 1, 0, 0, -1, -3, -2, -1, 0, 0, 1, 1, 1, 1, 0, 0, 0, -2, -2, -1, 1, 1, 0, 0, 0, 0, 1, 0, 0, -2, -4, -3, -2, -2, 0, 1, 1, 2, 0, 0, 0, 0, -2, -3, -3, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, -2, -3, -4, 0, 1, 3, 3, 1, 0, 0, 0, 0, -1, -4, -2, -1, 0, 0, 0, -1, -1, 0, 1, 0, -1, -2, -3, -2, -1, 0, 2, 3, 6, 4, 1, 0, 0, 0, 0, -3, -3, -2, 0, 0, 0, -1, -1, 0, 0, 0, 0, -2, -4, -3, -3, 0, 3, 6, 6, 5, 3, 1, 0, 0, -1, -2, -3, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, -2, -4, -3, -2, -1, 1, 4, 4, 3, 2, 1, 0, -1, 0, -2, -3, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -3, -3, -1, 2, 4, 4, 2, 2, -1, 0, -1, -1, -1, -1, -2, -1, 1, 1, 1, 0, 0, 0, 1, 0, -2, -3, -4, -2, -1, 0, 0, 1, 1, 0, -1, 0, 0, 0, -1, -1, -2, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, -3, -3, -3, -1, 1, 0, 2, 1, 0, -1, 0, -2, -1, -3, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, -2, -3, -2, 0, 0, 1, 1, 0, 0, -2, -1, -2, -1, -2, -2, -1, 1, 1, 1, 2, 3, 0, 0, 0, 0, -1, -4, -4, -3, -1, 1, 1, 0, 1, 0, -1, 0, -1, -2, -2, -1, -1, 0, 1, 1, 0, 2, 1, 2, 0, 0, 0, -2, -3, -2, -2, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -2, -3, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -2, -2, -2, -3, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, -2, -1, 1, 1, 0, 0, 0, -2, -2, -3, -1, -1, 0, 0, 0, 0, 1, 1, 1, 2, 0, 1, 0, 0, -2, -1, 0, -1, 1, 2, 3, 0, 0, 0, -1, -1, -2, -3, -1, -1, 0, 1, 1, 3, 3, 4, 3, 2, 2, 1, 1, 0, 0, 0, 1, 3, 4, 2, 1, 1, 1, 0, -2, -1, -1, 0, 2, 2, 4, 4, 5, 6, 5, 5, 5, 3, 3, 2, 3, 3, 6, 6, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 2, 0, 1, 0, 0, 1, 1, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 0, 2, 0, 0, 1, 2, 1, 2, 2, 2, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 0, 1, 1, 0, 0, 0, 1, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 3, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 2, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 2, 2, 1, 0, 1, 0, 0, 1, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 1, 1, 1, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 1, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 1, 1, -1, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, -1, -1, -1, -1, -1, 1, 1, 0, 1, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 2, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 1, 0, 2, 1, 0, 0, 0, 0, 1, 0, 0, -3, -1, 1, 1, 2, 3, 1, 2, 2, 4, 5, 5, 6, 6, 5, 3, 4, 2, 3, 2, 0, 0, 1, 2, 2, 3, -4, 0, 1, 3, 1, 0, 1, 1, 1, 0, 2, 4, 3, 5, 4, 4, 2, 1, 0, 0, -1, 0, -1, 0, 1, 2, -2, 0, 3, 2, 2, 0, -1, 0, 0, 0, 1, 2, 3, 6, 4, 5, 3, 1, 0, 0, 0, 0, -1, 0, 0, 1, -3, 0, 1, 0, 1, 1, -1, 0, 0, 1, 1, 2, 3, 3, 4, 4, 2, 2, 0, 0, -1, -1, 0, 0, 1, 2, -1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 2, 3, 3, 4, 1, 0, 0, -1, 0, -1, 0, 0, 0, 3, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 2, 0, 0, 0, 0, -1, 0, 0, 1, 2, -2, -2, 0, 0, 0, 0, 1, 1, 0, 0, -2, 0, 0, 1, 0, 1, 2, 0, 1, 0, 0, 0, 0, -1, 0, 1, -2, 0, 0, 0, 1, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, -1, 1, 1, 0, 1, 0, 0, -2, -3, -3, -3, -1, 0, 1, 1, 2, 1, 0, 2, 1, 0, 0, 1, 1, 0, 2, 0, 1, 1, 0, 0, -1, -2, -2, -3, -4, -2, 0, 0, 1, 1, 2, 0, 1, 2, 1, 1, 0, 0, 2, 1, 4, -1, 1, 0, 1, 0, -2, -3, -3, -5, -4, -3, -1, 2, 3, 3, 2, 1, 2, 2, 1, 1, 3, 2, 1, 2, 4, 0, 0, 0, -1, -1, -1, -3, -3, -4, -5, -1, -1, 1, 2, 1, 2, 0, 2, 1, 3, 2, 4, 2, 3, 3, 4, 0, -1, 0, -1, -1, -4, -6, -6, -7, -4, -4, 0, 0, 2, 1, 0, 0, 2, 3, 4, 5, 5, 5, 5, 4, 4, -2, -1, -1, -1, -4, -3, -6, -6, -7, -5, -3, -1, 0, 2, 3, 2, 2, 3, 5, 5, 5, 4, 5, 4, 5, 6, -1, -1, -1, -1, -4, -5, -5, -6, -7, -5, -4, 0, 0, 1, 2, 3, 3, 3, 4, 6, 6, 5, 6, 4, 5, 4, -2, 0, 0, -1, -3, -3, -4, -5, -5, -6, -3, -1, 0, 0, 2, 0, 0, 2, 3, 5, 5, 5, 5, 3, 5, 6, -1, -1, 0, -2, -2, -4, -3, -2, -3, -4, -3, -2, 0, 0, 0, 0, 1, 0, 3, 2, 4, 4, 4, 5, 3, 5, -1, 1, 0, -1, -1, -1, -2, -1, -2, -1, -1, 0, 0, 1, 1, -1, 0, 0, 1, 1, 1, 3, 3, 2, 3, 4, -1, 0, -1, -2, -1, 0, -1, 0, 0, 0, -2, 0, 0, 2, 1, 0, 0, 0, 0, 1, 1, 2, 1, 1, 2, 5, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 2, 1, 2, 1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 4, -2, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 2, 3, 1, 0, 2, 1, 0, 0, 0, 2, 0, 0, 3, 3, -4, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 1, 1, 0, 1, 0, 0, 1, 0, 2, 3, 4, -4, -2, 0, 1, 1, 1, 1, 0, 0, 1, 1, 1, 3, 2, 0, 0, 0, 1, 0, -1, 0, 1, 1, 1, 3, 4, -4, -2, 0, 0, 3, 1, 1, 0, 0, 2, 1, 3, 3, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 3, -4, -2, 0, 2, 2, 2, 1, 1, 1, 3, 2, 4, 4, 3, 2, 0, 2, 0, -1, -1, 0, 0, 1, 3, 3, 6, -5, 0, 1, 0, 0, 1, 1, 1, 3, 3, 4, 5, 3, 4, 1, 1, 2, 1, 1, 0, 0, 0, 1, 3, 3, 5, -5, -3, -3, -1, 0, 0, -1, 0, 0, 0, 0, 2, 1, 3, 3, 4, 3, 3, 4, 5, 3, 4, 4, 5, 6, 7, -4, -3, -2, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 1, 1, 2, 2, 2, 1, 1, 2, 3, 2, 2, 4, 6, -3, -2, -1, 0, -1, 0, -1, -1, 0, -2, 0, -1, 0, 0, 0, 0, 1, 1, 2, 1, 1, 0, 1, 2, 3, 3, -5, -2, 0, 0, -1, -1, 0, 0, -3, -2, -4, -2, -2, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 2, 2, -4, -1, -1, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, -1, 0, 1, 2, 0, 0, 1, 1, -1, 0, 0, 2, 4, -3, -1, 0, 0, 0, 1, 1, 0, 0, -2, -2, 0, 0, -1, -1, 0, 1, 1, 1, 1, 0, 0, 1, 0, 1, 2, -4, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, -2, -1, -2, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 3, -6, -4, -2, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, 0, -2, -1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 1, -5, -3, -1, 0, 0, 0, 0, 1, 0, -1, -1, -1, -2, -3, -3, -3, -2, 0, 0, 1, 1, 0, 0, 0, 0, 1, -5, -3, -2, -1, 0, 1, 0, 0, 0, 0, -1, -2, -2, -2, -3, -2, -1, 0, 1, 2, 0, 1, -1, 0, 0, 0, -3, -3, 0, 0, 1, 0, 0, -1, -1, -1, -1, 0, -2, -1, -2, 0, 0, 0, 2, 3, 2, 0, 0, 0, 1, 1, -2, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 1, 2, 1, 1, 1, 1, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, 0, 1, 2, 2, 3, 1, 0, 0, 1, 1, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -2, -2, 0, 2, 2, 2, 2, 0, 0, 0, 0, 2, -3, -2, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, -2, -1, -3, -2, -1, 2, 2, 2, 1, 1, 0, 0, 0, 1, -4, -3, -1, -2, -1, 0, -1, 0, -1, 0, -1, 0, -1, -3, -1, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -3, -2, -2, -1, -1, 0, 1, -1, -1, -2, 0, -1, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, -4, -2, -2, -1, -2, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 2, -5, -4, -2, -2, -1, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 2, 1, 2, 0, 0, 0, 1, 1, 1, -4, -4, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, -3, -3, -1, -2, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 2, 3, -2, -2, -3, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, -2, 0, -1, -1, -1, -2, 0, -2, -1, -1, 1, 2, 3, -3, -1, 0, 0, -2, -1, -1, -1, -2, -1, -1, -1, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 1, 1, 3, 4, -1, -1, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, -1, 1, 2, 2, 5, 5, -1, 0, 0, 0, 0, 0, -1, -2, -2, 0, -1, 0, 0, 0, 2, 1, 1, 2, 0, 1, 1, 1, 4, 4, 7, 8, -2, 0, 1, 1, 2, 1, 0, 0, 1, 2, 1, 3, 4, 4, 5, 4, 4, 3, 3, 4, 4, 6, 6, 8, 9, 11, 4, 3, 0, 0, 1, 3, 4, 1, 0, 0, 0, -1, -2, -3, -3, -2, -2, 0, -2, -1, -2, 0, 0, 0, 0, -2, 4, 1, 0, 0, 1, 3, 3, 2, 1, 1, 0, 0, -1, -2, -3, -3, -2, -3, -1, -3, -3, -1, -2, 0, 0, 0, 5, 1, 0, 0, 1, 3, 2, 1, 1, 1, 1, 0, -3, -2, -5, -4, -2, -3, -1, -3, -3, -1, -3, -2, -2, 0, 5, 3, 1, 2, 2, 3, 3, 2, 2, 2, 1, 0, -1, -3, -3, -4, -5, -2, -2, -1, -3, -1, -2, -2, -2, 0, 6, 3, 0, 2, 1, 2, 3, 2, 2, 2, 0, -1, -2, -2, -3, -3, -5, -3, -2, -2, -3, -2, -3, -2, -3, -1, 6, 4, 2, 2, 3, 3, 3, 3, 3, 0, 0, -1, -1, 0, -2, -3, -5, -3, -2, -3, -2, -1, -2, -2, -3, -1, 5, 4, 3, 2, 4, 3, 3, 3, 1, 1, 0, 0, 0, 0, 0, -2, -2, -4, -3, -2, -4, -2, -1, -1, -4, -3, 6, 4, 3, 2, 3, 1, 1, 2, 0, 0, 0, -1, 0, 1, 0, -1, -2, -1, -3, -4, -3, -3, -1, -1, -3, -4, 7, 5, 3, 2, 1, 2, 2, 1, 0, -2, -2, 0, 0, -1, 0, 0, -1, -2, -3, -4, -4, -2, -2, -1, -3, -2, 5, 3, 0, 0, 3, 4, 4, 1, 0, -1, -2, -2, -1, 0, 1, 0, 0, -1, -1, -2, -3, -2, -1, -1, -2, -2, 5, 1, -1, -1, 2, 4, 4, 2, 0, 0, -2, -2, 0, 0, 0, 1, 0, 0, -2, -3, -2, -1, -1, -2, -2, -3, 5, 1, -1, 0, 2, 5, 4, 3, 0, 0, -2, -1, 0, 0, 1, 1, 1, 0, 0, -1, -1, -2, -1, -2, -1, -2, 5, 1, 0, -1, 2, 5, 4, 4, 0, 0, -3, -2, -2, 0, 0, 1, 1, 1, -1, -1, -3, -1, -1, -1, -1, -1, 4, 2, 0, -1, 2, 4, 6, 3, 1, -1, -3, -1, 0, 0, 0, 1, 2, 1, -1, -3, -3, -1, 0, -2, -1, -1, 5, 1, -1, 0, 3, 3, 5, 2, -1, -2, -3, -1, 0, 0, 0, 1, 2, 0, 0, -3, -1, -1, -1, -1, -2, -2, 5, 0, 0, 0, 1, 2, 4, 0, 0, -3, -2, -2, -1, 0, 0, 2, 0, 0, -1, -2, -1, -1, -1, -1, -3, -1, 5, 1, 0, 2, 2, 3, 3, 0, -2, -1, -3, -3, 0, 0, 0, 0, 0, -1, 0, -1, -3, 0, -2, -4, -2, -1, 4, 3, 2, 1, 2, 2, 1, 1, -1, -1, -1, -2, -2, 0, -1, 0, 0, -1, -1, -3, -3, -2, 0, -2, -2, -2, 4, 3, 2, 2, 2, 3, 3, 0, 1, 0, 0, -4, -2, 0, -1, -2, 0, -1, -1, -3, -3, -2, -1, -3, -2, -1, 4, 2, 0, 2, 2, 3, 1, 2, 1, 0, -1, -3, -1, -1, -1, -2, -2, -2, -2, -3, -3, -1, -2, -3, -1, -1, 5, 2, 0, 1, 1, 1, 1, 1, 2, 3, 0, -1, -2, 0, -1, -1, -1, -1, -4, -2, -3, -1, -3, -1, -1, -2, 7, 2, -1, 1, 1, 2, 1, 2, 2, 1, 0, -1, 0, 0, 0, -2, -2, 0, -2, -2, -2, -2, -2, -1, -2, 0, 8, 1, 0, 1, 1, 1, 3, 3, 3, 2, 0, 0, 0, -1, -1, 0, -2, -2, -2, -2, -1, -1, -1, -2, 0, 0, 8, 2, 1, 2, 2, 1, 3, 2, 1, 1, 2, 0, -1, 0, -1, -1, -1, 0, 0, -2, -1, -1, 0, -1, -2, 0, 6, 4, 2, 1, 4, 3, 4, 3, 2, 2, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 8, 3, 2, 3, 3, 5, 2, 3, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 2, 1, 0, 0, 0, 1, 2, 0, 0, 2, 1, 2, 0, 0, 0, 0, -1, 0, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 2, 1, 0, 2, 1, 0, 0, 1, 0, 0, -1, 0, -2, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 1, 2, 0, 0, 1, 1, 0, 1, 2, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 3, 1, 1, 2, 1, 2, 1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, -1, -1, -2, 0, -1, 0, 0, 1, 2, 3, 1, 1, 2, 0, 1, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 0, 1, 2, 1, 2, 0, 2, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 2, 0, 2, 1, 0, 1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 2, 0, 0, 0, 0, 2, 0, 0, 0, 2, 2, 0, 0, -1, -1, -1, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, -1, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 1, 2, 0, 0, 0, 1, 2, 2, 2, 1, 2, 0, 0, 0, -1, 0, 1, 1, 0, 0, 1, 2, 0, 0, -1, 0, 2, 1, 1, 0, 2, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 3, 1, 2, 1, 2, 2, 3, 1, 0, 0, 0, 0, 0, -2, 0, 1, 1, 1, 0, 1, 1, 1, 2, 0, 0, 0, 2, 0, 2, 1, 2, 3, 2, 0, 0, 0, -1, 0, -2, -1, -1, 0, 0, 0, 1, 2, 2, 1, 1, 0, 1, 1, 0, 1, 1, 3, 3, 2, 2, 3, 1, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 1, 0, 2, 3, 2, 5, 3, 3, 2, 2, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 2, 3, 2, 3, 3, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 1, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, -1, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, -1, 1, 0, 1, 1, 1, 1, 2, 2, 3, 3, 2, 2, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, -1, 0, -1, 0, 1, 1, 2, 0, 1, 1, 1, 1, 2, 2, 2, 1, 2, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 1, 2, 0, 2, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, -1, 0, 0, -2, -2, -1, -2, -1, -3, 0, -2, 0, 0, 0, -1, -2, -1, -2, -1, -1, 0, 0, 0, 0, 0, 1, 2, 0, 1, 1, 2, 2, 2, 1, -3, -1, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 1, 1, 2, 0, 1, 0, 1, 2, 0, 0, 1, 0, 1, 0, -1, -1, 0, -2, -2, 0, 0, -2, 0, -1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 1, 0, 0, 0, -2, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -2, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, -2, -1, -1, 2, 1, 2, 1, 2, 1, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, -2, 0, 0, -1, 0, 0, -2, -1, 0, 0, 1, 2, 1, 2, 2, 0, 0, 0, -1, -1, 0, 0, -2, -2, -1, -1, -1, -2, -1, -1, 0, 0, -1, -1, 0, 0, 0, 3, 1, 2, 3, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -3, -2, -1, 0, 1, 0, 2, 3, 2, 3, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -2, 0, 0, 0, -2, -1, 0, -1, 0, 2, 0, 1, 1, 3, 3, 1, 1, 2, 1, 0, 1, 0, 0, -1, -2, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 2, 0, 2, 2, 3, 3, 3, 1, 2, 2, 1, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, -2, 0, 0, -1, 0, 1, 0, 2, 3, 3, 2, 1, 3, 1, 2, 1, 0, 0, -1, -2, 0, -1, -1, 0, 0, 0, -3, -2, -1, 0, 0, 0, 0, 2, 2, 2, 2, 3, 2, 1, 1, 2, 1, -1, -2, -2, -1, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 2, 2, 1, 2, 2, 3, 2, 1, 0, 0, 0, -2, -1, -2, -1, 0, 0, 1, -2, 0, -2, 0, 1, 0, 1, 2, 1, 1, 2, 1, 1, 0, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, -2, 0, 0, 1, 0, 2, 0, 0, 0, 0, 1, 2, 3, 0, 0, 0, -1, 0, -1, 0, 1, 0, 1, 0, -2, -1, 0, 0, 1, 0, 2, 2, 2, 2, 2, 0, 1, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -4, -1, -2, -1, 0, 1, 2, 3, 2, 1, 1, 0, 0, 0, 2, 0, 1, 1, 0, 0, 1, 1, -1, 0, 0, 1, -2, -3, 0, -1, 0, 2, 3, 3, 4, 3, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, -2, -3, 0, 0, 0, 2, 1, 4, 2, 2, 0, 0, 1, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, -2, -3, -1, 0, 0, 2, 3, 2, 3, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, -2, -3, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, -1, 0, 0, 0, 1, 2, 1, 1, 2, -2, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -2, 0, -2, -1, 0, 0, 0, 0, 0, 1, 0, 2, 1, 2, -1, -2, -1, 1, 2, 0, 0, -2, -2, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 2, 2, -1, -2, 0, 0, 0, 0, -1, 0, 0, -2, -1, -2, -1, 0, 0, 0, 0, 1, 1, 2, 2, 1, 2, 2, 3, 1, -3, -2, -2, -2, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 1, 3, 3, 2, 4, 4, 3, 4, 2, 2, 2, 0, 0, -3, -4, -2, -2, 0, 3, 5, 5, 6, 6, 7, 4, 3, 2, 2, 1, 0, 0, 1, 1, 0, 0, 1, 1, 0, -2, -2, -2, -2, 0, 0, 1, 3, 4, 4, 5, 2, 1, 2, 0, 1, 1, 0, 0, 0, 0, 0, -1, 2, 1, 0, -1, -2, -2, -2, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -1, 2, 1, 0, -1, -3, -2, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, 0, 0, 3, 0, 0, -1, -1, -2, -1, -2, -1, -2, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, -1, -1, -1, 3, 2, 2, -1, -1, -2, -3, -3, -3, -1, -1, -1, -2, 0, -1, 1, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 3, 0, 1, 0, 0, -1, 0, -2, -1, -1, 0, -1, 0, -2, -1, -1, 0, 1, 2, 0, 2, 0, 1, 0, 0, -1, 2, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, -1, -1, -4, -3, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, -2, 1, 1, 1, 2, 1, 2, 1, 3, 3, 2, 1, 0, -4, -4, -4, -4, -2, 0, 1, 1, -1, -1, -2, -1, -3, 0, 1, 0, 1, 2, 0, 0, 1, 2, 3, 5, 2, 0, -3, -6, -6, -5, -3, 0, 0, 1, 0, -2, 0, -3, -3, -2, 0, 0, 0, 2, 0, 0, 0, 0, 2, 3, 1, 0, -3, -7, -6, -6, -1, 0, 2, 2, 0, 0, -2, -3, -4, -4, -3, -2, 0, 1, 0, 0, 0, 0, 2, 2, 1, -1, -3, -6, -8, -5, -1, 3, 4, 3, 0, 0, -1, -4, -4, -4, -2, -3, 0, 0, 0, 0, 0, 1, 3, 4, 2, 0, -3, -4, -7, -4, 0, 3, 5, 4, 1, 0, -2, -2, -4, -4, -2, -1, -1, 1, 1, 0, 1, 2, 2, 4, 2, 0, -3, -5, -7, -4, -1, 3, 6, 4, 3, 0, -1, -3, -3, -4, -1, -1, 0, 2, 0, 0, 1, 1, 3, 3, 3, 0, -3, -6, -6, -5, -1, 3, 4, 3, 2, 0, -1, -2, -4, -3, 0, 0, 0, 1, 2, 2, 1, 1, 3, 2, 2, 0, -3, -6, -7, -3, -1, 0, 3, 2, 0, 0, -2, -4, -2, -3, 0, 0, 0, 2, 1, 1, 1, 2, 1, 0, 0, -2, -3, -7, -7, -5, 0, 0, 1, 2, 0, 0, -3, -2, -2, -3, 0, 0, 0, 1, 1, 2, 1, 1, 1, 0, -1, -1, -4, -4, -6, -3, -1, 1, 1, 2, 0, 0, 0, -1, -2, -3, 0, 0, 2, 0, 2, 2, 2, 0, 0, 0, 0, -2, -3, -5, -3, -2, -1, 0, 1, 2, 2, 0, -1, -2, -2, -3, 2, 0, 1, 1, 1, 2, 2, 0, -2, -1, -1, -1, -3, -4, -2, 0, 0, 1, 2, 2, 1, 0, 0, -1, 0, -2, 3, 0, 1, 0, 0, 0, 0, -1, -1, -1, -2, -2, -4, -3, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -3, 2, 0, 0, 0, 0, -1, 0, -1, -2, 0, -1, -2, -3, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, 1, 0, 0, 0, -2, -3, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, -2, -2, 0, 0, -1, -1, -2, 2, 0, 0, 0, -2, -1, -3, -1, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, -3, -2, -2, -1, -2, -1, -3, 2, 2, 1, -1, -3, -3, -2, -1, 0, 1, 0, 3, 4, 4, 5, 2, 1, 0, 0, -2, -2, -1, -2, -1, -3, -2, 6, 2, 3, 1, 0, 0, -2, -2, 0, 0, 4, 5, 6, 7, 6, 5, 4, 3, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 1, 1, -1, 0, 1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, -1, -2, -2, -3, -2, -3, -1, 0, 0, 0, 2, 1, 2, 2, 2, 1, 1, 0, 0, 2, 0, 1, 3, 4, 2, 1, -2, -1, -2, 0, 0, -1, -2, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 2, 1, 2, 1, -1, -2, 0, -2, -2, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -3, -1, 0, -1, 1, 1, 0, 2, 3, 2, 2, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -4, -1, 0, 0, 1, 2, 2, 1, 3, 2, 2, 1, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -3, -2, -2, 1, 1, 2, 2, 4, 2, 3, 4, 3, 1, 0, -1, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, -3, -3, 0, 0, 0, 1, 1, 1, 2, 4, 3, 1, 0, -1, -1, -1, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, -4, -4, 0, 0, 1, 0, 0, 1, 2, 2, 2, 2, 0, 0, -2, -1, -2, 0, 0, 0, 0, -1, 0, -1, -1, -2, -3, -4, -1, 0, 0, 1, 0, 1, 2, 3, 2, 2, 0, -1, -2, -3, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -3, -4, 0, 1, 0, 0, 1, 0, 1, 4, 3, 1, 0, -1, -2, -3, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, -3, -3, 0, 0, 2, 0, 1, 2, 3, 3, 2, 3, 0, 0, -1, -2, -2, 0, 0, 0, -1, -2, 0, 0, -2, -1, -2, 0, 0, 1, 1, 2, 2, 3, 3, 4, 2, 1, 0, 0, -2, -1, -2, -1, 1, 0, -1, -1, -2, -2, -1, -1, -2, -2, 0, 1, 3, 1, 2, 2, 3, 2, 3, 2, 1, 0, -2, -2, -1, -1, 0, 0, -1, -2, -2, -1, -1, -1, -3, 0, 0, 1, 2, 2, 2, 4, 3, 2, 1, 1, 0, 0, -1, -2, -1, -1, -1, -1, 0, -2, -2, -2, -2, -1, -2, -1, -1, 0, 1, 2, 4, 2, 3, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -2, 1, 1, 3, 3, 4, 2, 2, 0, 1, 0, -1, -2, -2, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, -1, -3, -2, 0, 2, 1, 4, 3, 4, 2, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -2, -2, 0, -2, -1, 0, 1, 1, 2, 1, 1, 2, 1, 1, 0, -1, -1, -2, -2, 0, -1, -1, 0, -2, 0, -2, 0, 0, 0, -1, 0, -1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, -2, -1, -1, -2, -1, -2, -2, -2, -2, -1, -1, 0, -1, -3, -1, 0, 0, 0, -1, -1, -1, -1, 1, -1, -1, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, 0, -1, -2, -2, 0, 0, 0, -2, 0, -2, -2, -2, -2, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, -2, 0, -2, -1, -1, 0, -1, 0, -1, -1, -2, -2, -2, -3, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, -1, -1, -2, 0, -2, -2, -2, -2, -2, -2, -2, -1, 1, 1, 2, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, -6, -4, -1, -2, -2, 0, -1, 0, -1, -1, 0, 2, 3, 3, 2, 2, 3, 3, 3, 3, 1, 2, 0, 1, 2, 5, -6, -3, 0, 0, 0, 0, -1, -1, -2, -1, 0, 2, 2, 3, 1, 3, 2, 0, 1, 1, 0, 0, 0, 1, 1, 3, -3, -1, 2, 1, 0, 0, -1, -2, -1, -2, 0, 2, 2, 2, 4, 2, 0, 1, 0, 0, 0, -2, -1, 0, 2, 2, -3, 0, 1, 2, 2, 1, -1, -2, 0, -2, -1, 0, 2, 4, 3, 2, 1, -1, -1, -2, -2, -1, -1, 0, 1, 2, -4, -1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, -2, -1, -2, -2, -1, 0, -1, 2, 2, -6, -2, 0, 1, 1, 0, 2, 0, 2, 1, 0, 1, 1, 1, 1, -2, -1, -1, -3, -2, -3, -2, -1, -1, 0, 2, -5, -2, -1, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, -1, -1, -3, -3, -2, -3, -4, -3, -2, 0, 1, -6, -3, -1, 0, 0, 0, 1, 3, 2, 2, 0, 0, 0, -1, -1, 0, -1, -2, -2, -2, -1, -2, -1, 0, -1, 0, -3, -3, -1, 0, 0, 0, 0, 0, 2, 1, 2, 3, 2, 2, 1, 0, 0, 0, 0, -1, -3, -2, -2, 0, 1, 0, -4, -1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 3, 5, 5, 4, 2, 1, 0, -2, -2, -2, -1, 0, 0, 1, 2, -4, 0, 0, -1, 0, -2, 0, -1, 0, 2, 1, 5, 6, 4, 4, 2, 1, -2, -1, 0, -1, -1, 0, 1, 2, 2, -2, 0, 0, -1, -1, -2, -1, 0, -1, 0, 3, 5, 6, 5, 5, 2, 0, -2, -1, -2, -2, 0, 1, 1, 3, 3, -2, -1, -1, -2, -1, -3, -3, -1, 0, 0, 1, 3, 5, 4, 5, 3, 0, -2, -3, -2, 0, -1, 2, 1, 1, 4, -4, -2, 0, 0, -2, -1, -3, -1, 0, 1, 1, 4, 5, 5, 5, 2, 1, 0, -3, -3, -2, 0, 1, 1, 3, 4, -3, -2, 0, -1, -2, 0, -2, -1, -2, 0, 2, 3, 4, 4, 4, 4, 2, 0, -1, -3, 0, 0, 1, 4, 4, 4, -4, -2, -1, -1, -1, -1, 0, 0, -1, 0, 1, 2, 2, 3, 4, 2, 2, 1, -1, 0, 1, 1, 3, 4, 4, 4, -5, -3, -1, -2, -2, 0, 0, 1, 0, 0, 2, 3, 3, 3, 3, 3, 1, 0, 1, 0, 2, 1, 2, 3, 3, 5, -5, -3, -2, -1, -1, 0, 1, 1, 3, 1, 1, 0, 3, 2, 2, 1, 0, 0, 0, 0, 1, 2, 0, 1, 2, 4, -6, -3, -3, -1, 0, 2, 1, 3, 3, 3, 3, 2, 2, 0, 1, 0, -1, -2, -2, 0, -1, 0, 0, 0, 2, 3, -5, -3, -1, -1, 1, 0, 1, 3, 2, 2, 2, 1, 2, 0, 0, 0, 0, -2, -1, -2, -2, 0, 0, 1, 0, 2, -4, -3, 0, 0, 0, 1, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, -2, -2, -2, -1, -1, 0, 1, 0, 2, -6, -3, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 2, -5, -4, 0, 0, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 1, 3, 2, -7, -3, -1, 1, 2, 1, -1, -3, -2, 0, 0, 2, 2, 2, 0, 1, 1, 1, 1, 1, 0, 0, 2, 3, 1, 2, -7, -4, -2, 1, 1, 0, 0, -2, 0, 0, 1, 2, 3, 2, 1, 1, 3, 2, 2, 3, 1, 3, 3, 4, 3, 2, -5, -3, -1, 0, 0, 0, 0, 0, -2, 0, 1, 3, 2, 3, 3, 3, 2, 1, 3, 3, 3, 5, 5, 5, 5, 3, -4, -1, -1, 0, 0, -1, 0, 1, 1, 2, 2, 2, 4, 3, 3, 2, 2, 1, 2, 3, 1, 2, 2, 3, 3, 6, -3, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 2, 0, 1, 1, 2, 0, 0, 0, 0, 1, 0, 1, 3, 3, -2, -2, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, 0, -1, 0, 1, 0, 1, 3, 2, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 3, -3, -2, -1, 0, 0, 0, 1, 0, -1, -2, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 2, -3, -1, 0, 0, 1, 0, 1, 0, -1, -1, -2, -1, -1, -1, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 1, -2, 0, 0, 0, 1, 1, 1, 1, 0, 0, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 1, -4, -1, 1, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -2, -1, -1, -1, -1, 0, 0, -2, 0, 0, 0, 0, 0, -3, -1, 0, 1, 0, 0, 1, 0, 0, -1, -2, -1, -1, -2, -2, -2, -1, 0, 1, 0, -1, -1, -1, 0, 0, 1, -3, -1, 0, 0, 0, 1, 0, 1, 0, 0, -1, -2, -2, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 1, 1, -1, -1, 0, 1, 0, -1, 0, 1, 0, -1, -1, -1, -2, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 1, 1, -3, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -1, 0, 0, 1, 2, 1, 2, 2, 0, 0, -1, -1, 0, 1, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 2, 3, 3, 2, 2, 0, 0, 0, 0, 0, 2, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 2, 1, 2, 4, 0, 0, 0, 0, -1, 0, 2, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 1, 1, 3, 2, 0, 0, 0, 0, -1, 0, -2, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 1, 1, 1, 2, 1, 0, 0, -1, -1, -1, 1, -2, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, -1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -2, -1, 0, 0, 1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -1, 0, 1, -2, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 3, -3, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, -1, 0, 0, -1, -1, -1, 1, 3, -1, -1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, -1, -1, -1, 0, 0, 1, -2, -1, -1, -1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -2, 0, 0, 0, 2, 2, -3, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 2, 3, 4, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 1, 2, 4, 5, -1, -1, 0, 1, 0, 1, 0, 0, 1, 1, 2, 2, 3, 2, 2, 2, 1, 1, 2, 1, 1, 3, 2, 4, 4, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 2, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, -1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 1, 0, -1, -1, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, 1, 0, 1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -3, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 1, 1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 1, -1, -2, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 1, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, -1, 0, 1, 0, 0, -1, -1, -2, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -2, -2, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, -1, -2, -1, -1, -1, -2, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, -1, -1, 1, 1, 1, 0, -1, -1, -2, 0, -1, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 1, 1, 0, 0, 0, 0, -1, -2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -2, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 1, 0, 0, 1, 0, 0, 0, -1, 2, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 2, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 2, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 0, 0, 0, 0, -1, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 2, 0, 2, 0, 0, 0, 0, 1, 0, 0, -1, -2, -1, -1, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, 1, 2, 1, 2, 0, 0, 0, -1, -1, 0, -2, -2, -2, -2, 3, 1, 1, 1, 0, -1, 0, 0, -1, 0, 0, 2, 1, 2, 2, 5, 3, 4, 2, 2, 1, 1, 2, 1, 1, 3, 4, 3, 0, -1, -2, 0, -2, -2, -2, -1, 0, 0, 2, 1, 1, 3, 1, 1, 0, 2, 0, 1, 2, 2, 1, 1, 4, 2, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 2, 1, 2, 0, 2, 3, 4, 0, -1, -2, -1, -2, -3, -1, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 1, 1, 0, 0, 1, 3, 0, 0, 0, -1, -2, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 1, 1, 0, 0, 2, 2, 0, -1, 0, 0, 0, -1, -2, -1, -2, -1, -2, 0, 0, 0, 0, 0, 1, 2, 1, 3, 1, 0, 0, 0, 2, 2, 1, -1, 0, 0, 0, 0, -2, -1, -3, -2, -2, 0, -1, 0, 0, 0, 0, 1, 1, 0, 2, 0, 0, 0, 1, 2, 0, 1, 0, 0, -1, -1, -1, -2, -1, -3, -1, 0, -1, 0, -2, 0, 0, 0, 1, 0, 1, 1, 0, 0, 2, 3, 2, 0, 0, -1, 0, 0, -1, -1, -2, -2, -1, 0, 0, -1, -2, -1, -1, 0, 1, 0, 1, 0, 0, 0, 0, 3, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -4, -3, -2, 0, 0, 1, 2, 0, 0, 0, 0, 3, 0, 0, -1, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, -4, -3, -2, -2, 1, 2, 2, 2, 2, 1, 1, 1, 2, 0, -2, -2, -1, 1, 0, 0, -1, -1, 0, 0, -2, -3, -4, -4, -2, 0, 2, 2, 3, 3, 1, 0, 1, 0, 1, 0, -2, -2, 0, 0, 0, 0, -1, -3, -1, -1, -2, -2, -2, -2, -2, 0, 2, 2, 6, 5, 3, 0, 0, 0, 2, 0, -3, -2, -2, -1, 0, 0, 0, -2, 0, 0, -1, -3, -3, -2, -2, 0, 2, 5, 5, 3, 4, 2, 1, 1, 0, 0, -3, -2, -1, -1, 0, 0, -1, -2, -1, 0, -2, -2, -4, -3, -2, 0, 2, 3, 4, 5, 2, 1, 1, 0, 2, 0, -1, -1, -1, 0, 1, 0, -2, -1, 0, -1, -1, -2, -4, -3, -2, 0, 2, 3, 2, 3, 2, 1, 0, 0, 1, 0, -1, -2, -1, -1, 0, -1, 0, -1, -1, 0, -2, -2, -2, -4, -2, -1, 0, 2, 2, 0, 1, 0, 0, 0, 2, 0, -1, -2, 0, -1, 0, -1, -2, -1, -1, -1, 0, -1, -3, -2, -1, -1, 0, 2, 1, 2, 1, 1, -1, 0, 3, 0, -2, -2, 0, 0, 0, -1, 0, -2, -1, -1, 0, -1, -1, -2, -1, 0, 1, 2, 2, 3, 1, 0, 1, 1, 3, 0, -2, -2, -1, 0, -1, 0, -1, -1, -1, -2, -1, -1, -1, -1, -1, 0, 2, 2, 2, 3, 2, 1, 0, 0, 2, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, -1, -2, -2, -1, 0, -1, 1, 1, 3, 2, 1, 0, 1, 2, 1, 2, 0, -1, -3, -1, -2, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 2, 2, 0, -2, -2, -3, -2, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 2, 2, 0, 0, -2, 0, -1, -2, 0, 0, 0, 1, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 4, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 2, 4, 1, 0, 0, 0, -1, -2, 0, 0, -1, 0, 0, 0, 0, 1, 2, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 3, 4, 3, 2, 3, 2, 1, -1, -1, -3, -1, -1, -3, -2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 3, 1, 3, 3, 2, 1, 0, 1, -1, -2, -3, -3, -4, -3, -1, 0, 0, 0, -2, -1, -1, 0, -2, 0, 0, 1, 0, 2, 2, 1, 2, 1, 1, 0, -1, -1, -2, -2, -2, -3, -2, 2, 0, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, -1, -1, 0, 0, 0, -3, -2, 1, 1, 0, -1, -1, -2, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -3, -2, -3, -3, -3, -4, -4, -3, -3, -2, 0, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, -1, 4, 0, 0, 0, -1, -2, -2, -4, -3, -4, -4, -4, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 3, 2, 2, 0, -1, -1, -1, -4, -3, -5, -5, -3, -3, -2, -1, 0, 1, 0, 0, 0, 0, 2, 0, 1, 0, 0, 2, 2, 0, 2, 0, -2, -3, -1, -2, -3, -4, -5, -3, -3, -1, -2, 0, 1, 2, 2, 1, 0, 1, 0, 0, 0, 3, 2, 1, 1, 0, -1, 0, -1, -3, -4, -4, -5, -5, -3, -3, -1, 0, 1, 1, 3, 1, 1, 0, 1, 1, 0, 2, 1, 0, 0, 0, -2, -1, -1, -1, -2, -3, -4, -6, -4, -3, -2, 0, 2, 4, 3, 3, 3, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, -3, -3, -3, -3, -5, -5, -4, -5, -4, -2, 0, 3, 4, 5, 4, 3, 1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -3, -3, -2, -4, -3, -3, -4, -4, -2, -2, 0, 4, 6, 6, 5, 2, 2, 2, 0, 0, -1, -1, 0, -2, -2, -2, -2, -4, -4, -3, -3, -5, -3, -5, -2, -2, 0, 3, 7, 5, 4, 3, 3, 2, 0, 0, 0, 0, 0, -1, -2, -3, -3, -3, -4, -3, -4, -3, -4, -4, -4, -1, 0, 4, 5, 5, 6, 3, 3, 0, 0, -1, 0, 1, 0, -1, 0, -3, -2, -2, -3, -4, -5, -4, -5, -6, -4, -2, 0, 1, 4, 5, 5, 2, 3, 1, 0, 0, 1, 0, 1, 0, -2, -1, -1, -2, -3, -3, -5, -4, -6, -4, -5, -3, -2, 0, 3, 2, 3, 3, 1, 1, 0, 0, 2, 1, 1, 0, 0, -1, 0, -2, -2, -4, -5, -6, -4, -5, -4, -2, -1, 1, 1, 2, 2, 2, 0, 2, 0, 0, 1, 1, 1, 0, 0, -1, -1, -1, -3, -3, -5, -3, -4, -3, -3, -1, -1, 1, 1, 3, 2, 1, 2, 0, 0, 0, 1, 1, 0, -1, 0, -1, -1, -1, -3, -4, -3, -3, -3, -2, -1, 0, 0, 0, 1, 4, 3, 1, 2, 1, 0, 0, 0, 0, 0, 0, -2, 0, -2, 0, -2, -4, -4, -3, -3, -1, 0, 0, 1, 2, 2, 3, 2, 3, 3, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, -2, -3, 0, -2, -1, 0, 2, 0, 1, 2, 2, 1, 1, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 2, 1, 2, 2, 1, 0, 1, 0, 0, 0, 0, 0, 2, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, -1, 0, -1, -1, -2, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 3, 3, 2, 0, 1, 0, 0, -1, -2, 0, -1, -1, -2, 0, 1, 2, 0, 1, 1, 0, 0, 0, 3, 2, 3, 4, 4, 4, 3, 3, 2, 1, 0, 0, 0, -1, -1, -1, -2, 0, 2, 1, 1, 0, 1, 1, 1, 0, 0, 0, 1, 2, 1, 1, 0, 1, 1, 1, -1, -1, -3, -3, -3, -3, -5, -4, 2, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 2, 0, 1, 0, -1, -1, 0, 0, 0, -1, -2, -3, -3, -3, -5, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, -3, -3, -4, 2, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, -2, -2, -2, -3, 2, 0, -2, 0, 0, -2, -1, -2, -1, -1, 0, -2, 0, -2, 0, -1, -1, -1, 1, 0, 0, 0, 0, -2, -3, -2, 0, 0, -1, 0, -1, -1, -2, 0, -3, -3, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -3, 2, 0, 1, 0, 0, 0, 0, -1, -2, -3, -3, -3, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -2, -1, 3, 3, 1, 0, 0, 0, 0, 0, -2, -2, -2, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 4, 3, 1, 1, 0, 0, -1, 0, -1, 0, -3, -2, -2, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 4, 2, 2, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, -3, -2, -2, 0, 0, 0, 0, 0, 0, 0, -2, 3, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, -1, -1, -1, -3, -2, 0, 0, 0, 0, 0, -1, -2, -1, 2, 0, 0, 0, 2, 0, 0, 1, 1, 1, 2, 0, 0, -1, -2, -2, -3, -2, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 0, -1, -2, -2, -1, -2, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, -1, -1, -2, -3, -1, 0, 1, 0, 1, 0, -1, -2, -2, 2, 1, -1, 0, 0, 1, 1, 0, 0, 2, 2, 1, 0, -1, -2, -2, -2, -1, -1, 0, 0, 1, 0, 0, 0, -1, 3, 1, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, -3, -3, -1, -3, 0, -1, 0, 0, 0, 0, 0, 0, 0, 3, 1, 1, 0, 0, 0, -2, -1, -2, 0, 0, 0, -1, -1, -2, -3, -3, -2, 0, 0, 0, -1, 0, 0, 0, 0, 5, 1, 0, 1, -1, -1, -3, -2, -3, 0, 0, -1, 0, -1, -2, -3, -2, -1, -2, -1, 0, 0, 0, 0, 0, -2, 6, 2, 2, 0, 0, -2, -1, -2, -1, 0, -1, 0, -1, -2, -1, -2, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 5, 4, 2, 0, -1, -2, -1, -2, -3, -2, -2, -2, -3, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 3, 1, 1, 0, -1, -3, -2, -2, -2, -1, -1, -2, -1, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, -1, 6, 2, 1, 0, 0, 0, 0, -3, 0, -1, -1, -2, -2, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 5, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -2, 0, -1, -1, -1, 0, 0, 0, -1, -1, 0, -1, -1, -3, -2, 4, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, -2, -1, -3, -4, 4, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, -2, -2, -3, -4, -4, 4, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, -1, -1, -2, -3, -3, -3, -5, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, -1, -1, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, -1, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, -1, 0, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 1, 0, -1, 0, 0, -1, -1, -2, -1, -1, -3, -2, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, -1, 0, 0, 0, -1, -3, -2, -2, -3, -1, -2, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -2, -3, -2, -1, -3, -2, 0, -1, -2, -1, 0, 0, -2, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 1, -1, -2, -2, -2, -2, 0, -1, -2, -2, -2, 0, 0, 0, -2, 0, -1, 0, 0, 0, -1, 0, 0, 2, 0, 2, 2, 0, 0, -1, -1, 0, -1, -1, -2, -1, 0, -2, -1, 0, 0, 0, 0, 0, -2, 0, 0, 0, 1, 0, 2, 2, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, 0, 0, -1, -1, -1, -1, -2, -1, -2, -1, 0, 1, 1, 0, 2, 2, 2, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, -1, -1, -1, -2, -2, 0, 0, -2, 0, -1, 1, 3, 2, 1, 1, 0, 0, -1, 0, 0, -2, -2, 0, -2, -1, -1, 0, 0, -2, -2, -1, -2, -1, 0, 0, 0, 2, 2, 1, 2, 1, 0, 0, 1, -1, -1, 0, -1, 0, -2, -2, -2, -1, 0, -2, 0, 0, -2, -1, -2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, -1, 0, 0, -1, -1, -2, -2, 0, 0, 0, 0, 0, 2, 2, 1, 2, 0, 1, 0, 0, 0, -1, -1, 0, -1, -1, -1, -2, 0, 0, 0, -2, -1, 0, 0, 0, 1, 1, 1, 1, 2, 1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 2, 0, 0, 0, 0, -1, 0, -1, -1, -2, 0, -1, -2, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 2, 2, 1, 0, 0, -1, 0, 0, -2, -1, -1, -1, 0, 0, 0, -2, -1, -2, 0, 0, -1, 0, -2, 0, 0, 0, 2, 2, 0, 1, 0, 0, -2, -2, -2, -2, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 1, 3, 3, 2, 0, 0, -1, -2, -2, 0, -1, -1, -1, -1, 0, -1, -1, -1, -1, -1, -2, -1, 0, 0, 1, 0, 2, 3, 2, 0, 0, 0, -2, -2, 0, -2, 0, -2, -2, -1, -1, 0, 0, -1, 0, 0, -1, -2, 0, 0, 1, 0, 1, 2, 0, 1, 0, 0, 0, -1, -2, 0, -2, 0, -2, -1, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -2, -1, -3, -1, -2, 0, 0, -1, -2, 0, -1, -1, 0, -1, -1, -1, -1, 1, 0, 0, 0, 0, -1, 0, -1, 0, -2, -1, -1, -2, 0, -1, -1, 0, 0, 0, -1, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, -3, -2, -2, 0, 0, -1, 0, 0, 0, 1, 1, 2, 2, 0, 2, 2, 1, 0, 0, 1, 0, 1, 1, 2, 2, 1, 1, 0, 2, 2, 0, 0, -1, -2, -2, -3, -5, -6, -7, -8, -8, 1, 2, 0, 0, 0, 0, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, -3, -2, -4, -5, -5, -6, -6, -9, 0, 1, 1, 0, -1, 0, 0, 1, 1, 1, 2, 1, 0, -1, -2, 0, -3, -3, -3, -2, -2, -3, -5, -5, -5, -7, 1, 0, 1, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, -1, -2, -3, -5, -3, -4, -2, -3, -3, -2, -4, -6, -7, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -3, -4, -3, -3, -6, -4, -3, -1, -1, -4, -3, -6, -5, 3, 1, 1, 0, 0, 0, -1, 0, 0, -2, -3, -3, -4, -5, -3, -4, -4, -5, -3, -2, -2, -3, -2, -2, -4, -5, 3, 3, 0, 0, 0, 1, 0, -1, -1, -3, -4, -3, -5, -3, -4, -3, -4, -3, -2, -3, -2, -1, -2, -1, -3, -5, 1, 2, 1, 1, 0, 0, 0, -2, -2, -1, -4, -2, -4, -3, -2, -4, -3, -3, -4, -2, -2, -3, -2, -3, -4, -5, 1, 2, 3, 2, 0, 0, -1, -1, -3, -2, -1, -3, -1, -2, -3, -1, -2, -2, -3, -2, -2, -1, -2, -2, -3, -3, 1, 2, 1, 2, 0, 0, -2, 0, -1, -1, -1, -2, -1, -2, -1, -2, -3, -4, -3, -2, -2, 0, -1, 0, -2, -3, 2, 2, 1, 1, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -3, -3, -3, -5, -5, -2, -1, -1, -1, 0, -3, -2, 2, 1, 1, 0, -1, -1, -2, -1, 0, 0, 0, 0, -1, -3, -3, -3, -2, -5, -3, -2, -1, -2, -2, 0, -3, -4, 0, 0, 1, 0, -1, -1, 0, 1, 0, 0, 1, 0, -1, -2, -3, -3, -3, -4, -2, -2, -2, -1, -1, -2, -1, -2, 0, 0, 1, 1, 0, 0, -1, 1, 1, 0, 1, 1, 0, 0, -2, -3, -4, -3, -3, -2, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 0, 0, 0, -2, -4, -3, -3, -3, -2, -2, 0, 0, -2, -2, -3, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, -1, -1, -2, -4, -4, -1, -3, -2, -1, -2, -1, -2, -2, -2, 1, 0, 0, 1, 0, 0, -1, -1, -1, -2, -1, -1, -1, -2, -2, -3, -4, -4, -2, -3, -2, -2, -3, -2, -3, -4, 1, 0, 0, 0, 1, 1, 0, -1, -2, -3, -3, -3, -4, -3, -3, -3, -4, -3, -5, -4, -3, -3, -2, -4, -3, -4, 0, 2, 0, 2, 0, 0, 1, -2, -3, -3, -4, -4, -4, -2, -3, -3, -3, -5, -3, -4, -3, -2, -3, -4, -4, -4, 0, 1, 2, 2, 0, 0, 0, -2, -2, -3, -3, -3, -2, -3, -3, -3, -4, -4, -4, -3, -3, -4, -3, -3, -4, -3, 0, 2, 1, 2, 0, 0, 0, -2, -2, -1, -1, -1, -2, -3, -3, -3, -4, -3, -2, -3, -2, -2, -1, -4, -3, -4, 1, 2, 2, 1, 1, 0, 0, 0, -1, -2, 0, -3, -2, -2, -3, -1, -3, -1, -1, -2, -2, -3, -3, -2, -3, -4, 0, 2, 1, 0, 0, -1, -1, -2, -1, -1, 0, -1, -1, 0, -1, -1, -1, -2, -1, -3, -2, -4, -2, -4, -6, -5, 1, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -2, -2, -1, -1, -2, -4, -5, -3, -3, -6, -5, 2, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, -1, -1, -2, -1, -2, -2, -1, -2, -2, -4, -6, -6, -6, -5, 1, 0, -1, -1, -3, 0, -2, -1, 0, 1, -1, 0, 0, -1, -1, -2, -3, -3, -2, -3, -4, -5, -5, -5, -6, -8, 3, 0, -1, -2, -3, -4, -3, -3, -2, -2, -2, 0, 0, 2, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -3, -1, -2, 0, -1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, -1, 0, 0, 1, 0, 0, -1, -2, -1, -2, -3, -1, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, -1, -3, -2, -2, -1, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, -1, -1, 0, -2, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 2, 0, 0, -1, 0, 1, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 2, 1, 3, 3, 3, 4, 2, 0, 0, -1, 0, -2, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, -1, -1, 1, 0, 2, 1, 2, 2, 3, 2, 2, 0, -1, -1, -2, -1, -2, -1, 0, -1, -1, 0, 0, 0, 0, -1, -2, -1, 0, 1, 3, 2, 1, 1, 3, 3, 2, 1, -1, -3, -2, -2, -2, -1, 0, 0, 0, 0, 0, -1, 0, -2, -2, -2, 0, 0, 1, 2, 0, 2, 2, 1, 0, 0, -1, -4, -3, -2, -2, 0, 0, 0, 1, 0, -1, -1, -1, -4, -3, -3, 0, 2, 2, 1, 1, 0, 0, 2, 1, 0, -3, -3, -3, -2, -2, 0, 2, 1, 1, 0, 0, 0, -2, -3, -3, -1, 0, 1, 3, 0, 1, 2, 2, 2, 0, 0, -2, -4, -3, -4, -2, 1, 2, 1, 0, 0, 0, -2, -2, -1, -3, -2, 0, 3, 3, 2, 2, 2, 2, 2, 1, -1, -1, -4, -4, -4, -2, 0, 1, 1, 0, 0, -1, 0, -3, 0, -2, 0, 1, 3, 2, 3, 2, 1, 3, 2, 2, 0, -1, -4, -3, -4, -2, 0, 0, 0, 0, 0, -2, 0, -3, 0, 0, -1, 0, 3, 3, 3, 2, 2, 1, 3, 1, 0, -2, -2, -3, -4, -2, 0, 0, -1, 0, 0, -1, -2, -3, 0, -1, 0, 0, 2, 2, 2, 3, 3, 2, 1, 0, 0, -1, -2, -2, -3, 0, 0, 0, 0, -1, -2, -1, -2, -1, 1, -1, -1, 1, 1, 1, 2, 2, 1, 0, 0, 0, -1, -1, -1, -1, -2, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, -1, 0, 1, 2, 3, 3, 1, 0, 0, 0, -2, -2, -1, -1, -1, -1, 0, 1, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 2, 1, 1, 1, -1, 0, -1, -1, -3, -1, -1, 0, 0, 1, 1, 2, 1, 0, 0, 0, -1, -1, -2, -1, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, -3, -2, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, -1, 0, -1, -1, 0, -1, 0, -1, -2, 0, -2, -1, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -2, -1, -2, 0, -1, 0, -2, 1, 0, 0, -1, -2, -2, -3, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, -1, 1, 0, 0, 0, 0, -2, -3, -2, -1, -2, -1, -1, 1, 0, 2, 2, 2, 0, 1, 0, -1, -1, -1, -1, 0, -1, 3, 1, 0, 0, -1, -1, -2, -1, -1, -2, -1, 1, 0, 3, 3, 3, 2, 2, 2, 1, 1, 0, 1, 0, 1, 0, -3, -1, 1, 1, 1, 1, 2, 2, 4, 4, 6, 4, 5, 6, 5, 6, 4, 4, 3, 3, 2, 1, 1, 3, 2, 4, -3, 0, 0, 0, 1, 0, 1, 3, 3, 1, 2, 4, 4, 4, 3, 4, 4, 3, 1, 2, 0, 0, 1, 0, 1, 3, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 3, 2, 3, 4, 3, 1, 0, 0, 0, 0, 0, 0, 2, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 2, 3, 2, 0, 0, 0, 0, 0, 0, 2, -2, 0, 1, 0, -1, -2, 0, 0, -1, 0, -1, 0, 0, 0, 1, 4, 3, 2, 2, 0, 0, 0, 1, 1, 1, 2, -2, 0, 0, -1, -1, -1, -2, -2, -3, -3, -1, -1, -1, 0, 1, 2, 3, 2, 1, 2, 0, 0, 1, 0, 0, 2, 0, 0, 0, -1, -1, -1, 0, -2, -3, -5, -2, -2, -2, -3, -1, 1, 1, 3, 2, 2, 1, 2, 1, 1, 0, 0, -1, 0, 0, 0, -1, -2, 0, -2, -3, -6, -6, -5, -6, -4, -3, -1, 0, 2, 2, 1, 2, 1, 2, 1, 1, 1, -3, 0, 1, 0, 0, -1, -1, -1, -3, -5, -6, -6, -7, -6, -4, 0, 1, 2, 2, 1, 2, 0, 2, 0, 1, 0, -1, 0, 1, 3, 0, 0, -2, -3, -3, -6, -5, -8, -7, -6, -2, 0, 2, 4, 5, 2, 2, 1, 0, 1, 0, 1, -1, 1, 1, 2, -1, -1, -3, -2, -5, -6, -5, -7, -7, -5, -2, 0, 3, 5, 7, 6, 2, 2, 1, 1, 2, 3, -1, 1, 2, 1, 0, -3, -2, -5, -6, -6, -7, -7, -6, -4, -2, 2, 3, 6, 8, 7, 4, 2, 3, 2, 2, 1, 0, 1, 1, 0, -1, -3, -2, -4, -6, -4, -5, -6, -7, -4, -2, 0, 5, 7, 10, 9, 5, 3, 1, 2, 1, 2, -1, 0, 1, 0, -1, -1, -3, -4, -6, -5, -8, -6, -6, -6, -3, 0, 3, 6, 10, 7, 5, 3, 2, 0, 2, 2, -1, 0, 1, 0, -1, -2, -3, -4, -5, -6, -7, -8, -8, -7, -5, 0, 4, 5, 7, 6, 4, 3, 2, 2, 1, 2, -1, 0, 0, 0, 0, -1, -3, -4, -3, -4, -6, -8, -8, -5, -5, -2, 3, 4, 5, 4, 3, 1, 1, 1, 3, 3, -2, 1, 0, 1, -1, -2, -3, -3, -4, -4, -6, -7, -6, -5, -4, 0, 0, 3, 4, 4, 2, 1, 1, 0, 3, 3, 0, 1, 0, 0, -2, -2, -3, -2, -3, -4, -5, -4, -5, -4, -3, 0, 2, 1, 2, 3, 2, 1, 1, 1, 1, 3, -2, 1, 1, 0, 0, 0, -2, -2, -5, -4, -5, -4, -4, -3, -1, 0, 2, 2, 3, 3, 1, 1, 0, 0, 2, 3, -1, 0, 0, -1, -1, 0, -1, -1, -5, -4, -4, -2, -2, -2, 0, 0, 2, 1, 0, 1, 0, 0, 1, -1, 0, 2, -1, 0, 0, 0, 0, 0, -1, -2, -3, -2, -4, -3, -2, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 3, -2, 0, 0, -1, 0, 0, 0, -1, 0, 0, -2, -2, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 1, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 2, -1, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, -2, 0, 1, 1, 2, 4, -3, 0, 0, 2, 0, 1, 0, 2, 2, 3, 1, 4, 2, 2, 3, 1, 1, -1, 0, -2, -1, 0, 1, 1, 2, 6, -2, 0, 1, 2, 2, 3, 2, 2, 4, 4, 7, 7, 6, 5, 5, 4, 2, 1, 1, 1, 1, 1, 2, 3, 5, 5, 5, 3, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 1, 1, 1, 0, 0, -1, -1, -3, -3, -3, -4, 3, 2, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, -2, -3, -3, -2, -3, 3, 2, 1, 0, 0, -2, 0, -2, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -3, -3, -4, 2, 1, 0, 0, -2, -2, -1, -2, -3, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, -1, -2, -2, -2, 4, 2, 0, 0, 0, -1, -2, -3, -2, -3, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -3, 4, 2, 0, 0, 0, 0, -2, -1, -2, -3, -3, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 5, 1, 2, 1, 0, 0, 0, -2, -1, -2, -3, -3, -2, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, -2, -3, 6, 4, 2, 1, 1, 0, 0, -1, -1, -3, -3, -3, -1, -2, -1, 0, 0, 0, 0, 1, 0, 1, 0, -1, -2, -2, 5, 4, 1, 2, 2, 0, 0, 0, -1, -2, -2, -2, -1, -1, -3, -3, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 4, 3, 1, 0, 2, 0, 0, 0, -2, -1, 0, 0, -1, -2, -3, -3, -3, 0, 0, 0, 1, 0, -1, -1, -1, -1, 2, 0, 1, 1, 1, 1, 0, -1, 0, 0, 0, 0, -1, -3, -3, -4, -3, -1, 0, 0, 0, 0, 0, -1, 0, -1, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, -1, -1, -2, -3, -3, -1, 0, 0, 1, 0, 0, -1, 0, -2, 1, -1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, -2, -1, -3, -2, -1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -3, -3, -1, -1, 0, 2, 2, 0, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, -1, -1, -3, -2, -2, 0, 0, 1, 1, 0, 1, 0, -1, -1, 4, 2, 0, 1, 0, -1, -2, -2, -2, -1, -1, 0, -1, -2, -4, -4, -1, -1, 0, 1, 1, 0, 0, 0, 0, -1, 6, 2, 0, 0, 0, -2, -3, -3, -2, -1, -1, 0, -2, -2, -4, -1, -1, 0, 0, 0, 1, 0, 1, 1, -1, -1, 7, 3, 1, 0, -2, -2, -3, -4, -3, -2, 0, -2, -1, -2, -3, -3, -1, 0, 0, 1, 1, 0, 1, 1, 0, -1, 6, 2, 2, 1, -1, -2, -3, -3, -2, -1, -2, -2, -1, -3, -3, 0, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, 8, 4, 2, 0, -1, -3, -3, -3, -3, -3, -3, -2, -1, -3, -3, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 7, 4, 0, 0, -1, -2, -3, -3, -2, -3, -1, -3, -2, -2, -2, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 6, 3, 1, -1, 0, -2, -2, -2, -2, -2, -1, -2, -1, -2, -1, 0, 0, 1, 0, -1, 0, -1, 0, -1, -1, -2, 6, 2, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, -1, -1, -2, 0, -2, -3, 6, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, -1, -2, 0, -2, -3, -3, -2, 5, 3, 0, 0, 2, 0, 0, -1, 0, 1, 2, 2, 2, 2, 1, 0, 1, 2, 0, 0, 0, -2, -1, -2, -3, -2, 7, 3, 1, 1, 2, 0, 0, 0, 1, 0, 1, 2, 3, 2, 2, 2, 1, 1, 0, -1, -1, -2, -2, -2, -3, -5,
    -- filter=0 channel=8
    1, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 2, 1, 1, 1, 1, 0, 1, 1, 2, 1, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 2, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 2, 1, 1, 0, 0, 0, 0, 1, 1, 2, 0, 0, 1, 0, 1, 0, -1, -1, 0, -2, -1, 0, 0, 0, 1, 0, 1, 2, 2, 1, 0, 0, 1, 0, 1, 2, 2, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 1, 0, 1, 1, 0, 2, 0, 0, 0, 0, 0, 1, 2, 0, 1, 1, 0, -1, -1, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 1, 1, -1, 0, 0, -1, 0, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 2, 1, 0, 2, 0, 0, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 1, 0, 2, 1, 0, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 1, 2, 0, 0, 0, 1, 0, 1, 0, 2, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 1, 0, 0, -1, 0, -1, 0, -1, -1, 0, 1, 0, 0, 0, -1, 0, 2, 0, 1, 2, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, -1, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 2, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, -1, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 2, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 2, 2, 0, 1, 1, 0, -1, 0, 0, 0, 0, 1, 1, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 0, 0, 0, -1, 0, -1, -1, -2, 0, -1, 1, 0, 2, 3, 2, 3, 3, 3, 4, 3, 5, 4, 4, 2, 3, 1, 2, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 1, 2, 2, 2, 3, 4, 3, 3, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 3, 1, 1, 1, -1, -1, 0, 1, 0, 0, 1, 0, 1, 0, 0, -1, -1, -2, -2, 0, 0, 0, 0, 1, 1, 0, 3, 1, 1, 0, -1, 0, 0, 0, 0, 2, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, -2, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, -1, -1, -1, -2, 0, 0, -1, 0, 0, -1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, -2, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 2, 1, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, -2, 1, 1, 0, 0, 0, 0, 1, 2, 2, 0, 0, 1, 0, 0, 0, -2, -1, -1, -1, -1, 0, -1, -1, -1, 0, -1, 1, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, 1, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, 1, -1, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, 2, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, -2, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, 2, 2, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -2, 2, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, 0, 0, 0, -1, -1, -1, -2, -2, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 1, 1, 0, 0, 0, 1, 0, -1, -1, -1, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, 0, 1, 0, -1, 0, -1, -1, -2, -1, -1, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, -1, 0, -1, -2, -1, -1, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, -1, -1, 0, -2, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 2, 0, 0, 1, 2, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 1, 1, 1, 3, 3, 3, 3, 3, 3, 2, 2, -3, -3, -3, -3, -2, -3, -2, -2, 0, -1, -2, -2, 0, -1, -1, -1, -1, -2, -4, -3, -3, -5, -6, -9, -10, -12, -4, -4, -3, -2, -2, -1, -1, -2, -1, -1, -1, 0, 0, 0, 1, 0, -1, 0, -2, 0, 0, -2, -4, -5, -7, -10, -5, -3, -3, -2, -2, -1, 0, -2, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -6, -8, -4, -3, -2, -1, -3, 0, -1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 1, 1, 0, 1, 0, -1, -5, -7, -4, -2, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 0, 0, -2, -3, -7, -4, -3, -3, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 2, 0, -1, -2, -1, -6, -3, -4, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 1, 2, 2, 0, 0, 0, -2, -6, -5, -4, -2, -2, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 1, 0, 0, -1, -7, -5, -5, -3, -1, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 2, 1, 2, 0, 0, -2, -7, -4, -4, -3, -1, -2, -2, 0, -1, -1, -1, -1, -1, -2, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, -1, -2, -7, -5, -2, -2, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -3, -7, -4, -4, -3, -1, -2, -2, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, -2, -5, -3, -4, -3, -2, 0, 0, 0, 0, 1, 0, 0, 0, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6, -4, -2, -1, -2, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, -5, -2, -4, -2, -1, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -2, -4, -3, -4, -4, -1, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 1, 1, 1, -1, -6, -4, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -2, -6, -3, -4, -3, -2, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 1, 0, 0, 1, 0, -1, 0, 1, 0, 0, -5, -8, -4, -2, -3, -1, -1, 0, 0, 0, 1, -1, 0, -1, 0, 1, 2, 0, 1, 0, 0, 1, 0, 0, 0, 0, -5, -8, -2, -2, -3, -1, -1, -1, -1, 0, -1, 0, -1, -1, -1, 0, 2, 0, 0, 1, 1, 1, 0, 1, 0, -1, -4, -9, -4, -3, -2, -2, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 2, 0, 0, 0, 1, -1, -4, -9, -3, -2, -2, -1, -3, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 2, 0, 1, 0, 0, 0, -3, -5, -10, -2, -3, -3, -2, -2, -1, 0, -1, 0, 0, -1, 0, -1, 0, 1, 2, 0, 0, 0, 0, 0, 0, -1, -5, -7, -9, -3, -4, -3, -3, -2, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, -1, -4, -5, -8, -10, -4, -3, -4, -4, -3, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -5, -6, -8, -9, -10, -13, -4, -5, -5, -5, -2, -1, -2, -2, -1, -1, -1, -2, -2, -3, -2, -3, -3, -3, -5, -6, -8, -8, -11, -12, -13, -14, 0, -1, 0, 0, -1, -1, -1, -1, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -2, -1, 0, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, -1, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -2, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -2, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, -2, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, 0, 0, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, 0, -1, -1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -2, 0, -1, -1, -1, 0, -1, 0, -2, -1, -1, -1, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -2, -2, -1, 0, 0, -2, 0, 0, 0, -2, -1, -1, 0, 0, 1, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -2, 0, -2, -2, -1, -2, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 3, 3, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 3, 1, 2, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, -1, -2, 0, -1, 0, 0, 0, 2, 0, 1, 2, 1, 1, 0, 1, 0, -2, -2, -3, -2, -3, -2, -3, -3, -3, -3, -3, -2, -2, -2, -1, 0, 0, 3, 1, 1, 2, 2, 2, 1, 0, 0, -1, -1, -2, -2, -3, -1, -2, -2, -1, -3, -3, -1, 0, -2, 0, 0, 0, 1, 1, 2, 1, 0, 1, 1, 0, 0, 0, -2, -2, -2, 0, -2, -2, -2, -1, -2, -3, -2, -2, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, -2, -2, 0, -2, -1, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, -2, -1, -1, -1, -1, 1, 1, 1, 2, -2, -1, 0, -2, -1, -2, -1, -1, -2, -1, 0, 0, -1, -1, -1, 0, -1, -2, -2, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, -1, -2, -2, -2, -1, 0, 0, 0, 0, -1, -1, 0, -1, -2, -1, -1, -1, 0, 0, 0, -1, -2, -1, -2, -2, -2, -1, -2, -1, -3, -1, -1, 0, 1, 1, -1, -1, -2, -1, 0, -2, -1, -1, 0, 0, 0, -2, 0, -2, -2, 0, -2, -2, -1, -1, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, -2, -1, 0, 0, -1, 0, -2, -2, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -2, -1, -1, -1, -1, -1, 0, -1, 0, -2, -2, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, -2, -1, -3, -3, -1, -3, -3, -1, -1, 0, -1, -1, -2, -2, -1, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, -1, -3, -3, -4, -2, -4, -2, -2, -1, -2, -1, 0, -2, 0, -2, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, -3, -3, -2, -3, -2, -2, -2, -1, -1, -1, 0, 0, -2, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -3, -4, -2, -2, -4, -2, -2, -2, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, -1, -2, -3, -2, -3, -2, -1, -2, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -3, -1, -2, -3, -3, -2, -1, -2, -1, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, -1, -1, -1, -2, -2, -1, 0, 0, -1, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, -2, 0, -1, -1, -2, -2, -1, -1, 0, -2, -2, -1, -1, -1, -1, 0, 0, 0, -1, -2, -1, -1, -1, -1, -2, -1, 0, 0, 0, -1, -1, -1, -2, -1, -1, -2, 0, -1, -1, -1, -2, -1, -2, 0, -1, -2, -2, -2, -1, -1, -1, 0, 0, -1, 0, -1, -1, -2, 0, 0, 0, -2, 0, -2, -1, 0, 0, 0, -1, -2, -2, 0, -2, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, -1, -1, -2, -1, -2, -1, 0, -2, -2, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, 0, -1, -1, -2, -2, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -2, 0, -1, -1, -2, -2, -2, -1, -2, -1, -1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, -2, -2, -1, 0, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 1, 1, 0, 0, -1, -1, 0, -1, -2, -1, -2, 0, -1, -2, 0, -2, 0, 0, 0, 0, 0, 1, 2, 2, 2, 0, 2, 1, 1, 0, -2, -2, 0, -2, -2, -1, -2, -2, -1, -2, -3, -2, -1, 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 1, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -2, -2, -1, -2, -2, -2, -1, -1, -2, -4, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -2, 0, 0, -1, -1, -1, -1, -1, -1, -1, 0, -1, 0, 0, -1, -2, -1, 0, -2, 0, -1, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, -2, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, -2, -1, -2, 0, 0, 0, 0, 1, 2, 0, 1, 0, -1, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, -2, -2, -2, -1, 0, 0, 1, 1, 2, 2, 1, 0, 2, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, -1, 0, 0, -2, -1, -1, 0, 0, -1, 0, 0, 1, 2, 2, 1, 0, 0, -1, -1, 0, -2, 0, 0, -1, -1, -1, 0, -1, 0, -2, -1, 0, 0, 0, 0, 1, 1, 3, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -1, -1, 0, 0, -2, -1, 0, -1, 1, 0, 0, 1, 1, 2, 2, 2, 2, 1, 0, -1, 0, -1, 0, 0, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 0, 0, 0, -1, -1, 0, -1, -2, -2, 0, -1, -1, -3, 0, -1, -1, -1, 0, 0, 1, 0, 1, 1, 1, 3, 3, 1, 0, -1, 0, 0, -2, -2, -2, -2, -2, 0, -1, -2, -3, -2, 0, -1, -1, 0, 0, 2, 1, 1, 2, 3, 1, 1, 1, -1, 0, -1, -2, -2, 0, 0, 0, -2, 0, -2, -2, -1, -1, 0, 0, 0, 0, 1, 3, 2, 1, 2, 1, 1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, -1, -2, -2, 0, -1, 0, 0, 0, 0, 1, 2, 2, 1, 2, 1, 1, 1, -1, 0, -1, 0, -2, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 0, -1, -1, 0, 0, -1, 0, 0, 0, -2, -1, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 2, 1, 2, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 2, 2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 2, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 1, 2, 0, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 1, 0, 1, 2, 1, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, 0, 2, 2, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, -1, 0, -1, -1, 0, 0, 1, 0, 1, 0, -1, -2, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, -1, 0, 1, 0, 1, 0, 0, -1, -1, 0, -1, -1, -2, -2, 0, 0, -1, 0, 0, 0, -2, -2, 0, -1, -1, 0, -2, -1, 0, 0, -1, -1, -2, -3, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, -1, -2, 0, -2, -2, -1, -2, -3, -3, -2, -1, -2, -1, -2, -4, -2, -2, -2, -1, 0, -2, 0, 0, -2, -2, -1, -4, -4, -4, -5, -6, -5, -7, -6, -6, -4, -6, -7, -9, -11, -15, -21, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, -3, -3, -3, -2, -3, -3, -3, -2, -2, -1, -3, -3, -6, -13, -19, -3, -2, 0, -1, 0, 0, 1, -1, -1, -1, -1, -3, -1, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, -3, -8, -14, -2, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, -1, -2, -5, -13, -2, -1, -2, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 1, 2, 1, 0, 0, 1, 3, 0, 1, -1, -5, -11, -3, -3, -2, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 2, 2, 1, 0, 3, 1, 1, 0, -1, -3, -9, -1, -2, -3, -3, -1, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 3, 2, 2, 2, 3, 3, 1, 2, 0, -2, -10, -1, -2, -2, -3, -2, -1, 0, 1, 0, -1, 0, 0, 0, 0, 2, 1, 3, 1, 1, 3, 3, 2, 0, 0, -2, -10, -2, -2, -4, -3, -2, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 2, 2, 2, 1, 2, 3, 1, 0, 0, -1, -9, -4, -2, -3, -2, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 3, 1, 2, 2, 2, 1, 1, -3, -7, -2, -3, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 3, 1, 2, 2, 3, 2, 1, -3, -8, -3, -2, -2, -2, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, 1, 1, 1, 1, 0, 1, 1, 1, 1, 0, -1, -7, -2, -2, -3, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 2, 0, -1, -6, -3, -2, -3, -1, -1, 0, 0, 1, 0, 0, 0, -2, -1, 0, 0, 2, 1, 1, 1, 0, 2, 2, 1, 2, 0, -7, -1, -3, -2, -2, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 3, 1, 2, 0, 0, 1, 3, 2, -2, -5, -1, -1, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 3, 1, 0, 0, 2, 2, 2, 1, -2, -7, -1, -3, -2, -2, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 1, 2, 3, 1, 1, 0, 2, 3, 0, -1, -6, -2, -2, 0, 0, 0, 1, 0, -2, -2, -2, 0, -1, 1, 2, 1, 3, 2, 2, 1, 1, 2, 3, 1, 1, -1, -7, -2, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 2, 3, 1, 0, 3, 1, 1, -2, -9, -1, -1, 0, 0, 1, 1, 0, -2, -1, 0, 0, 0, 2, 2, 2, 1, 2, 1, 3, 0, 0, 2, 1, 0, -4, -10, -1, -1, -2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 1, 1, 1, 0, 0, 1, 0, -3, -10, -3, -1, -2, 0, 0, 2, 0, 1, 0, 1, 1, 2, 1, 2, 1, 2, 2, 2, 2, 1, 0, 0, 0, -1, -7, -12, -2, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 3, 3, 2, 2, 0, 0, 0, 0, -4, -6, -13, 0, 0, -2, -2, 0, 1, 2, 0, -1, 1, 0, 0, 0, 0, 1, 1, 3, 3, 3, 0, -1, -1, -1, -6, -8, -15, -1, 0, 0, -2, -1, 0, 2, 0, 0, -1, 0, 0, -3, -2, -2, 0, 0, 3, 0, 0, -1, -3, -4, -7, -12, -17, -2, 0, -1, -1, -1, 1, 1, 1, -1, 0, -2, -2, -2, -2, -2, -3, -2, 0, -2, -3, -4, -5, -7, -11, -14, -19, 7, 5, 3, 0, 0, -1, 0, 0, 0, 0, 2, 2, 2, 2, 1, -1, 0, -1, 0, 2, 3, 3, 2, 2, 0, -1, 7, 6, 5, 2, 1, 0, 0, 1, 0, 2, 2, 3, 3, 1, 0, -2, -3, -3, -1, 0, 1, 0, 3, 2, 2, 0, 7, 8, 4, 3, 2, 0, 1, 0, 1, 3, 2, 2, 2, 0, 0, -3, -2, -3, -4, -2, -1, 0, 3, 3, 2, 0, 7, 6, 4, 1, 0, 1, 0, 2, 1, 2, 3, 2, 1, 0, 0, -2, -3, -5, -3, -3, 0, 0, 2, 1, 1, -1, 8, 7, 3, 1, 1, 1, 2, 0, 0, 2, 3, 4, 1, 2, 0, 0, -1, -4, -4, -2, -1, 0, 0, 1, 0, -1, 9, 7, 3, 1, 1, 2, 1, 3, 3, 2, 1, 4, 2, 0, 1, 1, -1, -1, -3, 0, 0, 0, 0, 0, 0, 0, 6, 6, 2, 2, 0, 0, 0, 3, 1, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 5, 4, 3, 0, 0, 0, 2, 3, 2, 2, 1, 0, 0, -1, 0, 0, -1, -1, 1, 2, 2, 2, 0, 1, 1, -1, 5, 4, 3, 0, 0, 2, 2, 2, 3, 2, 0, 0, -2, -1, 0, -1, -2, 0, 0, 3, 2, 2, 2, 0, 0, -1, 7, 5, 1, 0, 0, 1, 2, 2, 2, 0, 0, -1, -2, -1, 0, -1, -1, 0, 0, 1, 3, 2, 1, 2, 0, -1, 5, 4, 3, 1, 0, 0, 0, 1, 0, -1, -1, -3, -2, -1, 1, 0, -1, 0, 2, 1, 2, 3, 3, 3, 0, 0, 6, 4, 1, 1, 0, -1, 0, 0, 0, -3, -4, -5, -4, -1, 0, 0, 0, 0, 2, 2, 3, 4, 3, 3, 1, -1, 5, 4, 4, 1, 0, 0, 1, 0, -1, -3, -4, -4, -3, 0, -1, 0, 1, 2, 2, 4, 3, 4, 3, 1, 0, -3, 5, 4, 3, 2, 0, 0, 0, 1, 0, 0, -3, -4, -3, -1, 0, 0, 2, 1, 3, 3, 2, 3, 1, 1, 0, -3, 7, 4, 2, 1, 0, 1, 1, 0, 1, 0, -1, -3, -4, -2, 0, 0, 3, 2, 2, 3, 3, 3, 3, 0, 0, -2, 7, 5, 1, 0, 0, 0, 1, 0, 0, -1, 0, -2, -3, -1, 0, 1, 2, 2, 2, 3, 2, 1, 0, 2, 0, -2, 5, 3, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, -2, -1, -2, -1, 0, 0, 1, 0, 0, 0, 0, 2, 0, -1, 3, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, -2, -2, 0, 0, 0, 0, -1, 0, 0, 1, 1, 2, 0, 0, 3, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -2, -2, -1, 0, 0, 1, 1, -1, 3, 0, 0, 1, 0, 1, 1, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -1, 0, 0, -1, 2, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 0, 1, 0, -1, 0, -1, 0, -1, -1, -3, -1, -2, 0, 0, -1, 1, 1, 1, 1, 0, 0, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -3, -2, -2, -4, -3, -2, -1, -2, 3, 1, 0, 0, 0, -1, 0, 0, 2, 0, 0, 0, -1, 0, -2, -3, -1, -2, -2, -3, -2, -3, -2, 0, -1, -2, 3, 1, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, -3, -2, -1, 0, -1, -2, -1, 0, 0, 0, -2, 3, 3, 3, 1, 0, 0, 0, 1, 1, -1, 0, 0, 0, -1, -2, 0, 1, 0, 0, 0, 0, 0, 1, 3, 1, -1, 3, 4, 4, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 3, 2, 3, 4, 3, 4, 4, 4, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, -1, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, -2, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 1, 0, 1, -1, 0, -2, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 1, 1, 1, 1, 1, 2, 0, 0, -2, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, -2, 5, 3, 2, 0, 0, -2, -2, -4, -2, -3, 0, 2, 3, 1, 1, 0, 2, 2, 2, 5, 4, 5, 3, 1, 0, -5, 6, 6, 3, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -2, 0, -1, -1, 0, 2, 4, 3, 3, 0, -4, 8, 7, 5, 1, 0, 0, 0, 1, 1, 1, 2, 2, 2, 0, -1, 0, -2, -1, -3, -1, 0, 3, 3, 3, 0, -3, 7, 6, 4, 0, 1, 0, 0, 1, 3, 4, 4, 3, 2, 0, 0, -1, -2, -3, -4, -2, 0, 2, 3, 2, -1, -3, 7, 6, 4, 0, 0, 1, 0, 1, 1, 4, 5, 3, 2, 2, 1, 1, -2, -3, -3, -1, -2, 0, 1, 0, 0, -6, 7, 6, 3, 0, 0, 0, 2, 2, 2, 5, 5, 5, 3, 1, 1, 1, 0, 0, 0, -1, -1, 1, 1, 0, -2, -6, 6, 4, 2, 0, 0, 0, 0, 2, 2, 4, 4, 3, 2, 2, 2, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, -4, 5, 4, 0, -1, 0, 0, 3, 3, 3, 2, 3, 1, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 0, 0, -2, -7, 4, 3, 1, 0, 0, 2, 3, 5, 5, 3, 1, 1, 0, 0, 0, -1, 0, 0, 1, 2, 3, 1, 0, 0, -2, -6, 4, 2, 1, 1, 0, 0, 2, 5, 4, 3, 0, 0, 0, 1, 1, 1, 0, 0, 0, 2, 4, 3, 1, 0, -1, -7, 4, 2, 1, 0, 0, 1, 2, 4, 3, 2, 0, 0, -1, 1, 0, 1, 1, 0, 0, 1, 1, 3, 1, 2, -1, -6, 4, 4, 2, 0, 0, 0, 2, 1, 0, -1, -1, -2, -2, 0, 0, 0, 0, 1, 3, 2, 4, 1, 1, 2, 0, -6, 5, 4, 2, 1, 0, 0, 1, 1, 0, -2, -2, -2, -1, 0, 0, 1, 2, 1, 1, 2, 2, 2, 2, 0, 0, -6, 5, 4, 2, 1, 0, 2, 2, 3, 1, -1, -3, -2, 0, 0, 2, 1, 2, 3, 2, 3, 2, 1, 0, 0, -2, -8, 7, 4, 2, 1, 0, 1, 2, 2, 1, 0, -1, -1, -2, 0, 1, 2, 3, 3, 3, 4, 3, 1, 2, 0, -2, -8, 6, 3, 1, 0, 0, 2, 1, 2, 0, 0, -1, -1, 0, -1, 0, 2, 1, 4, 3, 4, 1, 1, 1, 0, -2, -6, 5, 3, 0, 0, 0, 0, 2, 2, 0, -1, -1, -2, 0, 0, 0, 0, 2, 1, 0, 0, 1, 1, 0, 1, 0, -5, 3, 1, 1, 0, 0, 2, 2, 1, 1, 0, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 2, 1, -3, 1, 1, 0, 0, 0, 2, 2, 2, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, -2, -1, 0, 0, 0, 1, -1, -4, 0, 0, 0, 1, 2, 2, 1, 2, 2, 1, 2, 1, 0, 0, 1, 0, 0, -2, -3, 0, 0, 0, 0, 0, -2, -6, 1, 0, 1, 0, 0, 2, 1, 1, 2, 2, 0, 1, 0, 0, 0, 0, -1, -1, -1, -2, -1, -2, 0, 0, -2, -5, 1, 0, 0, 0, 0, 0, 1, 2, 0, 2, 1, 2, 1, 1, 0, -1, -1, -2, -1, -2, -3, -2, -1, -2, -3, -8, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -2, -1, -2, -3, -3, -2, -2, -2, 0, -1, -2, -6, 2, 2, 0, 0, -1, -1, 0, 0, -1, 0, -2, -1, -1, -2, -2, -3, 0, -2, 0, 0, 0, 0, -1, -2, -2, -6, 3, 2, 1, 1, -1, 0, -1, 0, 0, -2, -2, -2, -2, -2, -3, -1, -1, 0, 2, 1, 1, 1, 2, 1, 0, -7, 5, 3, 4, 1, 0, -1, 0, 0, -1, -1, 0, -2, -1, -2, -1, 0, 1, 3, 3, 3, 4, 4, 3, 2, -1, -5, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, -1, 0, 0, -2, -2, -1, -2, 0, -1, 0, -1, -2, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 2, 1, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, 0, 0, 1, 1, 0, 0, 2, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 1, 0, 0, 0, 0, 1, 0, 2, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, 0, -2, -1, 1, 1, 0, 2, 0, 0, 1, 1, 1, 1, 1, 2, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, -2, 0, -1, 0, 0, 0, 2, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -2, -2, 0, -2, -1, -2, 0, -1, 0, 2, 2, 1, 2, 2, 2, 0, 0, 1, 1, 2, 0, 0, 0, -1, -1, -1, -2, -1, -2, -3, -1, 0, -1, 0, 1, 0, 2, 2, 2, 2, 1, 2, 1, 0, 0, 1, 0, 0, 0, 0, -1, -2, -1, -3, -1, -2, -2, -2, -1, 0, 0, 0, 0, 2, 1, 2, 1, 0, 0, 2, 0, 1, 0, 0, -1, -1, 0, -2, -2, 0, -1, -3, -2, -1, -1, -1, 0, 0, 0, 2, 1, 2, 2, 1, 1, 0, 0, 2, 0, 0, 0, 0, -2, 0, 0, -2, -1, -3, -2, -2, -1, -1, 0, 1, 0, 2, 3, 3, 4, 1, 1, 0, 1, 1, -1, 0, -1, 0, -1, 0, -1, -2, 0, -1, -2, -2, -1, 0, 0, 0, 0, 0, 1, 2, 3, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, -2, -1, -3, -1, -2, -2, 0, 0, 0, 0, 2, 1, 3, 3, 0, 1, 1, 2, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -2, -2, -3, -1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 1, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, -1, -1, -2, -2, -1, 0, 0, 1, 0, 2, 1, 1, 2, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -2, 0, -1, 0, -1, 0, 0, 0, 0, 2, 3, 2, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, -2, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 1, 2, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -2, 0, 0, 0, 1, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 3, 1, 1, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 0, 1, 0, 1, 1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 2, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 1, 1, 1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 3, 3, 2, 1, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, -1, 0, 0, -1, 1, 2, 1, 3, 3, 2, -2, 4, 3, 2, 1, 0, 1, 0, 1, 0, 0, 2, 1, 0, 0, 0, 0, -2, 0, -1, 0, 0, 2, 2, 1, 1, 0, 3, 2, 2, 1, 1, 1, -1, 0, 0, 0, 0, 1, 1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 1, 2, 1, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 1, 2, 1, 1, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 1, 0, -2, 2, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, 2, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -2, 2, 2, 0, 0, -1, 0, 1, 1, 1, 2, 0, -1, 0, 0, 1, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, -2, 0, 0, 0, -1, 0, 0, 1, 1, 2, 3, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 1, 0, 1, 1, 0, -2, 1, 0, 0, 0, 1, 1, 3, 3, 2, 1, 1, 0, 0, 0, 0, -2, -1, -1, 0, 0, 1, 2, 1, 1, 0, -2, 0, 1, 1, 0, 0, 2, 1, 2, 2, 0, 0, -1, 0, 0, 0, -1, -1, -2, -2, 0, 0, 1, 1, 1, 0, -1, 0, 1, 0, 1, 1, 0, 0, 2, 1, 0, -1, -2, -2, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 0, -2, -2, -1, 0, 0, 1, 0, 0, 1, 1, 0, 1, 2, 1, -2, 2, 1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, -1, -1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, -1, 1, 0, 1, 0, 0, -1, 0, 0, 1, 1, -1, -2, -1, -1, 0, 1, 0, 0, 1, 1, 1, 2, 0, 1, 0, -1, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, -1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 1, 1, 1, 1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, -1, -2, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 3, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 2, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, -1, -1, 0, -1, -2, 0, -1, -1, -1, 0, -2, -3, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -2, -2, -1, 0, 0, 0, -3, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -2, -1, -1, -1, -1, -1, 0, -1, 0, -1, -1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -2, -2, -1, -2, -1, 0, 0, 0, 0, 1, 0, 0, -1, -3, 2, 1, 1, 0, 1, 0, 0, 0, 0, -1, -2, -1, 0, -1, -1, -3, 0, -1, -1, 0, 1, 0, 0, 1, 0, -4, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, -4, 3, 2, 2, 1, 2, 1, -1, -1, -1, 0, -1, -1, 0, 0, -2, -3, -2, -2, -3, -2, -1, -3, -3, -2, -2, -6, 2, 4, 1, 2, 2, 0, -1, -1, -1, 0, -1, -1, 0, -1, -1, -2, -3, -2, -1, -2, -2, -1, 0, 0, -1, -3, 2, 2, 3, 2, 2, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -3, -1, -3, -3, 0, 0, 0, 0, 0, -4, 3, 3, 2, 3, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, -3, 3, 4, 3, 0, 1, 1, 0, 1, 2, 1, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, -2, -2, 3, 2, 1, 1, 0, 1, 2, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 2, 0, 0, 1, 0, 3, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 1, 0, 0, -1, 2, 0, 0, 0, 0, 0, 2, 2, 2, 1, 2, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 2, 2, 0, 0, -1, 1, 0, 1, 0, 0, 0, 1, 2, 3, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 1, 2, 2, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 2, 2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 2, 2, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, -2, 0, 0, 0, 0, 1, 0, 1, 2, 1, 3, 2, 3, 1, -1, 2, 0, 0, 0, 0, 1, 1, 1, 1, 0, -1, -1, -1, -1, 0, 0, 1, 0, 2, 2, 3, 1, 4, 3, 1, 0, 1, 1, 0, 2, 0, 0, 0, 3, 0, 0, 0, 0, 0, -2, 0, 0, 0, 2, 3, 3, 3, 2, 2, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 2, 1, 1, -1, 0, -1, -1, 0, 1, 2, 2, 3, 3, 3, 1, 2, 2, 0, -2, 3, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -1, 0, 1, 0, 1, 2, 0, 1, 1, 1, 1, 1, 0, 1, 2, 0, 1, 0, 0, 1, 0, 1, -1, -1, -1, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -3, 0, 0, 1, 1, 1, 1, 0, 2, 0, 0, 0, 0, 0, 1, -1, -2, 0, 0, -2, 0, 0, -1, -2, -1, -1, -2, 0, 1, 0, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, -1, -2, 0, 0, 0, -1, 0, -1, -1, 0, -1, -2, 0, 2, 1, 0, 2, 2, 1, 0, 0, 1, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, -1, -1, -1, 0, -2, -2, 1, 2, 1, 1, 1, 2, 2, 1, 1, 1, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, 3, 1, 1, 1, 1, 3, 0, 1, 1, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, -3, 5, 5, 4, 3, 1, 2, 2, 2, 5, 5, 6, 5, 4, 2, 2, 1, 0, 2, 4, 3, 4, 6, 8, 7, 9, 8, 5, 6, 3, 3, 1, 1, 0, 3, 3, 5, 5, 4, 2, 0, 0, -1, -1, 0, 0, 0, 0, 3, 4, 6, 5, 4, 6, 4, 4, 1, 2, 0, 1, 1, 2, 3, 1, 1, 0, -1, -2, -3, -3, -2, -2, -1, 0, 0, 2, 4, 3, 3, 6, 4, 2, 1, 0, 0, 0, 2, 2, 2, 1, 2, 0, -1, 0, -2, -3, -3, -2, -1, -1, 0, 1, 2, 2, 0, 4, 5, 1, 0, 0, 1, 1, 0, 2, 2, 0, 1, 0, 0, -2, -1, -3, -1, -1, -1, 0, 0, 1, 2, 2, 0, 6, 3, 1, 1, 0, 1, 0, 3, 2, 2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 6, 3, 3, 1, 0, 2, 3, 2, 3, 2, 0, 0, -3, -1, -2, -2, 0, 0, 1, 0, 1, 0, 1, 1, 2, 0, 4, 4, 2, 0, 2, 4, 3, 2, 2, 3, 0, -1, -1, -2, -3, -3, -2, 0, 1, 2, 1, 0, 0, 1, 1, 0, 4, 3, 2, 2, 2, 3, 3, 3, 2, 1, 0, -1, -2, -1, 0, 0, -2, 0, 2, 2, 2, 2, 2, 2, 1, 0, 3, 3, 1, 2, 1, 2, 3, 1, 2, 0, 0, -1, -1, 0, 0, -1, -1, 1, 1, 4, 2, 1, 2, 1, 2, 1, 4, 2, 2, 0, 0, 0, 0, 1, 0, -2, -2, -2, 0, 0, 0, 0, 1, 2, 4, 5, 4, 3, 3, 2, 0, 0, 4, 3, 2, 1, 0, 0, 1, 0, -1, -1, -1, -2, -2, 0, 0, 1, 3, 3, 3, 4, 4, 3, 3, 2, 2, 0, 4, 2, 2, 0, -1, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 2, 1, 3, 6, 4, 4, 3, 3, 2, 0, -1, 5, 2, 1, 0, 0, 0, 0, 0, -1, -3, -1, -2, -1, 0, 1, 2, 4, 3, 3, 5, 4, 3, 1, 1, 0, -3, 4, 1, 1, -1, -2, 0, 0, 0, -1, 0, -2, -1, 0, 0, 2, 3, 3, 3, 2, 3, 4, 3, 1, 1, 1, 0, 3, 2, -1, 0, -1, 0, 0, 1, 0, -2, 0, -1, 0, 0, 1, 2, 2, 0, 2, 1, 2, 2, 3, 3, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 0, 2, 1, 2, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 2, 2, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 2, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, -1, -2, -1, 0, -1, -2, -3, -1, -1, 0, 0, 1, -1, 1, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -2, -2, -1, -1, -2, -2, -3, -3, -1, -1, 0, 0, 0, 2, 1, 0, 0, -1, -1, 0, 1, 1, 0, 0, 0, 0, -1, -2, -4, -5, -4, -5, -3, -2, -1, 0, 1, 0, 0, 3, 1, 1, 0, 0, 0, 0, 1, 1, 0, -1, 0, -2, -4, -3, -4, -5, -5, -4, -2, -3, -2, 0, 3, 2, 2, 2, 1, 2, 0, 0, 0, 0, 0, 1, 1, -1, -1, -2, -2, -3, -2, -4, -4, -3, -1, -1, 0, 1, 3, 5, 2, 2, 2, 3, 2, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, -1, 0, 0, 2, 4, 5, 5, 6, 4, 5, 4, 3, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 5, 4, 6, 4, 4, 5, 6, 6, 6, 9, 8, 9, 7, 5, 4, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -4, -2, -3, -2, -2, -1, 0, 0, -2, -3, -4, -9, 5, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -2, -2, -2, -1, 1, 0, 0, 0, -4, -7, 5, 3, 1, 1, 0, 1, 0, 0, 1, 2, 1, 1, 0, -1, -1, -2, -2, -4, -2, 0, 0, 2, 2, 0, -3, -7, 3, 2, 1, 1, 0, 1, 0, 1, 1, 2, 2, 2, 1, 0, 0, -1, 0, -3, 0, 0, 0, 0, 0, 0, -1, -8, 2, 2, 0, 0, 0, 0, 2, 3, 2, 3, 1, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, -3, -6, 3, 3, 1, 0, 0, 0, 1, 1, 3, 2, 1, 2, 2, 0, 1, 2, 1, 0, 0, 1, 0, 0, 0, 0, -1, -7, 3, 1, 0, -1, 0, 0, 2, 3, 2, 3, 1, 1, 0, 1, 1, 0, 1, 2, 1, 2, 0, 0, 0, 0, -2, -8, 2, 0, -1, -1, -2, 1, 2, 1, 3, 1, 0, 0, 0, 0, 0, -1, 1, 1, 1, 4, 3, 1, 1, 0, -3, -7, 2, 0, 0, -2, 0, 0, 2, 1, 3, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 2, 3, 2, 2, 0, -1, -6, 1, 1, 0, -1, -1, 0, 1, 1, 3, 1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 2, 2, 2, 2, 0, -2, -6, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -2, 0, -1, 0, 0, 2, 0, 2, 1, 2, 2, 2, 2, 1, -2, -7, 2, 2, 0, 0, -1, 1, 0, 1, 0, -1, -1, -2, -1, 0, 0, 1, 1, 1, 0, 1, 3, 3, 3, 0, -1, -7, 1, 1, 2, 0, 0, 0, 1, 1, 0, -1, -1, -1, -2, 0, 0, 1, 1, 2, 2, 2, 3, 3, 0, 0, -3, -6, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, 1, 2, 3, 3, 3, 2, 2, 0, 2, 1, -3, -7, 3, 2, 1, 1, 1, 2, 2, 2, 0, 1, -1, -1, -1, 0, 1, 2, 2, 3, 3, 1, 1, 1, 1, 0, -2, -5, 1, 1, 1, 1, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 1, 1, 1, 0, -4, 2, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 1, 2, 2, 0, 0, -1, -5, 1, 1, 0, 1, 2, 1, 3, 2, 1, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, -5, 0, 0, 0, 1, 2, 2, 2, 3, 1, 1, 0, 1, 1, 1, 2, 0, 0, 0, -1, 0, 1, 1, 0, -1, -3, -6, 0, 0, 0, 0, 0, 2, 2, 3, 2, 2, 1, 1, 2, 1, 2, 0, 0, 0, -1, -1, -1, 0, 0, -1, -4, -7, 0, 0, 0, 0, 1, 1, 2, 2, 2, 2, 1, 2, 1, 2, 1, 0, -1, -1, 0, -1, 0, 0, -1, -1, -5, -9, 0, 0, 0, 1, 1, 2, 1, 1, 2, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, -2, -2, -1, -1, -2, -5, -7, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, 0, 0, -1, -2, 0, -1, -4, -9, 2, 1, 2, 0, 1, 1, 0, 0, -1, 0, -1, 0, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, -9, 3, 1, 1, 1, 1, 0, -1, -1, -2, -1, -1, -2, -1, -1, 0, -1, 0, 0, 1, 0, 2, 0, 0, -2, -5, -10, 3, 1, 0, 0, 1, 1, -1, 0, 0, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -5, -10, 0, 0, 0, 1, 0, 0, 1, 3, 5, 5, 5, 5, 5, 2, 2, 1, 2, 4, 3, 4, 4, 6, 5, 6, 6, 5, 0, 0, 0, 1, 1, 1, 0, 3, 5, 4, 5, 4, 2, 0, 0, 0, 0, 0, 1, 0, 1, 3, 3, 2, 4, 3, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 1, 0, 0, 0, 0, 0, -2, -1, 0, 1, 0, 2, 2, 1, 1, -1, 0, 0, -1, 0, 1, 2, 1, 2, 2, 1, 0, 0, -1, -1, 0, -3, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, 0, -1, 0, 0, -2, -2, -1, 0, -1, 0, 1, 0, -1, 0, -1, -1, -1, 0, 1, 2, 2, 3, 1, 2, 1, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, -2, 1, 1, 0, 0, 1, 3, 2, 1, 1, 2, 0, -1, -1, -2, -2, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 2, 3, 2, 2, 1, 1, 0, -2, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, 1, 0, 2, 2, 2, 3, 2, 3, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 0, -1, 0, -2, 1, 2, 1, 1, 1, 3, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 3, 2, 0, 0, 0, -1, -3, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 3, 2, 1, 1, 0, 1, 0, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -1, 0, 1, 1, 1, 1, 0, 1, 3, 3, 2, 2, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 1, 2, 2, 2, 2, 3, 2, 2, 2, 2, 1, 0, -2, 0, 0, 0, -1, -1, 0, 1, 0, 0, -2, -1, 0, 1, 3, 2, 1, 1, 2, 3, 2, 3, 2, 1, 0, 0, -2, 0, 0, -1, -1, 0, 0, 2, 0, 0, -1, -1, 1, 1, 4, 3, 1, 2, 3, 2, 1, 1, 1, 1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 1, 0, 2, 4, 2, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, -2, 0, 0, -1, -1, 0, 0, 2, 2, 2, 0, 1, 1, 2, 3, 1, 1, 0, 0, -1, -1, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 1, 0, 1, 2, 2, 1, 1, 0, 3, 2, 2, 0, -1, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 2, 1, 1, 1, 2, 2, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 1, 1, 2, 1, 1, 2, 1, 0, -1, -2, 0, -2, -1, 0, 0, 0, -1, -2, 0, 0, 0, 1, 1, 0, 0, 0, 1, 2, 2, 0, 0, 0, 1, -1, -1, -2, -2, -2, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, -2, -1, -3, -2, -3, 0, 0, 1, 0, -1, -2, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 2, 1, 0, -1, -1, -2, -3, -4, -3, -3, 0, 0, 1, 0, 0, -1, 0, -1, 1, 0, 1, 0, 0, 0, 1, 2, 1, 0, 0, 1, 1, 0, -2, -3, -3, 0, 0, 1, 1, 2, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 3, 1, 0, 1, 1, 2, 2, 1, 0, -1, 0, 0, 0, 2, 2, 3, 2, -1, 0, 0, 0, -1, 0, 0, 0, 2, 3, 2, 4, 4, 4, 6, 7, 3, 3, 2, 1, 4, 5, 6, 7, 5, 5, 5, 4, 5, 3, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, -2, -1, -1, 1, 1, 0, 1, 3, 1, 0, -2, 6, 4, 5, 2, 3, 0, 0, 0, 0, 0, 1, 1, 0, -1, -1, -1, -1, -2, 0, 0, 0, 1, 2, 2, 0, -1, 5, 6, 4, 2, 2, 1, 0, 0, 0, 0, 0, 2, 1, 0, -1, 0, 0, -1, -2, 0, 0, 1, 2, 1, 0, 0, 5, 5, 3, 2, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 5, 4, 3, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, -3, 4, 3, 2, 0, 0, 0, 1, 0, 2, 0, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 1, 1, 0, 1, 0, -1, 3, 3, 1, 0, -1, 0, 1, 2, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 2, 1, 2, 1, 2, 0, 0, -3, 3, 1, 0, 0, -1, 0, 1, 2, 2, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 2, 1, 0, 0, -3, 2, 3, 0, 0, -1, 0, 0, 3, 3, 2, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 1, 0, 2, 0, -2, 3, 1, 1, 0, 0, 0, 0, 2, 2, 2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 2, 2, 0, -3, 3, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, 0, 1, 1, 0, 1, 1, 1, 1, 2, 3, 1, 0, -2, 3, 2, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 1, 3, 2, 1, 1, 2, 1, 1, 0, 0, -1, 3, 2, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 2, 3, 1, 2, 2, 1, 1, 0, 0, -1, 2, 3, 2, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 2, 2, 1, 2, 1, 1, 0, -3, 2, 3, 2, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 1, 2, 1, 2, 2, 0, 0, 1, -1, 2, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 2, 0, 1, 1, 1, 1, 0, -1, 2, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, -2, 2, 2, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, -1, -3, 2, 1, 1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -2, 2, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, 0, 0, 0, -1, -1, -3, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -2, -1, -2, -1, 0, 0, -1, 0, 0, -1, 0, -3, 3, 2, 2, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, -2, 4, 3, 3, 1, 2, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, -2, 0, -1, 0, 1, 0, 0, 0, 1, 0, -2, 3, 4, 3, 3, 3, 0, 0, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 1, 1, 1, 2, 0, 1, 1, 1, -2, 4, 3, 4, 1, 1, 1, 0, -1, -1, 0, 0, -1, 0, 0, 1, 1, 1, 1, 1, 3, 3, 2, 2, 0, 0, -3, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, 0, -2, 0, 0, 1, 0, 2, 0, 2, 2, 1, 1, 1, 0, 0, 0, -1, 0, -2, -1, -1, 0, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, 0, 0, -2, -1, 0, 0, -1, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -2, 0, -1, -2, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, 0, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, -2, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, 0, -1, -2, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, -2, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, -1, 0, -2, 0, -1, -2, 0, -1, 0, 0, -2, -1, -1, -1, 0, -1, -1, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, -1, -1, -2, -1, 0, -2, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 1, 0, 1, 1, 0, 0, 0, 0, -2, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, -2, -2, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, -2, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -2, -3, -2, -3, -2, -1, -1, 0, -1, 0, -1, 0, -2, -2, 0, -2, 0, -2, -2, -4, -5, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -2, -2, -1, -2, -1, -2, -1, 0, -1, 0, 0, -2, -1, -2, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, 1, 0, 1, -1, -1, -2, 1, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 1, 0, -3, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 1, 1, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 2, 2, 2, 2, 1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 1, 2, 1, 2, 1, 1, 1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 1, 0, 1, 2, 1, 1, 2, 1, 2, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 2, 1, 0, 2, 1, 1, 1, 3, 2, 1, 0, -2, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 3, 1, 2, 1, 2, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, -2, 0, 0, 0, 1, 1, 1, 1, 0, 2, 2, 2, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -2, 0, -2, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, -1, -2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, -2, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 0, 2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, -3, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 2, 1, 2, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 2, 2, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 1, 0, 1, -1, -3, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 2, 0, 2, 1, 0, 0, -2, 0, -1, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 1, 1, 0, -3, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 2, 2, 2, 0, 0, -3, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, -3, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, -2, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, -2, -2, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -2, 0, -1, -1, -1, 0, -1, 0, 1, 1, 0, 0, 0, 0, -3, -4, -5, -5, -5, -6, -8, -7, -6, -5, -8, -6, -6, -4, -1, 2, 1, 3, 3, 0, 0, -1, -2, -5, -4, -4, -3, -5, -3, -4, -4, -6, -5, -5, -5, -5, -6, -6, -5, -3, 1, 3, 4, 4, 1, 0, 0, 0, -1, -1, -2, -1, -1, -3, -4, -4, -5, -3, -5, -3, -3, -5, -4, -4, -2, 0, 2, 2, 2, 1, 1, 2, 0, 0, 1, 1, 1, 2, 3, -4, -3, -4, -2, -5, -5, -5, -4, -5, -5, -4, -1, 0, 1, 2, 1, 0, 0, 0, 0, -1, 0, 2, 1, 1, 2, -3, -1, -3, -4, -4, -4, -4, -6, -4, -4, -3, -1, 0, 1, 3, 0, 0, 0, -1, 0, 0, 0, 2, 0, 0, 1, -3, -3, -2, -4, -3, -4, -4, -6, -5, -4, -1, -1, 1, 2, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, -3, -2, -4, -5, -5, -5, -6, -7, -4, -4, -2, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, -3, -3, -4, -5, -5, -8, -7, -7, -5, -2, -1, 0, 0, 2, 3, 3, 1, 0, 0, 0, 0, 0, 0, 0, 1, 3, -4, -3, -5, -5, -6, -6, -7, -5, -4, -3, 0, 0, 3, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, -5, -4, -4, -6, -4, -7, -7, -4, -3, 0, 0, 1, 1, 0, 0, 0, 2, 0, 0, 0, 0, 0, -1, -1, 0, 1, -4, -6, -4, -5, -7, -6, -7, -6, -3, -2, 0, 0, 0, -1, 0, 2, 2, 1, 0, 0, 0, 0, 0, -2, -2, 0, -5, -4, -5, -4, -6, -5, -6, -5, -3, -4, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -3, -1, 2, -5, -3, -3, -4, -5, -4, -5, -4, -5, -4, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, 0, 2, -5, -3, -3, -2, -2, -4, -4, -3, -3, -4, -2, -2, -1, 0, 0, 0, 0, -1, -1, -1, -2, -1, -2, 0, -1, 0, -3, -1, -3, -3, -4, -3, -5, -5, -3, -3, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, -2, 0, -2, -1, -1, 0, -2, -1, -1, -3, -4, -5, -4, -3, -4, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -2, 0, -1, -2, -2, -2, -3, -5, -4, -5, -5, -2, -1, 0, 0, 1, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, -2, -2, 0, -2, -3, -2, -5, -4, -3, -5, -3, -4, -4, -2, -1, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, -1, 0, -1, -2, -1, -3, -4, -3, -3, -4, -4, -4, -2, -1, -2, -1, 1, 1, 1, 1, 1, 0, 0, 1, 1, 1, 0, 0, -2, -2, -4, -4, -4, -4, -3, -3, -4, -4, -3, -3, 0, -2, 0, 0, 0, 2, 1, 1, 0, 1, 1, 2, 0, 1, -2, -3, -5, -5, -6, -5, -3, -3, -5, -3, -3, -3, -1, -1, 0, 1, 0, 2, 3, 3, 2, 2, 3, 0, 1, 0, -3, -4, -4, -3, -3, -5, -5, -4, -5, -2, -4, -2, 0, 0, 1, 0, 1, 1, 2, 2, 4, 3, 3, 2, 0, 1, -4, -4, -2, -3, -3, -3, -5, -5, -3, -2, -2, -3, -1, 0, 1, 1, 1, 0, 2, 2, 1, 3, 2, 3, 2, 2, -2, -4, -4, -4, -4, -4, -4, -4, -1, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 1, 0, -3, -3, -4, -3, -5, -5, -4, -2, -2, -1, -2, -4, -1, 0, 0, 0, 0, 0, 0, 1, 3, 3, 2, 1, 0, 0, -3, -3, -4, -3, -5, -5, -4, -3, -2, -3, -4, -4, -3, -2, -2, -2, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, -1, 1, 4, 2, 2, 3, 3, 1, 1, 0, 0, 0, 1, 1, 0, -1, -2, -3, -1, -1, -1, 0, 0, 0, 1, 2, 0, -4, 3, 2, 2, 2, 3, 2, 1, 0, 0, 1, 1, 1, 0, 0, -3, -2, -2, -2, -1, 0, 0, 1, 2, 0, 0, -2, 4, 4, 2, 3, 1, 0, 2, 2, 1, 1, 0, 0, -1, -2, -2, -2, -3, -2, -1, -1, 0, 1, 2, 2, 0, -3, 3, 3, 2, 1, 2, 0, 2, 0, 2, 0, 0, 0, 0, -2, -2, 0, 0, -3, -3, -2, 0, 0, 2, 1, 0, -3, 4, 3, 1, 1, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 1, 0, -1, 2, 2, 2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 0, 0, 1, 1, 3, 1, 1, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 1, 1, -1, 1, 0, 0, 0, 1, 0, 3, 2, 2, 1, 1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 2, 1, 0, 0, 0, -2, 1, 0, 0, 1, 0, 0, 2, 2, 3, 2, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 2, 2, 3, 1, -1, 0, 0, 0, 0, 1, 2, 3, 2, 2, 1, 1, -1, -1, 0, 0, -2, 0, -1, 0, 2, 1, 4, 3, 3, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 2, 3, 5, 4, 3, 0, 1, 0, 0, 0, 0, 1, 1, 3, 0, 0, 0, 0, -2, 0, 1, 1, 0, 2, 2, 3, 2, 5, 5, 5, 2, 0, 1, 1, 0, 0, 1, 0, 2, 1, 2, 0, -1, -2, -1, -1, 0, 1, 0, 1, 2, 4, 3, 3, 3, 4, 3, -1, 0, 0, 1, 1, 0, 0, 2, 2, 0, 0, 0, -2, -1, 0, 0, 2, 1, 1, 3, 3, 2, 2, 4, 4, 2, 0, 0, 1, 0, 0, 0, 1, 0, 2, 2, 0, 0, -2, -2, 0, 0, 3, 1, 3, 2, 4, 2, 2, 2, 4, 3, 0, 2, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -2, 0, -1, 0, 2, 2, 1, 1, 2, 3, 1, 3, 3, 1, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, -2, -3, -2, 0, 0, 0, 2, 2, 2, 2, 0, 0, 2, 4, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -2, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 2, 3, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -2, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 1, 1, 0, 0, 1, 2, 1, 0, 2, 0, 0, 0, 0, -1, -1, -2, -2, -1, -1, -2, -1, -2, -2, -1, 0, -2, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 0, -1, -1, -2, -1, -3, -1, -2, -3, -2, -2, -1, 0, -1, -1, -4, 0, 1, 1, 0, 1, 1, 1, 2, 0, 0, 0, -2, -2, -1, -3, -2, -1, -2, -2, -2, -2, 0, -1, 0, -1, -2, 0, 2, 1, 0, 1, 2, 1, 2, 1, 1, 0, -1, -2, -3, -1, -1, -1, 0, 0, -1, -1, -1, -1, 1, 0, -3, 1, 1, 1, 1, 2, 2, 2, 1, 0, 1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -4, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 1, 1, 2, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 3, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 1, 2, 1, 2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 2, 1, 1, 1, 1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 2, 1, 1, 2, 0, 2, 3, 3, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, 0, 1, 1, 1, 1, 2, 2, 2, 2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 3, 2, 1, 2, 2, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 0, 0, 0, 1, 2, 2, 3, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 2, 1, 0, -1, 1, 2, 2, 3, 2, 2, 2, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 1, 2, 2, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, -1, 1, 0, 2, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 1, 0, 0, 0, -1, 1, 1, 1, 1, 2, 1, 1, 1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 0, 0, -1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 2, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 3, 1, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -2, -1, -1, 0, -1, -1, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, -1, -2, -2, -2, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, -1, 0, -1, -2, -2, -4, -5, -6, -5, -7, -6, -4, -5, -5, -5, -5, -7, -12, -17, 0, 0, 0, 1, 2, 2, 1, 1, 0, 1, -1, -2, -3, -3, -4, -3, -4, -3, -1, -3, -2, -1, -2, -5, -8, -13, 0, 0, 1, 0, 1, 1, 1, 2, 0, 0, 0, 1, -1, 0, -1, 0, -2, -2, -1, 0, -1, -1, 0, -3, -5, -12, 0, 1, 0, 0, 1, 0, 0, 2, 2, 2, 2, 1, 2, 1, 0, 0, 1, 2, 0, 1, 0, 0, 0, -1, -3, -10, 0, 0, 0, -1, -1, 0, 0, 2, 2, 1, 1, 1, 3, 1, 2, 1, 3, 3, 1, 0, 1, 1, 0, 0, -3, -9, 0, 0, -1, -2, -1, -1, 1, 0, 1, 2, 1, 1, 2, 1, 1, 3, 2, 2, 2, 3, 2, 2, 1, 0, -2, -8, 0, -1, -2, -3, -2, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 1, 3, 4, 3, 3, 1, 3, 2, -1, -2, -10, -1, 0, -2, -2, -2, -1, 0, 1, 1, 1, 0, 1, 0, 0, 1, 1, 2, 2, 3, 3, 2, 1, 2, -1, -2, -7, -1, -1, -2, -1, -1, 0, 0, 2, 3, 1, 1, 0, 1, 1, 0, 0, 0, 3, 3, 2, 2, 2, 2, 1, -3, -8, -2, -1, -2, -2, -1, -1, 0, 1, 1, 1, -1, -1, 0, -1, 0, 1, 2, 2, 1, 2, 3, 3, 2, 0, -1, -8, -1, -1, -2, -1, -1, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 1, 0, 1, 0, 2, 3, 2, 3, 0, -1, -8, 0, 0, 0, -1, 0, 0, 0, 0, 1, -1, -1, -3, 0, -2, 0, 0, 0, 1, 0, 2, 3, 1, 2, 1, -1, -7, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -2, -2, -1, 0, 1, 2, 2, 2, 2, 1, 2, 0, -1, -5, 2, 0, 0, 0, 0, 2, 1, 2, 2, 0, 0, -2, -1, -1, -1, 0, 0, 1, 3, 0, 1, 2, 2, 1, 0, -7, 0, 1, 0, 1, 0, 0, 2, 2, 2, 1, 0, -1, -3, -2, -1, 0, 1, 3, 1, 1, 2, 1, 2, 0, -1, -7, 1, 1, 0, 0, 0, 2, 1, 0, 0, -1, -1, -3, -1, 0, 0, 2, 2, 1, 1, 2, 2, 3, 1, 0, -2, -6, 0, 0, 0, 1, 1, 2, 1, 0, -1, -1, -2, -1, 0, 0, 1, 2, 0, 0, 0, 2, 1, 1, 3, 1, 0, -7, 0, 0, 0, 1, 1, 3, 2, 0, 0, -1, -1, -1, 2, 2, 3, 2, 0, 0, 0, 1, 1, 1, 2, 0, -3, -7, -1, 0, 0, 1, 3, 2, 2, 0, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, -3, -8, 0, 0, 0, 1, 1, 2, 2, 1, 1, 1, 0, 0, 4, 4, 2, 1, 1, 0, 0, 0, 1, 0, 0, -1, -4, -8, -1, 0, 0, 1, 0, 1, 2, 2, 1, 1, 1, 1, 3, 3, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -4, -9, 0, 0, -1, 0, 2, 3, 2, 1, 1, 2, 2, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, -3, -7, -12, -1, 0, 0, 1, 0, 1, 2, 2, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4, -6, -14, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, -1, -2, -1, -6, -9, -15, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, -1, -2, -2, -2, -2, -1, -1, 0, -1, -3, -3, -4, -8, -10, -16, 0, 0, 0, -1, 0, 0, 0, 0, 1, -1, -1, -3, -3, -4, -4, -4, -3, -3, -4, -4, -6, -8, -10, -12, -15, -21, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 1, -1, 1, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, -3, -3, -2, 0, 1, 0, 0, 2, 1, 2, 1, 1, 4, 2, 2, 0, 0, -3, -3, -4, -4, -5, -6, -5, -4, -7, -5, -3, -1, 0, 1, 2, 1, 1, 0, 0, 0, 3, 3, 3, 2, 1, -1, -2, -3, -1, -2, -2, -4, -4, -5, -5, -4, -2, -1, 0, 0, 1, 0, 1, 0, 2, 2, 3, 4, 2, 2, 0, -1, 0, -1, -1, 1, 0, -2, -4, -4, -4, -2, -2, 0, 0, 0, 0, 1, 3, 1, 3, 2, 3, 3, 0, 0, 0, -1, -1, 0, 1, 0, 0, -1, -2, -2, -4, -3, -2, 0, 2, 2, 2, 3, 3, 2, 1, 2, 1, 2, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -3, -3, 0, 1, 2, 1, 2, 2, 3, 3, 3, 2, 0, 0, -1, -1, -2, -1, -1, 1, 0, 3, 1, 0, 0, 0, -2, -2, -1, 0, 1, 1, 3, 2, 2, 2, 2, 2, 1, -1, -2, -2, -2, -2, -1, 0, 1, 1, 0, 0, 0, 0, 0, -3, 0, 0, 0, 2, 4, 2, 2, 1, 1, 0, -1, -1, -2, -3, -1, -2, -2, -1, 0, 0, 1, 0, 2, 0, -1, -3, -2, -1, 2, 2, 2, 3, 0, 0, 1, -1, 0, -4, -4, -4, -1, -2, -2, -2, 0, 0, 2, 2, 2, 1, -1, -1, 0, 0, 0, 0, 2, 1, 0, 0, 0, -2, -2, -3, -4, -3, -1, -2, -2, -2, 0, 1, 0, 1, 3, 1, 0, -1, -1, 0, 1, 0, 1, 1, 0, -1, 0, -1, -3, -3, -2, -1, -3, -2, -1, -1, -1, 0, 1, 3, 4, 3, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -3, -2, -2, -1, -1, -3, -2, 0, 0, 2, 4, 4, 3, 0, -2, -1, 0, 1, 1, 0, 0, 0, -1, 0, -1, -2, -2, -3, -1, 0, -1, -2, -3, 0, 2, 3, 4, 5, 4, 0, -2, -1, 0, 2, 0, 0, 0, 1, 0, -1, 0, -3, -4, -3, 0, -1, -2, -1, -1, -1, 1, 2, 4, 4, 4, 1, -2, -1, 0, 1, 0, 2, 1, 2, 0, 0, -1, -4, -4, -3, -2, 0, -2, -3, -2, 0, 1, 2, 5, 4, 3, 1, -2, -1, 0, 1, 1, 1, 1, 1, 0, 0, -2, -2, -4, -2, -1, -2, 0, 0, -2, 0, 0, 2, 4, 5, 4, 0, -1, 0, 0, 0, 3, 2, 2, 0, 0, -1, -2, -2, -3, -1, 0, -1, -2, -1, -1, -1, 2, 3, 5, 4, 1, 0, 0, 0, 1, 0, 1, 0, 2, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 2, 4, 4, 1, -1, -2, 0, 0, 2, 3, 2, 2, 2, 1, 0, -2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 2, 2, 3, 2, 1, -1, 0, 0, 0, 2, 2, 3, 2, 3, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 2, 2, 3, 0, -2, -1, -1, 0, 2, 2, 2, 1, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 3, 3, 3, 0, -2, -2, -2, 0, 1, 2, 3, 3, 3, 3, 1, 1, 0, 1, 2, 0, 0, 0, 0, -2, -2, 0, 2, 3, 1, 0, -4, -2, -1, 0, 1, 1, 1, 2, 2, 4, 2, 2, 0, 2, 0, 1, 1, 1, 0, -1, -1, 0, 1, 1, 0, -2, -5, -2, -1, -2, 0, 1, 1, 3, 3, 4, 2, 2, 2, 2, 0, 0, 1, 1, 0, 0, -1, 0, -1, -1, -3, -3, -4, -2, -1, 0, -1, 1, 3, 4, 2, 3, 2, 3, 3, 3, 0, 2, 1, 2, 1, -1, -2, -4, -4, -4, -3, -5, -7, -2, -2, -1, -2, 1, 2, 3, 3, 3, 3, 4, 4, 2, 2, 0, 0, 0, 0, -1, -3, -4, -5, -5, -4, -4, -6, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, -1, 0, -2, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, -1, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, -2, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, -2, -1, -1, -1, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 1, 2, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, -1, 0, 1, 0, -1, 0, 1, 1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 2, 1, 1, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 1, 0, -1, 0, 1, 0, 0, -1, 0, 0, -1, 0, -1, 1, 0, 0, -1, 0, 0, 1, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, -1, 0, 0, 1, 1, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 3, 2, 2, 2, 2, 3, 3, 1, 0, 1, 2, 1, 1, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, -1, 0, 2, 2, 2, 2, 3, 3, 4, 3, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 3, 3, 2, 2, 3, 0, 1, 0, 0, -1, -1, -1, -2, -1, 0, 0, 1, 2, 0, 2, 2, 0, 0, 1, 1, 3, 3, 2, 4, 2, 3, 1, 0, 0, -1, 0, 0, -2, 0, 0, 0, 0, 1, 1, 1, 1, 2, 0, 0, 0, 2, 2, 2, 2, 2, 2, 4, 1, 2, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 2, 0, 0, 1, 0, 2, 2, 4, 2, 2, 2, 4, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 0, 2, 1, 0, 0, 1, 1, 2, 3, 4, 3, 3, 3, 2, 0, 0, 0, -2, -1, -2, 0, -1, 0, 1, 2, 2, 1, 2, 1, 0, 1, 2, 1, 3, 3, 4, 2, 4, 3, 2, 1, 0, -1, -1, -1, -3, -1, 0, 0, 0, 0, 2, 2, 3, 2, 0, 0, 1, 2, 2, 4, 3, 3, 3, 1, 0, 0, -2, -3, -3, 0, -1, -1, 0, 0, 0, 2, 2, 2, 3, 3, 0, 1, 1, 3, 4, 2, 4, 4, 3, 0, 0, 0, 0, -1, -1, -2, 0, -1, 0, 0, 0, 2, 1, 3, 4, 2, 1, 0, 0, 2, 2, 3, 4, 3, 2, 0, 0, 0, -1, -1, -2, -2, 0, 0, 0, 0, 1, 2, 3, 4, 6, 3, 2, 0, 1, 2, 1, 2, 2, 3, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 3, 4, 6, 5, 3, 3, 0, 0, 0, 1, 3, 1, 1, 1, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 1, 1, 3, 6, 6, 7, 5, 3, 0, 0, 2, 1, 1, 2, 2, 2, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 2, 4, 5, 6, 5, 3, 1, 0, 0, 1, 1, 3, 3, 1, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 1, 2, 3, 5, 6, 6, 6, 3, 0, 0, 0, 2, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 4, 5, 5, 5, 3, 0, 1, 0, 1, 1, 1, 2, 2, 0, 0, -2, -2, 0, 0, 0, 0, -1, 0, 0, 1, 3, 2, 5, 5, 5, 4, 0, 0, 2, 1, 2, 2, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, 0, 0, 1, 1, 3, 5, 3, 4, 2, 1, 2, 3, 3, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 1, 0, 1, 1, 4, 3, 5, 3, 2, 0, 2, 2, 3, 1, 3, 3, 2, 1, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 1, 4, 3, 3, 4, 1, 0, 2, 2, 3, 2, 1, 2, 3, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, 1, 2, 2, 2, 1, 2, 1, 0, 2, 3, 3, 2, 3, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 2, 3, 2, 1, 0, 0, 0, 0, 1, 3, 2, 3, 4, 3, 2, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, 0, 2, 1, 1, 0, 1, 0, 1, 0, 2, 3, 4, 2, 3, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 0, 0, 1, 0, 1, 1, 3, 4, 3, 3, 2, 2, 1, 1, 1, -1, 0, 0, 0, -1, -2, 0, 0, 0, 1, 1, 1, 0, 0, 2, 2, 2, 4, 5, 4, 3, 3, 3, 3, 2, 0, 0, 1, 0, 1, 0, -1, 0, 0, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 3, 4, 2, 3, 2, 2, 1, -1, -2, -2, -4, -4, -5, -4, -5, -5, -6, -4, -3, -2, -1, -2, -1, -4, -7, -14, 4, 4, 3, 3, 2, 2, 0, 0, 0, 0, -2, -2, -2, -3, -2, -4, -3, -2, -2, 0, 0, 1, 1, 0, -4, -10, 5, 4, 4, 3, 1, 3, 2, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -2, 0, 0, 0, 2, 2, 0, -2, -9, 4, 3, 2, 0, 0, 2, 1, 2, 1, 1, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 2, 3, 2, 2, -2, -9, 5, 1, 0, 0, 0, 0, 0, 0, 1, 3, 2, 2, 2, 0, 2, 2, 2, 1, 1, 1, 2, 2, 3, 3, 0, -7, 3, 1, 0, 0, -1, 0, 0, 1, 2, 3, 3, 1, 3, 1, 2, 3, 2, 2, 3, 1, 2, 3, 3, 1, -1, -6, 3, 1, -2, -3, -3, -1, 1, 1, 0, 2, 2, 2, 2, 1, 2, 4, 3, 4, 5, 4, 4, 2, 3, 0, -2, -6, 1, 0, -3, -3, -4, -1, 0, 0, 2, 0, 1, 0, 0, 0, 1, 3, 3, 3, 3, 4, 5, 4, 3, 1, -1, -7, 0, 0, -3, -4, -2, -1, 1, 2, 1, 1, 0, -1, 0, 0, 2, 3, 3, 3, 5, 4, 5, 5, 3, 3, -2, -7, 1, -1, -2, -3, -1, 0, 1, 0, 1, 0, -1, 0, 0, 1, 1, 1, 1, 2, 4, 4, 4, 5, 5, 3, -1, -6, 0, 0, -2, -3, -2, -2, 0, 1, 1, 0, -1, -2, -1, 2, 0, 1, 2, 1, 2, 5, 3, 4, 3, 2, 0, -5, 1, 0, 0, -1, -2, 0, 0, 1, 0, -2, -2, -2, 0, 0, 0, 1, 2, 4, 2, 4, 4, 3, 3, 2, -1, -7, 2, 0, 0, -2, -1, 0, 0, 2, 0, 0, -3, -3, -1, -1, 0, 0, 1, 2, 4, 4, 3, 3, 3, 1, 0, -4, 4, 0, 0, -1, 0, 0, 1, 1, 1, -1, -4, -3, -3, -1, 0, 1, 4, 4, 3, 3, 3, 2, 1, 1, 0, -5, 3, 2, 0, -1, 0, 0, 1, 0, 2, -1, -3, -3, -3, -1, 1, 3, 4, 4, 4, 2, 1, 3, 3, 2, -1, -5, 3, 1, 1, -1, 0, 0, 0, 0, 0, 0, -3, -4, -2, 0, 1, 2, 4, 5, 3, 2, 2, 2, 2, 1, 0, -3, 3, 2, 1, -1, 0, 0, -1, 0, 0, -1, -2, -3, 0, 0, 2, 3, 3, 5, 4, 4, 2, 2, 4, 3, 1, -4, 1, 1, 0, 0, 0, 1, 0, 0, -1, -2, 0, -1, 0, 1, 1, 3, 3, 3, 2, 2, 2, 2, 2, 2, 0, -3, 1, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 1, 2, 3, 3, 1, 1, 2, 1, 2, 3, 3, 1, 0, -6, 1, 0, 0, 0, 2, 1, 0, 0, 0, 2, 0, 1, 2, 3, 1, 0, 1, 1, 1, 0, 2, 2, 0, 0, 0, -7, 0, 0, 0, 0, 0, 2, 1, 2, 0, 1, 0, 1, 2, 2, 1, 1, 0, 0, 2, 0, 1, 0, 0, -1, -2, -8, 0, 1, 1, -1, 0, 2, 1, 1, 0, 1, 1, 1, 0, 2, 2, 0, 0, 1, 1, 1, 0, 0, -1, 0, -4, -10, 1, 2, 1, 1, 0, 2, 1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, -2, -5, -10, 2, 2, 1, 1, 1, 1, 2, 0, 0, -2, -2, -1, -2, -3, -1, -1, 0, 0, 1, 0, 0, -2, 0, -3, -7, -12, 3, 3, 1, 0, 0, 0, 2, 1, 0, -2, -2, -4, -3, -5, -4, -2, -1, 0, 0, 0, -2, -2, -2, -3, -8, -14, 2, 3, 1, 0, 0, 0, 1, 0, -2, -3, -2, -3, -4, -4, -5, -4, -2, -1, -1, 0, -3, -3, -4, -7, -12, -16, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, -1, 0, -1, -1, -1, 0, 1, 0, 0, 2, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 2, 2, 2, 1, 1, 1, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 2, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 2, 1, 1, 2, 1, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 1, 1, 2, 2, 2, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 2, 1, 2, 2, 1, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 1, 2, 1, 3, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 2, 2, 2, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 2, 2, 0, 0, 0, 1, 1, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 2, 0, 2, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 1, 2, 2, 1, 1, 1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 2, 2, 2, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 2, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 1, 1, 1, 2, 2, 1, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, -1, -2, -3, -3, -3, -2, -2, -4, -4, -3, -3, -2, -3, -2, -2, 0, 0, 0, 0, 2, 1, 0, 1, 0, 0, -1, -1, -1, 0, -2, -2, -2, -2, -2, -3, -2, -2, -3, -4, -3, -2, 0, 0, 1, 1, 2, 2, 1, 0, 1, 0, 0, 0, 0, -1, -3, -2, -2, -2, -3, -3, -2, -2, -2, -3, -3, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 2, 0, 1, 0, -2, -3, -1, -2, -1, -3, -2, -1, -1, -1, -2, -2, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -2, 0, 0, -1, -2, -3, -1, -1, -2, -2, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -2, 0, -2, -2, -2, -1, -2, -2, -2, -1, -2, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 1, 0, -1, 0, -1, 0, 0, -1, -3, -3, -3, -3, -2, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, -2, -3, -3, -3, -3, -3, -3, -3, -2, -1, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 1, 1, 1, 0, 0, -1, -2, -3, -2, -3, -2, -3, -3, -2, -1, -1, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -2, -2, -2, -3, -2, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -2, -2, -2, -2, -2, -1, 0, -1, 0, -2, 0, 0, -1, 0, 0, -1, 0, 0, 0, -2, 0, 0, -1, -1, -2, -1, -3, -2, -1, -1, -2, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, -2, 0, -1, -2, -2, -1, -2, -2, -2, -2, -2, -2, -1, -1, 0, 0, -2, -1, -1, -1, -1, -1, -2, -1, 0, -1, -1, -2, -2, 0, 0, 0, -2, -2, -1, -2, -1, -1, 0, 0, 0, 0, -1, -1, -2, -2, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, -2, -2, -1, -2, -2, -2, 0, 0, 0, -1, 0, -2, -2, -1, -2, 0, -1, -1, 0, -1, 0, 0, 0, -2, 0, -2, -2, 0, -1, -1, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, -2, 0, -1, -1, -2, -2, -2, 0, -1, -1, 0, -1, 0, 0, -1, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, 0, -1, -1, -1, 0, -2, -1, -2, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -2, -1, -2, 0, -1, -2, -2, -2, 0, -1, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, -2, -2, -1, -2, -3, -2, -1, -2, -1, -2, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, -2, -3, -3, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, -2, -3, -2, -1, 0, -3, -2, -2, -3, -1, -2, -2, -2, -1, 0, 0, 0, 0, 2, 1, 2, 0, 1, 1, 0, 0, -2, -2, -2, -1, -1, -3, -2, -1, -3, -1, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, -1, -1, -3, -1, -1, -3, -3, -1, -2, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, -2, -3, -2, -1, -3, -3, -2, -2, -2, -3, -2, 0, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -2, -1, -1, -4, -3, -2, -1, -1, -2, -1, -2, -2, -2, -3, -2, -2, -1, -2, -1, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 2, 2, 1, 0, 1, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 2, 1, 1, 2, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 1, 0, -1, -1, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -2, 0, -1, -1, 0, -1, 0, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, -2, -1, -1, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -2, -1, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, -1, 0, -1, 0, -1, 0, -1, -1, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, -2, 0, 0, -1, -1, 0, 0, 0, 0, -1, -2, -2, -2, 0, 0, -1, 0, 0, 0, 1, -1, 0, 0, 0, 0, -2, 0, -2, -1, 0, -2, -1, 0, -1, -1, -2, -1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -2, -1, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, 0, -1, -2, -2, -3, -2, -2, -2, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, 0, -1, -2, -1, -1, -1, -1, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, -1, 0, 0, -1, -2, -2, -2, -2, -1, -1, -2, -1, 0, 0, 1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, -2, 0, -1, -1, -3, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -2, -2, -1, -1, 0, 0, -1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -2, 0, -1, 0, 0, 0, 0, 1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 1, 1, 0, 1, 0, 1, 0, 0, 1, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, -1, 0, 0, -1, -1, 0, 0, -1, -2, -1, -2, -3, -1, -1, -1, -2, 0, -1, 1, 0, 2, 0, 0, -1, 0, -2, -3, -1, -3, 0, -1, -2, -1, 0, 0, -1, 0, 0, -1, 0, -2, 0, -1, 0, 1, 0, 2, 0, 2, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, 0, 0, 0, 1, 0, 0, 1, 0, 0, 2, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 2, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 1, 0, -1, -1, 0, -1, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, -1, 0, -1, -1, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, -2, 0, 0, -2, -2, -3, -2, -1, -2, -1, 0, -1, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -1, -1, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, -1, -1, -1, -1, -2, 0, -2, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, -1, -1, -2, -2, 0, -2, -2, 0, -2, -2, -1, -2, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -2, 0, 0, 0, -1, -2, -1, -1, -1, -2, -2, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, -3, -1, -2, -2, -1, 0, -2, -2, -2, -1, -3, -2, -1, -1, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, -1, -3, -3, -1, -2, -1, -2, -2, -3, -1, -1, 0, -2, -2, 0, -1, -1, 0, 1, 0, 1, 1, 0, 0, -1, -1, -1, -2, -2, -3, -1, -2, -1, -3, -3, -2, -3, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, -1, -2, -2, -2, -2, -3, -2, -3, -3, -3, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -3, -2, -2, -1, -3, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -1, -1, -2, -2, -1, -1, -2, -1, 0, -2, -1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -2, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 1, 0, 1, 1, 2, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 2, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 2, 3, 2, 2, 2, 1, 1, 0, 1, -1, 0, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 2, 1, 2, 1, 1, 3, 1, 0, 1, 1, 0, 0, 1, 1, 4, 3, 1, 2, 2, 1, 1, 0, 2, 0, 1, 0, 1, 0, 0, -1, -2, 0, 0, 1, 1, 1, 3, 1, 0, -3, 3, 3, 2, 1, 1, 0, 0, 1, 0, 1, 2, 1, 0, 0, -2, -2, -2, -3, 0, 0, 0, 0, 2, 2, 1, -3, 3, 4, 2, 1, 0, 1, 0, 2, 2, 0, 0, 0, 0, 0, -1, 0, -2, -2, 0, -2, 0, 0, 1, 0, -1, -2, 4, 3, 2, 2, 1, 1, 1, 0, 2, 1, 0, 1, 0, 0, 0, -1, 0, -2, -1, -1, 0, 1, 1, 0, 0, -4, 2, 1, 2, 1, 1, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 1, 0, 0, -2, 3, 1, 0, 0, 1, 1, 1, 2, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -3, 3, 1, 0, -1, 0, 1, 3, 2, 2, 3, 2, 0, 0, 0, 0, 0, -1, 1, 0, 0, 2, 0, 1, 0, 0, -4, 2, 0, 0, 0, 1, 2, 2, 3, 4, 2, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 2, 1, 0, 0, -4, 2, 0, 1, 0, 1, 2, 3, 4, 3, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 2, 1, 3, 2, 0, -4, 1, 1, 0, 0, 2, 1, 2, 2, 1, 2, 0, -1, 0, 0, 0, 0, 0, -1, 1, 1, 2, 1, 2, 3, 0, -3, 2, 2, 1, 0, 0, 2, 1, 2, 1, 0, 0, -2, 0, 0, 0, -1, 0, 0, 0, 1, 3, 4, 2, 2, 2, -2, 2, 2, 0, 0, 2, 1, 0, 3, 2, 1, 0, -3, -2, 0, 1, 1, 0, 2, 1, 2, 2, 4, 3, 4, 2, -3, 2, 0, 0, 0, 0, 1, 2, 1, 2, 0, -1, -1, -1, 0, 0, 2, 2, 3, 3, 2, 3, 3, 4, 4, 1, -2, 1, 1, 0, 0, 1, 0, 0, 2, 1, 1, -2, -1, -1, 0, 1, 2, 1, 3, 3, 4, 3, 3, 3, 1, 2, -2, 1, 2, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 3, 2, 2, 3, 2, 3, 3, 3, 2, 1, -2, 1, 2, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 2, 0, 2, 2, 3, 2, 0, 2, 4, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 2, 1, 3, 0, -1, 1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 3, 1, 0, -2, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, -1, -1, -1, 0, 0, -2, -1, 0, 0, 0, -1, -2, 1, 0, 1, 0, 0, 2, 2, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -2, -3, -1, -1, -1, -1, 0, -1, -4, 1, 0, 1, 0, 2, 1, 2, 1, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, -1, -1, -1, -1, 0, 0, -1, -3, 2, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, -1, -2, -2, -2, 0, -2, -2, -1, 0, 0, 0, -1, -2, -4, 2, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -3, -1, -2, 0, 0, 0, -1, 0, 0, 0, 0, -1, -5, 3, 1, 2, 1, 0, 2, 0, 0, 0, 1, 1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -6, 2, 2, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -3, -5, 0, 1, 0, 0, 0, 1, 1, 0, 2, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 3, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, -1, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 1, 0, 1, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -2, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, -1, 0, -2, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, -2, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, -1, 0, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, -2, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, -1, -2, -1, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, -2, -1, -2, -1, -3, -4, -3, -4, -5, -3, -4, -1, -3, 0, 0, -3, -3, -7, 2, 3, 1, 1, 0, 1, 1, 0, -1, 0, 0, -1, -1, -3, -3, -3, -1, -3, -2, 0, 0, 0, 1, 0, -2, -5, 2, 2, 2, 1, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, -2, -4, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, -1, -4, 2, 2, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 2, 2, 0, 2, 1, 1, 1, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 2, 2, 1, 2, 2, 3, 2, 1, 3, 1, 2, 1, 0, -2, 0, 1, 0, -2, -1, -2, 0, 1, 0, 1, 1, 0, 1, 0, 1, 1, 2, 3, 3, 3, 2, 3, 2, 0, 0, -3, 0, 1, 0, -2, -2, -1, 0, 0, 2, 1, 2, 0, 1, 1, 0, 1, 1, 3, 3, 2, 3, 2, 2, 1, 0, -3, 0, 0, 0, -1, -1, -1, 0, 0, 0, 2, 1, 1, 0, 1, 0, 1, 1, 1, 3, 2, 3, 4, 4, 2, 1, -1, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, 1, 2, 2, 2, 0, 1, 1, 3, 4, 3, 2, 0, -2, 0, 0, 0, 0, -2, -1, 0, 0, 0, 1, 0, -1, -2, 0, 2, 0, 1, 2, 1, 2, 2, 3, 3, 2, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, -2, -2, -1, 1, 2, 1, 1, 0, 1, 3, 3, 2, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, 1, 0, 0, 2, 1, 1, 1, 2, 0, 1, 0, -2, 2, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, -1, -1, -1, 0, 0, 1, 2, 2, 2, 1, 1, 1, 1, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 2, 1, 3, 2, 1, 1, 1, 2, 1, -2, 1, 2, 0, 0, 0, 0, 0, 1, 1, 0, -1, -1, 0, 0, -1, 1, 1, 2, 2, 2, 2, 2, 1, 1, 1, 0, 2, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, 0, 1, 1, 0, 1, 2, 2, 1, 3, 1, 3, 0, 0, 0, 0, 1, 0, 1, 2, 2, 2, -1, -1, 0, 0, 0, 0, 1, 0, 1, 2, 2, 2, 3, 2, 2, 2, 0, -1, 0, 1, 0, -1, 1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 2, 1, 1, 0, 0, 1, 1, 2, 1, 0, 0, -3, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 1, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 0, 1, 0, 1, 1, 1, 1, 0, 0, 1, 2, 1, 0, 0, -1, -4, 0, 0, 1, -1, 0, 0, 2, 2, 1, 1, 0, 0, 0, 2, 0, 0, 1, 1, 1, 1, 0, 1, 0, -2, -2, -4, 0, 0, 1, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, -2, -5, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 2, 2, 0, 0, 0, -2, -5, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -2, -1, -2, -2, -2, -1, -1, 0, 0, 1, 1, 0, -1, -3, -5, -7, 0, 0, 1, 1, -1, 0, 0, 0, 0, -2, -1, -1, -1, -3, -1, -2, -2, -2, 0, 0, 0, -4, -2, -5, -6, -10, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 1, 0, 1, 1, 1, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -2, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, -1, -1, -1, -1, 0, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -2, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 1, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, -2, -1, 0, -1, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -2, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, -2, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, -2, -1, 0, -1, -1, -2, -2, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -5, -6, -4, -3, -3, -1, -1, -2, 0, -2, -1, -1, -2, -3, -4, -5, -7, -9, -10, -10, -9, -10, -10, -10, -12, -12, -5, -5, -4, -3, -2, -2, -1, -2, -1, -1, -1, -2, -2, -2, -4, -4, -4, -5, -5, -6, -5, -7, -7, -8, -9, -9, -4, -5, -3, -1, -3, -1, 0, 0, 0, -1, -2, 0, -1, 0, -1, -1, -2, -3, -2, -1, -1, -2, -4, -5, -6, -7, -5, -3, -2, -3, -1, -2, 0, -1, 0, 0, 0, 0, -1, -2, -2, -2, 0, 0, 0, 0, 0, -1, -2, -4, -4, -4, -4, -3, -2, -3, -2, -3, -2, -1, -2, -1, 0, -1, 0, -2, -1, -1, -1, 0, 1, 0, 0, 0, 0, -3, -2, -2, -3, -2, -2, -2, -2, -1, -2, -1, 0, 0, -2, -3, -1, -2, -2, -2, -1, 0, 0, 2, 1, 0, 0, -1, -3, -2, -3, -3, -1, -3, -2, -2, -4, -1, -2, -2, -3, -2, -4, -4, -3, -2, -1, 0, 2, 1, 0, 0, -1, 0, -2, -2, -3, -4, -3, -3, -1, -2, -3, -4, -2, -2, -3, -3, -4, -2, -2, -1, 0, -1, 1, 1, 0, 1, 0, 0, -1, -1, -2, -3, -3, -2, -3, -2, -4, -4, -3, -3, -4, -5, -5, -4, -2, -1, -2, -1, 0, 1, 2, 0, 0, 0, 0, -2, -3, -4, -4, -2, -3, -3, -4, -5, -4, -3, -4, -5, -5, -5, -4, -2, 0, 0, 0, 1, 0, 0, 1, 1, 0, -2, -3, -3, -3, -3, -4, -4, -3, -4, -4, -4, -4, -3, -5, -4, -3, -2, -2, 0, 0, 1, 2, 1, 0, 0, 0, -1, -2, -3, -3, -2, -3, -3, -5, -4, -3, -4, -4, -5, -3, -4, -3, -3, -1, -1, 0, 0, 1, 2, 2, 1, 0, -1, -3, -2, -4, -2, -1, -2, -4, -2, -2, -3, -2, -3, -4, -3, -4, -3, -2, -3, -2, 0, 1, 3, 3, 1, 0, 0, -2, -3, -4, -2, -1, -1, -1, -2, -2, -4, -3, -5, -4, -3, -2, -1, -2, -2, 0, 0, 0, 2, 1, 1, 2, 0, -4, -4, -3, -2, -1, 0, -1, -3, -2, -2, -3, -5, -3, -3, -4, -2, -2, -1, -1, 0, 0, 2, 2, 3, 2, 0, -4, -2, -4, -2, -2, -1, 0, -3, -1, -2, -3, -4, -4, -2, -3, -1, -2, -2, -1, 0, 0, 1, 2, 2, 1, -2, -4, -2, -2, -2, -1, -1, -2, -1, -2, -2, -3, -3, -2, -3, -1, -2, -1, -2, -2, -2, 0, 0, 1, 0, 0, -2, -2, -4, -3, -3, -1, -1, -2, -3, -3, -4, -3, -3, -4, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -4, -4, -3, -3, -2, -2, -1, -1, -1, -2, -3, -3, -3, -1, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, -1, -4, -4, -4, -2, -2, -1, -2, -2, -1, -3, -1, -3, -4, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -2, -3, -4, -3, -4, -2, -3, -2, -1, -2, -2, -2, -1, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, -2, -2, -4, -3, -5, -5, -5, -4, -2, -2, -2, -2, 0, -1, -1, -1, -2, -1, 0, -1, 0, 0, 0, -1, 0, -1, -2, -3, -4, -4, -4, -4, -4, -3, -3, -1, -2, -1, 0, -2, 0, -1, -2, -1, -1, -1, -1, -1, -3, -1, -1, -2, -4, -5, -7, -6, -5, -6, -3, -3, -2, -1, -2, 0, 0, 0, -1, -1, 0, 0, -2, -1, -1, -2, -4, -4, -5, -4, -6, -8, -8, -9, -5, -5, -4, -5, -3, -3, 0, 0, -1, -1, -2, -1, -2, -3, -1, -2, -2, -3, -6, -6, -8, -8, -11, -11, -10, -10, -7, -6, -5, -4, -2, -3, -1, -1, 0, -2, -2, -2, -2, -4, -3, -4, -5, -8, -8, -10, -11, -12, -12, -13, -13, -14, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -2, -3, -2, -4, -2, -3, -1, -1, -1, -3, -4, -5, -8, -1, -1, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, -4, -5, 0, 0, -2, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, -4, -2, -2, -2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -4, -2, 0, -1, -1, -1, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 2, 2, 2, 1, 2, 1, 0, 0, -1, -3, -2, -2, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 2, 2, 2, 2, 0, 1, 0, -2, -1, 0, -2, 0, -1, -2, -1, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 3, 3, 3, 3, 1, 0, 0, -2, -1, 0, -1, 0, -2, -1, -1, 0, 1, 0, 0, 1, 1, 0, 2, 1, 3, 1, 2, 3, 4, 4, 2, 2, 1, -2, -3, -2, -2, -1, -1, -1, 0, -1, -1, 1, 1, 0, 0, 0, 2, 3, 2, 3, 2, 3, 4, 4, 3, 1, 1, -2, -2, -2, -2, -1, -2, -2, -1, -2, 0, 0, 0, -1, 0, 0, 0, 1, 1, 2, 1, 3, 4, 2, 3, 3, 1, -2, -2, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, -2, -1, -1, 1, 2, 0, 0, 2, 1, 2, 3, 1, 0, 1, 0, -1, 0, -2, -1, -2, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 1, 2, 1, 3, 1, 2, 1, -2, -2, -2, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 3, 3, 1, 1, 1, 0, -1, 0, -2, -2, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 1, 1, 2, 1, 2, 1, 1, 3, 1, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 2, 1, 3, 0, 0, 0, -1, 0, 0, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 1, 1, 0, 2, 2, 3, 0, 1, -1, -1, 0, -2, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 2, 2, 2, 0, 0, 0, 0, 1, 1, 3, 2, 0, -3, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 0, 1, 1, 1, 1, 2, 0, 0, -2, -2, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 2, 1, 1, 0, -4, -2, -1, -2, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 1, 0, -1, -2, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 1, 1, 1, 0, -4, -1, 0, -2, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 1, 1, 1, 2, 1, 2, 0, 1, -1, -3, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, -1, -5, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -2, -1, -3, -7, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, -1, 0, -2, -2, -2, -2, -2, -4, -5, -5, -7, -1, 0, -2, -1, -1, 0, -1, -1, -1, -1, -1, -2, -3, -1, -3, -3, -2, -3, -3, -4, -4, -5, -6, -8, -10, -9, 1, 1, 2, 1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 2, 1, 0, 1, 0, 1, 0, 0, 1, 2, 3, 2, 2, 1, 2, 0, 1, -1, -2, -2, -2, -1, 0, -1, -1, 0, 1, 2, 1, 3, 2, 0, 0, -1, 1, 3, 2, 4, 2, 1, 0, 2, 1, 0, 0, -2, -1, -3, -2, -1, 0, 0, 0, 3, 3, 5, 4, 2, 1, -1, 0, 2, 2, 3, 2, 0, 0, 1, 0, 0, -2, -1, -2, -2, -2, -2, -1, 0, 1, 2, 2, 3, 5, 2, 0, -1, 0, 1, 2, 3, 3, 0, 0, 0, 1, 0, -1, 0, -2, -2, -4, -4, -1, 1, 1, 0, 2, 3, 3, 3, 2, 1, 0, 1, 2, 3, 3, 0, 0, 1, 0, 0, 0, -2, -2, -3, -3, -4, -3, 0, 1, 1, 1, 1, 3, 4, 1, 0, 3, 3, 2, 2, 4, 0, 0, 0, 0, 0, -1, -2, -3, -2, -3, -2, -1, -1, 0, 0, 1, 1, 1, 1, 2, 0, 3, 2, 2, 3, 5, 0, 0, 0, 0, -2, -3, -3, -2, -3, -3, -2, -2, 0, 0, 0, 1, 3, 2, 0, 1, 1, 2, 3, 3, 4, 6, 0, 0, 0, 0, -3, -4, -2, -4, -2, -2, -2, 0, -1, 1, 2, 3, 4, 1, 1, 0, 1, 0, 1, 2, 5, 5, -1, 0, 0, 0, -3, -5, -3, -2, -2, -1, -2, -2, 0, 0, 1, 2, 5, 1, 0, 2, 0, 1, 0, 1, 4, 4, 0, 0, -1, 0, -3, -3, -3, -2, -1, -1, 0, 0, -1, -1, 1, 1, 3, 3, 1, 3, 1, 1, 0, 1, 2, 4, -2, 0, -1, -3, -3, -4, -3, -3, -1, 0, 0, 1, 0, -1, 0, 1, 2, 2, 3, 3, 2, 0, 0, 0, 1, 5, -2, -2, -2, -1, -2, -3, -3, -4, -1, 0, 0, 2, 1, 0, 0, 0, 2, 3, 2, 2, 1, 0, 0, 0, 1, 5, -2, -1, -1, -1, -2, -4, -4, -3, -2, -1, 0, 3, 1, 0, 0, 0, 3, 4, 2, 2, 2, 2, 0, 1, 2, 3, -2, 0, -2, -2, -2, -4, -5, -3, -1, -2, 0, 2, 2, 0, 1, 1, 2, 3, 4, 3, 2, 2, 0, 1, 2, 3, -1, -1, 0, -1, -4, -4, -3, -2, -2, -1, 0, 1, 2, 0, 1, 0, 2, 3, 2, 3, 2, 1, 0, 0, 0, 3, 0, 0, -2, -2, -2, -3, -3, -2, -3, -1, 0, 2, 1, 1, 1, 2, 2, 3, 3, 4, 2, 1, 0, 0, 1, 3, -1, 0, -1, -3, -4, -3, -2, -1, -2, -2, 1, 2, 0, 0, 0, 2, 2, 3, 4, 3, 3, 2, 0, 0, 1, 0, -1, 0, -2, -2, -4, -3, -2, -1, -2, -3, 1, 1, 2, 0, 0, 2, 3, 5, 4, 4, 2, 0, 2, 0, 0, 0, -1, 0, -2, -3, -2, -4, -3, -1, -3, -3, 0, 2, 0, 0, 1, 1, 3, 5, 3, 3, 3, 3, 2, 0, -1, 0, 0, 0, -1, -3, -1, -3, -3, -3, -3, -1, 0, 0, 1, 1, 0, 2, 3, 4, 4, 4, 2, 3, 1, 1, 0, 2, 1, 0, 0, -2, -2, -3, -2, -2, -2, 0, 0, 0, 0, 0, 1, 3, 3, 5, 5, 3, 3, 2, 3, 2, 0, 2, 1, 0, 0, 0, -2, -2, -2, -3, -1, 1, 0, 0, 0, 1, 0, 1, 3, 5, 4, 3, 1, 2, 2, 2, 1, 2, 0, 0, 0, 0, 0, -1, -3, -1, -1, 0, -1, 0, 1, 2, 3, 1, 2, 4, 3, 3, 1, 2, 2, 3, 1, 3, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 3, 1, 2, 3, 1, 2, 2, 2, 2, 1, 1, 0, 3, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -3, -1, 0, 2, 1, 2, 2, 1, 1, 0, 1, 2, 0, 0, 1, 3, -1, -1, -2, -2, -3, -2, -2, -3, -4, -4, -2, -3, -2, -1, 2, 2, 2, 4, 2, 1, 2, 2, 1, 0, 0, 2, -1, -1, -2, -2, -1, -2, -1, -1, -2, -3, -1, -1, 0, -1, 0, 1, 1, 1, 1, 0, 2, 2, 0, 1, 1, 0, 0, -1, -2, -1, 0, -2, 0, -2, -3, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 0, -1, 0, -1, -1, -1, -1, -1, -3, -2, -1, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 1, 0, 1, 1, 0, 0, -1, -1, -2, 0, -2, -2, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -3, -2, -2, -2, -1, -1, 0, 0, 1, 0, 0, -1, 0, -2, -1, 0, 0, -1, -1, 0, 0, -1, 0, -2, -1, -1, -3, -3, -3, -3, -1, 0, 0, 0, 0, 0, -1, -1, -3, -1, -1, -1, -1, -1, 0, 0, 0, -1, -2, 0, 0, -3, -2, -1, -3, -1, -2, 0, 0, 0, 1, 0, 0, -2, -1, -2, -1, -1, -1, 0, -1, 0, 0, -1, 0, -1, 0, -2, -2, -2, -1, -2, 0, 0, 0, 0, 0, 0, -2, -1, -1, -2, -2, -1, -1, -1, -2, -1, 0, -2, 0, -1, -1, -2, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, -2, -1, -2, -1, -1, -2, -3, -3, -3, -1, -1, -1, 0, -1, -1, -1, -1, -2, 0, 0, -1, -1, 0, -2, 0, 0, -2, -3, -3, -2, -3, -3, -3, -4, -1, -1, 0, -2, 0, 0, 0, -1, -1, -1, -2, 0, -1, -2, 0, -1, 0, -1, -1, -3, -3, -1, -1, -3, -3, -2, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, -3, -1, -2, 0, -2, -1, -2, -1, -2, -3, -4, -4, -4, -3, -1, 0, 0, -1, -1, 0, -1, -1, -1, -2, 0, 0, 0, -2, -2, -1, 0, -1, -2, -3, -2, -3, -2, -3, -3, -2, -2, 0, 0, -1, 0, 0, 0, -2, -1, -1, -2, -1, -1, 0, 0, -1, -2, -1, -1, -3, -3, -2, -2, -1, -2, -2, -2, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, -2, -1, 0, -1, -2, -2, -1, -2, -2, -1, -1, -3, 0, 0, 0, -1, 0, -2, -1, -1, -2, 0, -1, 0, 0, 0, -1, -2, -1, 0, -1, 0, 0, -2, 0, -1, -1, -1, -1, 0, 0, 0, -2, 0, -2, -1, -1, 0, -1, -1, 0, -1, -1, -1, -1, 0, -1, 0, -1, -2, -2, 0, -2, -1, 1, -1, 0, -2, 0, -1, -1, -2, -1, -1, -1, 0, 0, 0, -2, 0, -2, -1, -1, -2, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -2, -2, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, -2, -1, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -2, -1, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, -1, 0, 0, -1, -2, -2, 0, 0, -1, -1, 0, 0, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, -2, -1, -2, -1, -1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -1, -2, -2, -2, -2, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 2, 2, 2, 1, 1, 0, 1, 1, -1, -2, 0, 0, -2, -1, -2, 0, -1, -2, -1, -1, 0, -1, -1, 0, 0, 0, 2, 2, 2, 3, 0, 1, 0, 0, -2, -2, -2, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, -2, -2, -2, -1, -1, -2, -2, -2, -1, -1, -1, -1, -2, -1, -2, -1, -2, 0, 0, -2, 0, 0, -1, 0, -1, -1, -2, -1, -1, -2, -2, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, -2, 0, 0, -1, -1, -1, 0, 1, 0, -1, 0, -1, -1, -2, -1, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 2, 1, 1, 0, 0, 0, -1, 0, 0, 0, -2, 0, 0, -1, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 1, 0, 0, 0, 0, -2, 0, -1, -1, -2, -1, -1, -1, 0, -1, 0, 0, 1, 1, 0, 1, 0, 2, 1, 2, 2, 2, 1, 0, 0, -1, 0, -1, -1, -1, -2, 0, -2, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 2, 2, 1, 3, 1, 0, 0, -2, 0, 0, -2, -2, -2, -2, -1, -1, 0, -2, 0, 0, 0, 1, 0, 1, 1, 3, 3, 2, 1, 3, 2, 1, 0, -1, -1, -1, 0, -1, -1, -2, -2, -1, 0, 0, 0, -1, 0, 0, 0, 2, 2, 2, 3, 2, 2, 2, 1, 2, 0, -2, -2, 0, -1, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, 0, 1, 0, 0, 3, 3, 2, 2, 2, 1, 2, 0, -1, -1, -2, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 2, 1, 2, 1, 2, 2, 1, 0, -1, -2, -1, 0, 0, -1, -2, 0, 0, -1, -1, -1, 0, 0, 1, 2, 0, 0, 0, 2, 1, 2, 3, 2, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -2, -1, 0, 0, 1, 1, 0, 0, 0, 1, 2, 1, 1, 2, 0, 1, 0, -1, 0, 0, -2, -1, 0, -1, 0, -1, -1, -1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 2, 3, 1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 1, 2, 1, 0, 0, 1, 0, 3, 2, 1, 1, 1, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, 2, 1, 2, 2, 2, 0, -1, -2, 0, -2, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 1, 2, 2, 0, 1, -1, -1, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 2, 2, 2, 0, -1, -2, -1, -1, -2, -2, 0, 0, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 2, 1, 1, 2, 0, 0, -1, -1, 0, -1, -1, -2, -2, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, -2, -2, -2, -2, -2, -2, -2, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, -2, 0, -1, 0, -1, 0, 0, 0, -2, -1, -2, -1, -2, -2, -2, -1, -2, 0, -1, -2, -1, 0, -3, -1, -2, 0, -3, -3, -2, -3, -1, -2, -2, -2, -2, -2, -3, -2, -2, -2, -1, -2, -1, -1, -2, -1, -1, 0, -1, -2, -2, -2, -2, -2, -3, -3, -3, -3, -2, -4, -3, -4, 4, 3, 1, 1, 0, 0, -1, -1, -1, 1, 0, 0, 0, -3, -3, -3, 0, 0, 1, 2, 0, 1, 0, -3, -7, -15, 6, 4, 2, 2, 2, 0, 1, 0, 0, 2, 0, 0, 0, -2, -1, -1, -2, -1, 0, 1, 3, 3, 2, 0, -5, -13, 6, 5, 4, 1, 0, 1, 1, 3, 3, 2, 3, 0, 0, 0, 0, -1, -3, -1, 0, 1, 2, 4, 3, 0, -4, -13, 6, 4, 2, 0, 0, 1, 3, 4, 3, 5, 4, 2, 2, 2, 1, 0, -1, -1, -1, 0, 1, 2, 2, 0, -3, -13, 5, 2, 2, 0, 0, 1, 2, 4, 3, 6, 5, 3, 1, 3, 0, 0, -1, 0, 0, 0, 1, 2, 2, 0, -4, -12, 4, 2, 0, -1, 0, 2, 2, 4, 5, 4, 3, 3, 3, 1, 1, 2, 0, 1, 0, 1, 1, 2, 3, 0, -5, -12, 3, 0, -1, -1, 0, 2, 3, 4, 4, 5, 3, 3, 2, 2, 2, 1, 3, 2, 2, 2, 3, 3, 2, 0, -5, -11, 1, 1, -2, 0, 0, 2, 3, 4, 4, 2, 2, 1, 1, 1, 1, 0, 2, 2, 4, 3, 3, 2, 1, 0, -4, -12, 1, -1, -1, -1, 0, 1, 2, 4, 2, 2, 1, 0, 2, 0, 1, 1, 1, 2, 3, 5, 4, 5, 1, 0, -3, -13, 0, 0, -2, 0, 0, 1, 2, 2, 2, 2, 1, 1, 0, 0, 1, 1, 1, 2, 4, 5, 4, 5, 2, 0, -4, -11, 1, 1, 0, 0, 0, 0, 3, 3, 1, 0, -1, 1, 0, 0, 0, 1, 2, 3, 3, 4, 5, 5, 4, 1, -4, -13, 2, 0, 1, 0, 0, 1, 1, 2, 0, -1, 0, 0, 0, 1, 1, 2, 2, 4, 4, 5, 5, 5, 3, 0, -4, -11, 3, 2, 0, 0, 0, 0, 2, 1, 0, -2, -3, -1, -1, 0, 2, 3, 2, 4, 3, 4, 4, 3, 4, 0, -5, -12, 2, 1, 0, 0, 0, 2, 3, 4, 2, -1, -1, -3, 0, 1, 3, 5, 5, 6, 4, 5, 2, 3, 2, 0, -5, -11, 3, 2, 0, 0, 0, 2, 1, 3, 1, 0, -3, -3, -1, 0, 4, 5, 6, 5, 5, 4, 3, 2, 1, 0, -3, -12, 3, 2, 0, 0, 1, 2, 2, 3, 2, 0, -1, -3, 0, 1, 3, 5, 6, 4, 4, 4, 2, 3, 2, 0, -2, -9, 2, 1, 0, 0, 1, 1, 2, 2, 2, 0, -2, -1, 0, 3, 3, 3, 4, 3, 3, 2, 4, 3, 3, 1, -2, -10, 1, 1, 0, 2, 0, 2, 2, 2, 0, 0, -1, -1, 2, 3, 2, 2, 2, 1, 3, 2, 3, 3, 3, 1, -2, -9, 1, 0, 0, 2, 2, 3, 3, 3, 3, 1, 0, 1, 2, 4, 2, 2, 0, 1, 2, 3, 2, 1, 1, 0, -2, -9, 1, 1, 0, 2, 2, 1, 2, 3, 1, 1, 0, 2, 3, 3, 2, 1, 0, 0, 1, 0, 1, 1, 0, 0, -4, -12, 0, 1, 1, 1, 1, 2, 2, 3, 2, 2, 1, 2, 1, 1, 1, 1, -1, 0, 1, 0, 0, 0, 0, -1, -4, -14, 1, 1, 0, 2, 1, 2, 3, 2, 2, 1, 2, 1, 1, 0, 0, 0, 0, -1, 0, -1, -2, 0, 0, -2, -6, -14, 3, 1, 1, 2, 2, 2, 2, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 2, 0, 0, 0, 0, -1, -6, -14, 4, 2, 2, 1, 1, 2, 2, 1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 1, 1, 1, 0, 0, 0, -1, -7, -14, 3, 5, 3, 1, 0, 0, 2, 0, 0, 0, 0, -1, -3, -1, 0, 0, 2, 3, 3, 2, 0, 0, 0, -3, -6, -15, 4, 4, 3, 1, 0, 1, 2, 0, 0, -1, 0, -1, 0, 0, 1, 1, 2, 2, 3, 3, 1, 2, 0, -4, -9, -17, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 2, 1, 0, 0, 1, 0, -1, -1, -1, -1, 0, 0, -2, -3, -3, -2, -4, -3, -3, -3, -1, -1, 0, -3, -5, -5, 3, 3, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -3, -2, -1, -2, -2, -1, 0, -1, 0, 0, -1, -3, -5, 1, 2, 1, 2, 1, 1, 0, 1, 0, 0, 1, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -5, 3, 2, 1, 0, 0, 0, 1, 2, 2, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, -1, -1, -3, 2, 1, 1, -1, -1, 0, 0, 1, 1, 1, 1, 0, 2, 0, 0, 0, 0, 0, 2, 1, 0, 0, 1, 1, 0, -3, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 0, 0, 2, 2, 3, 0, 0, 1, 0, 0, -2, 1, 0, 0, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 2, 3, 3, 3, 2, 1, 0, -1, -3, 0, 0, 0, -1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 4, 3, 3, 2, 1, 1, 0, -4, 0, -1, -1, -2, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 4, 3, 2, 0, 0, 0, -3, 0, 0, -2, -2, -2, -1, 0, 0, 0, -2, 0, -1, -1, 1, 0, 0, 0, 3, 3, 2, 2, 1, 2, 0, -1, -4, 0, -1, -1, 0, -2, 0, -1, 0, 0, -1, -3, -2, -1, 0, 0, 0, 1, 1, 3, 3, 1, 1, 2, 0, -1, -4, 2, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -2, 0, 0, -1, 1, 0, 1, 3, 2, 2, 2, 2, 0, 0, -5, 2, 1, -1, -1, -1, -1, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 1, 3, 1, 2, 2, 1, 0, -2, -2, 1, 1, 0, -1, 0, 0, 0, 0, 0, -1, -3, -2, -1, 0, 0, 0, 0, 1, 3, 2, 2, 0, 1, 0, -1, -2, 0, 0, 1, 0, 0, -1, 0, 0, -1, -2, -1, -2, 0, 0, 1, 0, 1, 1, 3, 2, 2, 1, 2, 1, 0, -1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, 0, 0, 0, 1, 0, 2, 2, 2, 2, 1, 3, 1, 0, -3, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 1, 2, 3, 2, 2, 1, 3, 0, 0, 0, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 3, 3, 2, 2, 1, 0, -2, 1, 0, 1, 0, 1, 0, 1, 1, 1, 0, -1, 0, 0, 2, 1, 1, 1, 0, 2, 2, 2, 1, 1, 0, -1, -2, 1, 0, 1, 0, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, 2, 1, 0, 2, 3, 0, 1, 0, 0, 0, -1, -3, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 0, 1, 2, 2, 0, 1, -1, 0, -2, -3, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, -1, -2, -3, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 0, 0, 0, 0, -1, -2, -5, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 2, 1, 0, 0, 0, 0, -2, -4, 1, 2, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, -6, 0, 1, 0, 0, 0, 1, 0, 0, 0, -2, -1, -1, 0, -1, 0, -1, 0, 1, 0, 1, 0, 0, -1, -2, -4, -6, -7, -7, -6, -6, -5, -4, -5, -3, -2, -3, -3, -4, -4, -4, -5, -4, -6, -9, -9, -9, -9, -11, -12, -11, -12, -13, -6, -6, -4, -5, -5, -4, -4, -3, -1, -1, -2, -1, -3, -4, -4, -4, -3, -4, -4, -4, -6, -5, -7, -9, -9, -9, -6, -5, -5, -5, -5, -2, -2, -1, 0, -1, -1, -1, -2, -2, -2, -2, -2, -2, 0, -2, -2, -3, -4, -5, -8, -7, -6, -5, -5, -5, -5, -3, -2, -2, 0, -1, 0, -1, -3, -3, -1, 0, -1, 0, 1, 1, 0, -2, -3, -4, -4, -5, -5, -4, -4, -4, -4, -3, -1, -2, 0, 0, -1, -2, -2, -3, -2, -1, -1, 1, 3, 3, 1, 0, 0, -2, -4, -4, -3, -5, -4, -4, -3, -4, -3, -1, -2, 0, -1, -1, -3, -1, -1, -1, 0, 0, 3, 3, 1, 0, 0, 0, -2, -1, -4, -5, -4, -3, -2, -4, -4, -3, -3, -2, -2, -2, -2, -2, -1, -2, 0, 2, 3, 3, 2, 0, 1, 0, -1, -1, -3, -5, -5, -3, -4, -4, -4, -5, -4, -3, -5, -3, -4, -4, -1, -1, 0, 2, 3, 4, 3, 1, 1, 1, 0, 0, -5, -4, -5, -5, -3, -6, -5, -4, -5, -5, -4, -5, -4, -3, -3, -2, 0, 2, 3, 5, 3, 3, 3, 2, 0, -1, -4, -4, -5, -5, -5, -6, -6, -6, -5, -6, -4, -4, -4, -2, -1, -1, 1, 1, 5, 4, 5, 2, 1, 0, 0, -1, -4, -5, -5, -5, -4, -5, -5, -6, -5, -5, -5, -4, -5, -4, -1, 0, 1, 2, 5, 6, 4, 4, 4, 2, 0, -1, -4, -3, -4, -3, -4, -5, -5, -6, -5, -4, -4, -3, -3, -4, -1, -1, 1, 2, 3, 4, 6, 5, 3, 1, 0, -1, -4, -3, -3, -4, -2, -3, -4, -3, -3, -3, -4, -5, -4, -4, -1, -1, 0, 1, 2, 4, 6, 5, 2, 1, 1, -1, -3, -4, -2, -4, -3, -2, -1, -3, -4, -5, -5, -4, -4, -3, -2, 0, 0, 0, 2, 4, 4, 4, 3, 2, 1, -1, -5, -3, -3, -2, -3, -2, -1, -3, -2, -4, -5, -5, -3, -3, -1, 0, -1, -1, 2, 3, 5, 4, 4, 1, 0, 0, -4, -3, -3, -3, -2, -2, -1, -3, -3, -4, -3, -4, -3, -2, -1, -1, 0, 0, 0, 4, 5, 3, 2, 1, -1, 0, -4, -4, -3, -3, -3, -2, -3, -3, -2, -2, -2, -2, -2, -1, -1, 0, -1, -1, 1, 3, 4, 4, 2, 2, 0, -1, -5, -4, -3, -2, -2, -1, -2, -3, -2, -2, -2, -4, -2, 0, 0, 0, 1, -1, 0, 0, 4, 5, 4, 0, -1, -4, -5, -4, -5, -4, -4, -2, -4, -2, -3, -3, -1, -2, -2, -1, 0, 0, 0, 0, 0, 1, 4, 4, 1, 0, -1, -4, -4, -3, -4, -4, -3, -4, -2, -2, -1, -2, -3, -2, -2, -1, 0, 0, 0, 0, 1, 2, 4, 3, 2, 0, -3, -3, -5, -4, -6, -3, -5, -2, -2, -2, -1, -3, -2, -2, -2, 0, 0, 0, 0, 0, 2, 3, 1, 3, 0, -1, -4, -5, -4, -4, -4, -5, -4, -3, -3, -2, -1, -1, -1, -1, 0, 0, -1, -1, -1, 0, 0, 1, 0, 1, -1, -3, -4, -5, -4, -6, -5, -5, -4, -4, -2, -2, -1, 0, -1, -1, -1, -2, -2, -2, 0, 0, 0, 0, -1, 0, -3, -4, -5, -6, -6, -5, -5, -5, -4, -4, -2, -2, -1, -1, -2, 0, 0, -2, -3, -2, -1, -2, 0, 0, -2, -5, -5, -6, -8, -8, -6, -5, -6, -6, -6, -4, -2, -1, -2, -1, 0, -1, -2, -1, -2, -1, -3, -3, -5, -6, -6, -9, -9, -10, -11, -11, -7, -7, -6, -7, -5, -4, -3, -2, -1, -1, -2, -3, -4, -3, -3, -4, -7, -8, -8, -8, -10, -12, -13, -14, -13, -14, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -2, -2, -2, -2, -1, -2, -1, -2, -3, -1, -2, -4, -5, -7, -2, -1, -2, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, -1, -1, -2, -1, -1, -1, 0, -2, -2, -3, -4, -5, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -3, -4, -2, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -4, 0, -2, 0, -1, 0, 0, 0, -1, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, -2, -3, 0, 0, -2, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 2, 1, 1, 0, 1, -1, -4, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 2, 0, 1, 0, 0, -1, -2, -1, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 2, 2, 2, 2, 0, 0, -1, -2, -2, 0, -2, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 2, 0, 2, 1, 1, -2, -2, 0, 0, -2, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 1, 2, 2, 2, 2, 1, 0, -2, -4, -2, -1, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, 1, 0, 1, 1, 1, 1, 2, 1, 0, -2, -1, -1, -2, -2, -2, -1, -1, -2, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 2, 1, 1, 2, 0, 0, 0, -1, -3, -1, -1, -1, -1, -1, 0, -1, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 2, 2, 0, 0, -2, -2, -2, -2, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 2, 0, 0, -1, -2, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 1, 0, 0, -3, -1, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, -1, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -2, -1, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, -3, -1, -1, -2, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, -1, -3, -1, -1, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 2, 1, -1, -2, -4, -1, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -2, -4, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 1, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, -3, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, -2, -5, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, -2, -3, -5, -2, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, -2, -4, -4, -5, 0, 0, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -2, -1, -3, -4, -3, -4, -5, -8, 2, 2, 0, 1, 0, 0, 1, 1, 2, 2, 2, 3, 2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 2, 2, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 0, 1, 0, 0, -1, -1, -1, 0, 0, -2, -1, 0, 0, -1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 2, 2, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 3, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, -1, 0, -1, 2, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -2, -1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 2, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, -1, -1, -1, 0, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, -2, -2, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 3, 2, 2, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 2, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, 1, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, -1, -1, 1, 1, 1, -1, -1, 0, 0, 0, -1, 0, -1, -1, -1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, -1, 0, 0, -1, 0, -1, -1, -1, 1, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -2, -1, -2, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 2, 1, 3, 3, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 1, 0, 1, 0, 0, 0, 0, 2, 1, 2, 2, 1, 0, 0, 0, -1, 0, 0, 0, 1, 2, 1, 1, 0, 0, 2, 0, 0, 0, 0, 0, 1, 1, 2, 2, 0, 2, 1, 1, 0, 0, -1, -2, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 2, 1, 1, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 1, 0, 0, -2, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 1, 1, 0, -2, 2, 1, 0, -1, 0, 0, 2, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 2, 0, 0, 0, 1, 1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 2, 1, 0, 0, 0, 0, -3, 1, 0, 0, 1, 0, 0, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 0, -1, -1, 0, 0, 0, 1, 0, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 1, 1, -1, -3, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 1, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 1, 1, 0, -2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 1, 0, 2, 1, 2, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 0, 2, 0, 0, 0, -2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 1, 1, 1, 1, 2, 1, 2, 0, 2, 0, 1, 0, -1, -2, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -3, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, -1, 0, -1, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, -1, -2, 0, -1, 0, 0, -3, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, 0, -1, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 1, 2, 1, 0, 0, 1, 0, 2, 0, 0, -1, 0, 2, 0, 2, 1, 0, 1, -1, -2, -2, -3, -3, -3, -2, -2, -3, -2, -1, -1, -2, 0, 0, -1, -1, -3, -4, 1, 3, 1, 2, 2, 0, 0, 0, 0, -2, -2, -2, -2, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, -2, -2, 0, 2, 1, 0, 0, 2, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 1, 0, 0, -1, 2, 2, 3, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, -1, -1, -1, -1, 0, 0, -2, 2, 2, 2, 2, 1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 0, 1, 1, 0, -1, -2, 0, 0, 0, -1, -2, 1, 2, 2, 1, 0, -1, 0, 0, 1, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, -1, -2, 2, 2, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, -1, 0, 0, -1, 0, 1, 0, 0, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, 0, -1, -1, 0, 1, 1, 2, 2, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, -2, 0, 1, 0, 0, 1, -1, 0, 1, 2, 0, 0, 0, -1, -1, 1, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, -2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -2, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 1, 2, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, -1, 1, 0, 1, 0, 0, 1, 1, -1, 0, -2, 0, 2, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -2, 0, 2, 0, 0, 0, 1, 1, 1, 0, -2, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -3, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -3, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -2, -1, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -2, -4, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -4, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, -2, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, 1, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, -3, -2, -3, -3, -3, -2, -1, 0, 0, 0, 0, 0, 0, -3, -3, 1, 1, 1, 2, 1, 0, 0, 0, 1, 1, 1, 1, 1, -1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, -4, 1, 0, 2, 1, 0, 0, 1, 1, 2, 0, 1, 1, 0, 0, -1, -2, -1, -1, 0, 0, 1, 2, 0, 2, 0, -3, 1, 0, 1, 0, 0, 1, 1, 2, 1, 2, 0, -1, 0, -1, 0, -1, -1, -2, 0, 1, 2, 2, 2, 1, 0, -1, 1, 0, 0, 0, 1, 1, 2, 1, 2, 0, 1, 0, 0, -1, -1, -2, -1, -1, -1, 1, 2, 1, 1, 1, 0, -1, 1, 0, 1, 1, 0, 2, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 2, 1, -1, 2, 0, 1, 0, 1, 0, 2, 3, 2, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 2, 2, 1, 0, 1, -1, 0, 0, 0, 0, 0, 2, 1, 3, 2, 1, 1, 1, -1, -1, -1, 0, 0, -1, 0, 0, 2, 1, 2, 1, 1, -2, 0, 0, 1, 0, 1, 2, 1, 2, 3, 1, 1, 0, 0, 0, -2, 0, -1, 0, 1, 2, 2, 1, 1, 3, 0, -1, 0, 0, -1, 1, 0, 1, 1, 2, 2, 2, 1, 0, 0, 0, -1, 0, -2, -1, 1, 1, 2, 3, 3, 1, 1, -1, 0, 0, -1, 0, 0, 1, 2, 3, 2, 0, 0, 0, 0, -1, -1, -2, 0, 0, 1, 0, 2, 4, 2, 2, 1, -1, -1, -1, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 2, 3, 5, 3, 2, 2, -2, 0, 0, 0, 0, 1, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 3, 4, 5, 4, 2, 0, -1, -1, 0, 0, 0, 1, 2, 1, 2, 1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 3, 4, 3, 5, 4, 1, 0, 0, -1, 0, 0, 0, 1, 2, 2, 0, 0, 0, -2, 0, 0, 1, 1, 1, 1, 1, 2, 3, 5, 5, 3, 3, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 1, 1, 2, 1, 1, 0, 1, 3, 4, 3, 2, 0, -1, -1, -1, 0, 0, 0, 1, 1, 1, 0, -1, -2, 0, 1, 0, 2, 2, 0, 1, 0, 2, 3, 4, 3, 3, 0, 0, -1, 0, 0, 0, 0, 1, 2, 0, -1, -1, -2, 0, 0, 2, 0, 2, 1, 0, 1, 0, 3, 3, 3, 2, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, -1, -2, 0, 0, 1, 1, 0, 0, 2, 0, 0, 1, 1, 2, 4, 2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, -1, -1, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 1, 1, 4, 1, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 0, 0, -1, 1, 1, 0, -1, -2, 0, 0, 0, 1, 1, 1, 1, 2, -2, 0, 0, -1, 0, 1, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, -1, 0, -1, -2, -1, -1, 1, 0, 2, 0, 0, -1, 0, 0, 1, 1, 2, 0, 2, 1, 1, 0, 0, -1, 0, -1, -1, 0, -1, -2, -2, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 2, 1, 1, 0, 1, 1, 1, -1, -1, 0, 0, -1, -2, -1, -3, -2, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, -3, -2, -3, 0, -1, 0, 0, -3, 0, -1, -1, 0, 1, 1, 2, 1, 2, 0, 2, 1, -1, 0, -1, -1, 0, 0, -2, -1, -1, 0, -1, 0, -1, -5, 1, 0, 0, 0, 1, 0, 0, 1, 2, 2, 0, 0, 1, -1, -1, -1, 0, 0, -1, -2, -1, 0, 0, -1, -1, -3, 1, 0, 2, 0, 0, 0, 0, 1, 4, 4, 3, 4, 4, 4, 3, 1, 2, 4, 4, 3, 2, 5, 5, 9, 12, 14, 1, 2, 0, 0, 0, -1, 0, 2, 3, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 5, 7, 11, 0, 0, 1, 1, 0, 0, 0, 2, 2, 1, 0, 0, -1, 0, -1, -1, -2, -1, 0, 0, -1, 0, 1, 2, 5, 10, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, -1, -1, -1, -1, -1, -2, -1, -1, -1, -1, 0, -1, 0, 3, 4, 7, 0, 1, 0, 0, 3, 1, 1, -1, 0, 0, -1, -1, -2, -2, -2, 0, -1, -2, -1, -1, -1, 0, 1, 2, 3, 5, 0, 1, 2, 1, 2, 1, 1, 1, 0, -2, -1, -3, -1, -1, -1, 0, -1, -1, -1, -1, -1, 0, 0, 1, 1, 2, 1, 2, 1, 3, 1, 2, 1, 0, -1, -2, -2, -4, -3, -2, -2, -2, 0, -1, 0, 0, -1, 0, 0, 0, 1, 4, 3, 1, 2, 2, 1, 2, 1, 2, 0, 0, -1, -4, -3, -3, -2, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 3, 2, 3, 1, 0, 2, 1, 0, 0, 1, -1, 0, -2, -2, 0, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, 2, 3, 2, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 2, 2, 0, 0, 1, 1, 4, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 2, 0, 0, 0, 0, 3, 3, 1, 1, 0, 0, 3, 2, 0, 1, 0, 0, -2, -1, -1, -2, -4, -2, -1, 0, 0, 2, 0, 2, 0, 1, 2, 2, 1, 0, 0, 0, 1, 2, 0, 0, 0, 0, -1, -1, -1, -3, -4, -3, -1, 0, 1, 1, 0, 0, 1, 2, 2, 3, 2, 0, 0, 0, 3, 3, 0, 0, 0, -2, 0, -1, 0, -3, -4, -2, -2, 0, 0, 1, 1, 1, 0, 3, 2, 2, 1, 1, 0, 2, 1, 4, 0, 1, 0, -1, -1, -1, 0, -1, -2, -2, 0, 1, 1, 1, 0, 1, 1, 1, 3, 1, 1, 1, 0, 1, 2, 3, 1, 0, -1, 0, -2, -1, 1, 0, -1, -1, 0, 2, 1, 0, 0, 1, 1, 0, 0, 2, 0, 1, 1, 2, 3, 4, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 2, 2, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 1, 4, 1, 1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -2, -1, -1, 0, 1, 3, 5, 1, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, 0, -1, -1, -2, 0, 0, 2, 1, 4, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, -1, -1, -1, -1, 0, -1, 0, -2, -2, -1, -3, -1, 0, 2, 3, 5, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -2, -1, -3, -2, -2, 0, 1, 2, 3, 6, -1, 0, 0, 0, -1, -1, 0, 0, 1, 2, 1, 0, 0, 0, -1, 0, -2, -2, -3, -2, -1, 0, 2, 2, 6, 8, 0, 0, 1, 0, -1, -1, 0, 0, 2, 2, 1, 1, 0, 0, 1, 0, -1, -4, -3, -3, -1, 0, 2, 4, 6, 11, 0, 0, 0, 0, 0, -1, -1, 1, 3, 3, 1, 1, 3, 4, 4, 2, -1, -2, -2, 0, 1, 3, 5, 7, 9, 13, 0, 0, 1, 0, -1, -1, 0, 0, 3, 4, 4, 4, 6, 8, 9, 5, 4, 2, 4, 6, 6, 9, 11, 11, 15, 16, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 2, 1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 1, 0, 0, -1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 2, 2, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 2, 1, 2, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 2, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 1, 2, 2, 2, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 2, 1, 2, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 2, 1, 2, 0, 0, 1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 1, 1, 2, 1, 2, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 2, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 1, 1, 1, 2, 1, 1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, -1, 0, -1, -1, -1, 0, 1, 2, 1, 0, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 1, 1, 1, 1, 1, 2, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, -3, -2, 1, 2, 3, 3, 4, 4, 4, 5, 5, 4, 2, 1, 1, 0, 1, 0, 0, 1, 1, 1, 4, 7, 11, 16, -4, -2, 0, 2, 2, 4, 5, 4, 3, 2, 2, 0, 0, -2, -2, -2, 0, -1, -1, 0, 0, -2, 0, 4, 7, 13, -4, -2, 0, 2, 2, 4, 5, 5, 3, 0, 0, 0, -1, -4, -2, -3, -1, 0, 0, 0, -1, -1, 0, 2, 7, 10, -3, -2, 0, 0, 2, 3, 4, 2, 2, 0, 0, -1, -5, -3, -3, -1, 0, 0, 0, 0, -1, -1, 0, 1, 6, 9, -2, -1, 0, 2, 2, 3, 4, 3, 2, 0, -3, -4, -4, -4, -2, -1, 1, 0, 0, 0, 0, -1, 0, 1, 5, 7, -2, 0, 1, 2, 3, 4, 4, 3, 0, -2, -2, -5, -3, -2, -1, 0, 1, 1, 1, 0, 0, 0, 0, 2, 3, 8, -1, 0, 1, 1, 3, 2, 2, 1, 0, -2, -3, -4, -6, -3, -2, 0, 0, 0, 2, 1, 0, -1, 0, 1, 2, 6, -1, 0, 2, 2, 1, 3, 2, 1, -1, -3, -3, -4, -5, -2, -1, -1, 0, 1, 0, 0, 1, 0, 0, 0, 2, 7, 0, 1, 1, 3, 2, 1, 1, 0, -2, -1, -4, -4, -2, -1, -2, 0, 0, 0, 2, 2, 1, 0, 0, 0, 1, 7, 0, 1, 1, 0, 0, 0, 0, 0, -2, -3, -2, -1, -1, -1, 0, 0, 0, 2, 2, 2, 0, 1, 0, 0, 3, 7, -2, 0, 0, 0, 1, 0, -1, -2, -1, -1, -2, -1, 0, 0, 0, 1, 2, 1, 3, 3, 4, 3, 2, 2, 4, 6, -2, -1, -2, -1, 0, -1, -1, -2, -2, -4, -3, -2, 1, 1, 0, 0, 1, 0, 2, 3, 3, 3, 3, 3, 4, 6, -1, -2, -2, -2, 0, -1, -2, -3, -5, -3, -4, -3, 0, 1, 2, 1, 1, 1, 2, 2, 3, 3, 3, 2, 3, 8, -3, -1, -1, -1, 0, -1, -3, -3, -3, -3, -4, -2, 0, 1, 0, 0, 1, 2, 1, 4, 4, 3, 4, 4, 5, 8, -1, -2, -1, -2, -1, 0, -2, -2, -3, -4, -2, -1, 0, 0, 0, -1, 0, 0, 2, 3, 3, 3, 1, 3, 6, 9, -1, -1, 0, 0, -1, 0, -1, -3, -3, -4, 0, 0, 1, 1, 0, -1, 0, 1, 2, 1, 2, 2, 2, 4, 5, 10, 0, 0, 0, 0, 0, 0, -1, -1, -3, -3, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 3, 1, 2, 4, 5, 10, -1, 0, 0, 0, 0, 0, 0, 0, -3, -1, 1, 2, 2, 0, 0, 0, -1, 0, 0, 2, 2, 3, 2, 3, 5, 9, 0, 0, 0, 1, 0, 0, 0, -1, -3, -1, 0, 2, 3, 0, 0, -2, 0, -1, 0, 1, 1, 2, 1, 3, 4, 8, 0, 0, 1, 0, 2, 2, 0, -1, 0, -1, 0, 2, 2, 0, 0, -2, 0, 0, 0, 2, 1, 1, 0, 3, 5, 8, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -2, 0, 0, 1, 0, 1, 2, 6, 10, -2, -1, 0, 0, 1, 1, 1, 1, 3, 2, 2, 1, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 2, 5, 9, -1, 0, 0, 0, 1, 1, 1, 2, 2, 1, 2, 2, 1, 2, 2, 0, -1, -1, -1, -1, -1, -1, 0, 1, 6, 11, -2, -2, 0, 0, 0, 2, 0, 2, 2, 3, 1, 2, 3, 2, 1, 1, -2, -2, -2, 0, -1, -2, 0, 3, 6, 12, -3, -1, 0, 0, 0, 0, 2, 3, 4, 3, 4, 3, 3, 2, 2, 1, 0, -2, -1, -1, -2, 0, 3, 5, 9, 15, -5, -4, -1, 0, 0, 1, 2, 3, 3, 4, 6, 4, 5, 6, 4, 4, 1, 0, 0, 1, 1, 3, 7, 10, 13, 18, 5, 3, 2, 2, 1, 1, 0, -1, -2, 0, -1, 0, -1, -2, -3, -2, -4, -3, -1, 0, -1, 0, 0, -1, -3, -6, 4, 5, 3, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -3, -1, -2, -2, 0, 1, 0, 1, 1, -2, -4, 4, 4, 4, 2, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -3, -1, 0, 1, 1, 0, -1, -3, 3, 3, 1, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 2, 0, 0, 0, -1, -2, -1, 0, 2, 1, 0, -1, -5, 3, 4, 2, 0, 0, 0, 1, 0, 2, 3, 3, 4, 3, 2, 2, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, -4, 3, 2, 0, 0, -2, 0, 1, 0, 2, 3, 1, 3, 1, 3, 2, 2, 1, 0, 0, 2, 1, 2, 1, 0, -2, -3, 2, 3, 0, 0, -1, -1, 0, 0, 1, 1, 1, 1, 1, 2, 2, 1, 0, 0, 0, 3, 2, 2, 1, 1, -1, -3, 2, 1, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 3, 2, 2, 0, -1, -4, 1, 1, 0, -1, -2, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 3, 3, 1, 0, -3, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, -1, 0, 1, 0, 1, 0, 2, 2, 2, 3, 4, 2, 2, 1, -3, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 3, 2, 4, 1, 1, 0, -5, 3, 2, 0, 0, -1, -1, 0, 1, 0, 0, -1, -1, -2, 0, 0, 0, 1, 1, 2, 1, 1, 1, 2, 0, -2, -3, 2, 4, 2, 0, 0, 0, 0, 0, 1, 0, -1, -2, -2, 0, 0, 1, 2, 1, 2, 1, 0, 0, 0, 0, -1, -5, 2, 2, 2, 0, 0, 1, 1, 0, 1, 1, 0, -1, -3, -1, 0, 0, 2, 2, 2, 1, 2, 1, 1, 0, -1, -3, 4, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 1, 1, 3, 3, 1, 0, 1, 1, 0, -1, -3, 3, 1, 2, 1, 0, 0, 0, 0, 1, 1, 0, -2, -1, -1, 1, 0, 0, 1, 1, 1, 2, 1, 1, 1, 0, -1, 3, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 2, 1, 0, 2, 2, 2, 0, -3, 3, 2, 1, 1, 1, 1, 2, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 1, 0, 0, 0, 1, 1, 0, -1, -2, 0, 1, 0, 2, 2, 2, 1, 2, 2, 2, 0, 0, 2, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -5, 1, 0, 0, 1, 1, 2, 2, 3, 1, 2, 1, 1, 1, 2, 2, 1, 0, 0, -1, 0, 0, 0, 0, -2, -2, -5, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, -1, 1, 0, 0, -1, -1, -2, -5, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -4, -5, 1, 2, 1, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, -2, -2, 0, -1, 0, 0, 1, 0, 0, -1, -2, -2, -5, 3, 3, 3, 0, 1, 0, 0, 1, 0, -1, -1, 0, -1, -2, -3, -1, -1, 0, 1, 1, 0, 1, 1, -1, -3, -6, 4, 3, 1, 2, 1, 1, 0, 0, -1, -2, -1, 0, -2, -2, -1, -2, 0, 0, 1, 0, 1, 0, 0, 0, -3, -6, 3, 2, 1, 2, 0, 0, 0, 0, -1, -2, -1, 0, -2, 0, 0, -1, 0, 0, 0, 1, 1, 0, -1, -3, -5, -7, -5, -3, -3, -1, -1, -2, -2, 0, 0, 0, -2, -1, 0, -2, -2, -3, -2, -3, -4, -6, -5, -6, -8, -8, -11, -13, -4, -4, -3, -2, -2, -2, -1, -1, 0, -1, 0, 0, 0, 1, 1, 0, -1, -2, -2, -2, -3, -3, -4, -7, -7, -13, -5, -2, -1, -2, 0, 0, 0, -1, 0, 0, 1, 1, 2, 0, 1, 1, 0, -1, -1, -1, -1, -2, -3, -4, -7, -11, -3, -4, -1, -1, -1, 0, -1, 0, 0, 1, 0, 1, 1, 2, 0, 2, 0, 0, 0, 0, 1, 1, 0, -1, -4, -8, -4, -3, -2, -2, -2, 0, 0, 0, 0, 1, 1, 2, 2, 2, 2, 1, 0, 1, 0, 0, 1, 0, -1, -3, -4, -6, -2, -3, -2, -2, -1, 0, 0, 1, 0, 0, 1, 1, 0, 1, 2, 0, 0, 1, 0, 0, 1, 0, -2, -2, -4, -7, -2, -2, -2, -1, -1, 0, 0, 0, 2, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, 0, -2, -7, -3, -3, -2, -1, -1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, -3, -7, -3, -2, -2, -1, -1, -1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -2, -6, -4, -2, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -2, -5, -3, -4, -2, -1, -1, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -6, -4, -4, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, -1, 0, -1, 0, 1, 1, 0, -3, -3, -3, -1, -2, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, -2, 0, 0, 0, 0, 0, 0, -5, -3, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, -4, -2, -2, -2, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 2, 1, 0, -4, -3, -1, -3, -1, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, -1, 1, 0, 0, 0, -1, 0, 0, 2, 2, -1, -4, -1, -1, -3, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, 1, 0, -1, 0, 0, 1, 0, 2, -1, -5, -3, -2, -2, 0, 0, 1, 1, 0, 0, -1, -1, -1, -1, 0, 2, 1, 0, 0, -1, 0, 0, 0, 1, 0, -1, -6, -3, -3, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -7, -3, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, -2, -7, -2, -3, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, -1, 1, 0, -1, -4, -9, -3, -3, -2, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, 0, 0, -1, 0, 0, -1, -5, -9, -2, -3, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -1, 0, -2, -5, -7, -10, -3, -2, -3, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, -1, -2, -2, -3, -5, -10, -11, -1, -3, -3, -3, -1, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, -2, -1, -3, -5, -6, -7, -10, -11, -15, -2, -4, -3, -3, -2, 0, 1, 0, -1, -1, -2, 0, 0, -2, -3, -3, -3, -2, -4, -5, -7, -8, -11, -11, -15, -17, 2, 2, 3, 1, 0, 0, 1, 5, 6, 8, 8, 8, 6, 5, 5, 2, 1, 0, 3, 2, 1, 2, 4, 4, 6, 7, 2, 2, 2, 2, 0, 0, 0, 4, 5, 6, 6, 7, 4, 2, 1, 1, 0, -1, 0, 0, -1, 0, 1, 4, 3, 6, 1, 3, 1, 1, 0, 0, 1, 1, 3, 4, 4, 3, 2, 2, 2, 0, -1, -1, -1, -4, -3, -2, 0, 2, 3, 2, 1, 0, 0, 1, 1, 1, 1, 2, 2, 1, 3, 3, 1, 2, 1, 0, -1, -1, -2, -2, -2, 0, 1, 1, 1, 1, 3, 2, 1, 0, 1, 1, 1, 2, 3, 0, 0, 0, 1, 0, 1, 0, 0, -1, -1, -3, 0, 0, 0, 0, 2, 0, 2, 2, 0, 1, 1, 3, 2, 1, 3, 1, 1, 0, 0, 0, 0, 0, -2, -1, -2, -1, 0, 0, 1, 0, 0, 0, 3, 3, 1, 2, 3, 3, 3, 2, 3, 2, 0, -1, 0, -1, 0, -2, 0, -2, 0, 0, 0, 0, 0, 0, 1, 0, 3, 4, 2, 2, 3, 2, 2, 2, 3, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 3, 3, 3, 2, 1, 2, 3, 2, 2, 0, -1, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 1, -1, 3, 4, 2, 1, 1, 2, 2, 3, 1, 1, 0, 0, 0, 0, 0, 2, 1, 1, 1, 1, 1, 0, 1, 1, 1, 0, 2, 3, 1, 2, 1, 0, 1, 1, 0, 1, 0, -1, 0, 1, 2, 1, 2, 3, 4, 2, 2, 0, 0, 0, 0, 0, 3, 1, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 4, 2, 3, 2, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 2, 2, 2, 2, 4, 3, 4, 3, 3, 0, 0, 1, 0, 3, 2, 1, 0, 0, 0, 1, 0, -1, 0, 1, 2, 1, 2, 1, 2, 2, 4, 4, 4, 2, 3, 0, 0, 0, -1, 2, 3, 1, -1, 0, 0, 1, 2, 2, 0, 1, 2, 2, 0, 1, 3, 3, 3, 4, 1, 2, 0, 0, 1, 1, -1, 3, 1, 0, 0, 0, 1, 2, 2, 3, 1, 1, 2, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, -1, 3, 2, 0, -1, 0, 2, 3, 2, 3, 2, 2, 1, 0, 1, 0, 0, 0, -1, -1, 0, -1, -2, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 3, 1, 2, 4, 3, 2, 0, 0, 0, 1, 0, -1, -1, -3, -3, -1, -1, 0, 1, -1, 0, 1, -1, -1, 0, 1, 1, 1, 3, 3, 3, 2, 0, 1, 0, 0, -1, -1, -2, -3, -3, -2, -1, 0, -1, -1, 0, 0, -1, 0, 0, 1, 0, 2, 1, 4, 2, 1, 0, 0, 0, 0, -1, -2, -1, -3, -3, -3, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 1, 2, 0, -1, -1, -1, -1, -2, -2, -2, -5, -4, -3, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 2, 2, 1, 1, 0, 0, -1, -1, -4, -3, -3, -5, -4, -3, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 2, 2, 1, 0, 0, -1, -2, -3, -4, -5, -3, -4, -4, -1, 0, 1, 2, 0, 0, 2, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -3, -4, -4, -2, -2, -2, 0, 0, 3, 1, 1, 0, 1, 0, -1, 0, 0, 0, 1, 2, 1, 2, 3, 3, 2, 2, 0, -1, -3, -1, -1, 1, 1, 3, 4, 4, 0, 0, 0, 0, -1, -2, -1, -1, 1, 2, 3, 3, 6, 7, 8, 6, 3, 1, 2, 2, 1, 2, 5, 4, 5, 5,
    -- filter=0 channel=9
    3, 4, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 3, 3, 2, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, -1, 3, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 4, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 1, 1, 1, 1, 1, 1, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, -1, -1, -1, -1, -2, 0, 0, 0, 1, 0, 1, 2, 0, 0, 1, 1, 0, 0, 2, 0, 0, 0, 1, 0, 1, 0, 1, 0, -1, -1, 0, -1, 0, 0, 1, 1, 1, 0, 0, 2, 0, 1, 1, 1, 0, -1, 0, 0, 2, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, -1, 1, 2, 1, 2, 0, 1, 0, 1, 1, 1, 2, 0, -1, 0, 1, 1, 0, -1, -1, -2, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 2, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -1, 0, -1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 0, 0, -1, -1, 0, -2, -3, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 2, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, -2, 0, 0, -2, 0, 1, 1, 0, 0, 0, 1, 2, 0, 0, 3, 1, 0, 1, 0, -1, 0, 0, 0, 0, -2, -1, -3, -1, -1, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, -1, -1, 0, 0, 0, -2, -2, -2, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -2, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, -1, 0, 0, 0, -2, -2, -1, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, -1, 0, 0, -1, -1, 0, -1, -1, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, -2, -2, -2, -1, 0, 0, 0, 0, 1, 0, 1, 2, 0, 1, 0, 3, 0, -1, 0, 0, 0, -1, 0, 0, 0, -2, -3, -1, 0, 0, 1, 0, 0, 1, 0, 2, 3, 0, 1, 2, 0, 2, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, -2, -1, 0, 0, 2, 0, 0, 0, 2, 2, 2, 0, 1, 2, 1, 1, 1, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 2, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 2, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 2, 0, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 0, 2, 2, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 2, 0, 0, 1, 0, 0, 1, 2, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 2, 2, 1, 1, 1, 0, 0, 3, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 2, 0, 2, 2, 1, 1, 0, 10, 5, 2, 2, 0, 0, 0, 0, -1, -1, -1, -3, -4, -3, -4, -6, -6, -6, -7, -7, -6, -6, -5, -3, -2, -2, 8, 5, 1, 1, 0, -1, 0, 0, 1, 1, 0, 0, -2, 0, -1, -1, -2, -5, -5, -5, -4, -3, -2, -3, -2, 0, 7, 4, 2, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, -2, -3, -1, -2, -2, -1, -3, -1, -3, -2, 6, 3, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 2, 1, 0, 0, -1, 0, -2, -2, -1, -1, -2, -2, 5, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 2, 1, 0, -2, -1, -2, -2, 0, -1, -2, -2, -2, 4, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 1, -1, 0, -1, -1, -1, -1, -2, 0, -1, -2, -2, 0, -1, 0, 0, 0, 1, 1, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -2, -2, -2, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 2, 3, 1, 2, 0, 0, 0, 0, -1, -2, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 3, 2, 0, 0, 0, 1, 0, -1, -2, -2, 0, -1, -2, -2, 2, -1, -2, 0, -1, 0, 0, 0, 2, 0, 2, 2, 1, 0, 1, 1, 0, 1, -1, 0, -1, -1, -2, -1, -2, -2, 2, 1, 0, 0, 0, 2, 2, 3, 2, 1, 2, 1, 0, 1, 2, 3, 3, 2, 0, -1, -2, -1, -1, 0, -2, -1, 2, 0, 0, 0, 0, 2, 2, 2, 4, 1, 2, 1, 0, 2, 1, 2, 4, 3, 0, -1, 0, -1, 0, 0, -1, -1, 2, 0, -1, 0, 2, 1, 1, 2, 4, 3, 2, 2, 1, 3, 1, 2, 2, 3, 0, 0, 0, 0, -1, 0, 0, 0, 2, 0, -1, 0, 0, 0, 2, 2, 2, 2, 2, 1, 2, 3, 2, 2, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 2, 0, -1, -2, 0, 0, 0, 2, 1, 3, 2, 2, 1, 0, 1, 1, 0, 1, -1, -2, -1, -2, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 2, 2, 3, 1, 2, 0, 1, 0, 0, 1, 0, -1, -2, -1, -1, -1, -2, -1, 0, 0, 0, 0, -2, 0, 0, 1, 1, 3, 3, 1, 1, 2, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -2, 1, -1, 0, 0, 1, 0, 2, 1, 1, 0, 1, 2, 1, 1, 2, 2, 1, 0, 1, 0, 0, -1, -1, -1, 0, -2, 3, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 1, 0, 1, 0, 2, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 2, 0, 1, 0, 0, 2, 1, 3, 1, 1, 0, 1, 1, 0, 0, 1, -1, -1, -1, 0, -2, 0, -1, -1, 0, 0, 5, 3, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 1, 1, -1, 0, 0, -1, -1, -2, -2, 0, -2, -1, 5, 2, 2, 1, 0, -1, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, -1, -3, 0, -2, -2, 0, 4, 2, 1, 0, 1, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, -2, -2, -2, -1, -1, -1, -2, 0, -1, 0, 6, 2, 1, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, -2, -2, -1, -3, -1, -3, -3, -2, -2, 0, -1, 0, 5, 3, 1, 2, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -2, -3, -3, -4, -3, -3, -2, -1, -2, -2, -2, -2, 0, 0, 0, 2, 4, 3, 1, 2, 1, 0, 1, 2, 3, 4, 2, 1, 1, 2, 3, 3, 2, 2, 2, 1, 2, 5, 0, 2, 0, 2, 3, 2, 1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 3, 4, 0, 0, 2, 1, 2, 3, 1, 0, -1, -1, -1, -2, -1, 0, 0, -2, 0, -1, 0, -1, -2, 0, -1, 1, 2, 4, 2, 2, 0, 2, 2, 2, 0, -1, -3, -3, -1, -2, -1, -1, 0, -1, -1, -1, -2, 0, -2, -1, -1, 1, 2, 5, 0, 2, 0, 1, 0, 0, 0, 0, -2, 0, 0, 0, -2, 0, 0, 0, 0, -1, 0, -2, -3, -3, -1, 0, 0, 4, 0, 2, 0, 0, 0, -1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 1, 0, -1, -1, -2, -1, -2, -1, -2, 1, 4, 0, 2, 1, 0, -1, 0, 0, -1, -2, -1, 0, -2, -1, 0, 0, 0, 1, 0, 0, -2, -1, -2, -2, 0, 0, 4, 1, 2, 1, 0, 0, -1, -1, -2, -2, -1, -2, -1, 0, 1, 1, 0, 1, -1, -1, -1, -1, -1, -3, -1, 1, 4, 0, 3, 0, 1, 0, -1, -2, -1, -2, -1, -1, 0, 1, 0, 0, 0, 0, 0, -2, 0, -1, -1, -2, -1, 1, 4, 1, 1, 0, 0, 1, 0, -2, -2, -3, -1, 0, 0, 0, 1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, 2, 1, 1, 0, 0, 0, -1, -1, -2, -2, 0, -1, 1, 2, 0, 0, 0, -2, -2, -2, -1, 0, 0, 0, 0, -1, 2, 0, 2, 0, 0, -1, 0, -2, -2, -4, -1, 0, 0, 1, 0, 0, 0, -1, -4, -2, -1, 0, 0, -1, -2, -2, 0, 0, 2, 0, -1, 0, -1, -4, -2, -2, -2, -2, 0, 0, 0, 0, -1, -3, -4, -3, 0, 0, 1, 0, 0, -1, 0, 0, 2, 0, 0, -1, -1, -4, -4, 0, 0, -1, -1, 0, 0, 0, -1, -2, -4, -4, -1, 1, 0, 0, -2, -1, 0, 1, 2, 1, -1, -1, -3, -2, -2, -2, 0, 0, 0, 1, 1, 0, 0, -2, -1, -2, -1, 0, 0, -2, -3, -2, 1, 0, 2, 3, 0, 0, -1, -2, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, -2, -1, 0, -2, -4, -1, 3, 2, 2, 2, 1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 1, 1, -1, -2, -1, -2, -2, -1, -3, -3, -2, 0, 3, 0, 1, 1, 0, -2, -1, -3, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, -2, -1, -2, -3, -3, -3, -3, 1, 4, 0, 2, 1, 0, 0, -2, -3, -2, -2, -1, 0, 1, 1, 0, 0, -1, -1, -1, -2, -1, -1, -2, -4, -3, -1, 4, 0, 1, 0, 1, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -3, -2, -2, 0, 3, 1, 1, 2, 2, 1, -1, -1, -1, -1, 0, 1, 1, 2, 1, 0, -1, -1, -1, 0, -1, -1, -1, -2, -1, 1, 4, 1, 2, 1, 1, 1, 0, 0, -1, 0, 0, 0, 1, 2, 1, 0, 0, -1, 0, -1, -1, 0, -1, -2, -2, 0, 7, 1, 1, 1, 2, 3, 0, 0, 0, 0, 1, 1, 0, 2, 1, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 2, 6, 0, 1, 3, 3, 4, 1, 0, 1, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 2, 6, 0, 0, 1, 3, 4, 1, 2, 0, 1, 0, -1, 0, 0, 3, 2, 0, 0, 2, 1, 2, 3, 0, 0, 1, 2, 6, 0, 1, 2, 3, 4, 2, 2, 1, 0, 0, 0, 0, 1, 4, 4, 1, 2, 4, 5, 5, 3, 3, 2, 3, 5, 5, 0, 0, 0, 0, 0, 1, 2, 2, 1, 2, 2, 1, 0, 1, 2, 2, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 1, 1, 0, 0, 1, 1, 1, 1, 1, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 1, 1, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 1, 1, 0, 2, 2, 2, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 1, 0, 1, 0, 0, 1, 0, 2, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 1, 0, 2, 2, 0, 2, 2, 1, 1, 1, 2, 1, 2, 1, 2, 3, 2, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 1, 3, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 2, 1, 2, 0, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 2, 1, 2, 2, 2, 1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 1, 2, 1, 2, 2, 1, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -2, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, -2, -1, -2, 0, 0, 0, 0, -1, 0, 1, 1, 2, 3, 2, 0, 0, 1, 1, 1, -1, -1, -1, -3, 0, -1, -1, -2, -3, -1, -2, 0, -1, -1, 0, 0, 0, 2, 2, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -2, -2, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 1, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 2, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 2, 2, 1, 0, 0, 0, -1, -1, -1, -1, -1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -2, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 2, 2, 2, 2, 0, 0, 1, 2, 1, 2, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 2, 1, 1, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 1, 2, 2, 2, 0, 0, 0, 0, -1, -1, -1, -1, 0, 1, 2, 2, 1, 0, 0, 0, 0, -1, 1, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 2, 1, 2, 1, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 1, 1, 1, 0, 2, 1, 1, 0, 0, 1, 0, 0, -1, 1, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 1, 1, 2, 1, 2, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 2, 0, 2, 0, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 1, 1, 0, 1, 2, 3, 2, 3, 2, 3, 2, 2, 2, 1, 1, 2, 2, 0, 0, 1, 0, 1, 0, 0, 0, -3, 0, -2, -1, 0, 0, 0, 0, 0, 2, 1, 2, 5, 5, 5, 5, 1, 0, 0, -1, -1, -1, 0, -1, -2, -2, -2, -1, 0, -1, -1, 0, 0, 0, 1, 0, 1, 2, 4, 5, 3, 4, 1, 0, 0, -1, -2, -2, -1, -1, -2, -2, -3, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 2, 3, 3, 2, 2, 0, -2, -1, -3, -4, -3, -2, -2, -2, -2, -1, -2, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 3, 3, 4, 1, 1, 0, -1, -3, -4, -2, -4, -4, -2, -3, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, 1, 2, 3, 3, 2, 2, 1, 0, -1, -2, -3, -3, -4, -3, -3, -3, -2, 0, 0, -2, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 0, 0, 0, 0, -2, -1, -3, -2, -2, -3, -2, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 2, 0, 0, -2, -2, -3, -3, -3, -3, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 3, 2, 3, 1, 1, 0, 0, -2, -1, -1, -3, -4, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 4, 2, 3, 3, 1, 1, 2, 1, 0, -2, -1, -2, -3, -4, -5, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 3, 4, 2, 3, 4, 3, 3, 0, 0, 0, 0, -2, -2, -2, -3, -3, 0, 1, 1, 1, 0, 0, 0, 2, 2, 0, 2, 4, 4, 4, 3, 3, 1, 0, 0, 0, -2, -2, -2, -2, -3, -3, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 3, 4, 3, 2, 3, 4, 3, 0, 0, 0, -2, 0, -2, -1, -3, -4, -1, 0, 0, 2, 1, 2, 0, 0, 1, 1, 2, 3, 2, 3, 2, 3, 3, 2, 0, -1, 0, -2, -2, -2, -2, -2, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 3, 2, 3, 4, 4, 4, 4, 1, 0, -1, -2, -2, 0, -1, -1, -4, 0, 0, 2, 3, 2, 0, 0, 0, 0, 0, 1, 2, 3, 3, 3, 3, 1, 1, -1, 0, -2, -2, -2, -1, -3, -3, 1, 0, 1, 2, 2, 1, 1, 1, 1, 1, 2, 2, 3, 3, 3, 2, 0, 0, 0, -3, -2, -1, -2, -2, -3, -4, 0, 1, 1, 1, 0, 0, 0, 1, 1, 2, 1, 3, 2, 1, 2, 2, 0, 0, -1, -2, -2, -3, -3, -3, -3, -5, -1, 0, 1, 2, 0, 1, 0, 1, 0, 0, 1, 2, 1, 2, 2, 0, 1, 0, -2, -1, -2, -3, -4, -2, -2, -4, -1, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -3, -3, -2, -4, -2, -2, -4, -4, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -2, -1, -2, -3, -3, -4, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -2, -1, -2, -4, -3, -3, -4, -2, -4, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 0, 1, 2, 0, 0, 0, -2, -2, -4, -3, -3, -3, -2, -2, 0, -1, 0, 0, 1, 0, 0, 0, 1, 1, 2, 3, 1, 2, 1, 0, 1, 0, -2, -1, -1, -2, -3, -3, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 3, 2, 2, 2, 2, 1, 0, 0, 0, -2, -2, -2, -1, -1, -3, -2, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 2, 2, 3, 1, 2, 2, 0, 0, 0, -1, 0, 0, -1, -2, -1, -3, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 1, 1, 3, 2, 1, 1, 0, 2, 2, 0, 0, 0, -2, 0, -1, -1, -2, -1, -1, -2, -1, 0, 0, -1, -1, -1, 0, 0, 2, 2, 1, 0, -1, -1, 1, 2, 3, 7, 8, 10, 12, 15, -2, 0, -2, -2, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 2, 1, -1, -4, -3, 0, 0, 1, 3, 7, 7, 12, 0, 0, -1, -2, 0, 0, -1, -2, -2, 0, -2, -2, 0, 1, 0, 0, -2, -4, -4, -4, -3, -2, -1, 1, 5, 9, -1, 1, -1, -1, 0, 1, 0, -1, 0, -2, -1, -1, 0, 0, 1, 0, -2, -4, -6, -5, -7, -7, -4, -1, 0, 6, -1, 0, 1, 0, 2, 2, 1, 0, 0, -1, 0, -1, -1, -1, 1, -1, -3, -6, -6, -7, -6, -8, -5, -4, 0, 4, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, -1, -5, -5, -5, -7, -7, -6, -5, -1, 5, -1, 0, 1, 1, 0, 2, 2, 0, 1, 0, -1, -1, 0, 1, 1, 0, 0, -4, -4, -6, -4, -6, -8, -6, -1, 5, -3, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 0, -1, -4, -5, -4, -5, -6, -6, -2, 5, -3, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 2, 1, -1, -3, -4, -3, -3, -2, -4, -4, -1, 4, -1, -2, -1, -1, -2, 0, 1, 0, 0, 0, 0, 1, 1, 4, 4, 1, 0, -2, -5, -3, -3, -1, -3, -3, -4, 3, -1, -2, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 3, 3, 4, 3, 0, -2, -5, -4, -1, -2, -2, -2, -3, 2, -2, -1, 0, 0, 0, 2, 1, 2, 1, 2, 0, 1, 2, 4, 4, 3, 0, -3, -6, -5, -2, 0, -1, -2, -3, 2, -2, 0, 2, 0, 0, 0, 0, 2, 2, 1, 1, 0, 1, 5, 4, 4, 1, -3, -4, -3, -1, -1, -2, -3, -2, 1, -2, 1, 1, 0, 0, 0, 1, 2, 1, 3, 3, 3, 4, 5, 4, 2, 0, -1, -3, -3, -1, 0, -1, -2, 0, 1, -2, 1, 1, 0, -1, -1, 0, 2, 1, 1, 1, 4, 4, 4, 4, 2, 0, 0, -1, -2, 0, 0, 0, 0, -1, 2, -2, 0, 0, 0, 0, -2, -1, 0, 1, 2, 1, 2, 4, 4, 4, 1, 0, -1, -2, -2, 0, -1, 0, -1, -1, 1, -2, -1, 1, 0, 0, -1, -2, 0, 1, 3, 2, 2, 2, 3, 2, 0, -2, -3, -4, -3, -1, -2, -3, -4, -2, 2, -1, 0, 0, 0, 0, 0, -2, -1, 0, 1, 2, 3, 3, 1, 2, -1, -2, -3, -4, -2, -3, -3, -2, -3, -3, 2, -1, -1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 4, 2, 0, 0, -2, -5, -5, -5, -5, -3, -4, -3, -3, 1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, -1, -4, -3, -5, -4, -4, -5, -4, -2, 2, -1, -1, -1, 0, 1, 0, 1, 2, 1, 0, 1, 1, 1, 1, 1, 0, -1, -4, -4, -3, -2, -3, -4, -3, -4, 3, -1, -1, -1, 0, 0, 0, 1, 0, 2, 1, 0, 0, 1, 1, 1, 0, -1, -4, -2, -5, -4, -4, -4, -5, -3, 2, -2, -2, 0, 0, 1, 0, -1, 2, 2, 1, 0, 1, 2, 2, 0, 0, -3, -3, -4, -3, -4, -2, -2, -4, 0, 5, 0, -1, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 2, 2, 3, 0, -2, -3, -4, -3, -2, 0, -1, -1, 0, 5, -2, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 3, 1, 0, -3, -4, -3, -2, 0, 1, 0, 1, 3, 8, -2, -2, 0, 0, 1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, -2, -2, -1, 0, 2, 3, 5, 5, 8, 11, 19, 12, 6, 1, 1, 0, 2, 0, 0, -1, -2, -4, -6, -6, -4, -6, -6, -8, -9, -6, -5, -5, -6, -3, -1, 0, 15, 8, 4, 1, 2, 3, 1, 2, 1, 0, 0, -1, 0, -2, -1, -2, -2, -4, -3, -5, -4, -5, -3, -2, -1, -1, 12, 8, 3, 2, 1, 3, 1, 2, 1, 2, 0, 0, 0, 0, 1, 0, 0, 0, -2, -2, -3, -2, -3, -3, -4, -1, 11, 4, 3, 2, 0, 1, 3, 2, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, -1, -2, -3, -3, -2, -3, -3, 8, 2, 1, 1, 0, 1, 1, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -2, 0, -1, -2, -1, -2, -3, -3, 4, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, -1, -2, -2, -1, -3, -2, -4, 1, -2, 0, 0, 0, 0, 4, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -3, -3, -2, -2, -2, -2, -2, -1, -5, -2, -1, 0, 0, 1, 1, 0, -2, 0, 2, 0, 0, 1, 0, 3, 0, 0, 0, -2, -2, 0, -1, -2, -1, 0, -2, -3, 0, 0, 0, 0, -1, -1, -3, 0, 1, 1, 0, 1, 2, 1, 0, 0, 0, -1, -2, 0, 0, -1, -2, 1, -3, -3, 0, -1, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -2, 1, 0, 0, 0, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, -3, -1, 0, 0, 0, 0, 4, 0, 0, 2, 0, 2, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 3, 4, 1, -1, -1, -1, 0, 0, 0, 0, 6, 3, 2, 2, 3, 2, 2, 1, 0, 0, -2, -3, -1, 0, 1, 2, 4, 2, 1, 0, -1, -2, 0, 0, 0, 0, 5, 0, 1, 1, 1, 2, 3, 1, 0, 0, -2, -1, 0, 0, 1, 2, 2, 3, 1, 0, 0, -1, 0, 0, 0, 0, 3, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 0, 2, 0, -1, -2, -1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -2, -1, -2, 0, 1, 0, 0, 1, -2, -3, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 0, 2, 2, 1, -2, -2, -1, -1, 0, 0, -1, 2, -1, -3, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 2, 0, -3, -2, 0, 0, 1, 3, 0, 0, 0, 0, 2, 1, 3, 2, 2, 1, 0, 0, -2, -2, 0, 0, -2, -1, 4, 0, -2, -2, 0, 2, 2, 2, 1, 0, 0, -1, 1, 3, 2, 3, 3, 0, 0, 0, -2, -2, 0, -2, -3, -2, 6, 3, 0, -1, 0, 1, 3, 4, 1, 0, 0, 0, 0, 2, 1, 1, 1, 2, 1, -1, -2, -1, -2, -1, -1, -1, 7, 5, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 2, 0, -2, -2, -2, -1, -2, -3, 9, 6, 2, 2, 0, 1, 0, 0, 0, 1, 2, 0, 1, 1, 3, 3, 2, 1, 0, -2, -3, -3, -3, -1, -3, -2, 11, 6, 3, 4, 3, 2, 0, 1, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, 0, -2, -4, -2, -1, -1, -2, -2, 13, 8, 4, 3, 3, 1, 2, 0, -1, 0, 0, -1, 0, -1, 0, 0, -2, -2, -3, -4, -6, -3, -2, 0, -1, -2, 17, 10, 5, 5, 2, 1, 2, 0, -1, -3, -3, -2, -4, -1, -2, -3, -4, -4, -6, -5, -6, -5, -3, -2, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, 0, 0, 0, 0, -1, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 2, 1, 1, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 1, 1, 1, 1, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 1, 0, 1, 1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 2, 25, 15, 9, 4, 1, 0, 1, -1, 0, -3, -4, -8, -9, -10, -9, -10, -10, -11, -13, -12, -10, -7, -4, -4, 0, 5, 21, 11, 5, 2, 3, 2, 0, 1, 1, 1, 0, -1, -3, -3, -3, -5, -4, -7, -7, -7, -6, -6, -4, -2, 0, 1, 18, 11, 5, 1, 1, 1, 3, 2, 3, 2, 1, 0, 0, 0, 0, 0, -3, -3, -5, -5, -5, -4, -5, -4, -2, -1, 14, 8, 5, 3, 0, 0, 2, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -3, -5, -3, -4, -6, -5, -3, 0, 11, 5, 2, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -4, -4, -5, -5, -4, -3, 8, 1, 0, 0, 0, 2, 0, 0, 0, -1, -1, 0, 0, -1, -2, -1, -1, -2, -3, -3, -2, -3, -4, -4, -6, -3, 2, 0, -1, 0, 0, 1, 2, 1, 0, -1, 0, -2, -1, -1, 0, -1, -1, 0, -3, -4, -4, -4, -4, -5, -5, -3, 1, -2, -3, -1, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 1, 2, 1, 0, -3, -2, -2, -3, -3, -3, -2, 0, -2, -2, -2, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 2, 2, 1, 0, -1, -2, -2, -2, -2, -3, -3, -2, 2, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 1, 2, 1, 1, 2, 0, 0, 0, -2, -2, -3, -1, -2, -3, 0, 4, 0, -1, -1, -1, 0, 0, 1, 0, -1, 0, 0, 0, 1, 2, 4, 2, 0, -2, -4, -3, -2, -1, -2, 0, 0, 7, 1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, -1, 1, 2, 3, 4, 2, 0, -3, -2, -2, -1, -1, 0, 1, 7, 1, 0, 1, 2, 2, 2, 3, 3, 0, 0, -1, 0, 1, 4, 4, 4, 5, 1, -2, -3, -1, -3, -1, 0, 1, 8, 0, 0, 0, 3, 3, 3, 3, 1, 0, 0, 0, 0, 2, 4, 5, 4, 2, 1, -2, -3, -3, 0, 0, 0, 3, 4, 0, -1, 0, 1, 1, 2, 0, 0, 1, 0, 0, 1, 1, 3, 2, 1, 1, -2, -2, -2, -3, -1, 0, 0, 2, 4, -3, -4, -2, -1, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 2, 1, -1, -2, -2, -2, -3, -2, 0, 0, 2, 1, -2, -4, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -3, -2, -3, -2, -1, 0, 1, 0, -3, -2, -2, 0, 0, 0, 0, 0, 1, 2, 2, 0, 2, 1, 1, 1, 0, 0, -2, -1, -1, -2, 0, -1, -1, 4, -2, -3, -1, 0, 2, 2, 0, 0, 0, 1, 1, 2, 4, 4, 2, 2, 0, 0, -1, -3, -1, -3, -3, -2, 0, 4, 0, -1, 0, 0, 2, 2, 2, 1, 1, 0, 0, 2, 3, 4, 3, 2, 0, 0, -1, -1, -3, -1, -3, -2, 0, 8, 4, 1, 0, 1, 3, 4, 2, 2, 0, 0, 0, 1, 3, 3, 3, 1, 0, -1, 0, -2, -3, -2, -4, -4, -1, 10, 5, 3, 0, 1, 0, 2, 1, 1, 0, 1, 0, 2, 3, 1, 1, 0, 1, 0, -2, -4, -4, -4, -3, -3, -2, 12, 6, 3, 1, 2, 1, 0, 1, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, -1, -3, -4, -3, -4, -4, -4, -2, 14, 7, 5, 2, 2, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, -2, -1, -3, -3, -5, -5, -4, -3, -2, 0, 15, 10, 6, 4, 3, 1, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, -3, -4, -5, -7, -5, -4, -3, -1, -1, 1, 20, 13, 6, 5, 3, 3, 1, 1, 0, -1, -2, -1, -3, -3, -2, -3, -5, -6, -8, -7, -6, -4, -2, 0, 1, 3, -1, -2, 0, 0, 0, -1, 0, -1, 0, -1, -2, -1, 0, 0, 1, 2, 3, 1, 1, 1, -1, -2, -2, -2, -2, -4, -2, -1, -1, 0, -1, -1, -1, 0, -2, -2, -3, -2, -1, 0, 0, 2, 0, 0, 0, 0, -1, -2, -2, 0, 0, -2, -2, 0, -1, -1, -1, 0, -2, -2, -1, -2, -2, -1, -2, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 1, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, -1, -3, -2, -2, -2, 0, 0, 1, 0, 2, 0, 0, 0, 1, 0, 1, 0, -1, -1, 0, -1, 0, -2, 0, -1, -1, -2, -1, 0, -1, -1, -1, 0, 0, 2, 0, 1, 0, 0, 0, 2, 1, 1, 0, 0, -2, -1, 0, 0, 0, 0, -1, -2, -3, -1, 0, 0, 0, 0, 2, 1, 0, 1, 0, 0, 1, 0, 1, 0, -1, -1, 0, 0, -1, -1, -2, -1, -2, -3, -2, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 1, -1, 0, -1, -1, 0, -2, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, -2, -2, 0, 1, 0, -2, -2, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, -2, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -3, 0, -1, -1, 0, 0, -1, 0, -2, -1, -1, -1, -2, -1, 0, 1, 1, 1, 0, 0, 0, -1, 1, 1, 0, 0, -3, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 1, 1, 2, 0, -1, -1, -1, 1, 0, 1, 0, -2, 0, 0, 1, 0, -1, -1, 0, -1, -2, -2, -1, 0, 0, 0, 1, 2, 2, 1, -1, -1, -1, 0, 1, 2, -1, 0, 0, -1, -1, 0, 0, 0, -2, -1, -2, 0, -2, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 2, 1, 1, -1, -1, 0, 0, -2, -1, -1, 0, -1, -2, -1, -1, -2, -1, 1, 0, 2, 0, 0, -1, 0, -1, 0, 1, 2, 2, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -2, -1, 0, 0, 1, 1, 3, 2, 0, -1, -1, 0, 0, 1, 2, 0, -1, 0, 0, -1, -2, 0, -1, 0, -1, 0, -1, -2, -1, -1, 0, 0, 2, 2, 0, 0, 0, 0, 0, 1, 1, 0, -2, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 2, 2, 0, 0, 0, 1, 2, 2, 1, -2, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 2, 1, 3, 2, 0, 0, -1, 0, 2, 0, 1, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, -1, 0, 0, 1, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, -2, -2, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 2, 1, 2, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, -1, -1, -2, -1, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -2, 10, 4, 3, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, -2, -2, -3, -4, -4, -4, -4, -5, -3, -2, -1, 1, 7, 4, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -1, -1, -3, -3, -5, -4, -4, -4, -2, -2, 0, 6, 4, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, -1, 0, -2, -3, -3, -3, -3, -4, -4, -3, -2, 5, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, -3, -4, -4, -3, -5, -5, -3, -1, 3, 1, 1, 1, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -3, -4, -3, -4, -4, -4, -1, 1, 0, 0, 1, 1, 0, 2, 2, 1, 1, 1, 1, 1, 2, 0, 0, 0, 0, -2, -4, -4, -3, -2, -3, -2, -2, 2, 0, -1, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 0, 1, 0, 1, 0, -2, -3, -3, -2, -2, -2, -3, -2, 0, -1, -2, -1, -1, -1, 0, 1, 0, 0, 0, 1, 1, 1, 2, 2, 0, 0, -2, -3, -3, -4, -3, -3, -4, -2, 1, 0, -2, -3, 0, -1, -1, 1, 0, 0, 0, 0, 0, 2, 2, 2, 0, -1, -2, -3, -4, -2, -2, -2, -3, -2, 3, 0, -2, -2, -2, -1, 0, 1, 2, 1, 0, 0, 2, 4, 2, 4, 3, 1, 0, -2, -2, -1, -1, 0, -2, -1, 5, 2, 0, 0, 0, 0, 2, 3, 2, 2, 1, 1, 1, 4, 4, 5, 4, 2, 0, -1, -1, -2, -2, -1, -1, 0, 5, 0, 1, 0, 0, 1, 0, 3, 2, 2, 1, 1, 3, 4, 5, 5, 5, 3, 0, 0, -1, -2, -1, -1, -1, -1, 3, 1, 0, 1, 1, 0, 1, 1, 1, 1, 1, 2, 3, 5, 5, 5, 4, 2, 0, 0, -3, -3, -3, 0, -1, -1, 3, 0, 0, -1, -1, 1, 0, 1, 2, 1, 2, 3, 2, 4, 3, 3, 2, 0, 0, 0, -3, -3, -2, -2, -2, 0, 1, -1, -3, -1, 0, -1, -1, 0, 0, 1, 0, 1, 3, 2, 3, 2, 0, 0, -1, -1, -2, -2, -1, -1, -2, -1, 1, -1, -4, -2, -2, 0, 0, 0, 0, 1, 1, 1, 0, 1, 2, 2, 0, 0, -1, -1, -2, -2, -2, -2, -1, -1, 2, -2, -2, -3, -2, -1, 0, 0, 1, 2, 1, 0, 2, 2, 2, 2, 1, 0, 0, -2, -2, -3, -2, -2, -2, 0, 3, 0, -1, -1, 0, 0, 0, 1, 0, 1, 1, 1, 2, 2, 3, 2, 0, 0, -2, -3, -2, -3, -3, -3, -3, -2, 4, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 1, 2, 2, 2, 2, 1, 0, -2, -1, -2, -2, -3, -4, -2, -2, 4, 1, 0, -1, 0, 0, 0, 3, 1, 0, 1, 2, 0, 1, 2, 1, 0, -1, -1, -2, -3, -4, -3, -4, -3, -1, 5, 3, 0, -1, -1, 0, 0, 1, 1, 1, 1, 2, 2, 0, 0, 0, -1, -2, -3, -4, -1, -2, -4, -2, -3, -1, 5, 2, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 2, 1, 2, 1, 0, -2, -2, -2, -4, -4, -3, -3, -3, -1, 7, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 0, 0, -2, -3, -3, -3, -3, -3, -3, -2, -1, 7, 5, 2, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -3, -3, -4, -4, -2, -1, 0, -1, 0, 9, 6, 4, 1, 0, 0, 1, 0, 0, 0, 0, -2, 0, -1, -2, -3, -4, -5, -4, -4, -4, -2, -1, 0, 1, 2, 11, 7, 5, 3, 0, 0, 1, 0, -1, -2, -2, -3, -3, -4, -3, -4, -5, -7, -4, -5, -5, -1, 0, 0, 4, 5, 11, 8, 3, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -3, -2, -2, -4, -4, -2, 0, 0, 2, 4, 6, 10, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -3, -2, -3, -1, -1, 0, 2, 4, 7, 5, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, -1, -2, -1, -3, -2, -3, -1, -1, -1, 0, 1, 8, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -2, -3, -1, -1, 0, 0, 1, 6, 3, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, -1, -2, -4, -4, -3, -3, -2, -1, 5, 0, -1, 0, 0, 1, 0, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, -2, -1, -3, -3, -4, -2, -3, -1, 0, 2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, -1, -2, -4, -2, -4, -2, -1, 0, 3, -1, -2, -2, -1, -1, -1, 0, 1, 0, 0, 0, 1, 1, 2, 0, 0, 0, -2, -3, -4, -4, -2, -3, -2, -1, 3, -1, -2, 0, -2, 0, -1, -1, 0, 0, -1, 0, 1, 3, 0, 1, 1, 0, 0, -2, -3, -2, -2, -1, -1, 0, 3, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 2, 1, 2, 2, 3, 2, 1, 0, -1, -1, -1, -2, -1, 0, -1, 5, 0, -1, -2, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 2, 1, 0, -1, -2, -2, -2, -2, -2, 0, 5, 0, -1, -2, -1, 0, 0, 0, 0, 1, 1, 0, 1, 2, 3, 1, 3, 2, 0, -1, -1, -1, -2, -1, -2, 0, 4, 2, -1, -1, -1, 0, 2, 2, 1, 1, 0, 0, 1, 1, 2, 4, 3, 1, 0, 0, -1, -3, -3, -1, 0, -1, 4, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 2, 3, 4, 3, 0, -1, 0, 0, -1, -1, -1, 0, 1, 4, 1, 0, -2, 0, 0, 0, 1, 0, 0, 0, 2, 2, 3, 4, 3, 0, 1, -1, 0, -1, 0, -2, 0, 0, 0, 2, 0, -2, -1, 0, -2, -1, 0, 0, 1, 1, 1, 1, 1, 2, 0, 2, 1, -1, 0, -1, -1, 0, -1, 0, 0, 3, 0, -3, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, 0, 0, -2, -2, -2, -2, -1, -2, -1, 4, 0, -1, -3, -2, 0, 0, 1, 1, 0, 0, 1, 0, 2, 1, 1, 0, 0, 0, -1, -1, -3, -3, -2, -2, -1, 3, 1, -1, -1, -1, -1, 0, 1, 2, 1, 1, 0, 1, 2, 1, 0, 0, 0, -2, -1, -1, -2, -2, -2, -3, -1, 3, 0, -1, -2, -1, -1, 0, 2, 1, 1, 1, 1, 2, 0, 1, 0, 0, -2, -1, -2, -2, -2, -3, -4, -2, -1, 4, 1, 1, 0, 0, 0, 0, 2, 1, 2, 0, 0, 2, 0, 1, 0, 0, 0, 0, -1, -3, -2, -4, -3, -1, -1, 4, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 2, 1, 0, 0, 0, -2, -3, -3, -2, -3, -2, -1, 0, 6, 2, 2, 0, 0, 0, 0, 1, 0, 0, 1, 2, 2, 2, 0, 1, 0, -1, -2, -3, -4, -2, -4, -3, -1, -1, 8, 4, 2, 2, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, -2, -2, -4, -3, -3, -2, -2, 0, 0, 8, 5, 3, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -3, -4, -3, -5, -4, -4, -2, -2, 0, 1, 8, 6, 2, 2, 0, 0, 1, 0, -1, -1, -2, 0, 0, 0, -2, -2, -5, -4, -5, -5, -3, -4, -2, -1, 0, 1, 13, 6, 0, -3, -1, -2, -1, 0, -1, -3, -3, -1, -2, -4, -6, -5, -6, -8, -10, -8, -9, -6, -7, -6, -6, -6, 11, 5, 1, -1, -1, 0, 2, 2, 0, 0, 0, 0, 2, 0, 0, -3, -2, -4, -7, -6, -4, -5, -6, -6, -6, -5, 9, 4, 0, -2, 0, 1, 2, 2, 1, 1, 0, 1, 3, 2, 0, -1, -3, -4, -4, -5, -3, -4, -5, -5, -5, -5, 6, 2, 0, -1, -1, 0, 1, 2, 0, 0, 1, 1, 3, 3, 2, 0, -2, -3, -2, -2, -3, -3, -4, -4, -4, -5, 3, 1, 0, -1, -1, 0, 1, 2, 0, 1, 0, 2, 3, 1, 1, 0, -1, -1, -2, -2, -2, -2, -2, -4, -4, -5, 2, -2, -2, 0, 0, 1, 2, 2, 0, 2, 1, 2, 1, 1, 1, 0, 0, 0, -2, -4, -4, -2, -3, -4, -4, -6, 0, -2, 0, 0, 0, 0, 2, 1, 0, 2, 0, 3, 3, 2, 2, 0, 0, 0, -1, -3, -3, -2, -1, -2, -3, -6, -1, -2, -2, 0, -1, 0, 1, 0, 0, 0, 2, 3, 2, 1, 3, 1, 1, 0, -1, -3, -3, -4, -3, -4, -3, -5, 2, 0, 0, -1, -1, -1, 0, 0, 0, 0, 2, 2, 2, 1, 2, 2, 2, 1, -1, -3, -4, -3, -2, -3, -2, -3, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 2, 4, 4, 1, 0, -2, -3, -2, -2, -2, -3, -3, 4, 2, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 3, 4, 3, 2, 1, -1, -1, -3, -1, -3, -1, -2, 5, 2, 0, 1, 3, 3, 1, 2, 2, 1, 0, 0, 0, 3, 4, 4, 6, 4, 0, 0, -1, -2, -2, -1, -2, 0, 5, 2, 0, 1, 2, 4, 3, 2, 3, 1, 1, 1, 1, 2, 4, 5, 4, 4, 0, 0, -2, -1, -2, -1, -3, -2, 4, 1, 0, 0, 0, 1, 1, 2, 1, 1, 0, 2, 2, 3, 3, 4, 3, 1, 0, -2, -3, -3, -2, -2, -1, 0, 2, -1, 0, 0, 0, 1, 2, 1, 0, 0, 1, 0, 2, 2, 3, 2, 1, 1, -1, -2, -3, -1, 0, 0, -2, -3, 1, 0, -1, -1, 0, 0, 2, 2, 0, 0, 2, 1, 2, 1, 3, 2, 1, 0, 0, -1, -1, -1, -1, -1, -3, -3, 0, -1, -1, 0, 0, 0, 1, 2, 1, 3, 3, 2, 1, 2, 1, 2, 2, 0, 0, 0, 0, -2, -1, -1, -2, -3, 2, -1, -1, -1, 1, 2, 3, 3, 2, 0, 1, 1, 2, 3, 3, 3, 1, 0, 0, 0, 0, -2, -2, -3, -4, -3, 2, 0, -2, -1, 1, 2, 2, 4, 2, 0, 0, 1, 1, 3, 4, 2, 1, 0, -1, 0, -2, -1, -3, -2, -3, -5, 5, 0, -1, -1, 0, 1, 3, 3, 2, 0, 0, 0, 2, 2, 3, 2, 0, 0, -1, -2, -2, -3, -3, -2, -2, -4, 6, 2, 0, 0, 0, 0, 3, 3, 1, 0, 1, 0, 2, 1, 1, 1, 1, 0, 0, -2, -3, -1, -2, -2, -3, -4, 7, 3, 1, 0, -1, 0, 1, 1, 1, 2, 2, 3, 2, 1, 1, 2, 0, 0, -2, -4, -4, -3, -2, -3, -4, -4, 7, 5, 3, 1, 0, 0, 0, 0, 0, 1, 3, 3, 3, 2, 1, 0, -1, -1, -3, -4, -5, -3, -4, -3, -4, -4, 8, 6, 3, 1, 0, 0, 0, 0, 0, 0, 2, 1, 2, 0, 0, 0, -3, -4, -5, -5, -4, -5, -3, -2, -4, -4, 11, 7, 4, 2, 0, 0, 0, 0, 0, -1, 1, 1, -1, -2, -2, -5, -4, -7, -7, -6, -7, -5, -5, -4, -6, -5, 13, 9, 4, 3, 3, 0, -1, -2, -2, -2, -2, -1, -3, -4, -8, -8, -8, -10, -9, -11, -9, -7, -7, -5, -6, -6, 10, 7, 2, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -2, -4, -4, -5, -3, -2, 0, 0, 1, 4, 10, 4, 3, 0, 0, 0, 0, 0, 1, 0, 2, 2, 1, 1, 1, 0, 0, -1, -3, -3, -4, -3, -1, 0, 0, 3, 8, 5, 2, 1, 0, 1, 0, -1, 0, 0, 1, 1, 1, 1, 1, 1, -1, -2, -2, -4, -3, -4, -4, -3, -1, 1, 5, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -3, -4, -4, -3, -4, -5, -3, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, -3, 0, 0, -1, 0, -1, 0, 0, -1, -2, -3, -3, -3, -6, -6, -4, 0, 1, 0, 0, -1, 1, 1, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, -2, -3, -4, -4, -4, -5, -3, -1, 0, -1, -2, 0, 0, 0, 0, 0, -2, -1, -2, 0, -1, 0, 1, 1, 0, 0, -1, -3, -3, -4, -3, -4, -3, -1, 1, -2, -2, -2, -3, -1, -1, -2, -2, -2, 0, 0, 0, 1, 0, 0, 0, -1, -2, -1, -3, -2, -2, -2, -3, 0, 1, -2, -3, -2, -2, -2, 0, -3, -2, -3, 0, 0, -1, 0, 2, 1, 1, -1, -1, -1, -3, -1, -1, -3, -3, 0, 2, 0, -2, -2, -1, -1, -1, -1, -1, -1, -2, 0, 0, 1, 2, 1, 1, 1, -1, -2, -2, -1, -3, -2, -1, 0, 4, 1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -1, 2, 2, 3, 3, 0, -1, -2, -3, -1, -3, -1, -1, 0, 4, 1, 0, 0, 2, 1, 2, 1, 0, 0, -1, 0, 0, 2, 3, 5, 2, 2, 0, -1, -1, -2, -2, -1, 0, 1, 6, 3, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 1, 3, 3, 4, 2, 3, 0, -1, -1, -3, -2, 0, 0, 1, 4, 1, 0, 0, 1, 2, 1, 0, -1, 0, 0, 0, 2, 3, 4, 4, 3, 1, 1, -1, 0, -2, -1, -1, 0, 2, 3, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 1, 2, 4, 3, 3, 2, 0, 0, -2, 0, -1, -1, 0, 0, 3, 1, -1, -2, -1, -1, 0, -1, -2, -2, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, -2, 0, 0, 0, -1, 0, 1, 2, -2, -3, -2, 0, -1, -1, -1, -2, 0, 0, 0, 0, 3, 1, 3, 1, 0, 0, 0, 0, -1, -1, -2, 0, 1, 3, 0, -1, -1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 3, 3, 0, 1, 0, -2, -2, -3, -2, -2, -1, 0, 3, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 3, 1, 0, -1, -1, -1, -3, -2, -3, -2, 0, 4, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 3, 1, 2, 0, 0, -1, -1, -2, -3, -4, -3, 0, 6, 3, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 2, 1, 0, 0, -2, -3, -2, -4, -2, -2, 1, 7, 3, 2, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 2, 2, 2, 0, 0, -2, -4, -4, -4, -3, -3, -3, -1, 8, 5, 1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 2, 2, 2, 2, 0, 0, -2, -3, -5, -3, -4, -3, -1, 0, 7, 4, 2, 0, 2, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, -1, -1, -5, -4, -5, -2, -2, -2, 0, 2, 10, 5, 3, 2, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -2, -3, -3, -4, -4, -3, -1, -1, 0, 2, 4, 12, 7, 4, 2, 1, 0, 0, 0, -1, -2, -3, -1, -3, -2, -2, -3, -4, -5, -5, -5, -3, -1, 0, 1, 4, 6, 6, 2, 0, -1, -2, -1, -1, -2, -4, -4, -5, -4, -3, -4, -5, -5, -6, -7, -8, -8, -7, -6, -4, -5, -6, -3, 6, 3, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, -3, -4, -5, -5, -3, -3, -4, -5, -4, -3, 7, 2, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 3, 4, 1, 0, -2, -4, -3, -3, -3, -2, -3, -3, -3, -2, 6, 4, 2, 2, 0, 1, 0, 1, 0, 1, 2, 2, 2, 4, 3, 1, -2, -1, -2, -3, -2, -1, -2, -3, -3, -3, 4, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 2, 2, 0, -2, -2, -2, -1, -2, -3, -2, -3, -3, 2, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 3, 2, 1, 1, 0, -1, -2, -1, -2, -3, -2, -2, -2, -2, 0, 2, 1, -1, 0, 0, 1, -1, 0, 1, 1, 1, 4, 3, 3, 1, 0, 0, -1, -1, -2, -2, -1, -2, -1, -2, 1, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 2, 2, 3, 4, 1, 0, 0, -2, -2, 0, -2, -2, -1, -2, -2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 3, 4, 2, 1, 0, -1, 0, -2, -2, 0, -3, -4, -4, 3, 0, 0, -2, -2, 0, 0, 0, 0, 0, 1, 2, 3, 2, 3, 5, 2, 2, 0, 0, -1, 0, -2, -2, -2, -4, 4, 0, -1, -1, -3, -2, -1, -1, 0, 0, 0, 2, 2, 5, 3, 4, 4, 1, 1, 0, 0, -1, 0, -2, -1, -1, 4, 1, 1, -1, -1, 0, 0, 0, 1, 2, 0, 1, 2, 3, 4, 5, 5, 3, 1, 2, 0, 0, 0, 0, -1, -1, 5, 2, 0, 0, -1, 0, 1, 2, 2, 1, 0, 1, 3, 3, 4, 5, 5, 4, 2, 0, 2, 1, -1, -1, -1, -1, 5, 2, 0, 0, 0, 1, 0, 0, 0, 1, 1, 3, 2, 4, 5, 6, 6, 4, 0, 1, 2, 0, 0, 0, -2, -1, 3, 1, 0, -1, 0, 0, 0, 0, 0, 1, 4, 3, 4, 4, 4, 4, 4, 3, 1, 0, 1, 0, 1, -1, -1, -1, 2, 1, 0, 0, 0, 1, 0, 1, 1, 3, 4, 4, 3, 4, 3, 4, 3, 2, 2, 1, 1, 2, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 1, 3, 2, 3, 3, 3, 3, 4, 3, 3, 3, 1, 2, 0, 0, 1, 0, -1, -1, -2, 1, -1, 0, 0, 0, 0, 1, 2, 1, 2, 3, 2, 3, 3, 4, 3, 3, 2, 1, 0, 0, 1, 0, -1, 0, -2, 1, 0, -1, 0, 0, 0, 1, 1, 3, 1, 2, 2, 4, 2, 2, 3, 2, 1, 0, 0, 0, 0, 0, -1, 0, -2, 3, 1, 0, 1, 2, 1, 3, 2, 0, 2, 2, 3, 2, 4, 2, 2, 2, 0, 0, -1, 0, 0, 0, -1, 0, -1, 3, 2, 0, 1, 1, 2, 1, 0, 1, 2, 1, 2, 2, 2, 3, 2, 1, 0, -1, -2, -1, -1, 0, -1, -1, -1, 5, 3, 2, 1, 0, 0, -1, 1, 1, 0, 1, 1, 2, 0, 2, 1, 0, -1, -2, -1, -1, -2, -1, 0, -3, -1, 6, 2, 3, 2, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -2, -3, -1, -1, -1, -2, -1, -2, 4, 3, 2, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, -2, -2, -3, -3, -3, -2, -1, -2, -2, -3, 6, 5, 2, 2, 1, 1, 0, 0, -1, -1, 0, 0, 0, -1, -2, -2, -2, -3, -4, -4, -3, -2, -3, -3, -4, -3, 7, 4, 3, 1, 0, 1, 0, -1, 0, -1, -3, -1, -3, -1, -4, -5, -6, -5, -7, -6, -3, -4, -5, -6, -5, -4, 10, 6, 4, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -3, -1, -2, -4, -6, -4, -4, -3, 0, 0, 0, 2, 10, 6, 3, 0, -1, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, -2, 0, -2, -4, -5, -3, -3, -1, -1, -1, 1, 8, 4, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, -2, -1, -2, -1, -2, -4, -4, -2, -3, -3, -1, 0, 6, 2, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, -2, 0, 0, -1, -2, -3, -3, -2, -4, -3, -3, -1, 4, 0, 0, 0, 1, 0, 1, 1, 1, 0, -1, -1, -1, -1, -1, 0, -2, 0, -1, -4, -3, -3, -3, -3, -4, 0, 2, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, -2, -2, -1, 0, -1, -3, -3, -3, -3, -4, -4, 0, 3, -2, -3, 0, -1, -1, 1, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, -1, -1, -4, -4, -3, -1, -2, -1, 0, 2, -1, -2, -1, -1, 0, 0, 1, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, -2, -4, -3, -2, -3, -2, 0, 1, -2, -2, -1, 0, -2, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, -1, -3, -4, -3, -2, 0, 0, -1, 4, 0, -3, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, -2, -2, -3, -3, -1, -1, 0, 3, 1, 0, -1, -1, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 2, 1, 2, 0, -1, -3, -2, -1, -2, -1, 2, 6, 2, 1, -1, 0, 0, 1, 1, 2, 1, 0, -1, -1, 0, 1, 2, 2, 2, 2, 0, -1, -3, -3, -2, 0, 1, 5, 1, -1, 0, 1, 1, 1, 2, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, -1, -3, -2, -2, 0, 1, 2, 4, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, -2, -2, -1, -1, 0, 0, 2, 4, -1, -3, -3, -2, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 1, 3, -2, -4, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, -1, 0, 0, -1, -3, -2, -1, 0, 0, 0, 2, -2, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, -1, -3, -2, -2, 0, 0, 3, -2, -3, -2, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 2, 1, 0, 0, 0, -1, -1, -3, -2, -1, -1, 0, 5, 0, -3, 0, -1, 0, 2, 2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, -1, -3, -2, -1, -2, -2, -1, 6, 1, -1, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -3, -1, -2, -2, 0, 0, 6, 3, 0, -1, -1, 0, 0, 2, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, -1, -3, -3, -3, -1, -1, 0, 7, 3, 1, -1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 2, 0, 1, -1, -3, -2, -2, -2, -2, -3, -1, 0, 7, 4, 1, 0, 0, 0, 1, 0, 2, 2, 2, 0, 0, 0, 1, 1, 0, -1, -2, -2, -3, -3, -3, 0, 0, 0, 10, 5, 2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -3, -4, -3, -3, -3, -2, -1, 1, 0, 11, 6, 3, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, -1, -3, -5, -5, -6, -4, -4, -2, 0, 2, 3, 12, 9, 4, 2, 0, 0, 0, -1, -1, -2, -4, -3, -4, -4, -4, -6, -5, -6, -8, -7, -5, -3, -1, 0, 1, 4, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, 1, 1, 0, 0, -1, -1, 0, -1, -1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, -1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 3, 2, 0, 0, 1, 1, 0, 0, -1, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 2, 1, 1, 0, 2, 0, 1, 0, -1, -1, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 1, -1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 1, 1, 1, 0, 0, -1, 2, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, -1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 2, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 2, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, -1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 1, 0, 1, 0, 0, 1, 1, 0, 2, 0, 1, 1, 0, 0, 1, 0, 1, 1, 1, 0, 0, -1, 2, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 3, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 3, 2, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 3, 1, 2, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, 1, 2, 1, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 1, 1, 0, 0, 0, -1, 1, 0, 0, 1, 0, 2, 2, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 3, 1, 2, 1, 0, 0, 0, -1, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 3, 1, 0, 0, 0, -1, 0, 0, 0, -2, -1, -1, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 2, 0, 0, -1, -1, 0, -1, -2, -3, -1, -1, -1, 1, 1, 1, 0, 0, 0, 0, -2, -1, -1, -2, 0, 0, 1, 0, 1, 0, 0, -1, -2, -2, -2, -3, -3, -1, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -1, -2, -1, 0, -1, -1, 0, 0, 0, 0, -1, -2, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, -3, -3, -2, -1, -2, -2, -1, 0, 0, 0, 0, -2, 0, 0, 0, 1, 0, 1, 2, 1, 2, 2, 0, 1, 0, -1, -1, -3, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, -2, -1, -2, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 1, 1, 3, 1, 2, 0, 0, 0, 0, 0, -3, -2, -1, -1, -1, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 2, 3, 2, 1, 2, 0, 1, 1, 0, -1, -2, -1, -3, -1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 2, 2, 2, 3, 2, 2, 1, 1, 0, 0, -1, 0, -2, -2, -1, 0, 0, 1, 2, 1, 2, 0, 1, 0, 0, 0, 0, 1, 2, 3, 2, 3, 1, 1, 0, -1, 0, 0, -1, 0, -1, 1, 1, 2, 0, 1, 1, 1, 1, 0, 1, 2, 2, 1, 3, 3, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 0, 2, 2, 1, 1, 0, 0, 1, 1, 1, 2, 3, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 2, 0, 1, 0, 0, 0, 0, 2, 2, 1, 2, 3, 2, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 1, 2, 3, 1, 3, 2, 1, 0, -2, -1, -1, 0, 0, 0, -2, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 2, 1, 1, 0, 0, -1, -1, 0, -2, 0, 0, 0, -1, -1, 0, -1, 0, 1, 1, 1, -1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, -1, -1, -2, -2, -2, -1, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, -1, -2, 0, -1, 0, 0, 2, 2, 0, 0, 0, 0, -2, -2, -3, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, -2, -2, -2, -3, -2, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, -1, -1, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, -2, -1, -1, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 3, 1, 0, 0, 0, -1, 0, -1, -1, -1, -2, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, 1, 0, 1, 2, 1, 2, 2, 0, 0, 0, 0, -1, -1, -2, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 1, 3, 2, 1, 1, 0, 0, 0, 0, 0, 0, -2, 0, -1, 6, 7, 8, 5, 2, 2, 0, 1, 0, -2, -3, -5, -4, 0, 1, 2, 1, 0, -1, 0, -1, -3, -3, -1, 0, 0, 5, 6, 5, 1, 0, 0, 0, 0, -1, -1, -3, -3, -1, 1, 2, 1, 0, 0, 0, 0, -1, -1, -1, -1, 2, 2, 3, 5, 3, 0, 0, 0, 3, 3, 1, 0, 0, 0, 1, 2, 1, 2, 2, 2, 2, 1, 0, 0, 0, 0, 0, 1, 5, 3, 2, 2, 2, 3, 3, 3, 1, 0, 0, 1, 2, 1, 1, 3, 3, 2, 3, 1, 0, 0, 0, 1, 0, -1, 5, 5, 2, 1, 2, 3, 3, 3, 1, 0, -2, 0, 1, 2, 2, 3, 3, 2, 2, 1, 0, 0, 0, 0, 2, 0, 7, 2, 2, 1, 0, 1, 2, 0, 0, -2, -2, 0, 0, 1, 3, 2, 0, 2, 1, 1, 2, 1, 1, 0, 1, 0, 5, 1, 1, 1, 0, 2, 2, 1, 0, 0, -2, -2, 0, 0, 1, 0, 0, 3, 4, 3, 4, 2, 1, 0, 2, -1, 3, 0, 1, 2, 1, 3, 3, 3, 1, 0, -1, -1, 1, 1, 1, 2, 4, 6, 7, 5, 4, 1, 1, 1, 1, -1, 1, 0, 3, 2, 3, 4, 3, 2, 1, 0, 1, 1, 3, 2, 3, 4, 6, 7, 7, 5, 3, 1, 0, 0, 0, 0, 0, 1, 3, 2, 4, 2, 1, 3, 2, 2, 2, 4, 4, 5, 6, 5, 3, 4, 5, 4, 2, 0, -1, 0, 3, 0, 1, 3, 2, 1, 2, 0, 1, 1, 3, 3, 4, 5, 4, 4, 4, 3, 2, 4, 5, 4, 1, 0, -2, 0, 0, -1, 2, 0, 3, 0, 0, 0, 0, 3, 4, 3, 4, 3, 2, 2, 4, 3, 4, 5, 6, 4, 2, 1, 1, 1, 1, 0, 4, 1, 2, 0, 1, 1, 1, 2, 3, 3, 3, 2, 1, 1, 4, 3, 6, 5, 5, 2, 2, 2, 1, 3, 2, -1, 3, 1, 4, 2, 2, 3, 4, 3, 4, 4, 1, 1, 2, 1, 4, 5, 7, 6, 4, 3, 2, 0, 2, 2, 2, 0, 6, 5, 6, 3, 3, 3, 4, 3, 2, 2, 3, 3, 3, 4, 6, 8, 7, 6, 3, 1, 0, 0, 0, 3, 0, -1, 6, 3, 4, 4, 1, 3, 3, 2, 1, 2, 3, 4, 4, 6, 5, 7, 5, 1, 0, 0, -3, 0, 1, 3, 1, 0, 5, 2, 1, 0, 1, 2, 1, 0, 0, 2, 3, 4, 4, 3, 4, 3, 1, 0, -2, -3, -3, 0, 2, 3, 2, 1, 4, 2, 0, 0, 0, 1, 2, 1, 1, 1, 3, 1, 0, 1, 3, 3, 2, 0, -1, -1, -1, 0, 1, 2, 1, 0, 4, 0, 1, 0, 0, 2, 2, 2, 1, 2, 2, 1, -1, 0, 4, 4, 3, 2, 1, 1, 1, 0, 0, 2, 0, -1, 2, 2, 1, 1, 1, 3, 3, 3, 0, 2, 1, -3, -3, 0, 2, 3, 3, 2, 2, 1, 1, 3, 2, 1, 2, 0, 3, 1, 1, 0, 1, 2, 2, 1, 2, 1, -1, -1, 0, 1, 2, 3, 2, 1, 1, 2, 1, 1, 1, 3, 1, 0, 2, 1, 0, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 2, 1, 1, 0, 1, 2, 0, 1, 3, 1, 0, 0, 2, 1, 0, -2, -1, -1, 1, 0, 0, 1, 1, 2, 3, 2, 2, 0, 0, 1, 0, 0, 0, 1, 3, 2, 0, 0, 1, 1, -2, -2, -3, 0, 2, 0, 0, 0, 1, 0, 2, 2, 1, 0, -1, 0, 0, 0, -2, 2, 2, 1, 0, 2, 1, 0, -1, -1, 0, 3, 3, 3, 0, 0, 1, 2, 2, 2, 1, 0, 0, -1, 0, -3, -3, 1, 0, 1, 0, 1, 3, 0, 1, 0, 2, 4, 5, 5, 4, 3, 2, 4, 4, 2, 3, 2, 0, 0, -1, -4, -6, 0, 1, 1, 0, 0, 0, 0, 1, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -1, 0, 1, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 7, 5, 2, -1, 0, 0, 0, -1, -1, -1, -4, -4, -3, -2, -3, -5, -4, -6, -7, -5, -3, -3, -1, 1, 1, 3, 6, 2, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -2, -3, -5, -6, -4, -4, -4, -1, 0, 1, 2, 7, 3, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, -1, -1, -3, -5, -5, -4, -4, -4, -2, -1, 1, 3, 1, 1, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 2, 0, -1, -2, -3, -3, -3, -4, -4, -4, -4, -2, -1, 2, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 0, -2, -2, -3, -5, -4, -4, -4, -4, -3, -1, 1, 0, 0, 0, 0, 1, 1, 2, 2, 0, 1, 1, 1, 2, 1, 1, -1, -3, -3, -4, -3, -5, -6, -5, -4, -2, 2, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 2, 2, 2, 3, 1, -1, -1, -3, -4, -4, -5, -3, -5, -3, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 2, 3, 0, -2, -3, -4, -4, -4, -3, -3, -2, -2, 1, 0, 0, -2, -1, 0, 0, 0, 0, 1, 0, 1, 2, 3, 2, 4, 1, -1, -1, -4, -3, -4, -4, -3, -3, -1, 2, 0, 0, -1, -1, -2, 0, 0, 0, 0, 1, 1, 4, 4, 2, 4, 2, 1, -1, -2, -2, -3, -3, -3, -3, -2, 3, 0, 0, 0, -1, 0, -1, 0, 1, 1, 2, 3, 1, 4, 3, 3, 2, 0, 0, -2, -2, -2, -2, -2, -2, 0, 2, 1, 0, 0, 0, 0, 0, 0, 1, 3, 2, 2, 1, 4, 5, 5, 4, 2, 0, 0, -3, -3, -1, -3, -2, 0, 2, 2, 0, -1, 0, 0, 0, 2, 1, 2, 0, 1, 2, 5, 6, 6, 4, 1, 0, -1, -1, -1, -2, -1, -2, 0, 3, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 2, 3, 4, 5, 4, 2, 2, 0, 0, -3, -1, -2, -2, -2, -1, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 3, 4, 4, 3, 3, 1, -1, -1, -2, -2, -1, -1, -2, 0, 1, 0, -1, -1, -1, -1, -1, 1, 1, 0, 0, 2, 2, 3, 3, 2, 1, -1, -2, -3, -3, -1, -1, -2, -1, 0, 1, -1, -2, -1, -2, -1, 0, 0, 2, 2, 2, 2, 1, 3, 2, 2, 0, -1, 0, -1, -3, -3, -1, -1, -4, -1, 0, -1, -1, -2, -1, 0, 0, 0, 2, 2, 1, 2, 2, 1, 2, 0, 0, -2, -1, -4, -2, -3, -2, -3, -3, -2, 1, 0, -2, 0, -1, 0, 1, 2, 1, 1, 2, 1, 3, 2, 1, 0, 0, -2, -4, -4, -5, -3, -2, -4, -2, -3, 3, -1, -1, 0, 0, 0, 1, 2, 3, 0, 2, 2, 2, 2, 2, 1, 0, -1, -2, -3, -4, -4, -5, -4, -4, -1, 3, 0, 0, 0, 0, 1, 1, 2, 2, 2, 3, 2, 4, 2, 2, 0, 0, -2, -2, -4, -3, -4, -4, -3, -4, -2, 3, 2, 0, 0, 0, 0, 1, 2, 2, 3, 3, 2, 2, 2, 1, 0, -1, -1, -2, -4, -3, -5, -3, -3, -3, -2, 3, 2, 1, 0, 0, 0, 0, 1, 2, 1, 3, 3, 3, 2, 1, 2, 0, -1, -4, -4, -4, -4, -5, -4, -3, -1, 5, 2, 1, 0, 0, 0, 0, 2, 0, 1, 2, 3, 2, 2, 2, 0, -1, -3, -4, -4, -4, -4, -4, -2, -3, 0, 6, 2, 1, 1, 0, -1, 0, 0, 0, 1, 1, 1, 2, 1, 1, 0, -2, -3, -6, -6, -4, -4, -3, -2, -2, 0, 6, 4, 1, 1, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -2, -4, -3, -5, -5, -4, -3, -2, -2, 0, 1, 2, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 2, 1, 4, 3, 3, 4, 3, 1, 0, 0, -2, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 2, 3, 3, 2, 3, 3, 0, 0, 0, -2, -2, -2, -1, -2, -4, 0, -1, 1, 1, 0, 1, 0, 1, 1, 1, 0, 0, 3, 3, 1, 0, 1, 0, 0, -1, -1, -3, -1, -1, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 0, 2, 0, 0, 0, 0, -3, -2, -2, -1, -1, -2, -1, 0, 0, 1, -1, 0, 0, 0, -1, 0, -1, 1, 1, 2, 1, 0, 0, -1, 0, -1, -1, -1, 0, -2, -1, -2, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 2, 3, 3, 3, 0, 2, 0, 1, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 2, 4, 4, 2, 2, 1, 1, 0, 1, -1, 0, -1, 0, -2, -1, 0, 1, 2, 0, 0, 0, 2, 2, 0, 0, 2, 3, 5, 5, 3, 2, 1, 2, 2, 0, -1, -2, -2, 0, -1, -1, 0, 2, 2, 2, 2, 0, 1, 1, 1, 1, 3, 4, 3, 5, 5, 4, 3, 2, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 2, 3, 1, 2, 3, 2, 2, 3, 3, 4, 5, 4, 4, 4, 2, 2, 0, -1, 0, -2, -1, -1, 0, -1, 0, 2, 3, 3, 1, 2, 3, 1, 1, 2, 2, 3, 3, 4, 4, 4, 4, 1, 1, 0, -1, -1, -1, 0, 0, -1, 0, 1, 1, 1, 2, 2, 2, 1, 1, 2, 3, 2, 4, 3, 2, 5, 3, 3, 0, 0, -1, -1, 0, -1, 0, -2, 1, 1, 3, 3, 1, 3, 1, 0, 0, 1, 3, 3, 4, 4, 2, 3, 4, 0, 0, 0, 0, -1, 0, 0, -1, -2, 0, 1, 1, 1, 1, 3, 2, 0, 1, 0, 1, 3, 3, 3, 3, 4, 2, 1, -1, 0, -1, 0, -1, 1, 0, -2, 0, 1, 3, 2, 3, 2, 2, 0, 0, 0, 3, 3, 3, 4, 3, 4, 2, 1, -1, -2, 0, 0, -1, -1, 0, -1, 0, 0, 0, 2, 3, 3, 2, 0, 0, 1, 0, 2, 2, 1, 2, 2, 1, 0, 0, -1, -1, -2, -2, -2, -1, -2, 0, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 1, 1, 0, 1, 2, 1, 0, 0, -1, -2, -2, -2, 0, -2, -2, 0, 1, 0, 1, 0, 2, 2, 1, 0, -1, -1, 0, 1, 0, 1, 1, 1, 0, 0, -1, -1, -3, -1, -1, -3, -3, -1, 0, 1, 0, 1, 0, 2, 1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, -1, -2, -1, -1, -1, 0, 0, 1, 0, 0, 1, 0, 1, -1, 1, 0, 0, 1, 0, 2, 0, 0, -1, 0, 0, -2, -1, -2, -1, -2, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 1, 0, 2, 1, 2, 0, 0, 1, 0, -1, -2, -2, -1, -1, -1, -1, 0, 0, 1, 2, 0, 1, 1, 1, 0, 0, 2, 1, 3, 3, 2, 0, 1, 0, 0, 0, -1, -1, -1, -1, -2, -3, 0, 0, 0, 1, 1, 0, 1, 2, 0, 0, 1, 3, 2, 2, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -1, -1, 0, 1, 0, 1, 1, 2, 1, 0, 1, 3, 2, 3, 3, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -3, -3, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 2, 1, 1, 3, 3, 3, 1, 1, 0, 0, 0, 0, -2, -2, -3, 6, 2, 1, 0, -2, -3, -2, -3, -1, -2, 0, 0, 1, 1, 1, 0, 0, -3, -5, -2, -1, 0, 3, 5, 5, 11, 5, 1, 0, -1, 0, -1, -2, -3, -2, -1, 0, 0, 0, 1, 0, -1, -2, -4, -6, -6, -4, -2, -1, 0, 3, 7, 4, 1, 0, -1, -1, 0, -2, -2, -2, -1, -2, -1, -1, 0, 0, -2, -2, -3, -7, -7, -5, -6, -5, -3, 0, 3, 5, 1, 1, 0, 0, 0, -1, -1, -1, 0, -2, 0, 0, 0, 0, -2, -3, -5, -6, -8, -8, -9, -8, -5, -2, 1, 4, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -2, -4, -6, -8, -7, -8, -6, -6, -5, 1, 2, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, -3, -4, -6, -7, -8, -7, -7, -5, 0, 0, 0, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 2, 0, 1, -2, -3, -4, -6, -7, -6, -6, -7, -4, 0, 0, -1, -2, -3, -3, -1, -1, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, -3, -5, -6, -6, -5, -6, -5, -4, 0, 1, -1, -3, -4, -3, -1, 0, 1, 0, 0, 1, 1, 2, 1, 3, 1, 0, -2, -4, -5, -6, -5, -5, -5, -3, 1, 1, 0, -3, -2, -3, 0, 1, 2, 1, 0, 0, 1, 0, 4, 2, 3, 2, -2, -4, -5, -5, -4, -4, -4, -2, 0, 2, 0, -1, -2, 0, 1, 0, 1, 1, 2, 2, 1, 0, 4, 4, 5, 2, 1, -2, -4, -5, -4, -2, -2, -1, 2, 4, 0, 0, -1, 0, 0, 1, 1, 2, 3, 2, 1, 2, 5, 7, 5, 4, 0, -1, -3, -3, -3, -3, -3, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 3, 4, 5, 7, 4, 2, 1, -1, -3, -4, -2, -3, -2, -1, 3, 2, 0, -2, -2, -1, -1, 0, 0, 0, 1, 3, 2, 3, 4, 4, 3, 1, 0, -3, -3, -2, -3, -3, -2, -1, 3, 0, -2, -2, -2, -2, -1, -3, -1, 0, 0, 2, 2, 4, 4, 2, 0, 0, -2, -1, -2, -2, -4, -2, -3, 0, 2, 0, -2, -3, -3, -3, -4, -2, -1, 0, 1, 0, 3, 2, 3, 3, 1, 0, -1, -4, -3, -2, -5, -3, -4, -3, 0, 1, 0, -3, -1, -1, -2, -1, -1, 0, 2, 3, 3, 2, 2, 2, 1, -2, -3, -3, -5, -3, -4, -6, -4, -3, 0, 3, 0, -1, -3, -2, -1, 0, -1, 0, 1, 1, 1, 2, 1, 0, 0, -1, -3, -4, -5, -7, -5, -5, -4, -5, 0, 2, 1, -2, -2, 0, -1, 0, 0, 0, 0, 1, 0, 3, 1, 0, -1, -2, -2, -4, -7, -6, -6, -7, -6, -5, 0, 2, 1, -1, -1, -2, 0, -1, 0, 1, 0, 0, 1, 2, 0, 1, -1, -3, -3, -5, -5, -7, -7, -6, -6, -4, 1, 4, 1, 0, -2, -1, -1, 0, 0, 0, 2, 1, 2, 2, 0, 0, 0, -2, -2, -5, -6, -7, -6, -6, -6, -3, 0, 4, 2, 0, -1, 0, 0, 0, 0, 2, 2, 0, 1, 0, 0, 0, 0, -2, -3, -6, -5, -6, -7, -5, -4, -1, 0, 5, 3, 1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 2, 1, 1, 1, 0, -3, -6, -6, -6, -5, -4, -3, -2, 2, 6, 3, 2, 0, 0, 0, 0, 0, 0, 2, 2, 1, 1, 1, 2, 1, -2, -5, -6, -6, -5, -5, -2, -1, 1, 7, 8, 3, 3, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 1, 0, -1, -4, -6, -5, -3, -1, 1, 3, 5, 11, 10, 7, 3, 1, 0, 0, -2, -2, 0, -1, -3, -4, -4, -3, -1, -3, -3, -5, -4, -3, 0, 2, 3, 6, 10, 16, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, -1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, -1, 1, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 1, -1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 2, 3, 3, 0, 0, 0, 0, -1, 0, 0, 0, -2, 0, 3, 8, 6, 6, 5, 4, 2, 2, 2, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 2, 5, 4, 3, 3, 2, 0, 1, 4, 2, 2, 0, 0, 3, 2, 1, 0, 0, 0, -1, -1, -1, -1, -2, -1, -2, 0, 1, 3, 2, 1, 1, 1, 2, 5, 3, 3, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 1, 1, 1, 2, 3, 6, 1, 3, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 0, 0, 1, 0, 2, 5, 6, 0, 2, 2, 2, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 1, 0, 0, 1, 0, 2, 1, 0, 1, 3, 3, 4, 1, 3, 2, 2, 0, 1, 1, 0, -1, -1, -1, -2, -1, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, 1, 3, 7, 1, 2, 1, 2, 2, 1, -1, -1, -1, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 2, 1, 1, 1, 3, 6, 0, 2, 2, 0, 2, 0, -2, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 3, 4, 4, 0, 1, 2, 5, 0, 1, 0, 0, 1, -1, -2, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 2, 4, 5, 1, 0, 0, 3, -1, 0, 0, -1, -1, -1, -2, 0, -1, -2, 0, 0, -1, 0, -2, -1, -2, -2, 0, 2, 4, 4, 2, 0, 0, 0, -1, 0, 0, 0, -1, -2, -3, -2, -2, -3, -1, -2, 0, -1, -1, -3, -4, -4, -3, 0, 3, 3, 0, 0, -2, 0, -1, 0, 0, -2, -2, -3, -2, -1, -1, -3, -2, -3, -2, -1, -4, -4, -4, -6, -3, 0, 3, 4, 0, 0, -2, -1, -2, 0, -2, -3, -4, -2, -2, -2, -1, -2, -3, -3, -1, -2, -2, -5, -4, -5, -1, 1, 4, 2, 0, -3, -4, 0, -3, -1, 0, -1, -2, -3, -2, 0, -1, -2, -2, -2, -1, -3, -3, -3, -2, -3, -1, 2, 4, 3, 0, -2, -3, 0, -1, -1, 0, 0, -2, -1, -1, 0, 1, 0, 0, 0, -1, -1, -3, -2, -1, -1, 0, 1, 1, 1, -1, -3, -2, 2, -2, 0, 0, -1, -1, -2, -1, 0, 1, 0, 0, 0, 0, -1, -3, -2, -1, 0, 0, 1, 2, 0, -1, -1, 0, 4, 0, 1, 0, 0, -1, -3, 0, 0, 0, 1, 0, 0, 0, -2, -4, -2, -2, 1, 1, 1, 0, 0, 0, 0, 1, 5, 0, 0, 0, -1, 0, -2, -2, -2, 0, 0, 0, 1, 0, -2, -2, -2, -1, 1, 1, 1, 2, 1, 0, -1, 2, 5, -3, 0, 0, 0, -1, -3, -3, -2, -2, 0, 0, 1, 0, -1, -3, -3, -1, 0, 0, 1, 1, 0, -1, -2, 1, 5, -1, -1, 0, 1, 0, -2, -2, -1, -2, 0, 0, 0, 1, -2, -1, -2, -1, 0, 2, 3, 0, 0, 0, 0, 1, 5, -2, 0, -1, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, -2, -1, 1, 2, 3, 3, 1, -1, -2, 0, 7, -1, 0, 0, 3, 4, 2, -1, 0, 0, 0, 0, -1, 0, 0, -2, -2, 0, 0, 2, 5, 3, 1, -1, 0, 2, 7, 0, 0, 1, 2, 4, 3, 0, -1, 0, -1, -1, 0, -1, 0, 0, -3, 0, 0, 5, 6, 6, 3, -2, -1, 2, 7, -1, 0, 0, 4, 4, 2, 1, 0, 0, -3, -3, -4, -1, 0, -1, 0, 0, 1, 4, 5, 6, 2, 0, 0, 2, 6, -2, -1, 2, 4, 4, 1, 2, 1, -1, -3, -2, -4, -2, 0, 1, 1, 0, 2, 4, 6, 5, 2, 2, 1, 2, 5, 1, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -1, -1, -1, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 1, 1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 2, 2, 1, 1, 1, 1, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 2, 2, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, -1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 2, 0, 0, 2, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 1, 0, 2, 1, 1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 2, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, -1, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, 1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -1, -2, -2, -1, -1, -3, -3, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -2, 0, 0, -1, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, -2, -1, -2, -2, -2, -1, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, 1, 0, 1, 3, 1, 2, 2, 2, 1, 0, -2, -2, -1, -3, -1, -2, -1, 0, 1, 1, 2, 0, 1, 1, 1, 1, 0, 0, 1, 2, 1, 4, 3, 2, 0, 0, -1, -2, -1, -2, -1, -3, 0, -1, 0, 2, 1, 3, 2, 2, 1, 1, 0, 0, 1, 1, 3, 4, 4, 4, 1, 0, -2, -2, -2, -2, -2, -3, -2, 0, 0, 2, 2, 1, 1, 2, 0, 1, 0, 2, 3, 2, 3, 3, 5, 5, 4, 0, 0, 0, 0, 0, -3, -3, -1, 0, 0, 0, 1, 0, 1, 1, 2, 1, 0, 2, 3, 3, 4, 4, 6, 4, 4, 2, 0, 0, 0, -2, -1, -3, -1, -2, -1, 0, 1, 2, 1, 2, 0, 0, 0, 1, 2, 4, 6, 5, 5, 4, 4, 2, 0, 0, 1, 0, 0, 0, -2, -2, -2, 0, 1, 0, 0, 1, 0, 0, 2, 3, 4, 4, 3, 6, 5, 4, 3, 2, 1, 0, 0, 1, 1, 0, -2, -2, -2, 0, 1, -1, 0, 0, -1, 0, 2, 1, 3, 4, 4, 4, 6, 3, 3, 2, 1, 0, 1, 1, 1, 0, -2, -4, -2, 0, 0, 0, 0, -1, 0, 0, 2, 2, 3, 3, 5, 4, 4, 5, 5, 1, 1, 0, 0, 0, 0, -1, -4, -3, -3, 0, 0, 0, 0, -1, -2, 0, 1, 2, 3, 3, 4, 3, 4, 5, 3, 2, 1, 0, 0, 0, 0, -1, -2, -4, -3, -1, 0, 0, 0, -1, 0, 0, 2, 2, 4, 3, 4, 4, 5, 5, 5, 2, 0, 0, 0, 1, 0, -2, -2, -3, -2, -1, -1, 1, 0, 0, 0, 0, 3, 4, 3, 3, 6, 6, 4, 4, 4, 3, 2, 0, 0, 0, 0, -1, -3, -4, -1, -2, -1, 0, 1, 0, 1, 2, 3, 3, 3, 3, 6, 4, 4, 4, 3, 2, 1, 0, 0, -1, -1, -2, -3, -3, -2, 0, 0, -1, 0, 0, 0, 0, 3, 3, 4, 4, 5, 5, 5, 3, 1, 1, 1, 0, 0, -1, -2, -2, -1, -2, -1, -1, -1, 0, 0, 1, 0, 0, 3, 4, 5, 4, 5, 4, 2, 1, 1, 1, 0, 0, 0, 0, 0, -2, -3, -3, -1, 0, -2, 0, 0, 0, 0, 0, 2, 3, 3, 5, 4, 5, 4, 1, 1, 0, 0, 0, -1, 0, -2, -4, -2, -3, -2, 0, -1, -1, 0, 0, 1, 0, 0, 3, 2, 3, 5, 5, 4, 1, 2, 0, 0, -1, -2, 0, -2, -4, -4, -2, -1, 0, -1, 0, 0, 0, 1, 0, 1, 1, 2, 3, 5, 5, 3, 0, 2, 0, -1, -1, 0, 0, -2, -2, -5, -3, 0, -1, -1, 0, 0, 0, 0, 1, 0, 2, 2, 4, 5, 4, 4, 2, 0, 0, 0, -1, 0, 0, -1, -3, -5, -3, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 3, 3, 5, 2, 2, 0, 0, 0, -1, -1, -1, -3, -3, -4, -4, 0, -1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 3, 2, 2, 1, 0, 0, -1, -1, -1, -1, -2, -3, -3, -2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, -1, -2, -3, -1, -1, -2, -3, -4, -4, -2, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -2, -2, -1, -1, 0, -2, -1, -3, -2, -3, -1, -2, -2, -3, -1, -2, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 1, 0, 1, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, -1, 0, 1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 8, 3, 1, -1, -2, -2, -3, -2, -1, 0, 0, -1, -2, -3, -3, -2, -4, -5, -4, -3, -1, 0, 4, 5, 9, 14, 6, 2, 0, 0, -2, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, -4, -4, -4, -1, -1, 0, 2, 4, 9, 5, 1, 0, -1, -1, 0, -3, -1, -2, -1, -1, 0, -1, 0, 0, 0, -2, -3, -3, -5, -3, -4, -4, -2, 1, 6, 2, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, 0, -1, -2, 0, 0, -1, -3, -4, -5, -3, -5, -5, -3, -3, 3, 0, 0, 0, 0, 0, 1, 0, 0, -2, 0, -1, -1, 0, 0, -1, 0, 0, 0, -3, -4, -4, -6, -6, -5, -3, 2, -1, -2, -1, 0, 0, 1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 1, 1, 0, -3, -3, -3, -3, -7, -6, -4, 2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 2, 1, -1, -4, -3, -3, -5, -4, -4, -2, 2, -1, -2, -3, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 2, 0, -1, -3, -3, -3, -3, -4, -5, -3, 2, -2, -2, -2, -2, -3, 0, 2, 2, 1, 0, 0, 0, -2, 0, 0, 2, 1, -2, -4, -4, -4, -3, -3, -4, -2, 1, -1, -3, -3, -5, -2, 1, 2, 3, 0, 0, -1, -2, -1, 0, 0, 0, 0, -1, -3, -3, -3, -3, -4, -2, -2, 2, -1, -1, -3, -1, 0, 3, 4, 3, 0, 0, -1, -3, 0, 0, 3, 3, 3, -1, -3, -4, -3, -2, -2, 0, 0, 3, 0, -1, 0, -1, 1, 4, 6, 5, 2, 0, -1, -1, -1, 1, 4, 4, 4, 0, -1, -4, -4, -2, 0, 0, 2, 3, 0, 0, 0, 0, 2, 4, 4, 4, 1, 1, 0, -1, 0, 1, 5, 5, 2, 0, -1, -3, -3, -3, -1, 0, 1, 6, 0, 0, 0, -1, 0, 2, 3, 2, 0, 0, 0, 0, 2, 4, 3, 3, 0, 0, 0, -1, -1, -1, -1, 0, 2, 6, -3, -4, -2, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -2, -1, -2, -1, 0, 0, 1, 4, -3, -4, -3, -2, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, -2, -2, -2, -1, -2, -2, -1, 1, 3, -3, -4, -5, -3, -2, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -2, -2, -2, -3, -3, -2, -3, 0, 3, 0, -2, -3, -2, 0, 0, -1, 1, 0, 0, 0, 0, 0, 2, 1, 0, -1, 0, -2, -3, -2, -2, -2, -3, -1, 2, 0, -4, -3, 0, 0, 0, 2, 0, -1, -2, -1, 0, 0, 1, 1, 0, 0, -1, -4, -3, -5, -3, -2, -2, 0, 2, 0, -2, -1, -2, 0, 0, 1, 2, -1, -1, -1, -1, 1, 2, 1, 2, 1, 0, -2, -3, -5, -4, -3, -3, -1, 1, 2, -1, -2, -1, 0, 1, 2, 1, 1, 0, 0, -1, 1, 1, 1, 1, 0, 0, -1, -4, -5, -4, -5, -4, -2, 0, 2, -1, -1, -1, 0, 0, 2, 1, 2, 0, 0, 0, 1, 2, 2, 0, 0, -1, -4, -5, -6, -4, -4, -3, -2, 2, 3, 1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 1, 2, 3, 3, 0, -3, -3, -5, -5, -3, -3, -3, -1, 2, 5, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 2, 4, 3, 0, 0, -4, -4, -3, -2, 0, 0, 2, 4, 7, 3, 2, 0, 0, 2, 1, 1, 1, 0, 0, -1, 0, 1, 1, 1, 0, -1, -2, -4, -2, 0, 1, 5, 5, 9, 9, 3, 1, 0, 0, 0, 0, -1, -2, -1, -3, -2, -4, -2, -1, 0, -1, -1, -3, -4, 0, 2, 5, 9, 10, 15, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 3, 3, 3, 2, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 2, 2, 1, 1, 0, 0, -1, -1, -2, -2, -2, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 1, 0, 1, 0, -1, -1, -2, -2, -2, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, -1, -1, -1, 0, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 1, 0, 0, 1, -1, -1, 0, -2, -1, 0, 0, -2, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 2, 2, 0, 0, 0, 1, 1, 0, 0, -2, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 3, 2, 2, 0, 1, 0, 0, 0, -1, -1, 0, 0, -2, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 2, 3, 2, 3, 2, 1, 1, 0, 0, 0, 0, -1, -2, 0, -2, 0, 1, 1, 1, 0, 1, 0, 0, 2, 2, 2, 1, 4, 3, 3, 2, 2, 1, 0, 0, -1, -2, -1, -1, -2, -2, 0, 1, 0, 2, 1, 2, 0, 2, 2, 0, 1, 3, 3, 3, 3, 3, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 1, 1, 1, 2, 2, 0, 2, 2, 2, 3, 4, 3, 3, 2, 3, 2, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 1, 1, 2, 0, 1, 1, 2, 1, 2, 3, 4, 5, 4, 3, 2, 2, 1, 0, -1, -1, -2, -1, 0, -1, 0, 0, 0, 0, 2, 1, 1, 2, 1, 1, 2, 2, 3, 4, 4, 3, 1, 3, 0, -1, 0, -1, 0, 0, 0, -2, 0, 2, 2, 0, 2, 3, 1, 0, 0, 0, 1, 2, 2, 2, 3, 3, 3, 1, 0, 0, -1, -2, -1, 0, 0, 0, 0, 1, 2, 3, 2, 2, 0, 0, 0, 1, 1, 3, 3, 3, 3, 4, 1, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 1, 1, 0, 0, 1, 3, 3, 1, 1, 2, 2, 0, 0, 0, -3, 0, 0, -1, 0, -1, 0, 0, 2, 0, 0, 1, 1, 1, 0, 1, 0, 2, 2, 1, 2, 3, 0, 0, -1, -2, -1, -2, -2, -1, 0, 0, -1, 0, 2, 0, 0, 1, 0, 0, -1, -1, 0, 0, 1, 1, 1, 1, 1, 1, 0, -1, -2, -2, -2, -1, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, -2, -3, -2, -1, -2, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, -3, -3, -1, 0, -1, -2, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 1, 1, 2, 0, 0, 0, 0, -1, -2, -2, -1, -1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 1, 2, 0, 1, 1, 1, 0, 0, 0, -2, -2, -1, -2, -2, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 2, 2, 2, 2, 2, 0, 0, 0, 0, -1, -2, -2, -2, 0, -2, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 1, 0, 1, 3, 2, 1, 0, 0, 0, 0, -2, -2, -2, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 2, 3, 3, 2, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 2, 3, 1, 1, 0, 1, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, -1, -1, -2, -1, -2, -3, -3, -3, -2, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 1, 0, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -2, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 1, 0, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 2, 1, 3, 3, 3, 2, 0, 1, -1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 2, 2, 0, 2, 2, 0, 2, 3, 3, 0, -1, -2, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 2, 3, 3, 2, 1, 2, 0, 1, 1, 2, 0, -2, -1, -2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 1, 1, 1, 1, 1, 0, 0, -1, -2, -2, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 2, 2, 3, 1, 2, 2, 1, 1, 2, 0, 2, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 2, 1, 2, 1, 1, 3, 1, 2, 2, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 2, 2, 1, 0, 2, 1, 1, 1, 2, 4, 4, 3, 3, 2, 1, 1, 0, -1, 0, 0, 0, 3, 1, 1, 2, 2, 2, 2, 0, 1, 1, 1, 2, 1, 3, 3, 3, 2, 1, 1, 0, 0, 0, -1, 0, 0, -1, 1, 2, 1, 2, 0, 1, 0, 0, 0, 0, 1, 2, 3, 3, 3, 3, 2, 0, 0, 0, -3, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 1, 2, 2, 2, 3, 1, 2, 0, 0, 0, -2, -1, -2, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 2, 2, 1, 0, -1, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 2, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, -1, -1, 0, 0, -1, 1, 1, 1, 2, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 2, 0, 1, 0, 1, 0, 0, -1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, -2, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 3, 0, 0, 1, 3, 3, 3, 2, 3, 3, 3, 4, 3, 1, 2, 2, 0, 0, 0, 0, -3, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 2, 2, 1, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 2, 2, 1, 2, 0, 0, 1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 2, 2, 1, 1, 0, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, -1, 1, 2, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 2, 1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 1, 2, 1, 0, 0, 0, 1, 1, 3, 2, 1, 1, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 1, 3, 1, 2, 2, 2, 1, 2, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 2, 2, 1, 0, 1, 1, 2, 2, 2, 3, 3, 2, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 2, 2, 0, 0, 1, 0, 2, 1, 3, 3, 3, 2, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 2, 1, 1, 0, 1, 1, 2, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 2, 0, 1, 1, 2, 1, 2, 2, 2, 3, 2, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 0, 0, 0, 2, 2, 1, 2, 1, 3, 2, 2, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 2, 2, 1, 1, 2, 1, 0, 0, 2, 1, 0, 1, 2, 2, 2, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 1, 2, 1, 1, 1, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 2, 0, 1, 0, 1, 2, 0, 1, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 2, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 2, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 2, 0, 2, 1, 0, 0, 0, 1, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 1, 2, 1, 0, 1, 0, 0, 0, -1, -1, -1, -1, -2, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 2, 0, 0, -1, 0, -1, -1, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 1, 0, 1, 0, 1, 1, 0, 2, 1, -1, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 1, 0, -1, 0, 0, -1, 0, 0, -2, -1, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, -1, -1, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 2, 0, -1, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, -1, -1, 0, 1, 0, 2, 1, 0, 0, -1, 0, -2, -2, -1, -1, 0, -1, 0, 0, 1, 2, 1, 0, 0, 0, -1, -2, 0, -1, 0, 1, 1, 2, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 2, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, 2, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 2, 0, 1, 1, 1, 1, 1, 0, -1, -2, -1, 0, -2, -1, 0, 2, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, -1, 0, -2, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 1, 1, 1, 1, 1, 3, 3, 4, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 1, 3, 1, 3, 3, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 2, 1, 2, 3, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 2, 0, 1, 0, 0, -1, -2, -1, -1, -2, -1, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -3, -1, 0, 1, 0, 2, 1, 0, -1, 0, 0, 2, -2, -2, -2, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -2, -1, -2, -1, 1, 1, 0, -1, 0, -1, -1, -1, -1, -2, -1, -3, -1, 0, -2, 0, 1, 0, 0, 0, -1, 2, -3, -3, -2, -2, 0, 0, 0, -1, -2, -1, -2, -1, -1, 0, -2, -2, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, -3, -2, -3, -3, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 2, -4, -4, -1, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, -2, -1, -1, 1, 1, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, -1, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 2, -1, 0, -1, 0, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 3, 3, 4, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 3, 3, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, 2, 2, 0, 0, -1, 0, 1, 2, 1, 0, 0, 0, 2, 1, 1, 4, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 2, 0, -1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 2, 3, 0, 0, 0, 0, 1, 1, -1, -1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 1, 2, 1, 1, 1, 0, 1, 2, 3, -1, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 1, 0, 2, 1, 1, 2, 1, 1, 0, 3, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, -2, 0, 0, -1, -1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 1, 2, 0, 0, 0, 0, 2, 1, 0, 0, 0, -1, -2, -1, -2, -1, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 2, 2, 2, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 8, 6, 1, 0, 0, -1, 0, -1, -2, -1, 0, -1, -2, -4, -3, -4, -4, -4, -6, -5, -6, -4, -1, -1, 1, 4, 6, 3, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -3, -3, -3, -5, -6, -5, -3, -2, -1, 0, 1, 6, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, -1, -3, -4, -4, -4, -5, -5, -3, -2, -2, 2, 4, 1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -2, -4, -5, -5, -3, -4, -3, -1, 0, 4, 1, 0, 1, 0, 1, 1, 1, 1, 0, 0, 1, 1, 2, 0, -1, 0, -1, -3, -3, -3, -5, -5, -4, -3, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, -3, -4, -3, -4, -4, -4, -5, -3, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -2, -3, -4, -4, -4, -3, -4, -2, -1, 2, 0, -1, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, -2, -4, -3, -4, -4, -2, -3, -3, 0, 1, 0, -2, -2, -1, 0, 1, 1, 0, 0, 0, 1, 2, 2, 1, 1, 1, 0, -3, -4, -2, -2, -2, -1, -3, 0, 1, 0, 0, -2, 0, 0, 1, 1, 0, 0, 0, 0, 1, 2, 2, 3, 1, 1, -1, -1, -2, -1, -1, -1, 0, 1, 3, 0, 0, -1, 0, 0, 1, 2, 2, 0, 1, 1, 1, 3, 3, 4, 3, 0, 0, -1, -3, -2, -3, -1, -1, 0, 4, 1, 1, 0, -1, 0, 1, 0, 2, 0, 0, 0, 1, 3, 5, 5, 5, 1, -1, -1, -3, -2, -1, -1, -1, 1, 3, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 2, 2, 4, 3, 4, 2, 0, -1, -1, -2, -3, -2, 0, 0, 0, 2, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 1, 2, 3, 3, 3, 1, 0, -1, -2, -1, -1, -1, -1, 0, 1, 1, -1, -1, -2, -1, 0, -1, 0, 0, 1, 0, 0, 1, 3, 2, 1, 1, 0, 0, -3, -1, -2, -1, 0, -1, 0, 0, -3, -3, -2, 0, -2, 0, 0, 2, 0, 0, 0, 2, 2, 1, 0, 0, 0, -2, -2, -3, -2, -2, -1, -2, 0, 1, -1, -2, 0, -1, 0, 0, 1, 2, 0, 1, 1, 0, 0, 1, 1, 0, -2, -3, -1, -3, -2, -4, -3, -2, 0, 2, -1, -2, -1, 0, 0, 1, 2, 2, 0, 1, 1, 1, 2, 0, 0, 0, 0, -2, -4, -3, -4, -4, -3, -2, 0, 2, 0, -1, -2, 0, 0, 0, 2, 1, 1, 0, 2, 0, 0, 0, 0, 0, -2, -2, -2, -4, -4, -3, -3, -4, 0, 4, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 2, 2, 1, 2, 0, 0, -1, -1, -2, -4, -3, -4, -3, -4, 0, 4, 1, -1, 0, 0, 1, 0, 2, 1, 1, 0, 1, 2, 2, 2, 0, 0, -2, -1, -4, -3, -4, -3, -3, -3, 0, 6, 1, 1, 1, 1, 0, 1, 2, 2, 1, 2, 2, 3, 1, 1, 0, 0, -1, -4, -2, -2, -3, -2, -3, -2, 0, 6, 3, 2, 1, 1, 0, 0, 2, 0, 1, 2, 1, 2, 2, 2, 0, -2, -4, -4, -5, -3, -2, -3, -3, -1, 1, 6, 3, 2, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 1, 0, 0, -3, -4, -5, -4, -3, -4, -3, -3, 0, 1, 9, 4, 3, 1, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, -3, -5, -5, -6, -5, -3, -2, -1, -1, 1, 4, 10, 6, 3, 3, 0, 0, 0, -1, 0, -2, -2, -3, -3, -3, -4, -5, -7, -8, -8, -6, -4, -3, -2, 0, 3, 4, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, -1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, 1, 0, 0, 0, -1, 0, -1, -2, -2, 0, -1, 0, -2, -1, -1, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, 0, 1, 0, -1, -1, -2, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, -2, -1, -2, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, -1, 0, -1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 1, 0, -1, -1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 1, 0, 0, 0, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 1, 2, 2, 1, 0, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 1, 1, 2, 1, 2, 1, 2, 2, 2, 1, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 2, 2, 1, 1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 0, 0, -1, -1, -1, 0, 0, -2, -1, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 2, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 2, 0, 0, 0, 1, 1, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, -1, -2, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, 1, 0, 1, 0, 0, 0, 2, 1, 2, 2, 2, 0, 0, 2, 1, 1, 1, 0, 1, 0, 0, 0, 0, -1, 10, 6, 2, 0, -1, 0, 0, -1, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, -2, -3, -2, 0, 0, 0, 2, 3, 7, 4, 1, 0, 0, -2, -1, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, -4, -4, -3, -2, -1, -2, 0, 1, 7, 3, 1, 1, 0, -1, -2, -1, -2, -2, 0, -1, 0, 0, 0, 0, 0, -1, -2, -3, -4, -4, -2, -2, -1, 0, 4, 2, 1, 0, 0, -1, 0, -1, -2, -3, 0, 0, 0, 0, 0, 0, 0, -2, -2, -3, -3, -3, -3, -3, -3, -1, 5, 1, -1, -1, 0, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, -4, -4, -4, -4, -4, -3, -3, 2, 0, 0, -1, 0, 0, 1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -2, -3, -3, -2, -3, -4, -5, -3, 0, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, -2, -3, -4, -4, -4, -2, 1, 0, -3, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -4, -3, -3, -3, -4, -2, 2, 0, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, -3, -3, -1, -2, -2, -2, 4, 0, -2, -3, -2, 0, 1, 2, 0, 1, 0, 0, 0, 0, 1, 1, 2, 1, 0, -3, -4, -2, -2, -1, -3, -1, 3, 1, -1, -1, -2, 0, 2, 2, 1, 0, 0, 0, 0, 0, 2, 3, 2, 2, 0, -1, -4, -1, -3, -2, -1, 0, 3, 2, 0, -2, 0, 0, 3, 4, 2, 0, 0, -1, 0, 0, 3, 2, 4, 2, 1, -1, -2, -2, -1, -2, 0, 0, 4, 0, -1, 0, 0, 2, 2, 3, 2, 1, 1, 0, 0, 1, 4, 3, 2, 1, 1, -1, -1, -2, -3, -1, -1, 0, 3, 0, -1, -2, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 2, 3, 0, 0, 0, -1, -2, -2, 0, 0, 1, 3, 0, -3, -3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 3, 2, -1, 0, 0, -1, -2, -1, 0, -1, 0, 2, -2, -2, -4, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, -2, 0, 0, 0, -1, -1, 0, 3, 0, -3, -3, -2, -1, -2, -2, 0, 1, 1, 0, 0, 1, 0, 2, 0, 0, -1, -1, -3, -1, -2, -1, 0, -1, 4, -1, -1, -2, -2, 0, 0, 0, -1, 1, 0, 0, 0, 2, 2, 1, 0, 0, 0, -2, -1, -2, -2, -3, -2, 0, 4, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, 0, -2, -1, -2, -3, -3, -2, 0, 6, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, -1, 1, 1, 0, 1, -1, -1, -1, -2, -3, -3, -1, -2, 0, 5, 2, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, -1, -1, -2, -4, -3, -2, -1, -1, 6, 2, 1, 0, 1, 1, -1, 0, 1, 1, 0, 0, 0, 1, 1, 2, 0, -1, 0, -2, -3, -3, -2, -3, -1, -1, 8, 3, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 2, 0, 3, 0, 0, 0, -1, -3, -3, -1, -2, 0, 1, 9, 3, 2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 2, 0, 0, -2, -2, -3, -1, -1, -1, 0, 1, 9, 5, 3, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, 0, 1, 1, 0, 0, -3, -2, -3, -2, 0, 1, 2, 5, 12, 8, 3, 2, 0, 0, 0, 0, 0, 0, -2, -3, -3, -3, -2, 0, 0, -1, -2, -1, -2, -1, 1, 3, 5, 6, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 0, 1, 1, 1, 2, 2, 1, 0, -1, -1, 0, 0, -1, -2, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, 0, 1, 0, 0, 0, 1, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, -1, 0, 1, 1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -2, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 1, 0, -1, -1, 1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, 1, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 2, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, 1, 2, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 2, 1, 1, 0, 0, 0, 1, 0, -1, -1, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 2, 2, 2, 2, 2, 1, 2, 0, 0, 0, 1, -1, -1, -1, 0, -1, 0, 1, 0, 1, 0, 0, -1, -1, 0, 0, 1, 0, 2, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 2, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 2, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 1, 2, 1, 1, 2, 2, 2, 2, 1, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 1, 1, 3, 3, 1, 0, 2, 1, 0, -1, 0, 0, 0, -1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, -1, 3, 0, 0, 0, 1, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 1, 2, 1, 2, 0, 1, 0, 0, -1, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 1, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 2, 0, 0, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 3, 2, 2, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, -1, 0, 0, 3, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -2, -1, 0, 0, 3, 3, 3, 2, 0, 0, -2, 0, 1, 4, 3, 5, 4, 5, 5, 3, 3, 1, 2, 1, 0, 0, -1, 0, -1, 1, 1, 4, 1, 0, -2, -3, -4, 0, 0, 1, 2, 1, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 1, 2, 2, 1, -1, 0, -2, -3, -2, -2, 0, 0, 0, 0, 0, 0, -3, -3, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, -3, -2, 0, 0, 0, 0, 0, 0, -3, -3, -3, -1, -1, -1, 0, -1, 1, 0, -1, -1, 0, 0, 0, -1, -2, -3, -1, -2, 0, 0, 0, 0, -1, -2, -3, -4, -2, -3, -3, -2, -1, -1, 0, 1, 0, -2, -1, -1, -1, -2, -2, -1, -2, 0, 1, 2, 2, 1, 0, -3, -2, -4, -5, -2, -2, -2, -2, -2, 0, 1, 1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 2, 3, 3, 0, 0, -2, -4, -2, -4, -2, -2, -1, -2, -3, 0, 3, 3, 0, 0, -1, -1, -3, -2, 0, 0, 2, 3, 1, 1, 2, 0, 0, -1, -1, -1, 0, -3, -1, -1, -2, 0, 1, 2, 0, -1, -1, 0, -2, -1, 0, 0, 1, 2, 2, 1, 1, 0, 0, 0, -1, 0, -1, -2, -1, -2, -3, 0, 1, 1, 0, 0, -1, -3, -3, -2, 1, 0, 1, 1, 1, 1, 0, 0, -1, -1, 0, 0, -1, -2, -2, -3, -4, 0, 1, 1, 0, -2, -3, -3, -3, -3, -1, 1, 2, 0, 0, 1, -1, 0, -3, -1, -1, 0, 0, -2, -3, -2, -5, 0, 0, 1, 0, -2, -3, -3, -4, -1, 0, 1, 0, 0, 0, 0, 0, -1, -3, -3, -3, -1, 0, -1, -3, -3, -5, 0, 0, 0, 0, -3, -5, -5, -3, -2, 0, 0, 0, 1, 0, 0, 0, -1, -3, -2, -2, 0, 0, -2, -2, -3, -4, 0, 2, 0, -1, -1, -4, -4, -2, -1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -2, -2, -3, -1, -1, -3, -4, -3, 0, 0, 1, 0, -1, -3, -4, -2, 0, 0, 2, 1, 1, 1, 1, 2, 0, 0, -2, -3, -2, -3, -2, -3, -3, -3, 2, 3, 2, 1, -1, -1, -2, -2, 0, 0, 1, 2, 1, 3, 1, 2, 1, 0, -2, -3, -3, -2, -2, -4, -4, -2, 1, 3, 2, 0, 0, -3, -4, -1, 0, 0, 1, 2, 3, 3, 1, 0, -1, 0, -1, -2, -3, -1, -3, -4, -3, -4, 2, 3, 0, 1, -2, -2, -3, -2, -1, 0, 2, 2, 2, 2, 2, 0, 0, 0, -3, -2, -3, -2, -2, -3, -3, -3, 0, 2, 1, -1, -1, -2, -2, -3, -2, 0, 1, 2, 1, 3, 1, 0, -2, -2, -2, -2, -4, -4, -3, -2, -3, -3, 0, 0, 0, 0, -2, -2, -4, -2, 0, 0, 2, 1, 3, 0, 0, -1, 0, 0, 0, -4, -5, -3, -5, -4, -5, -3, 0, 0, 1, 0, 0, -3, -2, -2, 0, 1, 2, 3, 2, 2, 1, 0, 0, 0, 0, -2, -4, -2, -5, -3, -4, -3, 0, 1, 2, 0, 1, -2, -2, -1, 0, 2, 1, 3, 4, 1, 0, 0, 0, 1, 0, -1, -3, -3, -3, -2, -3, -2, 1, 2, 2, 3, 1, 0, 0, -1, -1, 2, 3, 2, 3, 3, 3, 0, 2, 0, 0, 0, -2, -2, -2, -2, -1, -2, 1, 2, 3, 4, 1, 1, 0, -1, 0, 0, 2, 1, 2, 3, 2, 2, 1, 3, 0, 0, -2, -2, -1, -1, -2, -2, 0, 3, 4, 4, 3, 1, 0, -1, -1, 0, 1, 1, 2, 4, 3, 3, 2, 2, 1, 0, 0, 0, 0, -1, -2, -3, 1, 1, 5, 5, 4, 3, 1, 1, 0, 0, 0, 0, 4, 5, 6, 4, 4, 3, 4, 3, 0, 1, 0, 0, -1, -2, 0, -1, -1, 0, -1, -2, -1, -1, 0, 0, 0, 1, 2, 5, 4, 2, 1, 0, -1, 0, -1, 0, 1, 1, 0, 1, -1, 0, -1, -1, 0, -1, -1, -2, 0, 0, 0, 1, 1, 1, 1, 1, 0, -1, -3, -3, -3, -3, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -2, -2, -2, -2, 0, 0, 0, 1, 0, -1, -2, -3, -4, -4, -2, -3, -1, -2, 0, 0, -1, 0, 0, 1, 0, 0, 0, -3, -2, -1, 0, 0, 0, 0, 1, 0, -2, -3, -4, -4, -4, -4, -3, -2, -1, 0, 0, 0, -1, -1, 0, 0, -2, -2, -2, 0, -1, 0, 0, 0, 0, 0, -2, -2, -3, -3, -3, -5, -3, -3, -2, 0, 0, 0, -1, 0, 0, 0, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -3, -2, -4, -4, -3, -3, -1, 0, -1, 0, -2, 0, 0, 0, -2, -2, -1, -1, 0, 1, 0, 0, 0, 1, 0, -1, -1, -3, -2, -3, -4, -4, -2, 0, 0, 0, -1, -1, -1, 0, 0, -2, 0, -1, 0, 1, 0, 2, 1, 0, 0, 0, -1, -2, -3, -3, -3, -3, -2, 2, 1, 0, -1, -2, -1, 0, -1, -1, -1, 0, 0, 0, 2, 2, 1, 1, 0, -1, -2, -3, -2, -3, -2, -4, -2, 3, 1, 0, 0, -1, -1, 1, 0, -1, 0, 0, 0, 0, 2, 1, 2, 2, 1, 0, -1, -1, -2, -2, -3, -2, -2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 3, 2, 2, 0, 0, 0, -1, -2, -2, -2, -1, -2, 1, 1, 2, 0, 0, 1, 0, -1, -1, 0, 1, 1, 2, 2, 3, 2, 1, 0, -1, -1, -1, -1, -1, -1, -3, -1, 1, 1, 0, 2, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 3, 2, 2, 0, 0, -1, 0, 0, -1, -2, -2, 0, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 3, 0, 0, -1, 0, 0, -1, 0, -1, -2, 0, 2, 1, 0, 2, 0, 0, -2, -1, 0, 0, 0, 0, 2, 3, 3, 0, 1, 0, 0, -2, 0, -1, -1, -2, -3, 0, 2, 2, 1, 1, 0, -1, -1, 0, 0, 0, 0, 2, 1, 2, 1, 1, 1, 0, -2, -2, -1, -2, -1, -2, -2, -3, 2, 1, 2, 0, 0, -1, -1, -2, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, -2, -2, -1, -3, -3, -3, -3, -3, 2, 1, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, -1, -1, -1, -2, -3, -2, -4, -4, -4, -2, 0, 1, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, -3, -3, -2, -4, -4, -5, -4, -2, 1, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -3, -3, -3, -3, -4, -2, -2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, -1, -4, -4, -4, -3, -4, -3, -1, 1, 1, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 2, 0, 0, -1, -2, -1, -2, -3, -2, -4, -4, -1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 2, 1, 2, 2, 2, 0, 0, 0, -3, -1, -3, -3, -3, -2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 2, 2, 1, -1, 0, -1, -1, -1, -1, 0, -1, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 1, 0, 1, 1, 2, 0, 1, 0, -1, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 1, 1, 2, 1, 2, 2, 1, 2, 1, 3, 4, 4, 3, 3, 5, 3, 1, 2, 1, 2, 0, 1, 0, 0, 0, 2, 4, 5, 6, 3, 3, 2, 2, 0, 0, -1, 0, 0, 4, 5, 3, 2, 0, 0, 0, 0, 0, -1, -2, -3, -2, 0, 3, 5, 5, 3, 4, 4, 2, 1, 1, 0, 0, 0, 3, 5, 3, 0, 0, 0, -1, 0, -1, -1, -4, -2, -2, 0, 1, 2, 2, 2, 4, 3, 3, 1, 2, 2, 1, 1, 4, 3, 2, 0, 0, 1, 0, 1, 0, 0, -3, -2, -2, -1, 1, 1, 3, 3, 3, 1, 2, 2, 3, 2, 2, 0, 3, 2, 1, 1, 1, 2, 1, 1, 0, -1, -3, -3, -2, -1, 0, 0, 2, 3, 3, 1, 0, 2, 4, 3, 3, 1, 4, 0, 0, 0, 0, 2, 3, 0, -1, -2, -2, -2, -3, -2, -1, 0, 2, 1, 1, 1, 1, 3, 5, 3, 3, 1, 5, 0, -2, -2, 1, 1, 0, 0, 0, -2, -2, -3, -3, -3, -1, -1, 1, 2, 3, 2, 2, 4, 5, 5, 3, 4, 4, 0, -2, 0, 1, 0, 1, 0, 0, -1, -4, -2, -1, -1, -1, -1, 0, 2, 4, 3, 1, 2, 4, 4, 2, 2, 3, 0, 0, 0, 1, 0, 0, 0, -1, -2, -3, -5, -4, -3, -2, 0, 0, 2, 4, 3, 1, 1, 3, 4, 2, 2, 5, 3, 2, 0, 0, 0, 0, 0, 0, 0, -4, -4, -6, -4, -3, -1, 0, 3, 3, 2, 0, 1, 1, 3, 2, 1, 5, 2, 4, 1, 0, 0, 0, -1, 0, -1, -2, -3, -5, -4, -5, -1, 0, 1, 4, 4, 1, 0, 0, 3, 2, 2, 6, 5, 2, 1, 0, -1, 0, 1, 0, 0, -2, -3, -5, -5, -3, -4, -1, 0, 4, 3, 1, 1, 0, 2, 3, 1, 6, 2, 2, 1, -1, -1, 0, 0, 0, -2, -4, -3, -5, -5, -4, -3, 0, 0, 1, 2, 2, 0, 2, 2, 3, 0, 6, 1, 1, 1, 0, -1, -2, 0, -1, -3, -5, -4, -6, -5, -3, 0, 0, 0, 2, 1, 1, 2, 2, 3, 2, 0, 4, 2, 0, 0, 0, 0, -2, -1, -2, -2, -5, -6, -5, -4, -2, 0, 1, 1, 0, 0, 1, 1, 3, 3, 1, 0, 5, 2, 1, 0, 0, -1, -2, -3, -2, -3, -4, -3, -5, -4, -2, 2, 1, 0, 1, 0, 1, 2, 3, 2, 1, 1, 4, 0, 0, -1, -1, 0, 0, -1, -1, -2, -2, -2, -4, -3, 0, 1, 1, 0, 0, 1, 1, 2, 4, 4, 1, 1, 4, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -4, -3, -3, 0, 2, 0, 1, 0, 1, 3, 3, 5, 5, 4, 1, 6, 1, 0, 0, 0, 0, 1, 0, -1, 0, -3, -3, -5, -2, 0, 1, 0, 1, 2, 3, 4, 4, 5, 3, 5, 1, 6, 3, 0, 0, -1, 0, 0, 0, 0, 0, -2, -3, -4, -1, 0, 2, 2, 0, 3, 3, 5, 4, 5, 4, 4, 3, 7, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -3, -4, 0, 2, 2, 0, 0, 2, 5, 6, 6, 4, 5, 5, 3, 4, 3, 0, 0, 1, 1, 1, 0, -1, -2, -2, -1, -1, 0, 1, 1, 1, 1, 1, 3, 4, 4, 3, 4, 3, 2, 6, 4, 1, -1, 0, 2, 2, 0, 0, -2, -2, -1, -1, -1, 0, 1, 0, 1, 2, 3, 4, 3, 3, 4, 4, 2, 7, 5, 1, 0, 0, 1, 1, 0, 0, -1, -1, 0, -2, -1, 0, 0, 0, 0, 3, 3, 3, 3, 2, 3, 3, 2, 7, 5, 3, 0, 0, 1, 2, 0, 1, 0, 0, 0, -1, -1, 0, 0, 1, 2, 1, 0, 2, 2, 4, 2, 3, 0, 8, 7, 4, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 2, 2, 2, 1, 0, -1, 2, 3, 3, 0, 1, 0, 0, 0, 0, 0, 0, -1, -3, -1, -1, -1, -2, -3, -1, 0, 0, -3, -3, 0, 0, 0, 2, 2, 2, 1, 0, -1, 1, 1, 1, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 1, 1, 0, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 1, 1, 2, 2, 0, 0, 0, 1, 0, 1, 1, 1, 1, 2, -1, 0, 0, 0, 0, 2, 0, 0, -1, 0, 0, 1, 0, 2, 1, 1, 1, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 2, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 2, 2, 1, 1, 2, 0, 0, 0, 0, 0, -3, -1, 0, 0, 1, 1, 1, 0, 1, 0, 1, 1, 0, 2, 1, 1, 0, 2, 0, 1, 0, 0, -1, 1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, -1, -2, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 2, 1, 3, 3, 2, 3, 0, 1, 0, 1, 1, 1, 2, 1, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, 1, 1, 1, 1, 1, 1, 3, 2, 2, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 2, 1, 1, 0, 0, 0, 0, -2, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 2, 2, 2, 1, -1, -1, -1, 0, 0, 2, 0, 2, 2, 0, 1, 0, 0, 1, 1, 1, 0, 0, 1, 1, 1, 2, 1, 1, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 2, 2, 0, 0, 0, 1, 0, 0, 1, 0, 2, 1, 1, 0, 0, 2, 0, 1, 0, 0, 0, 1, 1, 2, 1, 1, 1, 0, -1, 0, 0, 0, 0, 1, 0, 2, 0, 0, 1, 2, 2, 2, 1, 0, 0, 0, 2, 2, 2, 0, 2, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 2, 3, 2, 0, 1, 0, 0, 2, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 0, 0, 0, 2, 1, 0, 0, 2, 0, 1, 1, 1, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 1, 1, 0, 2, 0, 0, 1, 2, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -2, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 1, 0, 0, 2, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, -1, 1, 0, 0, 0, 1, 2, 1, 1, 3, 2, 2, 3, 1, 2, 1, 2, 2, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 3, 3, 4, 5, 4, 4, 1, 0, 0, 0, 0, -2, -3, -2, -3, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 3, 1, 2, 1, 1, 0, 0, 0, -2, -1, -1, -1, -3, -3, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 2, 1, 1, 0, 0, 0, -2, -3, -2, -1, -2, -1, -1, -1, 0, 0, 0, 0, -1, 1, 0, 0, -1, -1, 0, 0, 1, 2, 0, 0, 1, 0, -1, -1, -3, -1, -2, -2, -1, -3, 0, 0, -1, 0, -1, 0, -1, -1, 0, -1, -1, 1, 1, 2, 2, 1, 0, 0, -1, -1, -2, -2, -3, -2, -2, -2, -1, 0, 0, -1, 0, 0, 0, -1, -2, 0, -1, 1, 2, 1, 0, 0, 1, 0, 1, 0, -2, 0, -2, -1, -2, -1, -1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 2, 1, 2, 1, 1, 0, 0, 1, 0, -1, -1, -1, -1, -2, -3, 0, 0, 1, 1, 0, -1, 1, -1, 0, 0, 0, 1, 2, 1, 2, 3, 1, 0, 1, 0, -1, 0, -1, -2, -2, -1, 0, 2, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 2, 1, 1, 1, 2, 0, 0, 0, -1, -2, -1, -2, -2, -1, 0, 1, 3, 2, 1, 0, 1, 0, 0, 1, 3, 3, 3, 2, 2, 1, 1, 0, 0, -1, -2, -3, -3, -2, -1, -1, 2, 1, 3, 2, 0, 1, 1, 0, 1, 0, 2, 3, 3, 3, 3, 3, 2, 0, 0, -1, -1, -1, -1, -3, -1, -1, 2, 3, 1, 2, 1, 1, 0, 1, 0, 2, 2, 2, 3, 2, 4, 3, 2, 1, -1, 0, -2, -2, -2, -1, -1, -2, 0, 2, 1, 3, 2, 3, 0, 0, 0, 1, 1, 1, 2, 3, 2, 3, 1, 0, 0, 0, 0, -2, 0, 0, -1, -3, 2, 2, 2, 1, 2, 1, 0, 0, 0, 1, 1, 2, 3, 1, 3, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 3, 2, 2, 1, 1, 0, 0, 0, 1, 1, 2, 3, 3, 3, 2, 2, 1, -1, -2, -2, 0, -1, 0, -1, -3, 1, 1, 2, 1, 2, 2, 0, 0, 0, 0, 3, 2, 3, 4, 2, 3, 1, 1, -1, -1, -2, 0, 0, 0, -1, -3, 3, 1, 2, 2, 3, 0, 1, 0, -1, 1, 2, 1, 1, 3, 2, 1, 2, 0, -1, -2, -2, -3, -2, -1, -2, -1, 2, 2, 1, 2, 1, 2, 0, -1, 0, 0, 0, 1, 0, 2, 2, 1, 0, 0, 0, -1, -3, -3, -1, -1, -1, -2, 0, 0, 1, 2, 1, 1, 0, -1, 0, -2, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, -3, -2, -4, -3, -3, -1, 0, 1, 1, 2, 0, 2, 1, -1, -2, -1, 0, 0, -1, 1, 1, 0, 1, 0, 0, -2, -3, -4, -3, -3, -3, -3, 0, 1, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 2, 0, 0, -1, -2, -4, -2, -2, -3, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 2, 2, 2, 0, 2, 1, 0, 0, 0, -2, -2, -2, -3, 0, -2, 0, 0, 0, 1, 1, 2, 1, 1, 1, 2, 2, 2, 3, 1, 2, 1, 1, 1, -1, -2, 0, -2, -1, -1, -1, -2, 0, 0, 1, 0, 1, 1, 1, 0, 0, 1, 1, 1, 3, 1, 0, 0, 0, 0, 1, 0, 0, 0, -2, -1, -2, -1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 2, 1, 3, 2, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 1, 3, 3, 4, 3, 2, 2, 2, 1, 0, 0, 0, 0, 0, -3, -2, 13, 6, 3, 1, 0, 0, 0, 0, -1, -2, -3, -3, -5, -3, -5, -4, -6, -6, -6, -6, -2, 0, 1, 5, 7, 15, 11, 6, 2, 1, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, -2, -5, -6, -6, -3, -3, -3, 0, 0, 4, 9, 8, 5, 3, 2, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -2, -4, -5, -5, -3, -3, -3, -1, 2, 8, 6, 4, 0, 0, 2, 1, -1, -2, -3, 0, 0, 0, -1, 0, 0, 0, -1, -2, -4, -2, -4, -5, -3, -3, 0, 7, 3, 1, 0, 0, 2, 1, -1, -2, -1, -1, 0, 0, -2, -1, 0, 0, 0, -2, -3, -3, -5, -5, -5, -4, -1, 5, 0, 1, 0, 0, 2, 1, -1, -2, -3, -1, -1, -2, -3, 0, 0, 1, 1, -1, -2, -3, -4, -4, -5, -3, 0, 4, -1, -1, 0, 0, 0, 1, 0, -1, -2, 0, -1, -2, -2, -2, 0, 0, 0, 0, -4, -2, -3, -4, -5, -3, 0, 5, 0, -2, 0, 0, -1, 0, 0, -3, -1, -2, -3, -2, -2, -1, 0, 0, 0, -2, -4, -3, -3, -2, -3, -3, 0, 5, -1, -1, -3, -2, -1, -1, -1, -3, -1, -1, -3, -4, -2, -2, 1, 2, 0, -2, -2, -3, -3, -2, -4, -1, 1, 6, 0, -2, -2, -1, -1, 0, -1, -1, -2, -1, -3, -4, -2, 0, 2, 2, 1, -1, -2, -3, -2, -1, -1, -2, 0, 8, 1, 0, -1, -1, 1, 2, 0, -2, -2, -4, -3, -3, -1, 0, 3, 3, 2, 0, -2, -3, -3, -1, -1, 0, 1, 9, 2, 0, 0, 1, 2, 2, 1, 0, 0, -3, -4, -4, -1, 1, 4, 5, 3, 0, -1, -3, -1, 0, 0, 1, 4, 7, 2, 1, 2, 2, 2, 2, 2, 0, -1, -2, -2, -3, -1, 0, 3, 3, 2, 0, -1, -2, -3, 0, 0, 2, 3, 9, 1, 0, 0, 1, 3, 2, 0, -2, -2, -2, -2, -1, 0, 0, 2, 2, 2, -1, -1, -3, -2, 0, 1, 3, 4, 9, 0, -3, -1, 0, 1, 0, 0, 0, -3, -2, -1, 0, -1, 1, 0, 0, 0, -2, -1, -2, -1, 0, 0, 2, 1, 8, -2, -4, -2, 0, 0, 0, -2, 0, -2, 0, -3, -1, 0, 1, 0, 0, 0, -1, -1, -2, -2, 0, 1, 1, 1, 6, -3, -4, -2, 0, 0, -1, -2, -1, 0, -2, -1, -1, 0, 1, 0, 0, 0, -1, 0, -2, -3, -2, -1, 0, 0, 5, -3, -3, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 1, 0, -1, -3, -3, -2, -2, -2, 0, 1, 7, 0, -2, 0, 0, 1, 1, 0, 0, -2, -1, -2, 0, 0, 2, 0, 1, 0, -1, -3, -3, -3, -2, 0, -1, 0, 5, 0, -1, 0, 0, 2, 1, 1, 0, -2, -1, -1, 0, 2, 2, 2, 0, 1, -1, -1, -3, -4, -2, -2, -1, 0, 6, 2, 1, 0, 0, 3, 1, 1, 0, 0, -2, 0, 1, 3, 1, 1, 2, 0, -1, -2, -4, -5, -1, -1, -2, 0, 4, 5, 2, 0, 0, 0, 2, 0, 0, 0, -1, -1, 0, 1, 4, 2, 2, 0, -1, -2, -3, -3, -4, -4, -2, 0, 5, 5, 3, 2, 2, 1, 2, 1, 0, 0, 0, 0, 0, 2, 3, 3, 2, 0, -2, -5, -4, -4, -3, -3, -2, 0, 6, 8, 3, 3, 2, 2, 1, 0, 1, 0, 0, 0, 1, 3, 4, 2, 0, -3, -3, -6, -6, -3, 0, -2, -1, 0, 6, 8, 4, 3, 2, 1, 2, 1, 0, 0, -1, -1, 0, 0, 1, 0, 0, -4, -5, -7, -4, -2, 0, 0, 1, 3, 9, 11, 7, 5, 5, 3, 1, 0, -1, -1, -4, -3, -2, -2, -1, 0, -3, -6, -8, -8, -6, -2, 1, 3, 3, 5, 12, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, 2, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 2, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 2, 1, 0, 1, 0, 1, 0, 1, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, -1, 0, 1, 1, 0, 0, 1, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 2, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 2, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 2, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 1, 0, -1, 0, 0, -2, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 2, 2, 3, 2, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 3, 0, -1, 0, 0, 0, 0, -1, -1, -2, 0, 0, -1, 0, 0, 1, 2, 0, 1, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, -1, -1, -1, 0, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 1, 0, -2, 0, -1, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, 0, -1, 0, -2, -1, -1, 0, 0, 0, 0, -1, -2, -1, 0, 0, -1, 0, 0, 2, 1, 0, 0, 1, 0, -1, 0, -1, 0, 2, -2, -1, 0, -1, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 2, 1, 1, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, -2, -1, 0, -1, 0, -1, -1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 1, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -2, -1, 0, 0, 2, 2, 0, 0, -1, -1, 0, 0, -1, 1, 1, 0, -2, 0, 0, 1, 1, 3, 1, 0, 0, -1, -1, -2, 0, 0, 3, 2, 1, -1, 0, -1, 0, 0, 0, 1, 2, 0, 0, 0, 0, 2, 1, 2, 1, 0, 0, 0, -1, 0, 0, 2, 2, 1, 0, 0, 0, 0, -1, 0, 1, 2, 2, 0, -1, 1, 1, 1, 3, 2, 0, 0, -1, -1, -1, -1, 0, 2, 2, 2, 1, 0, 0, 0, 0, 0, 1, 0, 2, 0, -2, 0, 1, 2, 2, 0, 0, -1, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, -3, -3, 0, 0, 2, 0, 0, -1, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 2, 3, -2, -2, -1, -1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 3, -2, -3, -1, -1, 0, 1, 1, 0, 0, -2, -2, -2, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 1, 0, -2, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, -1, 0, 0, 0, 2, -2, -1, -2, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 1, 0, 2, 1, 0, -1, -2, 0, -1, 0, 0, 2, -1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -1, 2, 0, 2, 0, 0, 0, -1, 0, -2, -1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 1, 1, 2, 1, 1, 1, 0, 0, 0, -2, 0, -1, 0, 1, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 2, 1, 2, 1, -1, -1, 0, -2, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, -1, -2, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 0, 0, -1, -1, 0, 0, 0, 2, 0, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -1, 2, 1, 1, 2, 4, 4, 1, 1, 1, 0, 0, -1, 0, 0, -2, -1, 0, -1, 0, 0, 1, 0, 0, -2, 0, 0, 1, 3, 3, 3, 5, -4, -3, -1, 0, 3, 3, 2, 2, 2, 1, 2, 2, 5, 7, 7, 10, 9, 6, 4, 2, 2, 0, -2, -3, -3, -5, -2, -1, 0, 0, 1, 3, 3, 1, 0, 0, 0, 2, 3, 3, 4, 5, 6, 2, 2, 0, 0, -2, -2, -2, -1, -2, -3, -2, 0, 0, 0, 2, 0, 0, -1, -3, -2, 0, 2, 2, 0, 3, 1, 1, 0, -2, -1, -1, -2, 0, -2, -2, -2, 0, 0, 0, -1, 0, 0, -1, -3, -5, -2, -1, 2, 0, 0, 0, 2, 0, 0, -2, -2, -3, 0, 0, 0, -2, -1, -1, 0, -2, -3, -1, -2, -2, -4, -4, -2, -2, 0, 0, 0, 1, 0, 0, 0, -2, -1, -1, -1, 0, -1, -3, -2, -1, 0, -2, -3, -3, -2, -4, -5, -3, -3, 0, 0, 0, 0, 1, 1, 1, 0, -3, -4, -2, -1, -2, -1, -2, 0, 0, 1, 0, -1, -3, -2, -2, -3, -3, -1, 0, 3, 2, 1, 1, 2, 1, 0, -2, -3, -2, -2, -2, -2, -4, 0, 2, 2, 0, -2, -2, -2, -3, -4, -2, -1, 1, 3, 3, 2, 3, 4, 3, 1, 0, -2, 0, 0, -2, -3, -3, 1, 1, 3, 2, -1, -4, -3, -3, -2, 0, 1, 3, 3, 1, 3, 1, 1, 1, 0, 0, -1, -1, -2, -2, -3, -4, 0, 2, 2, 2, 0, -2, -4, -3, -3, 0, 2, 1, 2, 2, 2, 1, 1, 0, -1, -1, -3, -2, -2, -4, -3, -3, -1, 0, 3, 2, 0, -1, -3, -3, -2, 1, 1, 2, 2, 2, 2, 0, 0, -1, -1, -2, -1, -2, -3, -3, -2, -4, -1, 2, 3, 1, 0, -1, -2, -3, -1, -1, 1, 0, 1, 0, 0, 0, 0, -1, -4, -3, -4, -3, -3, -5, -3, -4, 0, 1, 1, 2, -1, -1, -2, -2, -3, -2, -1, 0, 0, 1, 0, 1, 0, -2, -3, -4, -3, -1, -3, -4, -4, -3, 0, 0, 2, 1, 0, -2, -3, -3, -4, -2, 0, 0, 1, 1, 1, 0, 0, 0, -3, -4, -3, -1, -2, -3, -3, -5, 0, 2, 3, 2, 1, -1, -3, -3, -2, -3, 0, 0, 0, 2, 1, 2, 1, 0, -4, -3, -3, -4, -4, -3, -3, -4, 0, 4, 5, 1, 1, -1, -1, -3, -2, 0, -1, 1, 0, 2, 3, 2, 1, 0, -2, -4, -5, -4, -5, -4, -4, -3, 1, 3, 5, 3, 0, 0, -3, -4, -3, -2, 0, 0, 1, 2, 2, 1, 0, 0, 0, -4, -5, -4, -4, -2, -2, -3, 2, 4, 3, 1, 0, -1, -3, -5, -5, -2, -1, 0, 0, 0, 2, 0, 0, -1, 0, -4, -5, -5, -4, -3, -1, -4, 0, 1, 3, 1, -1, -3, -3, -3, -4, -2, 0, -1, 0, 0, 3, 0, 1, -1, 0, -3, -4, -5, -5, -4, -3, -2, 0, 2, 1, 0, -1, -3, -3, -3, -2, -1, 0, 1, 0, 0, 1, 1, 1, 1, 0, -3, -4, -6, -6, -3, -4, -2, 0, 2, 1, 1, 0, -1, -2, -2, -1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, -1, -4, -5, -4, -2, -3, -4, -1, 2, 3, 1, 0, -1, -1, -1, -1, 0, 1, 1, 3, 2, 3, 3, 2, 3, 0, -1, -2, -4, -2, -1, -1, -2, 0, 3, 3, 4, 3, 0, 1, 0, 0, 1, 1, 3, 4, 3, 3, 1, 3, 2, 0, 0, -3, -3, -4, 0, -2, -3, 0, 4, 4, 3, 5, 2, 1, 0, 0, 1, 3, 4, 2, 1, 3, 2, 1, 2, 2, 0, -3, -2, -2, -1, -2, -2, 0, 3, 3, 3, 4, 2, 2, 1, 0, 0, 3, 3, 3, 5, 2, 4, 4, 3, 2, 2, -2, 0, -1, 0, -1, -4, 0, 2, 3, 3, 4, 3, 2, 3, 3, 2, 2, 4, 6, 5, 6, 6, 8, 7, 6, 3, 0, 0, 1, 0, -2, -4, -2, -1, -1, -2, -1, 0, 0, -1, -1, -1, 0, 0, 2, 2, 3, 2, 0, 0, 0, 2, 3, 2, 3, 2, 4, 4, -3, -1, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 3, 2, 3, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -2, 0, -1, 0, 1, 2, 4, -2, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 1, -1, -1, 0, -2, -1, -1, -1, 0, 0, 2, -2, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -1, -1, 0, 2, -2, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, 0, -1, -2, -3, -2, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, -2, -1, 0, -2, -2, -2, 0, 3, -1, 0, 0, -1, 0, 1, -1, 0, 0, 0, -1, 0, 1, 1, 1, 2, 0, -1, -1, -1, 0, 0, -1, -1, 0, 2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 3, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 2, 0, -1, -2, 0, -1, -1, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 2, 2, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 1, -1, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 1, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 2, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, -2, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -2, -2, -2, -1, -1, -1, 0, 0, 2, -1, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -2, -1, -2, -1, 0, -1, -1, 0, 1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, -2, -2, 0, -1, 2, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, 0, 2, -2, -1, 0, 1, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 4, -2, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 4, -1, -2, -1, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 2, 1, 0, 1, 2, 3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 1, 3, 3, 2, 3, 3, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -1, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -2, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 2, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 1, 0, 1, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 3, 1, 2, 2, 1, 0, 0, 0, 0, -1, 0, -2, 0, 0, -1, -1, -1, -1, 0, -1, -1, -1, 0, 0, 1, 0, 4, 1, 0, 0, 1, 0, 1, -1, -1, -1, 0, -1, -2, -1, 0, -2, -3, -4, -2, -1, -3, -1, 0, -1, -1, 0, 4, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -2, -1, -2, -2, -1, -1, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, -2, -1, -1, -1, 0, -1, -1, -1, 1, 0, 1, 0, 1, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, -2, 0, -2, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 2, 0, 0, 1, 0, 0, -1, -1, -1, -1, -1, 0, -1, 1, 1, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 2, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 1, 2, 2, 2, 1, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 0, 0, -1, -1, 0, 0, -1, 0, -2, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, 0, 1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 2, 1, 0, 1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, 0, 2, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -1, 0, -1, 0, 0, -1, -1, 4, 1, 0, 0, 0, 1, 0, -1, -1, 0, 0, -1, -2, 0, -1, -2, -1, -2, -3, -3, 0, -1, 0, 0, 0, -1, 9, 7, 5, 3, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -3, -3, -3, -3, -2, 0, 1, 2, 4, 7, 4, 3, 2, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, -1, -1, -2, -2, -3, -3, -1, 0, 0, 0, 0, 7, 4, 2, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -3, -2, -2, -1, -2, -2, -2, 0, 5, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -3, -3, -3, -2, 0, 5, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, -2, -1, -2, -4, -4, -2, -3, -2, -3, -1, 6, 1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, -2, -4, -4, -2, -2, -2, -3, 5, 0, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -3, -2, -3, -2, -3, -2, -4, 2, 0, -2, -1, -2, -1, -1, 0, -1, -1, -1, 0, 1, -1, 0, -1, -1, 0, -1, -1, -1, -2, -2, -3, -1, -2, 2, -1, -1, -2, 0, -2, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -3, -3, -1, -2, -2, 2, 0, -1, -1, -1, -3, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -3, -3, -3, -1, -1, -2, 5, 1, 0, 0, -1, -3, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, 0, 0, 0, 5, 2, 0, -1, 0, 0, 0, 1, 1, 1, 0, 1, 0, -1, 1, 0, 2, 0, 0, 0, -1, -1, -1, -1, 0, 0, 6, 2, 0, -1, 0, 0, 0, 1, 3, 2, 1, 0, 1, 1, 0, 2, 2, 1, 1, 0, -1, -2, -1, -2, -1, -1, 6, 1, 0, 0, 0, -1, 1, 1, 1, 1, 1, 0, 0, 1, 2, 3, 2, 2, 0, 1, -1, -2, -1, 0, -2, 0, 4, 2, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 1, 0, 0, -1, 0, 0, -3, 0, -2, -1, 0, 4, 0, -2, -2, -3, -1, -1, 0, 0, 1, 0, 2, 1, 1, 2, 2, 0, 0, -1, -1, -2, -1, -1, -2, -1, 0, 4, 0, -3, -2, -1, -1, -1, 0, 0, 0, 2, 2, 0, 1, 1, 2, 0, -1, -2, -2, -2, -1, -1, -1, -1, 0, 5, 0, -2, -2, -2, -1, -1, -1, 0, 1, 1, 0, 1, 1, 0, 2, 0, -1, -1, -1, -1, -2, -3, -1, -2, -2, 6, 0, 0, 0, -1, 0, 0, 1, 1, 2, 1, 1, 0, 1, 0, 0, 0, 0, -2, -2, 0, -2, -3, -1, -3, -2, 6, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 1, -2, 0, 0, -1, -2, -2, -3, -1, -1, 5, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, -2, -2, -2, -2, -1, -3, -1, -1, 6, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, -2, -2, 0, -2, -3, -3, -2, -1, 4, 4, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, -2, -2, 0, -1, -2, -3, -3, -2, -1, 6, 2, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -2, -3, -3, -2, -2, -2, 0, 6, 4, 1, 0, 0, -1, 0, 1, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -3, -1, 0, 0, 0, 0, 7, 5, 2, 0, 0, 0, 0, 2, 0, 1, 0, 1, 1, 0, 0, 1, 1, 0, -1, -3, -1, -2, 0, -1, 1, 2, 5, 2, 0, 0, -2, 0, -1, -2, -1, -4, -4, -4, -2, -2, -3, -5, -3, -6, -5, -3, -3, 0, 0, 2, 3, 4, 4, 1, -1, -1, -1, 0, -1, 0, -1, 0, -1, -1, -2, 0, -2, -2, -3, -3, -2, -4, -3, -1, 0, 0, 1, 2, 2, 2, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -3, -1, -3, -2, -3, -3, -1, -2, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 2, 0, 0, 0, -2, -2, -3, -3, -3, -3, -1, -1, 0, 3, 2, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 3, 2, 0, -1, -3, -2, -2, -2, -4, -4, -2, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 1, 0, 1, 1, 3, 3, 1, 0, -1, -3, -3, -3, -2, -4, -2, -2, -1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 3, 4, 1, 0, 0, -3, -3, -3, -2, -4, -3, -3, 0, 1, 2, 0, 1, 0, 1, 1, 0, 0, 1, 1, 1, 2, 3, 4, 3, 0, 0, -2, -1, -1, -2, -5, -4, -3, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 2, 2, 2, 4, 3, 1, 0, -1, -2, 0, -2, -2, -4, -2, -1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 2, 2, 2, 4, 5, 2, 2, 0, -1, -2, 0, 0, -1, -4, -3, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 4, 5, 4, 3, 1, 0, 0, -2, -1, 0, -1, -2, -2, -1, 0, 1, 0, 0, 0, 0, -1, 0, 1, 2, 2, 1, 4, 5, 6, 5, 3, 1, -1, 0, -1, 0, 0, -2, -2, -2, 1, 1, 0, 0, -1, -1, 0, 0, 1, 1, 1, 2, 2, 3, 5, 3, 2, 0, -2, -2, 0, 0, -2, -1, -1, -1, 1, 2, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 4, 4, 4, 5, 2, 1, 0, 0, -1, -1, -2, -2, -3, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 3, 4, 4, 3, 3, 1, 0, 0, -2, -2, -1, -2, -1, -2, -1, 1, -1, 0, -1, 0, 0, 0, 1, 0, 1, 1, 2, 3, 4, 4, 3, 1, 0, -1, -1, -2, -2, 0, -2, -3, -1, 0, 0, -1, 0, 0, 0, 1, 2, 1, 1, 2, 3, 2, 2, 3, 2, 1, 0, -1, -1, -2, -2, -2, -1, -2, 0, 1, -1, 0, -1, 0, 0, 0, 2, 2, 2, 3, 2, 3, 2, 2, 1, 0, -1, 0, -1, 0, -1, -3, -3, -2, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 3, 3, 2, 0, 1, 0, -1, -2, -2, -2, -2, -3, -2, -2, -1, 0, 0, -1, 0, 0, 1, 1, 1, 0, 1, 1, 2, 3, 2, 2, 0, -1, -1, -2, -2, -2, -3, -4, -3, -3, 0, 1, 0, -1, 0, 0, 2, 1, 0, 0, 1, 2, 3, 4, 3, 0, 0, 0, -1, -2, -1, -3, -1, -2, -5, -3, 0, 1, 1, 0, 1, 0, 0, 0, 0, 2, 2, 1, 2, 3, 2, 1, 1, 0, 0, -1, -2, -2, -3, -4, -4, -4, 0, 3, 1, 0, 2, 0, 1, 1, 1, 2, 0, 1, 2, 2, 2, 1, 0, 0, -2, -2, -1, -1, -3, -2, -2, -3, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 1, 1, 2, 0, 2, 1, 0, 0, -2, -4, -2, -2, -2, -3, -2, -1, 0, 2, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -3, -3, -5, -3, -1, -3, -1, -3, -1, 1, 3, 2, 3, 0, 1, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, -4, -5, -6, -4, -3, -2, -2, -1, -1, 0, 3, 8, 3, 0, -2, -2, -3, -3, -3, -3, -2, -4, -5, -5, -6, -6, -7, -8, -10, -10, -9, -9, -9, -7, -7, -7, -8, 7, 2, 0, -2, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -4, -5, -7, -7, -4, -3, -5, -4, -3, -5, -8, 8, 4, 0, 0, 0, 0, 1, 2, 3, 3, 2, 2, 3, 3, 3, 1, -2, -1, -2, -4, -3, -2, -2, -2, -4, -5, 6, 4, 1, 0, 0, 2, 1, 1, 2, 3, 3, 4, 4, 4, 2, 2, 0, 0, -2, 0, 0, -1, -3, -1, -5, -7, 5, 3, 1, 0, -1, 2, 1, 1, 3, 3, 1, 4, 3, 4, 3, 2, 0, 0, 0, 0, -1, -2, -2, -3, -4, -6, 5, 2, 0, -1, 0, 2, 2, 1, 1, 1, 3, 3, 3, 3, 1, 1, 0, 0, 0, -1, 0, -2, -2, -3, -4, -4, 3, 1, 0, 0, 1, 2, 1, 1, 1, 1, 4, 4, 2, 3, 2, 1, 1, 0, -1, -2, 0, -2, -1, -4, -4, -5, 1, 1, 0, 0, 1, 2, 1, 0, 0, 2, 3, 3, 3, 3, 1, 0, 1, 1, -1, -1, -2, -2, -3, -3, -4, -5, 0, 0, 0, -1, 0, 2, 1, 0, 0, 1, 2, 2, 2, 3, 3, 3, 3, 2, 0, -1, 0, -3, -3, -4, -6, -5, 2, -1, 0, -2, -1, 0, 0, 0, 0, 1, 2, 2, 2, 3, 3, 2, 4, 2, 1, 0, -1, -3, -3, -3, -4, -6, 1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 1, 1, 2, 2, 4, 5, 5, 3, 1, 0, -1, -3, -2, -2, -5, -5, 3, 1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 3, 4, 5, 4, 2, 1, 0, -1, -3, -3, -5, -4, 4, 1, 0, 0, 0, -1, -1, 2, 1, 1, 1, 2, 2, 1, 3, 4, 5, 6, 3, 3, 1, -1, -1, -3, -4, -5, 3, 2, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 1, 2, 4, 7, 5, 5, 1, 1, -1, 0, -1, -2, -5, 4, 1, 0, 0, 1, 2, 1, 3, 3, 4, 3, 3, 2, 2, 3, 3, 7, 5, 3, 2, 1, 0, -1, -1, -4, -4, 3, 2, 0, 0, 0, 3, 1, 4, 5, 3, 2, 3, 1, 2, 4, 5, 3, 4, 1, 0, 0, 0, 0, -2, -3, -4, 3, 1, 0, 0, 0, 3, 1, 4, 5, 4, 4, 3, 2, 2, 4, 4, 3, 3, 0, 1, 1, 0, 0, 0, -1, -3, 2, 0, 0, 0, 0, 1, 2, 4, 4, 4, 4, 3, 1, 1, 4, 4, 2, 2, 0, 0, 1, 0, 1, -1, -3, -5, 2, 0, 0, 0, 0, 0, 2, 2, 3, 2, 2, 0, 0, 2, 3, 4, 2, 2, -1, 0, 0, 0, 1, 0, -3, -4, 4, 0, 0, -2, 0, 1, 3, 3, 3, 3, 0, 0, 0, 1, 3, 2, 1, 0, 0, -1, -1, 0, -1, 0, -2, -5, 5, 0, 0, -2, -1, 0, 1, 2, 3, 2, 0, 0, 0, 1, 1, 0, 0, -2, -1, -2, 0, -2, 0, 0, -2, -5, 6, 2, 0, 0, -1, 0, 1, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, -1, -2, -2, -1, -1, 0, -1, -2, -6, 5, 4, 2, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, -1, -1, -2, -1, -2, -2, -3, -1, 0, -1, -6, 6, 2, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, -2, -1, -1, -3, -1, -1, -2, -3, -4, -1, -2, -4, -8, 5, 3, 1, -1, 0, 0, 0, -1, 0, -2, -1, -2, -3, -4, -3, -3, -4, -3, -5, -5, -5, -5, -3, -4, -6, -8, 5, 3, 1, 0, -1, -1, 0, -1, -2, -3, -3, -3, -4, -5, -8, -8, -7, -7, -7, -8, -7, -8, -7, -8, -7, -10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, 0, 0, 1, -1, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 2, 3, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 2, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 2, 2, 0, 1, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -2, 0, 0, -1, -1, 0, 0, 0, -1, -2, -1, -2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, -1, 0, 0, 0, -1, -2, -1, 0, 0, 0, 1, 1, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 1, 1, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 1, 1, 2, 0, 2, 2, 1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 2, 0, 1, 1, 2, 2, 0, -1, 0, -1, 0, 0, 0, 1, 2, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 1, 2, 2, 2, 1, 2, 1, 1, 0, 0, 0, 0, -1, 0, 1, 2, 2, 2, 2, 1, 1, 1, 1, 0, 2, 1, 0, 1, 2, 2, 2, 1, 1, 0, 1, 0, 0, 0, -1, 2, 2, 2, 2, 3, 2, 1, 0, 0, 0, 0, 2, 1, 2, 1, 2, 2, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 3, 1, -1, -1, 0, 1, 0, 0, 1, 2, 3, 2, 3, 2, 0, 0, 0, 1, 0, 0, -2, 0, 0, 2, 3, 3, 1, 0, -1, -1, 0, 0, 0, 2, 1, 1, 2, 3, 1, 2, 1, 0, 1, 1, 0, 0, 0, 2, 1, 3, 3, 3, 3, 1, 0, 0, 1, 0, 2, 2, 1, 3, 3, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 1, 2, 1, 1, -1, -1, 0, 1, 0, 0, 1, 3, 1, 1, 1, 1, 0, 0, 0, 1, 0, -1, -1, 2, 1, 2, 2, 1, 3, 2, 0, 0, 0, 2, 1, 1, 0, 2, 1, 1, 2, 1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 1, 1, 2, 2, 2, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, 2, 0, 2, 1, 0, 2, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 1, 1, 0, -1, -1, -1, 0, 0, -1, 0, 1, 0, 0, 1, 1, 0, 2, 1, 0, 0, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 1, 0, 1, 1, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, 0, -1, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 2, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 1, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, -4, -2, -6, -5, -5, -3, 0, 0, -1, 0, -1, -3, -3, -5, -5, -3, -4, -4, -3, -4, -5, -7, -8, -11, -1, -1, -2, -5, -3, -5, -2, 0, 0, 2, 1, 0, 0, 0, 0, 0, -2, -1, -2, -1, -1, 0, -3, -4, -5, -9, 0, 0, -2, -1, -2, -2, -1, 0, 0, 1, 3, 3, 3, 2, 2, 1, 0, 0, 0, 1, 0, 0, -1, -2, -4, -6, 0, 0, 0, -1, -2, -2, 0, -1, 1, 3, 3, 5, 5, 6, 4, 2, 1, 0, 1, 2, 2, 3, 0, -1, -2, -3, 1, 0, 0, -2, -3, -2, -1, -1, 0, 2, 3, 6, 8, 7, 5, 5, 4, 2, 1, 2, 3, 2, 1, 0, 0, -2, 0, 0, 0, -2, -1, 0, 0, 0, 1, 3, 3, 4, 6, 8, 5, 5, 3, 3, 2, 1, 2, 3, 1, 0, -1, -1, 1, 0, 0, -2, -2, 0, 0, -1, 0, 0, 3, 5, 6, 6, 6, 4, 3, 2, 1, 1, 0, 0, 1, -1, -1, -2, 0, 0, 0, -1, 0, 0, 0, 0, 2, 2, 4, 5, 6, 6, 3, 4, 4, 2, 2, 1, 1, 1, 0, 0, -1, -3, 0, 0, -1, 0, -2, 0, 0, 3, 4, 3, 3, 3, 4, 4, 3, 3, 3, 2, 4, 2, 1, -1, 0, -1, -2, -3, -2, -3, -3, -2, -3, -1, 2, 3, 3, 2, 4, 3, 1, 3, 3, 3, 2, 3, 1, 1, 0, -1, -1, -2, -4, -6, -1, -5, -5, -5, -3, 0, 0, 1, 1, 2, 2, 2, 2, 1, 3, 1, 2, 2, 3, 1, 0, -2, -3, -2, -3, -5, -2, -3, -5, -5, -3, -1, 0, 0, 0, 1, 3, 1, 0, 0, 1, 3, 2, 1, 3, 1, 0, -2, -3, -4, -4, -4, -2, -4, -4, -3, -3, -1, -1, 0, 1, 1, 1, 2, 1, 1, 1, 2, 3, 3, 2, 4, 1, -2, -2, -3, -2, -4, -5, -5, -5, -2, -1, 0, 0, 0, 2, 0, 1, 1, 1, 1, 1, 2, 2, 3, 4, 3, 1, 0, -3, 0, -3, -2, -5, -3, -3, -4, 0, -1, 0, 0, 1, 2, 2, 3, 2, 1, 2, 4, 6, 6, 5, 5, 2, 0, 0, 0, -1, -1, -3, -4, -4, -2, -2, 0, 0, 1, 4, 4, 3, 3, 0, 2, 4, 4, 6, 4, 6, 4, 2, 2, 1, 0, 0, -1, -4, -3, -4, -3, -1, 0, 1, 1, 4, 3, 3, 3, 2, 1, 2, 4, 5, 6, 3, 4, 3, 3, 1, 2, 0, 0, -2, -1, -3, -3, -1, -1, 2, 4, 4, 3, 2, 3, 1, 2, 1, 3, 4, 4, 4, 3, 3, 2, 1, 2, 1, 0, 0, -2, -2, -2, 0, 0, 1, 3, 2, 4, 3, 2, 1, 1, 2, 4, 4, 4, 1, 1, 1, 2, 3, 2, 3, 0, -2, 0, -2, -2, -2, -1, 0, 2, 2, 1, 1, 0, 1, 1, 2, 3, 3, 3, 2, 1, 1, 0, 2, 3, 2, 0, 0, 0, -1, -1, -3, -2, 0, 1, 2, 1, 0, 1, 0, 1, 2, 3, 2, 2, 1, 1, 0, 0, 2, 2, 1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 1, 1, 1, 2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 0, -1, 1, 0, 0, 0, -1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, -2, 0, 1, 1, 0, 0, 0, 1, 0, -1, -2, 0, 0, -2, -2, -1, 0, 0, 0, 0, -1, -2, -1, 0, 0, -1, -6, 0, 0, 1, -1, 0, 0, 0, -1, -4, -2, -1, -2, -1, -4, -2, -2, -1, 0, -1, -4, -3, -3, -2, -4, -5, -8, 10, 7, 3, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, -2, -3, -1, 0, 0, 1, 3, 7, 5, 3, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -2, -2, -2, -1, -2, 0, 0, 1, 6, 3, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -3, -3, -2, -3, 0, 6, 2, 1, 1, 0, 0, 0, 0, 0, -2, 0, -2, -1, 0, -1, 0, 0, 1, 0, 0, -2, -3, -3, -4, -4, -2, 2, 1, 0, 0, 0, 1, 0, -1, -1, -3, -2, -1, -2, -2, 0, 1, 1, 0, 0, 0, 0, -2, -2, -5, -2, -1, 0, -1, 0, 0, 2, 0, 1, 0, 0, -3, -2, -1, -2, -1, 0, 1, 1, 0, 1, 0, 0, 0, -3, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -3, -2, -1, -1, -3, -1, -1, 0, 1, 1, 0, -2, 0, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, -2, 0, 0, -1, -1, -2, 0, 0, 0, 1, -1, -1, -2, -1, -2, 0, -1, 0, 0, 1, 0, -1, 0, -1, -1, -2, -1, 1, 0, -1, -2, -1, 0, 0, 2, 0, 0, -2, -2, 0, -1, 0, 0, 1, 0, 1, 1, 0, -1, -1, -1, -1, 0, 1, 3, 0, 0, 0, 1, 1, 2, 1, 0, 0, -2, -2, -1, 0, 1, 1, 3, 2, 1, 0, -1, -1, 0, 0, -1, 0, 5, 0, 0, 1, 1, 4, 4, 1, 0, 0, -2, -1, 0, 0, 1, 2, 4, 3, 1, -1, 0, -1, 0, 0, 0, 2, 3, 0, 0, 0, 2, 3, 4, 1, 0, 0, -1, -2, 0, 0, 1, 2, 4, 2, 1, -1, -1, -1, 0, 0, 0, 1, 3, -1, -1, 0, 2, 3, 2, 2, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 3, 0, -1, -1, -2, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, -1, -3, -1, 0, 0, 1, 1, 0, -1, -1, 0, -1, 0, 2, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 2, -1, -1, 0, -1, 1, 0, 0, 0, 0, -1, 0, -1, 1, 2, 2, 2, 2, 0, 0, -1, -1, 0, 0, -1, 1, 1, -1, -2, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 2, 2, 3, 1, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, -1, -1, 1, 2, 1, 0, 1, 0, -2, 0, 0, 0, 2, 3, 3, 3, 1, 0, -2, -2, -1, -1, 0, 0, 4, 1, 0, 1, 0, 2, 1, 1, 0, -1, 0, 0, 0, 1, 3, 1, 1, 2, 2, 0, -2, -2, -1, -2, 0, -1, 5, 2, 0, 1, 1, 2, 1, 1, 0, 0, -1, 0, 1, 0, 1, 0, 0, 1, 1, 0, -1, -1, -1, -2, -2, 0, 6, 3, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 2, 2, 2, 0, 0, -1, -1, -3, -2, -1, 0, 0, 6, 4, 1, 2, 0, 1, 0, 0, -1, -1, 0, 0, 1, 0, 1, 1, 1, 0, 0, -1, -3, -1, -1, -2, 0, 1, 7, 4, 0, 0, 2, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -1, 0, 0, 2, 10, 4, 3, 1, 2, 2, 0, 0, 0, -1, -3, -2, -1, 0, -1, 0, 0, -1, -1, -3, -2, 0, 1, 1, 1, 3, 11, 6, 5, 2, 0, 0, 0, 0, -1, -1, -2, -4, -3, -3, -3, -3, -3, -4, -4, -2, -2, 0, 0, 3, 5, 6, -1, 0, 0, 0, 1, 1, 2, 0, 0, -1, 0, 0, 0, 2, 1, 0, 1, 2, 3, 4, 4, 4, 4, 5, 6, 8, 0, 0, 0, 0, 1, 3, 0, 0, -1, -2, -1, -3, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 3, 4, 7, 1, 1, 0, 2, 3, 3, 0, 1, 0, -2, -1, -2, 0, 0, -1, -2, -2, -1, -2, -1, -2, -1, 0, 0, 1, 6, 2, 1, 1, 2, 3, 2, 0, 0, 0, -1, -1, -1, -2, 0, 0, 0, -2, -2, -4, -3, -4, -3, -1, 0, 1, 6, 1, 2, 0, 1, 2, 1, 2, 1, -1, 0, 0, 0, -2, 0, 0, 0, -3, -3, -3, -3, -2, -3, -3, -1, 2, 4, 1, 2, 2, 1, 2, 1, 0, 1, 0, 0, -2, -1, -2, 0, 0, 0, -1, -2, -3, -2, -2, -2, -3, 0, 0, 6, 1, 1, 2, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -2, -4, -2, -1, -2, -3, -2, 0, 5, 0, 0, 1, 0, 1, 0, 0, 0, -1, -2, -1, -1, 0, 0, 1, 0, 0, -1, -4, -3, -1, -1, -1, 0, 0, 4, 0, 1, 1, 1, 1, 0, 0, -1, 0, -1, 0, -1, 1, 2, 1, 0, 0, -1, -3, -2, 0, 0, 0, -1, 0, 3, -1, 1, 1, 1, 0, 1, -1, 0, 0, -1, 0, 0, 0, 2, 2, 0, 0, -2, -2, -1, 0, 1, 0, 0, 0, 2, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 0, -1, -2, -1, -1, 1, 0, 0, -1, 0, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, -1, -3, -3, -1, -1, 0, 0, -1, 0, 2, 0, 0, 0, 0, -1, -1, 0, -2, 0, 0, 0, 1, 1, 2, 0, 0, -2, -4, -5, -3, 0, 0, 0, -1, -1, 2, -1, 0, 0, -2, -2, -1, -3, 0, 0, 0, 0, 0, 0, 0, 1, -1, -2, -2, -3, -3, 0, 0, 0, -1, -2, 1, 0, 1, 1, 0, -1, -3, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, -1, -3, -3, -1, 0, 0, 0, -1, -2, 2, 0, 1, 0, 0, -2, 0, -2, 0, 2, 1, 0, 0, 1, 1, -1, -2, -2, -3, -1, -1, 0, 0, -2, -3, -1, 3, 0, 2, 0, 1, -1, -2, -2, 0, 1, 2, 1, 0, 1, 0, 0, -1, -3, -4, -2, -3, -2, -3, -2, -4, -1, 2, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, -2, -3, -4, -2, -3, 0, -1, -3, -2, -2, 3, 0, 1, 0, 1, 0, -1, -2, 0, 0, 0, 0, 0, 1, 0, -2, -3, -3, -2, -2, -2, -1, -3, -3, -2, -1, 4, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -3, -2, -1, -2, -2, -1, -3, -3, 0, 2, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 1, 1, 1, 0, -1, -2, -2, -3, -1, -2, 0, -1, -1, -2, -2, 4, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, -2, -1, -2, -1, 0, -2, -1, -3, -2, -1, 4, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, -2, -2, -2, 0, 0, 0, -2, -2, 1, 7, 0, 0, 2, 0, 3, 2, 1, 0, 1, 0, -1, -1, 0, 0, 0, -2, -3, -3, 0, 0, 1, 1, 0, 1, 1, 8, -1, 0, 0, 2, 2, 2, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 1, 3, 3, 3, 3, 6, 8, 0, -1, 1, 3, 2, 0, 0, 0, 1, -1, -2, -3, 0, 1, 1, 0, 1, 0, 2, 2, 5, 5, 5, 6, 8, 10, 15, 8, 3, 0, 0, -1, 0, -1, -2, -5, -6, -6, -6, -4, -5, -5, -6, -6, -9, -8, -7, -6, -5, -7, -5, -5, 14, 6, 1, 0, 0, 0, 2, 0, -1, -2, -1, -2, -1, 0, 0, -2, -4, -3, -5, -6, -5, -4, -5, -5, -6, -6, 12, 7, 3, 0, 0, 1, 2, 1, 1, 0, -1, 0, 0, 1, 2, 0, -2, -2, -2, -4, -2, -3, -2, -4, -5, -6, 12, 6, 3, 1, 1, 1, 3, 2, 2, 0, 0, 0, 2, 1, 2, -1, 0, -2, -2, -2, -2, -1, -2, -4, -3, -5, 8, 4, 2, 0, 0, 2, 1, 1, 0, -1, 0, 0, 2, 1, 0, -1, -2, -2, -2, 0, -1, -1, -3, -3, -3, -4, 6, 3, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 2, 1, 0, 0, -1, -2, -2, -1, -3, -3, -2, -2, -3, 4, 0, -2, -1, 0, 0, 1, 0, -2, -1, -1, 0, 1, 1, 0, 0, 1, 0, 0, -3, -3, -1, -1, -3, -4, -4, 4, 0, -1, -1, -1, 0, 0, -1, -2, -1, 0, 0, 1, 1, 2, 0, 0, 1, 0, -1, -1, -3, -2, -3, -3, -3, 4, 0, -1, -2, -2, 0, -2, -2, -3, -3, 0, 0, 1, 2, 3, 1, 2, 1, 0, -1, -2, -1, -2, -1, -3, -2, 5, 0, 0, -1, -2, -1, -1, -3, -1, 0, 0, 0, 0, 3, 3, 3, 2, 1, 0, -1, -1, -1, 0, -2, -1, -2, 6, 2, 0, 0, -2, 0, -2, -1, -2, 0, 0, 0, 0, 2, 4, 5, 6, 4, 2, 0, -1, 0, 0, -1, -1, -3, 8, 2, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 2, 5, 5, 6, 4, 3, 0, 0, 0, -1, -1, -1, -2, 7, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 6, 5, 4, 2, 0, 0, -1, -1, -2, 0, -1, 6, 2, 0, -1, -2, -2, 0, 0, 0, 0, 1, 0, 1, 3, 5, 7, 6, 4, 2, 2, 0, 0, 0, -2, 0, 0, 5, 0, 0, -1, -1, 0, 0, 1, 0, 2, 2, 0, 2, 3, 4, 5, 5, 5, 2, 1, 0, -1, 0, -1, 0, -2, 5, 0, 0, -1, -1, -1, 0, 0, 1, 3, 4, 3, 3, 4, 6, 7, 4, 3, 3, 1, 1, -1, 0, -1, -1, -2, 5, 0, -1, 0, -1, 0, 1, 0, 2, 2, 4, 3, 4, 6, 5, 5, 6, 2, 2, 1, 0, 0, 0, 0, -2, -2, 3, 0, 0, -2, 0, 0, 0, 2, 2, 1, 2, 2, 4, 4, 5, 5, 5, 2, 0, 0, 1, 0, 0, -1, -2, -2, 6, 2, 0, 0, 0, 1, 2, 3, 1, 1, 2, 1, 3, 4, 5, 5, 4, 2, 0, 0, 0, 1, 0, 0, -2, -2, 9, 3, 0, -1, 0, 2, 1, 1, 2, 0, 0, 0, 2, 4, 5, 3, 2, 1, 0, 0, 0, 0, 0, -2, -2, -3, 8, 5, 0, 0, 0, 1, 1, 1, 2, 1, 0, 0, 1, 2, 2, 3, 2, 0, 0, -1, -1, -2, -1, 0, -3, -3, 10, 5, 1, 0, -1, 0, 0, 1, 0, 1, 1, 0, 1, 1, 2, 0, 1, -1, 0, -1, -3, -1, -2, -1, -3, -4, 11, 7, 2, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, 0, -2, -3, -2, -2, -2, -3, -3, 11, 8, 4, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -4, -4, -5, -3, -4, -2, -1, -2, -3, 12, 8, 3, 2, 1, 1, 0, -1, -1, -1, -1, -2, -2, -3, -3, -4, -5, -5, -4, -5, -6, -4, -4, -2, -4, -3, 15, 11, 5, 3, 1, 0, -1, 0, -3, -3, -4, -5, -6, -6, -7, -8, -8, -7, -7, -7, -6, -6, -6, -3, -5, -5,

    others => 0);
end iwght_package;
