library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    80, 84, 85, 85, 81, 81, 83, 87, 82, 64, 54, 60, 66, 66, 66, 
    80, 83, 85, 85, 88, 104, 62, 67, 40, 48, 26, 20, 35, 55, 66, 
    52, 66, 86, 87, 89, 84, 52, 24, 29, 56, 43, 37, 10, 25, 61, 
    6, 57, 72, 86, 72, 64, 51, 31, 28, 60, 46, 35, 25, 10, 45, 
    26, 58, 58, 91, 83, 57, 47, 34, 20, 60, 52, 23, 33, 10, 18, 
    44, 76, 66, 83, 109, 75, 66, 35, 11, 98, 55, 28, 36, 23, 10, 
    53, 46, 53, 56, 69, 97, 69, 54, 18, 86, 43, 29, 31, 42, 31, 
    65, 54, 24, 40, 59, 100, 56, 48, 42, 89, 60, 28, 37, 47, 57, 
    70, 68, 32, 58, 55, 46, 46, 46, 47, 29, 60, 20, 35, 59, 71, 
    93, 79, 32, 51, 32, 42, 60, 49, 40, 50, 8, 1, 26, 62, 61, 
    81, 73, 31, 120, 56, 30, 62, 50, 16, 0, 1, 3, 2, 8, 4, 
    28, 69, 54, 119, 42, 20, 12, 10, 6, 2, 2, 3, 9, 9, 6, 
    0, 29, 88, 87, 19, 8, 0, 2, 2, 4, 4, 8, 5, 5, 17, 
    0, 0, 58, 46, 19, 9, 2, 1, 4, 6, 4, 5, 0, 18, 0, 
    0, 0, 0, 4, 1, 9, 10, 8, 11, 11, 2, 6, 28, 12, 0, 
    
    -- channel=1
    54, 52, 56, 57, 56, 50, 57, 59, 55, 45, 37, 39, 46, 51, 52, 
    56, 55, 59, 57, 59, 45, 54, 41, 32, 24, 24, 17, 19, 42, 51, 
    24, 42, 58, 57, 58, 17, 22, 14, 29, 20, 20, 23, 23, 27, 40, 
    24, 37, 55, 55, 40, 38, 32, 32, 23, 22, 14, 17, 15, 23, 33, 
    33, 33, 55, 62, 46, 41, 12, 17, 9, 27, 23, 28, 20, 26, 24, 
    17, 8, 51, 27, 0, 18, 14, 26, 15, 30, 12, 14, 20, 23, 31, 
    27, 0, 32, 38, 12, 22, 11, 22, 18, 11, 11, 16, 16, 23, 31, 
    17, 2, 34, 35, 46, 20, 2, 2, 23, 14, 12, 10, 18, 20, 39, 
    5, 0, 11, 16, 27, 2, 14, 12, 32, 11, 9, 3, 14, 35, 53, 
    0, 4, 6, 4, 21, 22, 21, 21, 18, 15, 7, 17, 32, 40, 42, 
    0, 4, 0, 21, 37, 40, 14, 0, 12, 7, 14, 19, 5, 0, 2, 
    0, 0, 27, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    
    -- channel=2
    35, 39, 40, 37, 36, 39, 43, 43, 39, 35, 27, 28, 29, 26, 23, 
    33, 44, 47, 41, 45, 27, 36, 37, 38, 7, 0, 0, 1, 22, 22, 
    16, 41, 39, 40, 45, 61, 3, 0, 0, 15, 0, 0, 0, 0, 19, 
    0, 0, 35, 45, 27, 30, 9, 0, 0, 39, 0, 0, 0, 0, 26, 
    0, 16, 22, 81, 44, 41, 3, 0, 0, 18, 8, 0, 0, 0, 0, 
    0, 6, 11, 34, 49, 36, 0, 0, 0, 48, 2, 0, 0, 0, 0, 
    0, 0, 14, 14, 50, 29, 40, 0, 0, 56, 0, 0, 0, 0, 0, 
    0, 2, 0, 10, 50, 72, 0, 2, 0, 39, 0, 0, 0, 0, 0, 
    1, 23, 0, 9, 0, 25, 0, 0, 3, 9, 11, 0, 0, 0, 23, 
    13, 20, 0, 21, 0, 0, 14, 6, 0, 5, 0, 0, 0, 27, 29, 
    30, 22, 0, 46, 0, 0, 37, 19, 0, 0, 0, 0, 0, 0, 0, 
    10, 14, 10, 78, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 22, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=3
    47, 47, 44, 47, 49, 44, 48, 53, 54, 51, 43, 37, 36, 42, 45, 
    46, 47, 47, 50, 45, 30, 51, 50, 49, 24, 20, 26, 30, 36, 42, 
    52, 36, 50, 51, 52, 60, 49, 40, 16, 0, 10, 2, 19, 23, 29, 
    43, 1, 50, 49, 53, 29, 24, 10, 6, 0, 18, 17, 17, 16, 15, 
    16, 0, 45, 20, 7, 0, 22, 14, 16, 0, 17, 19, 7, 12, 12, 
    10, 6, 38, 39, 20, 12, 21, 19, 21, 0, 21, 22, 7, 7, 4, 
    0, 25, 35, 53, 15, 2, 29, 11, 27, 0, 28, 17, 7, 3, 10, 
    0, 12, 13, 37, 14, 3, 19, 19, 19, 0, 21, 25, 3, 8, 15, 
    4, 1, 17, 5, 17, 22, 28, 20, 2, 36, 35, 24, 6, 11, 28, 
    8, 2, 23, 0, 24, 0, 0, 15, 9, 21, 22, 9, 0, 19, 45, 
    1, 6, 28, 0, 0, 0, 0, 6, 10, 9, 0, 0, 0, 16, 26, 
    0, 0, 1, 0, 55, 21, 7, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 28, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=4
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=5
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 18, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 38, 0, 0, 0, 11, 1, 0, 
    31, 25, 0, 0, 0, 53, 21, 16, 0, 0, 0, 0, 0, 14, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 13, 6, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 14, 
    13, 0, 0, 41, 45, 14, 0, 0, 0, 0, 11, 14, 0, 0, 0, 
    0, 2, 9, 0, 15, 0, 2, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 49, 33, 0, 0, 6, 2, 0, 13, 0, 
    0, 0, 2, 0, 0, 53, 0, 0, 0, 18, 19, 50, 19, 0, 0, 
    3, 0, 0, 0, 0, 12, 0, 0, 2, 36, 47, 3, 0, 0, 0, 
    0, 0, 8, 0, 0, 0, 0, 34, 10, 0, 0, 0, 0, 9, 7, 
    61, 19, 0, 0, 97, 66, 45, 40, 9, 4, 0, 3, 0, 0, 0, 
    0, 47, 0, 27, 64, 0, 0, 0, 0, 0, 0, 0, 1, 6, 0, 
    0, 0, 36, 65, 10, 0, 0, 0, 0, 0, 6, 12, 3, 0, 49, 
    3, 0, 14, 48, 24, 20, 20, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=6
    11, 15, 12, 15, 13, 17, 15, 8, 11, 19, 18, 14, 16, 12, 7, 
    12, 15, 11, 18, 12, 62, 37, 28, 17, 23, 55, 37, 12, 9, 15, 
    31, 0, 15, 12, 9, 14, 27, 6, 14, 43, 66, 46, 50, 5, 14, 
    74, 18, 24, 14, 36, 20, 69, 42, 39, 16, 70, 33, 30, 19, 0, 
    94, 90, 45, 5, 139, 95, 82, 50, 32, 0, 74, 64, 36, 41, 0, 
    76, 91, 53, 16, 33, 52, 103, 57, 62, 21, 100, 48, 29, 43, 34, 
    72, 117, 26, 36, 18, 62, 105, 81, 65, 44, 87, 53, 30, 40, 46, 
    95, 109, 60, 62, 23, 84, 89, 44, 43, 31, 69, 48, 23, 40, 14, 
    118, 106, 93, 57, 61, 16, 37, 56, 35, 53, 23, 24, 1, 12, 25, 
    96, 95, 110, 53, 79, 30, 36, 109, 52, 31, 34, 6, 27, 35, 29, 
    91, 99, 101, 60, 183, 116, 101, 102, 88, 50, 40, 61, 63, 68, 69, 
    57, 85, 97, 125, 141, 46, 39, 36, 49, 53, 61, 62, 68, 70, 71, 
    86, 47, 56, 156, 68, 62, 62, 55, 54, 58, 65, 76, 79, 72, 85, 
    82, 71, 36, 134, 64, 61, 69, 59, 56, 64, 68, 67, 69, 79, 91, 
    89, 69, 65, 46, 49, 42, 51, 60, 68, 77, 72, 58, 76, 113, 85, 
    
    -- channel=7
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=8
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 6, 0, 0, 6, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 5, 26, 4, 3, 0, 3, 0, 
    0, 25, 0, 0, 0, 3, 0, 0, 0, 36, 0, 8, 0, 0, 15, 
    0, 20, 0, 20, 0, 15, 1, 0, 0, 48, 9, 0, 3, 0, 12, 
    16, 29, 0, 15, 59, 32, 4, 0, 0, 76, 3, 0, 10, 0, 0, 
    22, 9, 6, 0, 31, 44, 8, 3, 0, 65, 0, 0, 11, 13, 0, 
    32, 11, 7, 0, 15, 42, 0, 14, 0, 45, 5, 0, 17, 10, 0, 
    27, 38, 0, 25, 9, 24, 6, 5, 16, 0, 18, 0, 15, 8, 0, 
    33, 39, 0, 45, 0, 19, 32, 0, 17, 4, 0, 0, 11, 8, 0, 
    50, 37, 0, 87, 0, 3, 39, 18, 0, 0, 7, 11, 21, 14, 2, 
    53, 49, 13, 72, 1, 19, 33, 32, 17, 14, 16, 22, 23, 25, 21, 
    16, 54, 72, 33, 0, 20, 16, 18, 15, 18, 23, 25, 23, 26, 32, 
    15, 24, 88, 0, 7, 23, 15, 18, 21, 24, 25, 25, 22, 38, 19, 
    13, 26, 33, 14, 10, 25, 20, 17, 23, 23, 17, 24, 40, 20, 0, 
    
    -- channel=9
    74, 83, 78, 80, 80, 76, 84, 91, 85, 76, 66, 63, 66, 67, 69, 
    75, 85, 85, 86, 82, 59, 76, 79, 81, 26, 7, 6, 22, 52, 66, 
    65, 68, 80, 86, 83, 101, 54, 28, 0, 0, 9, 5, 11, 9, 51, 
    35, 0, 74, 84, 76, 49, 33, 8, 0, 12, 26, 14, 8, 0, 27, 
    24, 2, 66, 65, 61, 32, 37, 7, 3, 0, 21, 14, 1, 3, 0, 
    0, 10, 60, 46, 40, 35, 33, 23, 8, 0, 33, 17, 6, 5, 0, 
    0, 24, 36, 84, 41, 7, 63, 22, 30, 0, 31, 0, 0, 0, 0, 
    0, 30, 0, 55, 33, 44, 46, 24, 18, 13, 26, 7, 0, 12, 27, 
    3, 10, 0, 10, 5, 32, 20, 8, 2, 38, 21, 24, 0, 11, 44, 
    21, 9, 16, 0, 19, 0, 4, 29, 0, 37, 30, 0, 0, 39, 69, 
    6, 11, 24, 0, 13, 0, 2, 36, 15, 0, 0, 0, 0, 0, 0, 
    0, 0, 17, 12, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 41, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=10
    52, 53, 58, 58, 59, 52, 59, 65, 65, 46, 35, 39, 48, 53, 56, 
    62, 62, 58, 58, 58, 66, 61, 53, 30, 32, 26, 23, 22, 39, 51, 
    30, 30, 61, 64, 58, 0, 47, 28, 27, 0, 0, 2, 9, 10, 36, 
    28, 22, 56, 63, 61, 42, 24, 10, 1, 0, 11, 0, 11, 16, 11, 
    16, 0, 51, 40, 28, 11, 5, 18, 0, 5, 9, 18, 6, 18, 6, 
    0, 0, 53, 32, 0, 5, 22, 14, 17, 0, 0, 12, 0, 7, 23, 
    6, 0, 30, 61, 0, 17, 0, 12, 7, 0, 2, 15, 2, 4, 9, 
    2, 0, 14, 39, 2, 0, 0, 0, 10, 0, 4, 9, 0, 0, 24, 
    0, 0, 11, 0, 24, 0, 15, 12, 2, 10, 0, 0, 0, 18, 40, 
    0, 0, 5, 0, 0, 4, 8, 3, 0, 0, 0, 7, 0, 28, 47, 
    0, 0, 0, 0, 31, 3, 0, 0, 0, 7, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=11
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=12
    30, 30, 37, 33, 34, 34, 33, 34, 36, 25, 14, 21, 26, 26, 27, 
    37, 38, 40, 32, 41, 63, 13, 25, 2, 25, 11, 6, 14, 22, 27, 
    12, 25, 34, 33, 43, 33, 0, 0, 16, 56, 2, 0, 0, 16, 30, 
    0, 77, 26, 40, 29, 31, 22, 6, 11, 57, 0, 10, 0, 0, 47, 
    0, 61, 0, 65, 32, 28, 0, 0, 0, 69, 7, 0, 17, 0, 32, 
    0, 20, 0, 52, 41, 0, 0, 0, 0, 142, 0, 0, 20, 0, 1, 
    0, 0, 0, 0, 70, 58, 0, 0, 0, 120, 0, 0, 18, 27, 0, 
    0, 0, 0, 0, 58, 72, 0, 0, 0, 89, 0, 0, 25, 16, 1, 
    0, 7, 0, 29, 17, 0, 0, 21, 23, 5, 23, 0, 23, 28, 43, 
    2, 12, 0, 52, 0, 10, 27, 12, 13, 0, 0, 0, 39, 56, 18, 
    47, 7, 0, 123, 0, 10, 55, 0, 0, 0, 11, 25, 21, 1, 0, 
    24, 6, 0, 114, 0, 0, 0, 0, 0, 0, 0, 2, 1, 5, 0, 
    0, 29, 38, 16, 0, 0, 0, 0, 0, 6, 8, 9, 0, 0, 7, 
    0, 0, 71, 0, 0, 3, 0, 0, 2, 4, 2, 0, 0, 21, 0, 
    0, 0, 5, 0, 0, 6, 0, 0, 11, 5, 0, 1, 34, 0, 0, 
    
    -- channel=13
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 14, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 14, 15, 20, 6, 0, 
    29, 0, 0, 0, 0, 0, 0, 4, 10, 0, 14, 9, 20, 14, 0, 
    38, 0, 0, 0, 0, 0, 16, 9, 18, 0, 11, 13, 5, 14, 1, 
    46, 15, 0, 0, 7, 3, 0, 13, 19, 0, 23, 32, 11, 16, 9, 
    38, 32, 3, 0, 0, 0, 17, 10, 29, 0, 40, 22, 14, 5, 5, 
    26, 38, 29, 0, 0, 0, 36, 23, 12, 0, 18, 31, 11, 2, 0, 
    35, 33, 39, 6, 0, 30, 22, 6, 8, 15, 10, 35, 6, 0, 0, 
    23, 28, 47, 18, 33, 1, 5, 8, 15, 9, 35, 24, 0, 0, 0, 
    20, 27, 55, 0, 14, 15, 0, 45, 47, 42, 38, 27, 51, 68, 71, 
    82, 43, 33, 0, 89, 99, 81, 82, 75, 65, 67, 71, 69, 73, 74, 
    89, 69, 24, 34, 108, 62, 64, 63, 65, 65, 70, 70, 75, 79, 75, 
    98, 81, 44, 85, 64, 65, 66, 64, 63, 67, 77, 85, 87, 75, 94, 
    90, 81, 72, 104, 74, 68, 70, 63, 55, 65, 75, 74, 57, 83, 100, 
    
    -- channel=14
    57, 62, 56, 63, 64, 57, 64, 70, 70, 63, 54, 46, 48, 60, 63, 
    60, 64, 57, 67, 50, 47, 84, 73, 59, 17, 33, 48, 41, 34, 58, 
    87, 11, 63, 68, 62, 69, 79, 56, 11, 0, 31, 10, 47, 21, 28, 
    107, 0, 67, 58, 88, 17, 45, 26, 16, 0, 59, 28, 39, 39, 0, 
    44, 0, 79, 0, 20, 18, 69, 53, 45, 0, 34, 59, 17, 40, 12, 
    32, 7, 82, 64, 0, 9, 64, 46, 79, 0, 68, 61, 2, 21, 22, 
    14, 70, 42, 103, 0, 0, 45, 39, 74, 0, 71, 53, 11, 0, 35, 
    19, 39, 28, 67, 0, 0, 74, 32, 44, 0, 45, 68, 0, 17, 30, 
    30, 0, 78, 0, 49, 14, 48, 44, 0, 74, 35, 65, 3, 0, 33, 
    14, 0, 89, 0, 55, 5, 0, 41, 39, 29, 53, 7, 0, 17, 64, 
    0, 11, 90, 0, 46, 17, 0, 15, 40, 33, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 129, 43, 9, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 68, 81, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 88, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 13, 0, 0, 3, 9, 15, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 15, 25, 17, 0, 7, 
    40, 0, 0, 0, 0, 0, 26, 1, 11, 0, 31, 0, 22, 0, 0, 
    69, 18, 0, 0, 85, 0, 23, 7, 4, 0, 24, 12, 14, 30, 0, 
    0, 32, 0, 0, 19, 0, 54, 21, 31, 0, 12, 15, 9, 24, 5, 
    0, 42, 0, 20, 0, 0, 55, 27, 47, 0, 36, 7, 0, 16, 7, 
    0, 77, 0, 41, 0, 24, 19, 5, 31, 0, 31, 7, 1, 0, 2, 
    19, 35, 0, 40, 0, 0, 13, 12, 13, 0, 0, 10, 0, 8, 0, 
    36, 18, 60, 8, 27, 0, 3, 71, 0, 13, 30, 15, 18, 0, 0, 
    51, 14, 51, 0, 109, 20, 13, 58, 53, 21, 15, 27, 6, 17, 21, 
    0, 42, 58, 9, 39, 17, 0, 2, 26, 26, 32, 27, 36, 26, 33, 
    27, 0, 0, 30, 39, 31, 31, 26, 28, 29, 35, 31, 34, 39, 43, 
    47, 27, 0, 113, 40, 25, 32, 23, 31, 30, 26, 34, 40, 27, 32, 
    43, 38, 5, 48, 17, 14, 33, 38, 35, 35, 30, 29, 40, 48, 61, 
    
    -- channel=16
    84, 93, 87, 90, 87, 89, 92, 98, 96, 88, 78, 74, 77, 79, 81, 
    83, 98, 92, 95, 88, 75, 91, 97, 90, 41, 28, 34, 44, 61, 76, 
    88, 64, 91, 96, 93, 102, 76, 51, 26, 10, 26, 12, 24, 28, 57, 
    57, 0, 83, 93, 95, 57, 52, 26, 14, 13, 42, 34, 26, 14, 28, 
    31, 7, 76, 58, 63, 47, 57, 33, 25, 0, 37, 38, 17, 18, 15, 
    25, 15, 74, 93, 54, 55, 55, 37, 32, 0, 53, 38, 15, 18, 8, 
    14, 39, 51, 105, 42, 31, 64, 37, 43, 0, 48, 28, 9, 10, 19, 
    25, 31, 13, 65, 34, 44, 55, 37, 35, 19, 42, 34, 10, 26, 30, 
    31, 21, 30, 12, 47, 40, 39, 34, 4, 55, 50, 40, 14, 18, 56, 
    34, 19, 40, 0, 42, 20, 10, 39, 20, 49, 37, 12, 0, 45, 78, 
    12, 29, 43, 0, 21, 15, 11, 36, 24, 11, 0, 0, 0, 0, 5, 
    0, 0, 16, 11, 85, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 63, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=17
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    0, 5, 0, 0, 0, 9, 0, 7, 4, 22, 16, 12, 0, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 10, 46, 6, 23, 14, 3, 15, 
    0, 0, 0, 0, 0, 0, 9, 4, 15, 36, 3, 0, 7, 0, 16, 
    38, 30, 0, 8, 75, 45, 0, 0, 0, 38, 18, 15, 21, 5, 0, 
    31, 23, 11, 0, 34, 17, 22, 7, 0, 51, 18, 6, 18, 13, 3, 
    32, 22, 4, 0, 10, 41, 34, 38, 12, 39, 21, 10, 26, 27, 0, 
    34, 49, 14, 23, 0, 57, 16, 2, 14, 6, 29, 24, 34, 8, 0, 
    44, 49, 6, 45, 12, 24, 24, 0, 20, 27, 20, 17, 11, 0, 0, 
    54, 42, 19, 44, 0, 0, 45, 54, 21, 11, 12, 15, 33, 38, 28, 
    102, 75, 28, 46, 64, 73, 74, 74, 53, 50, 50, 58, 58, 57, 56, 
    56, 93, 70, 50, 55, 50, 51, 51, 47, 48, 53, 52, 60, 66, 56, 
    61, 60, 109, 55, 43, 54, 45, 50, 55, 56, 64, 70, 65, 64, 83, 
    59, 65, 70, 73, 53, 66, 65, 53, 50, 50, 55, 60, 56, 53, 51, 
    
    -- channel=18
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 17, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 16, 0, 0, 24, 28, 0, 
    0, 78, 0, 0, 0, 48, 0, 0, 0, 44, 0, 0, 0, 32, 34, 
    0, 64, 0, 0, 0, 9, 0, 0, 0, 96, 0, 0, 0, 0, 94, 
    0, 10, 0, 51, 0, 0, 0, 0, 0, 91, 0, 0, 0, 0, 29, 
    0, 27, 0, 0, 148, 0, 0, 0, 0, 160, 0, 0, 19, 0, 0, 
    0, 0, 18, 0, 96, 29, 0, 0, 0, 147, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 27, 87, 0, 9, 0, 91, 0, 0, 30, 10, 0, 
    0, 0, 0, 51, 0, 43, 0, 0, 31, 0, 45, 0, 38, 29, 0, 
    0, 0, 0, 58, 0, 0, 28, 0, 0, 21, 0, 9, 45, 28, 0, 
    96, 0, 0, 124, 0, 0, 39, 9, 0, 0, 0, 0, 10, 37, 2, 
    135, 76, 0, 79, 0, 0, 34, 32, 3, 6, 9, 10, 3, 1, 0, 
    0, 108, 94, 0, 0, 0, 0, 0, 0, 0, 3, 0, 2, 10, 2, 
    0, 7, 158, 0, 0, 4, 0, 0, 8, 4, 2, 17, 0, 20, 1, 
    0, 7, 14, 50, 0, 37, 29, 3, 0, 0, 0, 5, 21, 0, 0, 
    
    -- channel=19
    1, 0, 0, 0, 0, 0, 0, 0, 0, 7, 18, 16, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 27, 6, 0, 0, 26, 19, 0, 
    20, 45, 0, 0, 0, 51, 19, 26, 0, 0, 0, 0, 0, 26, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 6, 0, 0, 34, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 13, 0, 0, 0, 0, 18, 
    0, 0, 0, 8, 93, 12, 0, 0, 0, 1, 0, 0, 2, 0, 0, 
    0, 0, 31, 0, 33, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 24, 0, 12, 0, 0, 8, 1, 0, 
    0, 0, 0, 5, 0, 52, 10, 0, 0, 0, 46, 22, 23, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 15, 12, 0, 0, 0, 
    26, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 22, 16, 
    76, 31, 0, 0, 25, 63, 51, 49, 19, 0, 0, 0, 0, 0, 0, 
    0, 57, 22, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 64, 31, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 10, 
    0, 0, 6, 57, 9, 21, 14, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=20
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 19, 2, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 5, 1, 4, 38, 0, 12, 0, 0, 0, 
    0, 31, 0, 4, 16, 5, 3, 0, 0, 21, 15, 0, 4, 0, 0, 
    26, 41, 0, 0, 58, 13, 6, 0, 0, 69, 14, 0, 14, 0, 0, 
    20, 36, 0, 0, 25, 37, 40, 0, 0, 67, 7, 2, 7, 19, 0, 
    36, 26, 8, 0, 16, 75, 0, 15, 0, 40, 11, 1, 21, 10, 0, 
    43, 56, 9, 30, 9, 10, 3, 18, 14, 0, 40, 0, 0, 0, 0, 
    46, 54, 10, 42, 27, 0, 13, 23, 18, 17, 0, 0, 9, 0, 0, 
    72, 50, 7, 86, 17, 43, 70, 48, 13, 0, 25, 36, 46, 43, 36, 
    98, 62, 27, 97, 58, 37, 50, 48, 46, 47, 54, 56, 59, 65, 63, 
    64, 86, 64, 83, 17, 49, 48, 46, 48, 55, 61, 68, 68, 68, 72, 
    67, 63, 109, 44, 42, 54, 46, 52, 54, 60, 65, 72, 62, 91, 74, 
    60, 68, 62, 54, 46, 62, 59, 48, 55, 57, 60, 59, 78, 78, 49, 
    
    -- channel=21
    1, 8, 1, 9, 10, 4, 3, 8, 17, 20, 13, 0, 3, 10, 19, 
    3, 5, 0, 12, 0, 3, 39, 25, 29, 0, 28, 23, 0, 0, 13, 
    45, 0, 4, 11, 0, 0, 57, 31, 0, 0, 26, 11, 43, 0, 0, 
    123, 0, 8, 1, 42, 0, 34, 26, 8, 0, 58, 6, 39, 26, 0, 
    88, 0, 41, 0, 28, 7, 62, 51, 32, 0, 24, 65, 5, 47, 0, 
    49, 0, 49, 11, 0, 0, 64, 45, 83, 0, 68, 69, 0, 27, 22, 
    39, 47, 0, 82, 0, 0, 30, 42, 84, 0, 82, 54, 0, 0, 25, 
    33, 45, 17, 49, 0, 0, 79, 9, 42, 0, 46, 64, 0, 0, 1, 
    48, 0, 100, 0, 31, 0, 30, 30, 0, 37, 0, 63, 0, 0, 0, 
    10, 0, 120, 0, 57, 0, 0, 44, 10, 14, 56, 4, 0, 0, 18, 
    0, 0, 108, 0, 108, 39, 0, 19, 69, 46, 4, 0, 0, 0, 28, 
    0, 0, 18, 0, 138, 61, 0, 3, 15, 0, 0, 0, 0, 0, 4, 
    11, 0, 0, 39, 132, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 0, 0, 105, 35, 0, 12, 0, 0, 0, 0, 0, 0, 0, 11, 
    30, 0, 0, 10, 13, 0, 0, 0, 0, 0, 10, 0, 0, 22, 48, 
    
    -- channel=22
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 0, 0, 12, 0, 0, 
    19, 25, 0, 0, 0, 0, 9, 6, 1, 0, 0, 0, 0, 9, 0, 
    4, 31, 0, 0, 29, 28, 0, 5, 0, 0, 3, 12, 6, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 25, 15, 0, 0, 0, 4, 30, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 4, 6, 5, 
    7, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 16, 0, 14, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 17, 14, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 22, 66, 68, 3, 0, 0, 20, 48, 61, 47, 17, 18, 
    0, 0, 0, 1, 0, 0, 0, 0, 9, 24, 30, 28, 34, 34, 31, 
    49, 0, 0, 0, 0, 28, 27, 26, 29, 37, 42, 48, 28, 21, 49, 
    38, 43, 0, 0, 1, 28, 37, 32, 26, 34, 31, 20, 29, 54, 5, 
    39, 37, 31, 0, 12, 8, 0, 20, 37, 45, 36, 31, 53, 55, 37, 
    
    -- channel=23
    0, 0, 5, 8, 9, 6, 4, 1, 9, 0, 0, 0, 2, 10, 7, 
    10, 10, 6, 7, 5, 58, 38, 11, 0, 1, 45, 28, 0, 0, 8, 
    0, 0, 5, 6, 1, 0, 0, 0, 13, 3, 13, 12, 30, 0, 0, 
    62, 27, 12, 7, 27, 3, 46, 23, 7, 0, 13, 0, 0, 11, 0, 
    52, 56, 35, 0, 104, 80, 24, 23, 0, 0, 34, 45, 12, 31, 0, 
    9, 0, 31, 0, 0, 0, 41, 30, 47, 0, 20, 0, 0, 17, 44, 
    28, 12, 0, 18, 0, 10, 0, 27, 22, 0, 8, 25, 3, 9, 26, 
    34, 16, 49, 37, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 
    29, 0, 43, 0, 40, 0, 0, 21, 0, 16, 0, 0, 0, 0, 24, 
    0, 0, 37, 0, 19, 6, 0, 54, 23, 0, 0, 0, 7, 15, 7, 
    0, 0, 16, 3, 142, 104, 8, 0, 11, 27, 33, 48, 27, 2, 9, 
    0, 0, 14, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 8, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 5, 12, 0, 0, 9, 23, 6, 
    
    -- channel=24
    5, 14, 7, 12, 7, 10, 10, 4, 6, 13, 14, 8, 11, 10, 7, 
    5, 8, 6, 14, 5, 42, 31, 21, 18, 14, 44, 24, 0, 1, 11, 
    31, 0, 5, 9, 0, 6, 41, 4, 9, 21, 79, 58, 58, 0, 7, 
    93, 0, 13, 3, 29, 0, 65, 51, 42, 0, 91, 41, 51, 32, 0, 
    121, 58, 45, 0, 122, 76, 97, 69, 45, 0, 76, 80, 39, 57, 0, 
    93, 87, 65, 8, 38, 71, 121, 71, 79, 0, 115, 76, 30, 53, 39, 
    93, 123, 28, 52, 0, 45, 116, 89, 94, 0, 114, 69, 27, 39, 58, 
    107, 125, 54, 54, 3, 69, 117, 57, 68, 6, 93, 70, 24, 44, 32, 
    132, 103, 120, 53, 52, 21, 54, 59, 27, 34, 34, 56, 2, 18, 20, 
    109, 99, 150, 25, 103, 27, 22, 111, 49, 56, 57, 15, 15, 14, 25, 
    67, 96, 133, 14, 202, 111, 77, 118, 116, 48, 33, 49, 46, 36, 47, 
    34, 77, 113, 72, 179, 82, 43, 44, 65, 54, 63, 62, 71, 74, 81, 
    90, 26, 34, 150, 127, 70, 71, 62, 62, 62, 66, 76, 83, 77, 83, 
    100, 70, 0, 172, 86, 64, 78, 67, 64, 70, 72, 77, 78, 76, 103, 
    108, 79, 62, 60, 58, 49, 65, 71, 71, 80, 84, 65, 69, 121, 112, 
    
    -- channel=25
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 11, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 0, 0, 16, 6, 0, 
    20, 26, 0, 0, 0, 48, 13, 23, 0, 0, 0, 0, 0, 17, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 7, 3, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 3, 49, 1, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    0, 4, 19, 0, 8, 0, 7, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 23, 25, 1, 0, 0, 3, 0, 5, 0, 
    0, 0, 0, 0, 0, 45, 6, 0, 0, 7, 34, 36, 10, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 31, 32, 7, 0, 0, 0, 
    0, 0, 7, 0, 0, 0, 0, 28, 3, 0, 0, 0, 0, 22, 25, 
    66, 15, 0, 0, 78, 64, 46, 45, 19, 6, 0, 1, 0, 0, 0, 
    0, 44, 0, 19, 55, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 27, 68, 3, 0, 0, 0, 0, 0, 0, 12, 2, 0, 37, 
    0, 0, 7, 70, 18, 18, 17, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=26
    48, 48, 49, 54, 53, 45, 52, 56, 55, 46, 32, 27, 35, 46, 50, 
    48, 50, 51, 56, 48, 48, 67, 47, 32, 10, 25, 23, 11, 20, 46, 
    46, 1, 53, 55, 53, 34, 42, 20, 12, 0, 35, 19, 34, 3, 17, 
    75, 0, 51, 48, 60, 20, 46, 34, 16, 0, 43, 19, 23, 18, 0, 
    56, 14, 67, 5, 57, 50, 51, 39, 22, 0, 37, 52, 17, 31, 0, 
    42, 7, 67, 50, 0, 18, 54, 44, 52, 0, 59, 40, 6, 23, 21, 
    38, 39, 16, 74, 0, 5, 41, 41, 52, 0, 53, 39, 8, 7, 35, 
    37, 35, 30, 48, 9, 2, 56, 15, 32, 0, 36, 41, 0, 15, 28, 
    42, 14, 62, 0, 46, 0, 26, 32, 0, 42, 13, 28, 0, 6, 40, 
    22, 18, 65, 0, 44, 14, 0, 48, 32, 18, 23, 0, 0, 18, 44, 
    0, 21, 59, 0, 83, 54, 0, 14, 32, 19, 0, 0, 0, 0, 4, 
    0, 0, 28, 0, 74, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 50, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 40, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 4, 
    
    -- channel=27
    12, 0, 6, 5, 5, 1, 8, 6, 2, 7, 15, 11, 7, 10, 3, 
    6, 0, 2, 4, 3, 0, 33, 3, 14, 0, 0, 9, 11, 11, 3, 
    0, 12, 8, 3, 3, 0, 23, 16, 23, 0, 1, 6, 3, 27, 0, 
    0, 0, 12, 0, 0, 4, 0, 27, 3, 0, 6, 8, 7, 24, 0, 
    43, 0, 48, 20, 0, 35, 4, 17, 0, 8, 0, 31, 0, 4, 30, 
    104, 0, 67, 27, 0, 64, 0, 7, 0, 0, 36, 48, 0, 6, 25, 
    123, 0, 57, 0, 0, 0, 0, 25, 0, 0, 37, 23, 1, 0, 20, 
    92, 0, 82, 0, 0, 0, 46, 6, 16, 0, 11, 16, 0, 0, 25, 
    44, 0, 87, 0, 52, 16, 9, 0, 8, 0, 0, 33, 0, 0, 0, 
    0, 0, 23, 0, 33, 65, 13, 0, 45, 16, 20, 11, 0, 0, 16, 
    0, 9, 16, 0, 5, 30, 0, 0, 50, 14, 0, 0, 2, 0, 17, 
    0, 0, 38, 0, 14, 60, 0, 3, 14, 1, 0, 0, 0, 0, 0, 
    12, 0, 40, 0, 83, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 3, 17, 0, 25, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 8, 0, 6, 0, 0, 4, 0, 0, 0, 0, 0, 0, 17, 
    
    -- channel=28
    34, 41, 34, 38, 35, 34, 40, 36, 31, 38, 39, 35, 34, 32, 28, 
    34, 32, 34, 42, 32, 54, 48, 43, 40, 21, 39, 27, 19, 29, 35, 
    52, 30, 35, 37, 30, 48, 51, 12, 6, 27, 71, 57, 56, 14, 35, 
    76, 0, 42, 31, 47, 16, 59, 44, 44, 22, 87, 43, 47, 30, 6, 
    99, 68, 66, 0, 113, 65, 89, 57, 46, 0, 68, 65, 39, 49, 0, 
    76, 102, 81, 12, 64, 70, 108, 63, 67, 0, 110, 70, 37, 48, 30, 
    67, 124, 54, 57, 24, 46, 123, 84, 83, 17, 106, 56, 28, 34, 55, 
    82, 117, 53, 66, 13, 86, 124, 69, 67, 29, 90, 60, 28, 55, 48, 
    110, 101, 93, 66, 43, 41, 54, 51, 39, 46, 39, 62, 12, 33, 37, 
    107, 98, 126, 31, 90, 30, 30, 97, 46, 68, 67, 14, 27, 38, 48, 
    82, 92, 118, 17, 161, 80, 81, 126, 110, 42, 16, 30, 39, 49, 50, 
    60, 92, 106, 86, 173, 74, 39, 38, 52, 43, 52, 49, 55, 59, 62, 
    73, 43, 46, 152, 109, 54, 56, 50, 48, 46, 50, 57, 70, 63, 64, 
    79, 55, 16, 184, 70, 51, 58, 50, 49, 54, 57, 64, 62, 54, 96, 
    85, 60, 51, 71, 49, 43, 60, 59, 54, 60, 63, 50, 49, 95, 88, 
    
    -- channel=29
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 15, 16, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 20, 3, 4, 10, 2, 0, 
    4, 1, 0, 0, 0, 0, 0, 0, 12, 12, 0, 0, 8, 2, 0, 
    22, 32, 0, 0, 33, 0, 0, 0, 0, 21, 5, 7, 15, 9, 0, 
    19, 24, 0, 0, 0, 0, 8, 0, 3, 29, 10, 5, 12, 12, 3, 
    17, 29, 0, 0, 0, 17, 19, 18, 6, 16, 10, 8, 20, 13, 0, 
    27, 40, 14, 19, 0, 15, 1, 1, 10, 0, 6, 14, 14, 0, 0, 
    37, 41, 21, 31, 8, 1, 9, 1, 7, 9, 12, 12, 8, 0, 0, 
    48, 28, 23, 43, 3, 1, 33, 47, 27, 14, 30, 36, 43, 36, 25, 
    102, 68, 28, 32, 42, 75, 73, 73, 73, 71, 82, 86, 93, 94, 92, 
    103, 94, 59, 36, 67, 79, 78, 79, 80, 85, 92, 95, 97, 99, 104, 
    113, 96, 90, 76, 69, 84, 78, 79, 84, 91, 100, 108, 105, 113, 116, 
    109, 108, 91, 94, 80, 92, 94, 86, 81, 88, 92, 99, 100, 107, 103, 
    
    -- channel=30
    35, 38, 30, 31, 30, 31, 34, 39, 29, 25, 22, 24, 17, 17, 17, 
    26, 32, 32, 33, 32, 18, 5, 23, 25, 5, 0, 0, 14, 23, 16, 
    23, 51, 35, 36, 39, 104, 24, 13, 0, 8, 0, 0, 0, 4, 26, 
    0, 0, 29, 35, 18, 14, 0, 0, 0, 38, 0, 6, 0, 0, 31, 
    0, 0, 3, 22, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 
    0, 40, 2, 34, 136, 30, 5, 0, 0, 22, 3, 0, 1, 0, 0, 
    0, 33, 30, 12, 66, 22, 45, 0, 0, 52, 6, 0, 0, 0, 0, 
    0, 17, 0, 0, 12, 59, 20, 37, 0, 61, 20, 0, 2, 12, 9, 
    0, 30, 0, 22, 0, 60, 22, 0, 0, 18, 53, 6, 10, 20, 12, 
    49, 37, 0, 23, 0, 0, 4, 0, 0, 24, 0, 0, 0, 11, 17, 
    67, 27, 1, 28, 0, 0, 0, 32, 0, 0, 0, 0, 0, 0, 0, 
    66, 50, 0, 61, 68, 32, 29, 23, 0, 0, 0, 0, 0, 0, 0, 
    0, 43, 30, 74, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 46, 74, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=31
    3, 0, 0, 1, 7, 0, 0, 4, 9, 1, 0, 0, 0, 3, 7, 
    8, 2, 0, 0, 1, 6, 13, 0, 0, 17, 26, 25, 12, 2, 3, 
    0, 0, 6, 5, 6, 0, 19, 35, 15, 0, 0, 0, 8, 6, 0, 
    24, 19, 13, 7, 8, 21, 4, 0, 0, 0, 0, 0, 5, 8, 0, 
    10, 0, 11, 0, 0, 0, 0, 0, 0, 8, 7, 5, 0, 4, 5, 
    2, 0, 5, 7, 0, 0, 0, 4, 12, 0, 0, 3, 0, 0, 12, 
    9, 0, 6, 5, 0, 0, 0, 0, 0, 0, 4, 13, 12, 3, 0, 
    0, 0, 20, 19, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 
    0, 0, 14, 0, 12, 0, 18, 9, 0, 41, 0, 0, 0, 0, 0, 
    0, 0, 2, 9, 0, 0, 5, 0, 0, 0, 0, 5, 0, 0, 4, 
    0, 0, 9, 0, 8, 0, 0, 0, 0, 24, 25, 4, 5, 22, 33, 
    0, 0, 0, 0, 0, 20, 19, 18, 8, 2, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 6, 0, 0, 0, 3, 2, 2, 0, 0, 0, 0, 
    1, 4, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 4, 0, 0, 
    0, 0, 8, 1, 7, 0, 0, 0, 0, 3, 0, 1, 0, 0, 4, 
    
    -- channel=32
    107, 107, 107, 107, 108, 108, 108, 108, 109, 107, 106, 107, 108, 107, 108, 
    108, 108, 108, 108, 108, 108, 108, 107, 105, 84, 101, 109, 107, 108, 108, 
    107, 108, 109, 108, 109, 107, 106, 94, 81, 68, 81, 107, 108, 109, 109, 
    101, 101, 107, 110, 108, 96, 114, 93, 88, 73, 72, 101, 104, 107, 109, 
    64, 83, 120, 108, 108, 96, 104, 102, 105, 100, 84, 79, 77, 106, 111, 
    71, 81, 85, 89, 105, 73, 87, 93, 100, 93, 87, 79, 58, 100, 106, 
    47, 60, 83, 98, 67, 17, 27, 60, 101, 98, 91, 82, 87, 75, 95, 
    25, 69, 47, 89, 95, 83, 89, 63, 65, 56, 44, 46, 52, 64, 77, 
    86, 64, 74, 78, 88, 87, 96, 76, 72, 61, 69, 55, 57, 57, 60, 
    42, 50, 50, 48, 50, 49, 37, 37, 37, 30, 26, 22, 25, 31, 46, 
    0, 11, 0, 3, 12, 18, 14, 9, 12, 3, 3, 8, 25, 37, 50, 
    0, 15, 6, 0, 0, 0, 26, 0, 0, 5, 23, 41, 35, 44, 62, 
    0, 0, 0, 0, 0, 0, 63, 80, 73, 57, 34, 36, 49, 55, 79, 
    0, 0, 0, 0, 0, 0, 14, 16, 0, 7, 31, 46, 53, 68, 84, 
    0, 0, 0, 0, 0, 0, 0, 0, 23, 48, 53, 54, 63, 73, 88, 
    
    -- channel=33
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 10, 11, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 1, 2, 0, 0, 0, 0, 0, 0, 
    35, 32, 0, 0, 0, 0, 0, 0, 0, 0, 13, 23, 17, 13, 0, 
    0, 0, 0, 8, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 
    12, 14, 0, 0, 0, 33, 38, 0, 0, 0, 0, 0, 5, 11, 11, 
    26, 7, 28, 17, 0, 0, 0, 4, 10, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 8, 
    22, 26, 27, 25, 22, 18, 21, 22, 10, 13, 22, 25, 14, 1, 17, 
    29, 18, 2, 12, 23, 23, 5, 7, 15, 5, 0, 0, 17, 21, 17, 
    28, 26, 21, 22, 25, 25, 17, 0, 0, 0, 29, 32, 18, 18, 12, 
    28, 36, 34, 31, 30, 30, 21, 1, 37, 41, 25, 20, 22, 19, 13, 
    
    -- channel=34
    43, 44, 44, 44, 44, 44, 45, 44, 45, 42, 42, 44, 44, 44, 45, 
    44, 44, 44, 44, 44, 43, 44, 44, 41, 24, 38, 45, 44, 44, 44, 
    45, 46, 45, 44, 45, 42, 45, 32, 26, 2, 38, 52, 43, 44, 45, 
    39, 39, 43, 46, 47, 28, 45, 18, 14, 3, 2, 40, 39, 41, 43, 
    2, 21, 38, 47, 46, 31, 48, 39, 40, 27, 27, 18, 16, 48, 40, 
    11, 24, 46, 42, 34, 42, 42, 45, 53, 19, 1, 7, 0, 39, 45, 
    0, 25, 21, 25, 15, 0, 0, 0, 29, 41, 38, 31, 34, 32, 44, 
    0, 0, 0, 40, 15, 0, 21, 23, 15, 0, 0, 0, 0, 0, 17, 
    22, 37, 17, 47, 51, 34, 35, 9, 14, 24, 15, 11, 15, 8, 0, 
    49, 7, 9, 6, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 12, 
    0, 0, 0, 0, 0, 0, 58, 44, 52, 43, 31, 7, 0, 14, 20, 
    0, 0, 0, 0, 0, 0, 7, 78, 78, 29, 5, 15, 5, 11, 25, 
    0, 0, 0, 0, 0, 0, 0, 15, 2, 16, 12, 0, 6, 12, 23, 
    
    -- channel=35
    7, 6, 6, 6, 6, 6, 6, 6, 6, 7, 5, 6, 7, 6, 6, 
    7, 7, 7, 7, 7, 7, 7, 8, 11, 23, 7, 5, 7, 7, 7, 
    7, 7, 7, 7, 6, 8, 6, 18, 20, 15, 0, 0, 8, 7, 7, 
    6, 7, 8, 7, 6, 20, 3, 13, 0, 0, 0, 0, 8, 8, 7, 
    29, 19, 1, 7, 8, 13, 2, 7, 0, 3, 10, 17, 23, 0, 6, 
    0, 0, 0, 17, 12, 26, 11, 7, 0, 9, 0, 0, 0, 0, 4, 
    19, 12, 14, 0, 14, 18, 0, 0, 0, 5, 9, 12, 7, 11, 2, 
    0, 0, 5, 2, 5, 0, 0, 6, 20, 22, 17, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 9, 12, 4, 0, 0, 0, 0, 0, 7, 10, 
    0, 3, 4, 3, 2, 3, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 3, 10, 7, 7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 2, 10, 13, 4, 1, 0, 0, 0, 0, 1, 12, 6, 0, 0, 
    25, 4, 3, 6, 3, 3, 0, 2, 27, 23, 7, 1, 8, 3, 0, 
    27, 7, 6, 5, 3, 3, 2, 20, 8, 0, 9, 12, 6, 1, 0, 
    
    -- channel=36
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=37
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 17, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 13, 44, 22, 27, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    95, 76, 3, 0, 0, 0, 0, 0, 0, 0, 44, 76, 85, 36, 0, 
    0, 0, 0, 35, 29, 97, 105, 85, 48, 0, 0, 0, 0, 0, 0, 
    110, 99, 42, 0, 0, 8, 0, 0, 0, 12, 56, 82, 64, 81, 50, 
    0, 0, 18, 14, 0, 0, 0, 12, 61, 30, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 23, 35, 14, 0, 21, 14, 41, 65, 80, 46, 
    59, 90, 89, 81, 70, 49, 36, 14, 20, 14, 33, 22, 2, 7, 3, 
    63, 52, 70, 92, 107, 114, 106, 100, 84, 72, 50, 29, 0, 0, 0, 
    10, 5, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 17, 35, 20, 3, 1, 53, 17, 0, 16, 65, 33, 0, 0, 0, 
    0, 0, 1, 2, 0, 0, 5, 15, 52, 12, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=38
    140, 139, 139, 139, 138, 139, 139, 139, 136, 140, 139, 139, 139, 139, 139, 
    139, 138, 138, 139, 137, 138, 137, 138, 139, 137, 104, 126, 138, 138, 139, 
    136, 136, 137, 139, 138, 140, 135, 141, 111, 109, 96, 112, 139, 138, 140, 
    139, 143, 141, 139, 140, 147, 112, 139, 128, 137, 131, 125, 143, 142, 142, 
    47, 44, 107, 133, 135, 143, 137, 142, 142, 146, 130, 99, 77, 68, 139, 
    148, 152, 145, 108, 114, 96, 81, 90, 102, 141, 136, 143, 147, 119, 137, 
    39, 24, 72, 106, 154, 81, 43, 64, 101, 135, 117, 96, 87, 96, 75, 
    0, 100, 65, 56, 101, 139, 151, 143, 81, 75, 77, 78, 86, 107, 116, 
    17, 145, 145, 149, 143, 139, 125, 128, 126, 119, 118, 116, 89, 72, 68, 
    77, 63, 66, 69, 73, 80, 93, 80, 80, 76, 66, 59, 60, 63, 64, 
    0, 0, 0, 0, 0, 0, 1, 11, 25, 21, 21, 28, 38, 61, 59, 
    0, 0, 31, 15, 0, 0, 24, 71, 44, 42, 49, 68, 65, 48, 62, 
    10, 0, 0, 0, 0, 0, 0, 30, 35, 31, 15, 0, 35, 61, 81, 
    46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 55, 58, 63, 86, 
    29, 0, 0, 0, 0, 0, 0, 0, 10, 39, 54, 54, 62, 76, 96, 
    
    -- channel=39
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=40
    49, 49, 49, 49, 50, 49, 50, 49, 50, 49, 51, 49, 49, 49, 50, 
    49, 50, 50, 50, 50, 50, 51, 49, 48, 34, 58, 57, 50, 50, 51, 
    49, 51, 51, 49, 51, 49, 51, 41, 40, 28, 51, 62, 50, 50, 51, 
    53, 50, 50, 50, 52, 36, 60, 31, 38, 31, 39, 66, 48, 49, 50, 
    52, 62, 64, 50, 52, 34, 52, 42, 51, 44, 36, 39, 44, 68, 51, 
    23, 36, 44, 45, 50, 31, 45, 47, 53, 35, 31, 29, 17, 67, 52, 
    48, 65, 54, 48, 17, 0, 34, 56, 73, 44, 40, 39, 40, 38, 63, 
    38, 39, 26, 67, 43, 22, 38, 26, 44, 42, 34, 35, 38, 37, 46, 
    99, 23, 29, 39, 49, 41, 46, 18, 29, 26, 32, 24, 32, 38, 38, 
    47, 47, 53, 55, 56, 52, 41, 44, 43, 33, 36, 25, 30, 28, 37, 
    15, 33, 28, 33, 35, 41, 44, 42, 35, 32, 30, 31, 37, 30, 34, 
    0, 11, 0, 0, 0, 2, 32, 8, 17, 22, 27, 28, 23, 29, 36, 
    0, 0, 5, 0, 0, 0, 70, 41, 39, 35, 33, 36, 28, 25, 38, 
    0, 0, 0, 0, 0, 0, 38, 60, 47, 33, 19, 17, 16, 29, 38, 
    0, 0, 0, 0, 0, 0, 9, 19, 9, 15, 13, 11, 18, 27, 39, 
    
    -- channel=41
    26, 26, 26, 26, 26, 26, 26, 26, 27, 25, 23, 26, 27, 26, 26, 
    26, 26, 26, 26, 25, 25, 25, 26, 25, 31, 15, 18, 26, 25, 25, 
    28, 28, 26, 26, 25, 27, 25, 28, 23, 14, 9, 20, 25, 26, 25, 
    12, 17, 22, 27, 27, 33, 16, 26, 0, 0, 0, 0, 20, 21, 23, 
    0, 0, 11, 29, 27, 33, 17, 27, 14, 15, 24, 21, 17, 11, 19, 
    0, 0, 22, 30, 27, 48, 42, 40, 33, 20, 0, 0, 0, 0, 20, 
    0, 0, 6, 4, 25, 0, 0, 0, 0, 30, 38, 37, 37, 36, 15, 
    0, 0, 0, 0, 9, 0, 0, 17, 11, 0, 0, 0, 0, 0, 0, 
    0, 34, 0, 17, 23, 28, 25, 28, 7, 16, 10, 15, 13, 8, 0, 
    7, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 71, 71, 66, 50, 19, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 79, 90, 33, 0, 1, 9, 0, 3, 
    4, 0, 0, 0, 0, 0, 0, 17, 0, 2, 18, 7, 4, 1, 1, 
    
    -- channel=42
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 6, 14, 13, 4, 12, 21, 7, 8, 7, 0, 0, 0, 0, 
    25, 5, 3, 17, 19, 15, 0, 0, 2, 0, 0, 6, 18, 0, 0, 
    31, 19, 18, 21, 19, 19, 19, 76, 72, 57, 47, 3, 0, 0, 0, 
    24, 28, 24, 22, 25, 24, 28, 49, 54, 14, 0, 0, 0, 0, 0, 
    
    -- channel=43
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=44
    6, 8, 8, 8, 9, 8, 8, 7, 10, 9, 7, 8, 9, 8, 9, 
    5, 8, 8, 8, 8, 8, 9, 7, 6, 0, 14, 17, 8, 8, 9, 
    5, 7, 9, 7, 10, 7, 8, 0, 0, 0, 25, 24, 6, 9, 9, 
    12, 6, 8, 8, 8, 0, 26, 0, 12, 7, 22, 58, 5, 8, 8, 
    0, 0, 32, 7, 8, 0, 32, 2, 20, 2, 0, 0, 0, 21, 13, 
    25, 45, 31, 0, 5, 0, 0, 0, 2, 0, 3, 19, 1, 84, 17, 
    0, 0, 0, 18, 0, 0, 17, 47, 77, 8, 0, 0, 0, 0, 11, 
    26, 73, 0, 57, 3, 11, 62, 3, 0, 0, 0, 6, 25, 28, 44, 
    156, 11, 25, 36, 24, 0, 3, 0, 10, 0, 0, 0, 0, 0, 0, 
    59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 16, 
    0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 16, 27, 
    0, 43, 0, 0, 2, 19, 68, 16, 16, 20, 36, 43, 21, 4, 39, 
    0, 25, 2, 0, 1, 14, 96, 0, 9, 6, 0, 0, 22, 37, 50, 
    0, 11, 13, 2, 10, 12, 44, 0, 0, 0, 27, 48, 23, 37, 43, 
    0, 14, 20, 14, 17, 19, 32, 0, 21, 61, 36, 17, 29, 37, 43, 
    
    -- channel=45
    31, 30, 30, 30, 30, 30, 30, 29, 28, 31, 33, 31, 30, 30, 30, 
    32, 31, 31, 31, 32, 32, 31, 32, 34, 51, 41, 31, 31, 32, 31, 
    32, 31, 31, 31, 30, 32, 34, 44, 63, 65, 37, 30, 32, 31, 31, 
    39, 38, 34, 30, 30, 38, 27, 44, 32, 40, 34, 26, 40, 36, 34, 
    86, 72, 30, 31, 32, 42, 23, 35, 27, 37, 51, 66, 70, 48, 36, 
    9, 0, 29, 41, 35, 62, 54, 49, 45, 51, 41, 24, 28, 0, 38, 
    80, 74, 54, 25, 45, 76, 54, 38, 9, 35, 44, 51, 44, 51, 48, 
    30, 0, 44, 20, 44, 12, 0, 36, 65, 72, 65, 48, 38, 30, 22, 
    0, 36, 8, 7, 28, 48, 50, 52, 29, 39, 38, 47, 51, 67, 67, 
    18, 75, 81, 85, 82, 84, 85, 75, 68, 65, 67, 68, 49, 40, 35, 
    55, 46, 58, 57, 56, 60, 73, 72, 69, 70, 61, 52, 41, 26, 18, 
    16, 2, 2, 7, 10, 4, 0, 25, 32, 23, 6, 0, 0, 19, 8, 
    14, 4, 15, 15, 9, 4, 0, 0, 0, 0, 0, 16, 0, 5, 11, 
    28, 5, 4, 6, 5, 5, 0, 0, 0, 0, 0, 0, 12, 13, 20, 
    39, 0, 2, 5, 2, 4, 0, 0, 0, 0, 0, 17, 13, 15, 20, 
    
    -- channel=46
    10, 8, 8, 8, 7, 8, 7, 10, 8, 10, 6, 8, 8, 8, 7, 
    10, 9, 9, 10, 8, 10, 8, 10, 18, 54, 0, 0, 10, 9, 8, 
    8, 7, 8, 10, 7, 15, 2, 39, 25, 29, 0, 0, 10, 8, 8, 
    0, 6, 6, 8, 9, 50, 0, 37, 0, 3, 0, 0, 6, 6, 6, 
    27, 0, 0, 5, 9, 24, 0, 11, 0, 16, 18, 19, 27, 0, 0, 
    0, 0, 6, 20, 14, 32, 0, 0, 0, 15, 2, 0, 21, 0, 0, 
    22, 0, 0, 0, 42, 77, 0, 0, 0, 12, 16, 18, 0, 13, 0, 
    0, 0, 20, 0, 0, 0, 0, 35, 27, 33, 37, 12, 0, 0, 0, 
    0, 0, 0, 0, 0, 17, 8, 7, 0, 0, 0, 0, 0, 1, 9, 
    0, 0, 0, 0, 0, 0, 15, 9, 3, 12, 4, 7, 0, 0, 0, 
    37, 1, 32, 18, 9, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    21, 0, 5, 26, 17, 0, 0, 21, 0, 0, 0, 0, 0, 1, 0, 
    56, 4, 19, 34, 17, 9, 0, 23, 22, 37, 40, 22, 4, 0, 0, 
    91, 13, 9, 16, 12, 11, 0, 68, 84, 29, 0, 0, 5, 0, 0, 
    75, 20, 14, 12, 11, 8, 0, 18, 0, 0, 12, 7, 0, 0, 0, 
    
    -- channel=47
    29, 29, 29, 29, 28, 29, 29, 29, 27, 28, 30, 30, 30, 29, 29, 
    28, 28, 28, 28, 28, 27, 27, 29, 24, 29, 27, 26, 27, 28, 28, 
    28, 28, 28, 28, 27, 28, 28, 24, 21, 44, 7, 33, 28, 27, 28, 
    28, 28, 28, 28, 28, 38, 19, 45, 42, 44, 29, 0, 32, 30, 30, 
    0, 0, 37, 27, 26, 56, 18, 44, 27, 31, 29, 16, 0, 14, 32, 
    63, 49, 23, 6, 21, 10, 24, 30, 41, 59, 47, 47, 54, 0, 30, 
    0, 0, 14, 43, 59, 2, 0, 0, 0, 28, 25, 20, 38, 21, 10, 
    22, 10, 0, 0, 45, 67, 39, 13, 2, 11, 5, 11, 6, 29, 0, 
    0, 78, 58, 42, 34, 38, 30, 75, 48, 45, 60, 44, 33, 13, 18, 
    3, 17, 8, 14, 12, 22, 33, 15, 18, 18, 14, 29, 19, 20, 17, 
    0, 0, 0, 0, 0, 0, 0, 2, 12, 11, 11, 11, 14, 10, 9, 
    12, 0, 42, 12, 0, 0, 57, 2, 4, 6, 11, 9, 16, 13, 9, 
    0, 0, 0, 0, 0, 0, 0, 30, 18, 6, 0, 0, 0, 8, 7, 
    32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 3, 15, 
    33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 10, 12, 11, 15, 
    
    -- channel=48
    37, 36, 36, 36, 36, 37, 36, 38, 37, 37, 34, 35, 37, 36, 36, 
    37, 36, 36, 37, 36, 37, 36, 36, 40, 51, 24, 30, 37, 36, 36, 
    38, 38, 36, 37, 37, 39, 33, 45, 36, 25, 15, 18, 36, 37, 36, 
    26, 29, 33, 38, 39, 51, 25, 37, 6, 2, 0, 2, 29, 31, 33, 
    22, 14, 16, 39, 38, 36, 27, 35, 25, 31, 32, 28, 33, 7, 27, 
    0, 0, 25, 46, 39, 55, 38, 35, 23, 22, 2, 0, 7, 0, 24, 
    22, 16, 21, 7, 33, 13, 0, 0, 0, 36, 43, 44, 35, 38, 17, 
    0, 0, 9, 16, 14, 0, 0, 31, 31, 23, 9, 0, 0, 0, 0, 
    0, 19, 3, 20, 26, 33, 32, 26, 5, 12, 5, 17, 14, 14, 11, 
    6, 19, 13, 13, 10, 5, 6, 0, 2, 0, 0, 0, 0, 0, 0, 
    7, 0, 10, 6, 10, 9, 6, 2, 2, 1, 0, 0, 0, 0, 0, 
    4, 0, 6, 4, 2, 0, 0, 0, 0, 0, 0, 0, 18, 14, 3, 
    15, 0, 22, 21, 4, 2, 12, 90, 89, 86, 75, 43, 22, 11, 3, 
    28, 2, 6, 7, 3, 2, 22, 160, 159, 79, 29, 20, 18, 8, 6, 
    19, 1, 0, 0, 0, 0, 2, 62, 31, 17, 28, 16, 11, 6, 5, 
    
    -- channel=49
    52, 52, 52, 52, 53, 53, 53, 52, 52, 52, 55, 52, 52, 52, 53, 
    53, 53, 53, 53, 54, 53, 54, 52, 52, 59, 74, 59, 53, 53, 54, 
    56, 56, 54, 52, 53, 52, 57, 55, 73, 58, 73, 75, 54, 54, 54, 
    55, 54, 54, 53, 55, 50, 63, 41, 36, 28, 26, 51, 54, 54, 54, 
    103, 104, 71, 57, 56, 41, 47, 46, 50, 53, 73, 87, 93, 94, 57, 
    11, 16, 49, 68, 68, 88, 104, 98, 89, 51, 24, 14, 9, 43, 58, 
    109, 121, 85, 48, 34, 29, 45, 34, 43, 60, 78, 88, 83, 87, 95, 
    65, 13, 46, 75, 50, 0, 6, 47, 82, 69, 45, 31, 29, 22, 40, 
    38, 33, 9, 31, 58, 64, 71, 49, 43, 60, 63, 67, 83, 92, 77, 
    91, 108, 111, 112, 108, 96, 83, 72, 75, 63, 75, 63, 55, 54, 57, 
    61, 71, 78, 93, 100, 109, 113, 112, 96, 89, 78, 69, 57, 35, 44, 
    10, 29, 4, 0, 7, 21, 16, 0, 11, 15, 11, 11, 42, 42, 32, 
    0, 18, 33, 18, 6, 7, 86, 53, 38, 42, 63, 55, 19, 26, 33, 
    0, 2, 7, 6, 3, 3, 26, 44, 54, 37, 0, 8, 22, 31, 43, 
    0, 0, 0, 0, 0, 0, 5, 23, 0, 0, 14, 20, 22, 28, 39, 
    
    -- channel=50
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 53, 60, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 14, 0, 0, 0, 
    68, 99, 80, 0, 0, 0, 0, 0, 0, 0, 0, 25, 46, 109, 0, 
    0, 0, 0, 3, 25, 22, 94, 83, 68, 0, 0, 0, 0, 23, 3, 
    80, 123, 72, 19, 0, 0, 8, 6, 26, 0, 13, 30, 58, 37, 88, 
    94, 0, 0, 83, 6, 0, 0, 0, 22, 1, 0, 0, 0, 0, 0, 
    141, 0, 0, 0, 4, 0, 27, 0, 0, 0, 21, 1, 44, 49, 32, 
    98, 68, 73, 69, 58, 44, 10, 5, 19, 0, 19, 4, 13, 17, 29, 
    21, 67, 35, 70, 92, 106, 97, 89, 67, 49, 43, 37, 27, 0, 17, 
    0, 70, 0, 0, 0, 19, 44, 0, 0, 0, 0, 0, 0, 5, 17, 
    0, 26, 46, 3, 0, 6, 197, 10, 0, 0, 19, 38, 0, 7, 23, 
    0, 1, 12, 2, 3, 6, 87, 45, 13, 23, 0, 0, 0, 18, 31, 
    0, 0, 0, 0, 0, 0, 26, 36, 0, 3, 0, 0, 8, 9, 19, 
    
    -- channel=51
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 29, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 29, 14, 22, 16, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    100, 98, 31, 0, 0, 0, 0, 0, 0, 0, 9, 49, 73, 64, 0, 
    0, 0, 0, 21, 25, 60, 85, 69, 39, 0, 0, 0, 0, 0, 0, 
    107, 117, 66, 0, 0, 0, 2, 0, 0, 0, 25, 50, 53, 46, 60, 
    29, 0, 0, 37, 0, 0, 0, 0, 50, 41, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 24, 0, 0, 0, 0, 0, 34, 57, 48, 
    23, 79, 81, 80, 70, 57, 33, 22, 26, 9, 27, 22, 5, 3, 3, 
    61, 70, 71, 94, 108, 114, 106, 97, 78, 67, 53, 32, 6, 0, 0, 
    2, 16, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 17, 46, 24, 6, 2, 76, 9, 0, 0, 40, 52, 0, 0, 0, 
    0, 0, 6, 6, 1, 1, 32, 49, 67, 45, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 30, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=52
    72, 73, 73, 73, 73, 73, 73, 71, 72, 75, 74, 73, 73, 73, 73, 
    72, 73, 73, 73, 73, 73, 73, 72, 75, 67, 76, 79, 73, 73, 74, 
    72, 73, 73, 73, 74, 74, 74, 73, 72, 60, 81, 78, 73, 74, 75, 
    83, 76, 76, 74, 73, 64, 79, 58, 64, 60, 60, 94, 79, 78, 76, 
    71, 80, 89, 72, 74, 62, 78, 71, 78, 81, 79, 71, 71, 85, 80, 
    57, 63, 73, 69, 76, 79, 79, 80, 77, 64, 63, 60, 40, 93, 83, 
    62, 68, 78, 64, 60, 7, 36, 51, 97, 83, 78, 68, 71, 63, 82, 
    26, 60, 28, 72, 63, 50, 70, 61, 57, 48, 41, 45, 50, 58, 79, 
    82, 64, 61, 71, 82, 77, 93, 66, 66, 74, 74, 69, 68, 61, 56, 
    76, 67, 76, 76, 73, 74, 63, 61, 67, 50, 57, 43, 49, 47, 45, 
    9, 20, 22, 23, 30, 41, 52, 49, 46, 37, 36, 33, 33, 38, 40, 
    0, 13, 0, 0, 0, 0, 9, 5, 11, 12, 16, 35, 28, 17, 40, 
    0, 0, 0, 0, 0, 0, 41, 0, 0, 0, 0, 0, 20, 32, 58, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 24, 44, 64, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 20, 24, 36, 47, 66, 
    
    -- channel=53
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 44, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 28, 15, 34, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 40, 0, 42, 0, 17, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 25, 0, 7, 0, 15, 14, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 18, 0, 0, 0, 20, 18, 8, 43, 0, 0, 
    0, 0, 0, 0, 47, 109, 0, 0, 0, 0, 3, 3, 0, 0, 0, 
    0, 0, 2, 0, 0, 25, 0, 26, 2, 19, 31, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 0, 36, 0, 0, 0, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 16, 6, 0, 22, 0, 14, 0, 0, 0, 
    10, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 0, 21, 33, 13, 0, 0, 42, 10, 0, 0, 0, 0, 0, 0, 
    59, 0, 0, 22, 10, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    117, 3, 0, 8, 3, 1, 0, 0, 29, 2, 0, 0, 0, 0, 0, 
    95, 16, 7, 6, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=54
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 25, 42, 13, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    47, 51, 0, 0, 0, 0, 0, 0, 0, 0, 18, 44, 51, 34, 0, 
    0, 0, 0, 0, 0, 17, 24, 55, 36, 0, 0, 0, 0, 0, 0, 
    0, 69, 0, 0, 0, 48, 67, 0, 0, 0, 2, 28, 37, 41, 27, 
    80, 0, 39, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 26, 0, 
    0, 0, 15, 33, 20, 14, 61, 129, 94, 88, 85, 69, 0, 0, 0, 
    37, 7, 0, 0, 10, 15, 0, 0, 0, 0, 0, 0, 3, 1, 0, 
    26, 18, 15, 12, 17, 17, 0, 0, 0, 0, 27, 21, 0, 0, 0, 
    0, 32, 30, 28, 29, 32, 32, 0, 36, 27, 0, 0, 0, 0, 0, 
    
    -- channel=55
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 25, 47, 60, 18, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 10, 1, 9, 0, 0, 0, 0, 0, 0, 
    83, 84, 13, 0, 0, 0, 0, 0, 0, 0, 41, 73, 87, 34, 0, 
    0, 0, 0, 0, 23, 29, 0, 31, 27, 0, 0, 0, 0, 0, 0, 
    0, 63, 0, 0, 0, 86, 102, 20, 0, 0, 0, 24, 35, 50, 32, 
    33, 24, 76, 51, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 
    0, 0, 22, 34, 9, 0, 38, 126, 73, 68, 70, 66, 2, 0, 5, 
    44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 10, 4, 
    52, 5, 0, 0, 2, 2, 0, 0, 0, 0, 46, 38, 0, 0, 0, 
    20, 32, 23, 19, 20, 21, 22, 12, 54, 42, 11, 0, 0, 1, 0, 
    
    -- channel=56
    138, 135, 135, 135, 135, 136, 135, 137, 134, 137, 136, 135, 135, 135, 135, 
    137, 135, 135, 135, 134, 135, 134, 134, 136, 147, 99, 120, 135, 134, 134, 
    135, 134, 134, 136, 134, 139, 130, 145, 118, 126, 86, 99, 136, 134, 136, 
    128, 134, 133, 136, 137, 154, 105, 150, 127, 134, 116, 90, 137, 135, 136, 
    56, 50, 99, 130, 133, 148, 118, 142, 134, 152, 143, 112, 92, 62, 131, 
    141, 133, 123, 113, 119, 122, 99, 105, 104, 144, 135, 135, 144, 81, 127, 
    58, 30, 84, 104, 153, 107, 28, 31, 71, 140, 136, 120, 112, 108, 76, 
    0, 79, 64, 39, 108, 148, 130, 138, 86, 81, 79, 71, 67, 91, 96, 
    0, 139, 136, 126, 129, 140, 129, 157, 128, 130, 130, 133, 104, 82, 82, 
    54, 86, 82, 87, 87, 93, 103, 87, 87, 94, 77, 81, 69, 70, 63, 
    2, 0, 17, 9, 6, 11, 39, 45, 56, 53, 46, 42, 42, 67, 58, 
    20, 0, 55, 36, 4, 0, 8, 66, 41, 41, 46, 75, 78, 58, 52, 
    25, 0, 0, 3, 0, 0, 0, 102, 100, 91, 54, 20, 40, 48, 61, 
    79, 0, 0, 0, 0, 0, 0, 20, 13, 0, 13, 36, 52, 51, 69, 
    63, 0, 0, 0, 0, 0, 0, 0, 3, 19, 51, 50, 54, 63, 77, 
    
    -- channel=57
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 14, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 35, 23, 16, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    91, 76, 5, 0, 0, 0, 0, 0, 0, 0, 26, 58, 74, 34, 0, 
    0, 0, 0, 25, 19, 79, 83, 66, 32, 0, 0, 0, 0, 0, 0, 
    99, 92, 48, 0, 0, 0, 0, 0, 0, 3, 37, 60, 51, 56, 40, 
    0, 0, 4, 11, 0, 0, 0, 0, 48, 32, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 12, 26, 7, 0, 3, 0, 22, 44, 62, 43, 
    28, 79, 78, 77, 66, 52, 39, 20, 25, 12, 32, 25, 2, 3, 0, 
    59, 46, 66, 83, 94, 97, 93, 88, 73, 63, 45, 24, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 34, 21, 2, 0, 28, 4, 0, 0, 35, 27, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 13, 38, 10, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=58
    32, 30, 30, 30, 30, 30, 29, 30, 31, 31, 27, 30, 30, 30, 29, 
    31, 30, 30, 30, 29, 30, 29, 30, 33, 41, 0, 15, 30, 29, 29, 
    28, 28, 29, 31, 29, 33, 25, 41, 20, 22, 0, 0, 31, 30, 29, 
    20, 28, 28, 30, 29, 47, 8, 47, 28, 36, 27, 10, 28, 29, 29, 
    0, 0, 0, 26, 29, 39, 25, 33, 28, 38, 29, 11, 2, 0, 22, 
    34, 27, 27, 22, 17, 23, 0, 0, 0, 31, 37, 38, 50, 3, 20, 
    0, 0, 0, 1, 48, 52, 0, 0, 1, 29, 21, 12, 0, 7, 0, 
    0, 14, 14, 0, 12, 46, 34, 48, 3, 4, 15, 11, 10, 16, 21, 
    0, 27, 26, 24, 16, 26, 16, 28, 19, 16, 3, 16, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    7, 0, 14, 20, 4, 0, 0, 37, 9, 4, 2, 16, 7, 1, 2, 
    37, 0, 0, 1, 0, 0, 0, 8, 16, 18, 0, 0, 9, 9, 5, 
    61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 17, 17, 8, 5, 
    49, 17, 10, 6, 4, 4, 0, 0, 16, 12, 24, 17, 14, 13, 10, 
    
    -- channel=59
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 11, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 13, 0, 0, 0, 0, 0, 0, 0, 1, 10, 13, 14, 0, 0, 
    0, 0, 0, 21, 0, 42, 16, 14, 5, 0, 0, 0, 0, 0, 0, 
    16, 13, 0, 1, 0, 79, 0, 0, 0, 0, 15, 26, 9, 0, 7, 
    1, 0, 23, 0, 0, 4, 0, 0, 5, 6, 10, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 26, 3, 14, 0, 10, 10, 8, 6, 
    0, 15, 2, 10, 7, 2, 0, 4, 0, 24, 0, 9, 0, 4, 0, 
    22, 0, 10, 12, 10, 10, 8, 17, 10, 17, 12, 6, 0, 0, 0, 
    23, 0, 1, 8, 11, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 9, 0, 11, 12, 3, 0, 12, 6, 9, 17, 6, 2, 0, 0, 
    34, 4, 3, 7, 4, 2, 42, 10, 40, 15, 0, 0, 0, 0, 0, 
    41, 4, 0, 1, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=60
    135, 134, 134, 134, 133, 134, 134, 135, 132, 135, 135, 135, 134, 134, 134, 
    135, 133, 133, 134, 133, 133, 132, 133, 133, 146, 109, 120, 133, 132, 133, 
    135, 133, 133, 134, 132, 136, 131, 142, 124, 126, 99, 114, 135, 134, 134, 
    125, 132, 134, 134, 134, 151, 111, 141, 114, 115, 96, 87, 138, 135, 136, 
    73, 72, 114, 131, 132, 146, 117, 138, 128, 143, 149, 129, 110, 87, 135, 
    122, 116, 128, 118, 129, 139, 132, 134, 127, 143, 118, 113, 117, 73, 132, 
    75, 52, 95, 104, 147, 80, 18, 13, 54, 143, 146, 137, 130, 128, 95, 
    3, 60, 66, 50, 107, 115, 106, 134, 95, 77, 62, 52, 51, 71, 84, 
    0, 141, 118, 120, 131, 146, 139, 157, 126, 132, 134, 137, 118, 101, 88, 
    74, 96, 90, 91, 88, 91, 95, 72, 76, 75, 70, 70, 58, 64, 62, 
    0, 0, 8, 11, 15, 21, 42, 50, 57, 48, 40, 34, 31, 50, 55, 
    16, 0, 45, 21, 0, 0, 0, 14, 1, 3, 11, 41, 69, 57, 50, 
    12, 0, 0, 0, 0, 0, 0, 85, 75, 71, 52, 22, 28, 50, 65, 
    60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 57, 56, 79, 
    57, 0, 0, 0, 0, 0, 0, 0, 0, 17, 54, 59, 60, 69, 84, 
    
    -- channel=61
    38, 38, 38, 38, 39, 39, 39, 38, 38, 39, 42, 39, 38, 38, 39, 
    39, 39, 39, 39, 39, 39, 39, 38, 37, 43, 56, 44, 38, 39, 39, 
    40, 39, 39, 39, 38, 39, 42, 41, 56, 60, 57, 56, 39, 39, 40, 
    45, 43, 41, 38, 38, 37, 47, 42, 46, 45, 41, 46, 46, 43, 42, 
    77, 78, 63, 39, 39, 40, 35, 39, 42, 51, 63, 71, 70, 73, 49, 
    38, 33, 41, 40, 52, 58, 76, 73, 68, 55, 47, 36, 28, 39, 50, 
    81, 78, 67, 48, 40, 35, 48, 42, 41, 51, 60, 64, 67, 63, 69, 
    58, 36, 40, 45, 55, 31, 29, 39, 57, 52, 42, 37, 35, 37, 42, 
    38, 46, 28, 28, 46, 54, 64, 62, 57, 64, 73, 69, 75, 77, 70, 
    63, 85, 90, 90, 87, 84, 78, 71, 71, 65, 73, 70, 63, 57, 54, 
    44, 56, 57, 68, 73, 81, 92, 90, 85, 77, 73, 65, 60, 45, 40, 
    16, 28, 17, 8, 9, 17, 35, 18, 33, 34, 29, 27, 27, 30, 25, 
    0, 8, 11, 4, 6, 4, 32, 0, 0, 0, 0, 9, 4, 16, 32, 
    0, 1, 0, 1, 2, 3, 0, 0, 0, 0, 0, 0, 15, 26, 41, 
    6, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 18, 22, 29, 40, 
    
    -- channel=62
    56, 58, 58, 58, 58, 58, 58, 58, 58, 57, 58, 57, 58, 58, 58, 
    59, 59, 59, 59, 60, 59, 60, 60, 59, 65, 88, 69, 58, 59, 60, 
    62, 62, 61, 60, 59, 59, 61, 61, 75, 50, 60, 79, 60, 61, 61, 
    55, 53, 62, 61, 60, 62, 75, 44, 13, 0, 0, 40, 59, 60, 62, 
    115, 117, 98, 66, 63, 53, 48, 50, 41, 42, 61, 88, 102, 105, 68, 
    0, 0, 43, 71, 82, 86, 107, 100, 89, 55, 8, 0, 0, 17, 64, 
    98, 115, 90, 32, 29, 0, 6, 8, 24, 60, 73, 83, 84, 85, 95, 
    4, 0, 22, 81, 61, 0, 0, 20, 83, 64, 24, 2, 0, 0, 3, 
    0, 15, 0, 0, 34, 59, 77, 26, 0, 10, 20, 23, 48, 74, 65, 
    40, 77, 82, 79, 74, 63, 45, 27, 33, 3, 25, 11, 0, 0, 15, 
    20, 35, 31, 47, 63, 70, 62, 49, 40, 25, 11, 1, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 7, 
    0, 0, 0, 0, 0, 0, 69, 30, 0, 0, 28, 39, 0, 1, 21, 
    0, 0, 0, 0, 0, 0, 0, 12, 1, 0, 0, 0, 9, 18, 39, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 13, 18, 35, 
    
    -- channel=63
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 19, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 8, 0, 0, 
    0, 0, 0, 0, 0, 47, 55, 72, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 0, 0, 0, 0, 0, 0, 30, 51, 44, 37, 21, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 
    21, 14, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 1, 0, 15, 62, 51, 39, 22, 0, 0, 0, 0, 
    19, 7, 0, 0, 5, 4, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    20, 7, 5, 6, 6, 6, 0, 0, 0, 6, 17, 0, 0, 0, 0, 
    23, 21, 19, 19, 17, 19, 24, 23, 18, 0, 0, 0, 0, 0, 0, 
    
    -- channel=64
    61, 70, 89, 89, 98, 98, 106, 102, 107, 112, 105, 115, 107, 110, 110, 
    69, 78, 98, 96, 105, 100, 105, 107, 107, 82, 104, 115, 108, 111, 115, 
    75, 78, 102, 101, 107, 101, 94, 92, 107, 55, 98, 107, 106, 111, 116, 
    73, 82, 94, 103, 100, 104, 89, 79, 43, 31, 30, 47, 98, 97, 104, 
    43, 39, 42, 53, 60, 64, 62, 45, 36, 24, 25, 47, 52, 63, 57, 
    25, 30, 24, 29, 34, 32, 37, 24, 27, 30, 55, 72, 48, 70, 22, 
    22, 24, 18, 33, 46, 41, 37, 32, 37, 44, 73, 84, 64, 49, 26, 
    27, 33, 39, 43, 51, 57, 60, 57, 61, 43, 64, 77, 70, 26, 43, 
    33, 26, 54, 60, 53, 52, 56, 56, 61, 49, 59, 63, 63, 61, 55, 
    19, 39, 40, 42, 54, 56, 59, 54, 56, 65, 64, 58, 45, 33, 33, 
    45, 38, 43, 35, 43, 59, 38, 19, 48, 54, 43, 33, 24, 16, 8, 
    42, 42, 24, 18, 23, 48, 34, 25, 28, 30, 21, 14, 10, 4, 0, 
    33, 32, 25, 21, 21, 23, 22, 20, 16, 15, 14, 13, 0, 0, 0, 
    6, 8, 7, 11, 11, 10, 11, 9, 22, 0, 4, 0, 0, 0, 1, 
    0, 0, 1, 3, 6, 6, 6, 2, 24, 0, 0, 0, 0, 0, 0, 
    
    -- channel=65
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 1, 4, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 0, 0, 0, 3, 1, 2, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 21, 19, 0, 0, 
    6, 21, 7, 8, 9, 9, 0, 0, 3, 8, 27, 32, 16, 9, 19, 
    0, 2, 0, 0, 0, 0, 0, 6, 12, 13, 17, 0, 6, 4, 5, 
    6, 10, 19, 12, 1, 0, 0, 0, 0, 0, 0, 1, 3, 16, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 12, 20, 5, 1, 9, 0, 
    0, 9, 0, 0, 0, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 3, 8, 8, 
    0, 0, 0, 0, 0, 0, 0, 7, 2, 0, 5, 2, 7, 10, 11, 
    0, 0, 0, 0, 0, 0, 0, 9, 5, 0, 11, 12, 8, 12, 16, 
    0, 0, 5, 10, 11, 8, 3, 7, 20, 14, 9, 12, 13, 16, 16, 
    15, 17, 16, 16, 18, 20, 15, 12, 13, 11, 12, 12, 15, 16, 14, 
    
    -- channel=66
    0, 10, 19, 23, 26, 31, 39, 31, 44, 43, 46, 47, 40, 42, 49, 
    0, 17, 32, 26, 34, 33, 38, 40, 46, 19, 40, 55, 41, 45, 49, 
    5, 24, 40, 30, 41, 34, 27, 44, 45, 0, 43, 58, 33, 44, 54, 
    16, 20, 43, 47, 49, 44, 35, 15, 2, 0, 0, 0, 46, 45, 59, 
    0, 0, 0, 21, 19, 29, 19, 0, 0, 0, 0, 0, 26, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 33, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 32, 8, 27, 0, 
    0, 0, 0, 1, 2, 0, 0, 0, 1, 0, 11, 26, 20, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 17, 9, 0, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 3, 9, 4, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=67
    0, 0, 0, 0, 0, 0, 0, 6, 0, 2, 5, 3, 4, 5, 0, 
    1, 0, 0, 0, 1, 4, 7, 6, 3, 27, 1, 3, 8, 9, 1, 
    6, 0, 0, 6, 11, 8, 17, 13, 5, 37, 0, 1, 13, 14, 4, 
    9, 0, 3, 3, 15, 8, 17, 14, 28, 32, 14, 31, 13, 15, 9, 
    19, 14, 25, 23, 26, 24, 19, 24, 0, 0, 0, 0, 0, 23, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 13, 17, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 6, 20, 16, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 4, 9, 10, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 5, 6, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 14, 21, 13, 
    0, 0, 0, 0, 0, 0, 12, 13, 0, 6, 12, 18, 13, 8, 9, 
    0, 0, 4, 0, 0, 0, 4, 0, 0, 8, 11, 6, 8, 3, 6, 
    0, 0, 0, 0, 0, 9, 4, 0, 3, 5, 4, 0, 6, 0, 0, 
    4, 4, 2, 0, 0, 2, 3, 6, 0, 3, 0, 1, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 3, 0, 9, 0, 0, 0, 0, 11, 
    
    -- channel=68
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=69
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 32, 15, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 4, 32, 18, 42, 9, 28, 12, 6, 0, 
    21, 5, 24, 20, 16, 4, 5, 2, 77, 52, 42, 91, 55, 41, 43, 
    70, 58, 61, 71, 74, 74, 60, 50, 10, 4, 8, 0, 0, 12, 47, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 6, 
    0, 4, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 39, 46, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 37, 32, 3, 0, 0, 0, 
    12, 46, 13, 0, 14, 32, 24, 0, 0, 0, 0, 0, 0, 0, 34, 
    0, 0, 0, 18, 0, 0, 0, 27, 35, 0, 0, 12, 48, 55, 41, 
    0, 0, 2, 25, 49, 24, 21, 26, 0, 29, 56, 48, 29, 20, 26, 
    4, 7, 15, 6, 0, 0, 36, 17, 16, 16, 28, 28, 4, 14, 7, 
    24, 50, 51, 37, 45, 38, 9, 6, 34, 29, 5, 10, 17, 3, 0, 
    36, 30, 19, 11, 17, 25, 21, 12, 0, 3, 10, 6, 2, 0, 0, 
    2, 0, 0, 0, 0, 0, 3, 15, 10, 12, 4, 0, 0, 0, 18, 
    
    -- channel=70
    138, 99, 133, 137, 142, 134, 141, 149, 136, 145, 134, 139, 143, 150, 136, 
    132, 93, 122, 131, 135, 128, 132, 136, 132, 147, 77, 134, 140, 145, 131, 
    126, 82, 111, 124, 130, 122, 133, 98, 100, 136, 58, 109, 133, 126, 122, 
    109, 71, 100, 96, 110, 105, 113, 121, 80, 41, 38, 10, 31, 101, 77, 
    34, 32, 38, 36, 43, 47, 53, 80, 66, 70, 54, 53, 66, 89, 37, 
    47, 52, 79, 45, 85, 78, 90, 80, 67, 71, 60, 116, 123, 72, 65, 
    65, 55, 47, 51, 71, 94, 98, 98, 104, 101, 90, 94, 101, 64, 40, 
    86, 96, 106, 122, 122, 124, 124, 118, 100, 97, 47, 70, 88, 87, 76, 
    82, 67, 60, 99, 111, 100, 90, 89, 88, 108, 96, 96, 89, 86, 70, 
    75, 88, 107, 95, 84, 103, 109, 97, 67, 92, 95, 95, 70, 47, 25, 
    78, 96, 95, 86, 68, 70, 101, 45, 28, 72, 64, 48, 40, 28, 30, 
    55, 77, 90, 47, 55, 67, 75, 58, 47, 44, 41, 31, 27, 18, 8, 
    44, 56, 49, 42, 32, 22, 30, 40, 34, 25, 24, 20, 21, 8, 11, 
    2, 0, 7, 12, 21, 19, 17, 19, 18, 47, 14, 12, 9, 10, 13, 
    6, 4, 9, 12, 17, 23, 23, 18, 0, 30, 11, 5, 8, 9, 10, 
    
    -- channel=71
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=72
    31, 55, 57, 54, 56, 55, 54, 43, 56, 55, 49, 54, 50, 50, 57, 
    31, 53, 57, 48, 50, 49, 51, 48, 54, 30, 68, 60, 50, 50, 61, 
    28, 50, 54, 42, 43, 43, 35, 48, 57, 0, 73, 58, 43, 46, 58, 
    26, 51, 48, 51, 39, 45, 29, 25, 25, 21, 41, 53, 64, 39, 51, 
    32, 35, 34, 44, 39, 43, 42, 18, 17, 13, 20, 26, 32, 21, 41, 
    23, 21, 4, 26, 23, 23, 27, 16, 18, 13, 37, 30, 2, 22, 0, 
    24, 21, 16, 40, 43, 30, 32, 26, 25, 23, 47, 42, 9, 24, 0, 
    26, 24, 28, 37, 40, 40, 37, 33, 36, 15, 43, 42, 32, 0, 12, 
    33, 31, 57, 51, 42, 38, 36, 30, 36, 10, 33, 32, 31, 24, 22, 
    28, 39, 35, 38, 41, 34, 30, 25, 32, 33, 36, 26, 18, 12, 21, 
    41, 35, 35, 24, 35, 42, 15, 16, 45, 29, 22, 14, 5, 1, 0, 
    45, 35, 15, 23, 26, 42, 9, 9, 20, 16, 4, 2, 1, 0, 0, 
    32, 22, 11, 15, 18, 21, 14, 9, 5, 7, 0, 7, 0, 0, 0, 
    12, 12, 5, 7, 3, 3, 7, 2, 11, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 
    
    -- channel=73
    0, 0, 0, 0, 0, 4, 15, 23, 16, 20, 28, 24, 20, 24, 19, 
    0, 0, 0, 7, 16, 15, 23, 28, 20, 32, 2, 25, 24, 31, 19, 
    11, 0, 10, 19, 30, 23, 31, 30, 20, 40, 0, 29, 29, 36, 26, 
    29, 0, 31, 38, 51, 36, 45, 23, 14, 0, 0, 0, 19, 47, 43, 
    9, 0, 4, 11, 24, 27, 18, 22, 0, 0, 0, 0, 1, 15, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 40, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 41, 27, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 14, 18, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 5, 4, 34, 
    0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 10, 15, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=74
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 37, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=75
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=76
    0, 20, 22, 6, 9, 5, 11, 0, 20, 11, 0, 15, 2, 10, 12, 
    0, 19, 25, 2, 14, 3, 10, 8, 15, 0, 15, 21, 0, 7, 15, 
    0, 14, 27, 2, 17, 5, 0, 5, 14, 0, 60, 15, 0, 8, 20, 
    0, 13, 16, 8, 3, 13, 0, 4, 0, 0, 10, 0, 26, 3, 9, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 2, 15, 39, 0, 8, 
    24, 20, 0, 15, 23, 12, 13, 0, 1, 4, 42, 49, 0, 28, 0, 
    19, 0, 0, 34, 16, 0, 7, 3, 20, 20, 53, 17, 0, 3, 0, 
    8, 12, 26, 35, 18, 12, 5, 0, 0, 0, 13, 17, 1, 0, 32, 
    0, 0, 17, 10, 0, 0, 0, 0, 15, 0, 42, 16, 0, 0, 0, 
    0, 34, 18, 0, 0, 12, 11, 0, 0, 6, 8, 0, 0, 0, 0, 
    13, 2, 1, 0, 2, 8, 0, 0, 33, 11, 0, 0, 0, 0, 0, 
    43, 1, 0, 0, 8, 40, 0, 0, 10, 0, 0, 0, 0, 1, 0, 
    24, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 13, 0, 3, 3, 
    0, 0, 1, 10, 7, 5, 4, 0, 24, 0, 0, 4, 0, 10, 10, 
    5, 14, 14, 16, 15, 15, 12, 0, 41, 0, 8, 3, 8, 11, 0, 
    
    -- channel=77
    62, 45, 46, 50, 43, 41, 36, 39, 32, 34, 38, 31, 37, 34, 32, 
    58, 38, 38, 40, 34, 35, 33, 35, 33, 55, 40, 27, 35, 33, 28, 
    48, 34, 27, 31, 25, 31, 33, 40, 33, 70, 18, 32, 35, 28, 23, 
    38, 18, 14, 15, 18, 16, 33, 23, 66, 91, 61, 72, 36, 25, 19, 
    54, 43, 56, 44, 46, 42, 52, 66, 50, 43, 42, 18, 7, 27, 34, 
    34, 27, 35, 35, 31, 40, 42, 60, 43, 39, 15, 0, 13, 11, 38, 
    40, 41, 54, 35, 52, 52, 54, 51, 41, 37, 8, 22, 37, 25, 38, 
    45, 34, 22, 25, 41, 48, 52, 50, 49, 54, 35, 22, 26, 41, 0, 
    55, 64, 55, 54, 62, 67, 70, 61, 39, 37, 8, 24, 34, 24, 32, 
    67, 31, 43, 62, 61, 47, 40, 46, 48, 41, 35, 37, 44, 52, 41, 
    53, 60, 56, 57, 53, 54, 64, 70, 35, 40, 53, 61, 45, 42, 29, 
    42, 59, 70, 65, 50, 33, 56, 37, 37, 48, 46, 49, 39, 32, 33, 
    39, 51, 60, 44, 49, 57, 44, 33, 41, 46, 37, 29, 38, 28, 26, 
    40, 43, 38, 31, 31, 35, 41, 40, 24, 34, 33, 27, 29, 24, 19, 
    22, 20, 26, 26, 27, 25, 29, 31, 17, 48, 24, 25, 24, 22, 28, 
    
    -- channel=78
    7, 0, 0, 0, 0, 0, 0, 18, 0, 2, 4, 0, 8, 9, 0, 
    20, 0, 0, 2, 0, 7, 13, 5, 0, 68, 0, 0, 15, 14, 0, 
    25, 0, 0, 10, 13, 12, 38, 7, 0, 106, 0, 0, 25, 15, 0, 
    29, 0, 6, 1, 26, 9, 31, 36, 54, 57, 14, 36, 0, 15, 0, 
    21, 7, 31, 13, 28, 18, 13, 41, 4, 1, 0, 0, 0, 65, 28, 
    0, 0, 14, 0, 0, 0, 0, 5, 0, 0, 0, 0, 76, 0, 49, 
    0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 7, 47, 39, 59, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 0, 0, 17, 58, 17, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 17, 0, 7, 11, 19, 18, 
    2, 0, 0, 0, 0, 0, 0, 8, 0, 0, 1, 27, 26, 43, 16, 
    0, 0, 0, 0, 0, 0, 41, 35, 0, 0, 18, 35, 23, 12, 22, 
    0, 0, 31, 5, 0, 0, 19, 0, 0, 14, 16, 8, 22, 11, 21, 
    0, 0, 5, 0, 1, 11, 5, 0, 3, 9, 12, 0, 22, 4, 3, 
    12, 7, 2, 0, 0, 0, 2, 13, 0, 26, 5, 8, 6, 0, 6, 
    7, 0, 0, 0, 0, 0, 0, 15, 0, 38, 3, 7, 1, 0, 39, 
    
    -- channel=79
    57, 4, 39, 31, 37, 23, 32, 47, 26, 31, 27, 32, 26, 38, 23, 
    46, 0, 27, 24, 36, 18, 28, 46, 24, 33, 0, 27, 22, 38, 12, 
    45, 0, 17, 24, 31, 23, 37, 12, 6, 61, 0, 22, 25, 33, 15, 
    40, 0, 11, 20, 29, 20, 42, 29, 0, 20, 0, 0, 12, 29, 0, 
    5, 0, 0, 0, 0, 0, 0, 39, 34, 31, 22, 13, 0, 14, 0, 
    19, 5, 36, 9, 35, 10, 29, 36, 25, 35, 7, 49, 10, 73, 4, 
    19, 4, 17, 2, 13, 36, 33, 38, 31, 31, 0, 3, 66, 0, 10, 
    33, 39, 56, 38, 43, 41, 43, 28, 37, 26, 0, 9, 17, 39, 30, 
    19, 26, 0, 33, 29, 31, 26, 32, 14, 60, 14, 11, 17, 16, 21, 
    23, 31, 39, 19, 28, 32, 32, 23, 22, 33, 18, 26, 17, 9, 0, 
    40, 30, 24, 35, 15, 31, 36, 6, 0, 21, 17, 15, 16, 15, 13, 
    12, 23, 38, 10, 17, 0, 48, 32, 4, 11, 14, 18, 10, 7, 11, 
    7, 20, 37, 19, 5, 0, 14, 13, 9, 12, 14, 1, 19, 7, 10, 
    0, 0, 5, 4, 9, 9, 4, 8, 15, 12, 12, 5, 10, 7, 7, 
    9, 3, 4, 4, 10, 11, 9, 11, 0, 21, 8, 7, 5, 8, 12, 
    
    -- channel=80
    0, 0, 0, 4, 11, 16, 24, 32, 24, 32, 34, 31, 32, 33, 29, 
    8, 0, 6, 20, 24, 29, 36, 33, 29, 52, 15, 34, 38, 41, 32, 
    20, 4, 16, 30, 36, 35, 45, 38, 29, 55, 2, 28, 42, 44, 37, 
    38, 16, 44, 46, 56, 45, 47, 41, 38, 22, 0, 21, 25, 51, 47, 
    29, 21, 31, 36, 47, 47, 35, 35, 3, 0, 0, 0, 8, 42, 38, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 33, 32, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 46, 48, 35, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 11, 30, 36, 24, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 2, 23, 22, 25, 37, 
    0, 0, 0, 0, 0, 0, 0, 11, 1, 7, 14, 29, 29, 29, 16, 
    0, 0, 0, 0, 0, 0, 9, 1, 0, 13, 20, 16, 9, 1, 12, 
    0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    
    -- channel=81
    54, 69, 68, 69, 66, 65, 61, 52, 61, 60, 64, 57, 55, 54, 59, 
    52, 65, 67, 59, 58, 58, 60, 58, 59, 56, 78, 62, 56, 56, 61, 
    47, 63, 61, 49, 48, 50, 47, 71, 70, 39, 79, 80, 56, 56, 62, 
    52, 58, 63, 63, 51, 51, 43, 35, 71, 64, 69, 93, 95, 63, 72, 
    75, 71, 68, 78, 75, 78, 75, 60, 47, 43, 51, 23, 42, 31, 58, 
    32, 30, 26, 35, 23, 28, 46, 48, 42, 30, 30, 12, 0, 29, 20, 
    46, 42, 42, 54, 57, 43, 42, 31, 20, 24, 39, 53, 23, 44, 33, 
    39, 25, 24, 37, 50, 53, 54, 58, 66, 53, 66, 48, 40, 7, 0, 
    65, 78, 78, 73, 75, 80, 71, 50, 44, 18, 24, 37, 44, 34, 49, 
    43, 41, 58, 70, 60, 45, 47, 58, 69, 50, 48, 48, 58, 53, 51, 
    68, 60, 61, 63, 79, 75, 48, 51, 54, 60, 66, 55, 39, 32, 31, 
    69, 63, 51, 51, 41, 58, 55, 44, 46, 43, 40, 38, 25, 28, 20, 
    65, 70, 65, 58, 61, 57, 41, 35, 43, 43, 25, 30, 27, 23, 17, 
    48, 47, 37, 34, 33, 37, 38, 30, 22, 18, 27, 25, 21, 19, 16, 
    17, 18, 17, 18, 17, 17, 23, 24, 42, 19, 23, 22, 20, 20, 16, 
    
    -- channel=82
    0, 3, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 18, 0, 0, 0, 0, 2, 0, 0, 57, 10, 0, 0, 0, 
    0, 2, 21, 0, 0, 0, 0, 27, 33, 0, 108, 52, 0, 3, 9, 
    0, 5, 26, 29, 0, 2, 0, 0, 0, 9, 33, 68, 158, 39, 46, 
    57, 43, 48, 78, 64, 67, 51, 8, 0, 0, 11, 0, 14, 0, 33, 
    19, 0, 0, 11, 0, 0, 0, 0, 0, 0, 14, 0, 0, 55, 0, 
    14, 0, 0, 36, 23, 0, 0, 0, 0, 0, 14, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 60, 31, 0, 0, 0, 
    5, 27, 51, 23, 0, 10, 8, 0, 0, 0, 0, 0, 0, 0, 21, 
    0, 6, 2, 0, 3, 0, 0, 0, 34, 11, 0, 0, 2, 1, 26, 
    40, 0, 0, 0, 43, 55, 0, 0, 42, 38, 19, 6, 0, 2, 2, 
    70, 8, 0, 0, 0, 46, 0, 0, 11, 9, 1, 6, 0, 1, 0, 
    58, 30, 25, 22, 27, 30, 10, 5, 12, 18, 0, 14, 0, 5, 0, 
    23, 30, 19, 22, 17, 21, 18, 5, 22, 0, 7, 0, 0, 3, 0, 
    3, 7, 5, 4, 2, 0, 3, 0, 60, 0, 7, 2, 4, 10, 0, 
    
    -- channel=83
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 25, 20, 0, 42, 24, 0, 1, 0, 
    0, 1, 14, 17, 4, 0, 0, 0, 42, 67, 47, 105, 105, 30, 37, 
    74, 58, 70, 80, 82, 78, 65, 40, 4, 0, 0, 0, 0, 2, 54, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 
    0, 0, 8, 2, 5, 0, 0, 0, 0, 0, 0, 0, 0, 10, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 42, 19, 0, 0, 0, 
    4, 28, 27, 1, 0, 14, 14, 0, 0, 0, 0, 0, 0, 0, 19, 
    0, 0, 0, 0, 0, 0, 0, 1, 24, 0, 0, 0, 25, 40, 41, 
    3, 0, 0, 6, 32, 28, 0, 22, 20, 24, 37, 39, 22, 14, 12, 
    14, 3, 0, 10, 0, 6, 15, 0, 6, 17, 16, 17, 6, 7, 8, 
    21, 28, 34, 19, 31, 41, 17, 0, 16, 24, 6, 4, 7, 4, 0, 
    33, 37, 20, 12, 10, 16, 18, 12, 0, 0, 8, 3, 2, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 5, 19, 0, 2, 2, 0, 0, 2, 
    
    -- channel=84
    72, 78, 91, 87, 86, 79, 82, 74, 82, 84, 73, 80, 75, 79, 78, 
    68, 72, 85, 75, 78, 71, 76, 75, 78, 67, 75, 81, 72, 78, 77, 
    61, 62, 74, 62, 71, 63, 63, 67, 77, 31, 93, 78, 64, 68, 76, 
    49, 51, 62, 54, 52, 57, 51, 56, 45, 32, 43, 55, 82, 59, 55, 
    39, 36, 38, 48, 43, 49, 51, 48, 37, 39, 36, 32, 34, 24, 44, 
    34, 40, 28, 28, 42, 48, 57, 44, 41, 38, 44, 49, 16, 42, 11, 
    46, 36, 31, 51, 63, 53, 60, 49, 51, 51, 64, 53, 26, 36, 0, 
    50, 44, 56, 67, 72, 75, 76, 69, 67, 43, 45, 50, 41, 0, 15, 
    68, 50, 70, 81, 80, 72, 66, 57, 63, 34, 49, 46, 44, 41, 36, 
    42, 74, 67, 64, 64, 70, 68, 62, 53, 56, 55, 50, 39, 24, 21, 
    66, 67, 69, 58, 66, 64, 49, 24, 53, 62, 43, 29, 26, 13, 13, 
    72, 63, 46, 37, 42, 73, 43, 28, 32, 35, 31, 15, 17, 9, 0, 
    58, 50, 40, 35, 31, 31, 29, 30, 27, 18, 18, 19, 3, 4, 1, 
    15, 16, 15, 20, 20, 18, 18, 15, 24, 12, 7, 7, 2, 4, 3, 
    0, 1, 6, 9, 13, 14, 15, 4, 27, 0, 5, 1, 4, 4, 0, 
    
    -- channel=85
    25, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 2, 0, 0, 
    27, 0, 0, 0, 0, 0, 0, 0, 0, 58, 0, 0, 7, 0, 0, 
    29, 0, 0, 1, 0, 1, 23, 0, 0, 121, 0, 0, 13, 0, 0, 
    26, 0, 0, 0, 1, 0, 19, 31, 38, 48, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 37, 19, 11, 0, 0, 0, 38, 0, 
    0, 0, 23, 0, 0, 1, 0, 20, 0, 5, 0, 0, 78, 0, 61, 
    0, 1, 14, 0, 0, 8, 2, 7, 3, 0, 0, 0, 54, 6, 80, 
    0, 0, 0, 0, 0, 0, 0, 6, 0, 42, 0, 0, 7, 87, 19, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 36, 0, 0, 2, 15, 0, 
    19, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 21, 16, 33, 0, 
    0, 0, 0, 9, 0, 0, 45, 34, 0, 0, 9, 28, 22, 13, 14, 
    0, 0, 41, 8, 0, 0, 29, 7, 0, 6, 16, 8, 19, 7, 19, 
    0, 0, 10, 0, 0, 0, 5, 0, 1, 2, 13, 0, 25, 2, 6, 
    0, 0, 0, 0, 0, 0, 0, 7, 0, 29, 2, 5, 6, 0, 3, 
    3, 0, 0, 0, 0, 0, 0, 10, 0, 51, 0, 4, 0, 0, 34, 
    
    -- channel=86
    1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 24, 0, 0, 0, 
    25, 23, 12, 14, 36, 33, 17, 0, 2, 12, 31, 34, 37, 0, 0, 
    14, 8, 0, 15, 4, 22, 35, 47, 65, 46, 21, 0, 0, 0, 0, 
    36, 49, 54, 56, 28, 17, 10, 2, 0, 0, 0, 0, 0, 14, 75, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 12, 29, 0, 0, 0, 0, 
    34, 46, 14, 0, 0, 16, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 4, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 23, 5, 0, 0, 0, 0, 0, 0, 5, 1, 3, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 0, 10, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 15, 21, 1, 8, 10, 17, 18, 
    9, 15, 17, 19, 20, 21, 11, 0, 0, 2, 10, 11, 15, 15, 0, 
    
    -- channel=87
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 2, 0, 0, 
    6, 13, 14, 2, 37, 29, 8, 0, 0, 7, 24, 61, 76, 0, 19, 
    0, 0, 0, 0, 0, 16, 25, 44, 63, 46, 20, 0, 0, 0, 0, 
    27, 48, 59, 57, 28, 16, 10, 1, 0, 0, 0, 0, 0, 49, 89, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 41, 12, 0, 0, 0, 
    16, 30, 5, 0, 0, 9, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=88
    150, 91, 126, 137, 142, 134, 139, 153, 127, 143, 137, 136, 142, 146, 131, 
    143, 88, 114, 135, 134, 129, 134, 137, 126, 158, 70, 124, 142, 145, 124, 
    141, 78, 102, 127, 128, 123, 138, 99, 98, 171, 40, 103, 138, 127, 116, 
    128, 74, 106, 104, 119, 109, 126, 129, 88, 67, 23, 8, 38, 107, 80, 
    53, 40, 44, 34, 52, 53, 62, 98, 85, 82, 60, 60, 46, 92, 37, 
    38, 49, 86, 36, 73, 70, 84, 94, 71, 76, 44, 101, 127, 74, 84, 
    60, 62, 59, 37, 65, 96, 95, 97, 93, 93, 69, 89, 129, 64, 81, 
    85, 93, 102, 107, 115, 120, 125, 124, 110, 118, 46, 69, 92, 108, 67, 
    96, 77, 56, 102, 121, 110, 97, 95, 86, 122, 77, 87, 90, 99, 76, 
    82, 83, 100, 97, 90, 104, 112, 109, 75, 93, 94, 108, 87, 70, 35, 
    79, 98, 102, 105, 79, 74, 115, 62, 19, 78, 79, 68, 59, 42, 43, 
    44, 85, 106, 57, 55, 57, 108, 76, 47, 54, 58, 40, 42, 30, 25, 
    46, 75, 80, 61, 44, 35, 47, 50, 45, 36, 41, 27, 41, 20, 20, 
    18, 16, 22, 23, 32, 28, 23, 32, 21, 56, 26, 25, 22, 18, 23, 
    16, 9, 14, 15, 22, 28, 28, 32, 0, 56, 20, 19, 17, 15, 30, 
    
    -- channel=89
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 24, 9, 32, 5, 15, 0, 1, 0, 
    11, 0, 9, 7, 7, 0, 3, 0, 56, 67, 36, 88, 66, 31, 27, 
    65, 46, 59, 65, 68, 65, 52, 51, 8, 0, 1, 0, 0, 7, 36, 
    0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 26, 25, 2, 0, 0, 0, 
    9, 33, 8, 0, 6, 23, 19, 0, 0, 0, 0, 0, 0, 0, 26, 
    0, 0, 0, 9, 0, 0, 0, 15, 22, 0, 0, 9, 35, 48, 34, 
    0, 0, 0, 17, 36, 17, 16, 27, 0, 26, 44, 44, 27, 17, 21, 
    1, 3, 13, 9, 0, 0, 33, 5, 5, 18, 25, 20, 9, 10, 10, 
    16, 36, 45, 24, 34, 36, 12, 3, 22, 25, 7, 3, 15, 3, 0, 
    30, 30, 16, 7, 10, 18, 16, 14, 0, 0, 8, 4, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 12, 2, 11, 2, 1, 0, 0, 19, 
    
    -- channel=90
    24, 0, 4, 16, 17, 20, 23, 35, 19, 26, 28, 25, 33, 31, 23, 
    29, 1, 6, 26, 21, 27, 25, 22, 22, 49, 0, 18, 36, 30, 21, 
    34, 4, 9, 32, 31, 28, 38, 12, 8, 67, 0, 0, 35, 27, 18, 
    28, 4, 12, 9, 29, 23, 35, 40, 19, 2, 0, 0, 0, 14, 5, 
    0, 0, 0, 0, 0, 0, 0, 15, 7, 9, 0, 1, 2, 32, 1, 
    0, 1, 19, 0, 8, 13, 4, 9, 1, 8, 0, 18, 69, 1, 48, 
    0, 2, 2, 0, 0, 7, 8, 11, 18, 18, 0, 16, 39, 30, 36, 
    1, 8, 5, 6, 5, 10, 13, 18, 4, 28, 0, 3, 21, 48, 32, 
    0, 0, 0, 0, 5, 1, 2, 8, 9, 31, 12, 21, 17, 26, 13, 
    3, 0, 0, 2, 0, 9, 14, 16, 0, 6, 11, 24, 14, 13, 0, 
    0, 0, 3, 5, 0, 0, 24, 9, 0, 0, 4, 9, 9, 4, 7, 
    0, 0, 16, 0, 0, 0, 13, 4, 0, 4, 10, 0, 8, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 5, 0, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 21, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 2, 1, 3, 0, 19, 0, 0, 0, 0, 13, 
    
    -- channel=91
    0, 23, 0, 0, 0, 9, 0, 0, 0, 0, 15, 0, 11, 0, 8, 
    0, 30, 0, 10, 0, 9, 0, 0, 0, 0, 30, 0, 16, 0, 11, 
    0, 48, 0, 9, 0, 4, 0, 0, 10, 0, 0, 2, 13, 0, 0, 
    3, 57, 0, 5, 0, 0, 0, 0, 21, 9, 0, 34, 0, 0, 25, 
    8, 32, 3, 1, 9, 9, 16, 0, 17, 0, 6, 22, 8, 0, 25, 
    0, 18, 0, 6, 0, 3, 0, 9, 5, 0, 14, 0, 13, 0, 44, 
    0, 22, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 76, 
    1, 0, 0, 0, 0, 0, 0, 7, 0, 8, 0, 0, 7, 48, 0, 
    7, 5, 0, 0, 1, 3, 0, 0, 1, 0, 0, 0, 4, 20, 0, 
    9, 0, 0, 0, 0, 0, 0, 6, 23, 0, 0, 1, 15, 19, 18, 
    0, 0, 0, 9, 0, 0, 0, 24, 17, 0, 10, 10, 14, 14, 0, 
    0, 0, 0, 13, 0, 0, 7, 19, 5, 0, 10, 5, 2, 6, 10, 
    0, 8, 4, 12, 4, 0, 4, 2, 7, 0, 7, 7, 8, 3, 4, 
    2, 5, 1, 1, 1, 2, 0, 1, 0, 5, 2, 5, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 0, 29, 0, 4, 1, 0, 6, 
    
    -- channel=92
    135, 81, 119, 128, 134, 129, 137, 149, 127, 141, 139, 135, 137, 144, 128, 
    133, 82, 115, 129, 134, 126, 133, 140, 126, 156, 79, 127, 137, 145, 123, 
    134, 76, 108, 126, 132, 122, 138, 111, 108, 165, 51, 121, 141, 135, 120, 
    129, 70, 113, 114, 128, 114, 130, 124, 94, 67, 28, 21, 66, 127, 100, 
    65, 47, 56, 53, 71, 70, 75, 104, 76, 74, 57, 48, 54, 93, 42, 
    32, 40, 80, 33, 59, 56, 73, 85, 67, 69, 37, 90, 107, 86, 69, 
    55, 52, 52, 31, 57, 77, 74, 72, 69, 74, 64, 95, 123, 71, 73, 
    67, 71, 75, 84, 99, 105, 112, 113, 108, 117, 61, 73, 89, 84, 38, 
    82, 80, 51, 91, 110, 109, 99, 90, 78, 108, 70, 83, 87, 90, 90, 
    58, 60, 92, 90, 81, 91, 105, 110, 85, 94, 90, 104, 94, 76, 42, 
    75, 85, 90, 99, 85, 83, 107, 56, 16, 86, 88, 75, 61, 45, 45, 
    46, 77, 95, 45, 41, 55, 108, 75, 49, 54, 60, 47, 36, 28, 21, 
    50, 80, 86, 63, 51, 39, 41, 48, 50, 42, 37, 27, 38, 16, 15, 
    17, 16, 22, 23, 36, 34, 25, 32, 16, 50, 25, 19, 17, 13, 17, 
    14, 7, 12, 12, 18, 24, 28, 33, 2, 48, 16, 13, 13, 13, 28, 
    
    -- channel=93
    77, 71, 77, 71, 67, 58, 53, 49, 50, 50, 46, 45, 43, 46, 43, 
    67, 60, 64, 55, 54, 45, 46, 50, 45, 44, 52, 42, 39, 44, 41, 
    55, 48, 51, 40, 39, 36, 38, 46, 50, 42, 56, 55, 40, 39, 38, 
    43, 36, 34, 32, 24, 28, 31, 28, 44, 60, 50, 54, 63, 38, 32, 
    51, 39, 42, 40, 37, 37, 45, 53, 54, 55, 55, 38, 23, 22, 21, 
    46, 39, 40, 40, 33, 38, 54, 64, 56, 51, 45, 24, 2, 24, 11, 
    56, 48, 51, 53, 63, 59, 64, 58, 50, 49, 40, 32, 22, 14, 21, 
    59, 49, 47, 55, 66, 70, 73, 70, 72, 56, 47, 28, 23, 8, 2, 
    74, 76, 78, 80, 81, 85, 83, 68, 53, 39, 25, 27, 35, 30, 33, 
    67, 62, 70, 75, 79, 69, 63, 61, 62, 54, 43, 41, 43, 41, 36, 
    87, 78, 76, 73, 77, 81, 61, 53, 51, 56, 55, 53, 43, 39, 29, 
    78, 77, 70, 63, 57, 62, 64, 51, 48, 50, 47, 48, 37, 34, 28, 
    69, 73, 74, 63, 62, 59, 49, 46, 48, 50, 41, 39, 34, 31, 27, 
    47, 49, 46, 45, 44, 43, 45, 42, 40, 32, 36, 29, 31, 29, 27, 
    25, 25, 30, 30, 33, 34, 38, 34, 39, 35, 28, 27, 29, 30, 19, 
    
    -- channel=94
    15, 12, 41, 41, 49, 46, 57, 56, 61, 64, 62, 65, 52, 62, 56, 
    29, 22, 56, 46, 63, 54, 67, 72, 61, 68, 77, 70, 56, 71, 61, 
    36, 23, 60, 50, 69, 54, 64, 81, 75, 47, 67, 85, 65, 81, 71, 
    44, 20, 61, 69, 71, 62, 58, 31, 59, 62, 43, 93, 126, 86, 86, 
    66, 44, 68, 82, 86, 85, 70, 54, 1, 0, 0, 0, 1, 46, 53, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 0, 
    0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 3, 51, 29, 23, 0, 
    0, 0, 0, 0, 0, 0, 3, 6, 29, 29, 59, 50, 29, 0, 0, 
    1, 26, 33, 26, 22, 36, 42, 27, 12, 0, 0, 13, 25, 9, 47, 
    0, 0, 0, 20, 19, 0, 5, 23, 35, 33, 23, 26, 36, 36, 27, 
    10, 0, 6, 11, 37, 44, 23, 13, 11, 43, 45, 37, 8, 0, 0, 
    23, 14, 8, 0, 0, 17, 18, 0, 1, 14, 3, 3, 0, 0, 0, 
    12, 21, 22, 0, 19, 29, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    3, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=95
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 28, 39, 30, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 3, 
    7, 0, 0, 10, 13, 7, 0, 0, 0, 0, 0, 0, 12, 0, 0, 
    0, 0, 1, 4, 5, 11, 11, 18, 23, 11, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 43, 
    0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 
    23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 25, 10, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 21, 18, 0, 0, 0, 0, 1, 0, 7, 6, 1, 6, 
    0, 0, 0, 0, 0, 8, 1, 0, 0, 1, 1, 0, 0, 2, 5, 
    4, 3, 1, 0, 0, 0, 6, 8, 0, 0, 0, 0, 3, 2, 0, 
    1, 6, 10, 12, 7, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 
    
    -- channel=96
    79, 70, 57, 68, 73, 68, 70, 71, 71, 72, 73, 72, 80, 84, 87, 
    78, 75, 72, 43, 85, 91, 85, 92, 90, 93, 87, 87, 92, 86, 88, 
    75, 75, 79, 58, 51, 58, 53, 63, 56, 60, 68, 79, 88, 85, 88, 
    72, 74, 50, 42, 54, 51, 45, 51, 55, 48, 55, 55, 78, 84, 84, 
    74, 73, 70, 53, 59, 59, 64, 65, 64, 59, 63, 78, 74, 83, 82, 
    84, 74, 68, 80, 68, 69, 72, 71, 69, 70, 73, 76, 80, 81, 86, 
    90, 60, 43, 55, 85, 85, 82, 82, 83, 80, 82, 80, 81, 81, 83, 
    96, 87, 79, 41, 21, 72, 92, 89, 82, 79, 81, 80, 80, 78, 79, 
    100, 96, 91, 82, 11, 28, 47, 74, 88, 85, 85, 81, 80, 81, 82, 
    99, 93, 92, 86, 7, 10, 26, 30, 28, 29, 54, 76, 89, 88, 85, 
    99, 87, 91, 61, 52, 6, 13, 55, 44, 23, 30, 19, 66, 69, 79, 
    82, 70, 72, 71, 70, 59, 53, 60, 57, 55, 53, 54, 48, 52, 56, 
    45, 35, 32, 32, 35, 33, 30, 34, 34, 36, 34, 38, 40, 37, 34, 
    30, 24, 25, 26, 22, 20, 19, 22, 22, 17, 18, 18, 16, 14, 41, 
    21, 15, 14, 17, 16, 23, 18, 24, 22, 22, 18, 20, 21, 47, 27, 
    
    -- channel=97
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 8, 10, 6, 10, 11, 9, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 5, 2, 0, 1, 4, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 30, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 9, 11, 15, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 30, 35, 18, 32, 37, 32, 39, 25, 22, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 4, 7, 12, 16, 14, 12, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 4, 8, 6, 9, 12, 15, 17, 19, 20, 18, 20, 33, 
    23, 18, 18, 20, 22, 21, 24, 27, 26, 27, 28, 25, 28, 39, 20, 
    
    -- channel=98
    31, 24, 0, 13, 26, 18, 15, 19, 16, 18, 18, 19, 26, 36, 35, 
    25, 19, 7, 17, 50, 52, 44, 50, 51, 54, 53, 56, 42, 33, 36, 
    21, 13, 8, 50, 46, 63, 57, 75, 66, 61, 59, 59, 60, 30, 34, 
    18, 14, 1, 35, 42, 35, 33, 44, 37, 28, 43, 39, 54, 26, 30, 
    12, 13, 11, 12, 16, 16, 11, 18, 22, 12, 20, 34, 35, 25, 27, 
    22, 16, 20, 13, 16, 17, 23, 24, 21, 19, 21, 28, 23, 24, 26, 
    29, 0, 0, 18, 41, 28, 26, 27, 25, 23, 27, 25, 25, 26, 29, 
    35, 22, 12, 0, 0, 35, 49, 30, 27, 25, 26, 25, 24, 22, 25, 
    36, 32, 30, 25, 0, 0, 10, 31, 42, 35, 34, 26, 25, 23, 24, 
    40, 36, 33, 18, 0, 0, 0, 0, 0, 0, 15, 30, 41, 37, 30, 
    42, 32, 33, 7, 0, 0, 0, 11, 0, 0, 0, 0, 23, 25, 31, 
    47, 34, 31, 29, 32, 12, 23, 37, 22, 13, 23, 18, 25, 19, 22, 
    2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=99
    0, 0, 0, 1, 0, 1, 5, 2, 2, 2, 4, 4, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 3, 0, 0, 7, 7, 10, 0, 0, 0, 
    0, 0, 0, 2, 1, 1, 0, 0, 0, 2, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 16, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 27, 3, 12, 18, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 38, 12, 3, 1, 11, 29, 21, 16, 0, 0, 0, 
    0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 6, 11, 12, 11, 13, 0, 0, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    20, 15, 17, 14, 18, 14, 11, 11, 14, 13, 11, 11, 9, 10, 2, 
    13, 8, 8, 8, 10, 3, 6, 5, 8, 7, 8, 9, 3, 6, 17, 
    
    -- channel=100
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=101
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 16, 39, 38, 29, 34, 34, 29, 18, 0, 0, 0, 
    0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 2, 1, 0, 0, 0, 0, 0, 
    0, 2, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 74, 67, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 68, 44, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 60, 96, 82, 44, 4, 0, 0, 0, 0, 
    0, 0, 0, 13, 47, 21, 7, 0, 22, 75, 110, 114, 82, 30, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    81, 92, 103, 107, 113, 84, 59, 65, 73, 39, 48, 28, 46, 53, 47, 
    0, 0, 0, 0, 0, 0, 4, 26, 40, 47, 55, 59, 65, 69, 68, 
    38, 38, 34, 24, 23, 20, 15, 14, 9, 8, 4, 3, 2, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 
    
    -- channel=102
    97, 126, 126, 102, 95, 115, 113, 105, 111, 109, 113, 110, 111, 129, 126, 
    99, 118, 133, 97, 63, 55, 60, 57, 65, 67, 63, 60, 114, 124, 125, 
    93, 116, 133, 72, 101, 93, 90, 81, 105, 116, 105, 103, 98, 129, 128, 
    100, 115, 133, 84, 84, 85, 95, 89, 85, 90, 79, 100, 74, 122, 122, 
    115, 116, 123, 127, 98, 96, 94, 101, 102, 101, 97, 102, 128, 127, 124, 
    118, 122, 100, 115, 135, 133, 133, 136, 135, 133, 131, 129, 124, 125, 124, 
    119, 127, 106, 30, 42, 106, 124, 129, 129, 130, 123, 126, 125, 124, 121, 
    119, 132, 139, 157, 64, 19, 69, 120, 127, 124, 123, 125, 126, 127, 124, 
    119, 130, 133, 132, 122, 26, 12, 10, 47, 90, 106, 128, 126, 123, 122, 
    118, 127, 130, 137, 86, 2, 13, 27, 26, 7, 0, 16, 52, 95, 118, 
    113, 127, 127, 136, 119, 133, 61, 60, 135, 92, 101, 82, 78, 114, 107, 
    67, 75, 68, 63, 57, 63, 72, 74, 75, 84, 86, 92, 95, 84, 81, 
    56, 61, 64, 59, 56, 52, 51, 45, 43, 32, 31, 25, 24, 27, 11, 
    9, 5, 5, 3, 8, 5, 6, 6, 12, 11, 8, 13, 11, 11, 29, 
    15, 15, 16, 15, 14, 18, 24, 19, 25, 23, 20, 15, 14, 56, 50, 
    
    -- channel=103
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=104
    50, 49, 35, 40, 53, 47, 42, 46, 44, 47, 46, 45, 51, 49, 48, 
    52, 54, 43, 36, 64, 63, 54, 62, 56, 57, 57, 60, 62, 53, 54, 
    52, 51, 43, 48, 36, 48, 35, 53, 41, 37, 42, 49, 57, 51, 55, 
    50, 51, 38, 63, 61, 58, 52, 61, 68, 58, 65, 56, 78, 53, 57, 
    45, 51, 46, 34, 43, 43, 45, 49, 45, 41, 44, 57, 50, 50, 53, 
    43, 41, 41, 46, 40, 41, 46, 45, 42, 40, 42, 51, 51, 51, 53, 
    48, 33, 22, 51, 62, 57, 56, 55, 52, 48, 52, 49, 50, 52, 55, 
    53, 50, 28, 0, 18, 64, 62, 55, 52, 50, 51, 49, 50, 50, 53, 
    54, 51, 49, 37, 0, 18, 43, 57, 53, 49, 58, 53, 51, 50, 53, 
    52, 51, 52, 40, 0, 9, 14, 13, 20, 31, 61, 52, 50, 50, 55, 
    55, 53, 52, 23, 16, 0, 18, 46, 9, 5, 11, 12, 52, 50, 58, 
    44, 44, 40, 41, 44, 22, 26, 49, 47, 40, 44, 40, 49, 57, 56, 
    20, 25, 19, 14, 11, 10, 15, 28, 22, 25, 24, 29, 30, 27, 32, 
    12, 20, 16, 13, 5, 8, 9, 8, 2, 0, 1, 0, 0, 1, 10, 
    0, 1, 1, 1, 0, 5, 0, 2, 0, 0, 0, 0, 3, 2, 0, 
    
    -- channel=105
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 10, 12, 
    0, 0, 0, 28, 36, 48, 49, 44, 52, 51, 51, 41, 15, 10, 11, 
    0, 0, 0, 42, 42, 38, 47, 48, 42, 41, 39, 30, 31, 6, 8, 
    0, 0, 0, 13, 19, 14, 15, 14, 10, 18, 20, 21, 7, 5, 3, 
    0, 0, 0, 6, 0, 0, 0, 0, 3, 2, 2, 0, 8, 1, 1, 
    6, 3, 8, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 
    8, 0, 0, 0, 18, 7, 0, 1, 2, 4, 4, 5, 4, 4, 4, 
    7, 2, 12, 3, 0, 2, 22, 10, 7, 8, 4, 4, 2, 1, 0, 
    10, 12, 11, 22, 13, 0, 0, 15, 33, 27, 9, 3, 3, 2, 0, 
    16, 16, 13, 19, 35, 0, 0, 2, 0, 0, 0, 26, 35, 21, 6, 
    15, 10, 11, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 36, 38, 37, 36, 41, 29, 18, 19, 9, 13, 11, 8, 1, 6, 
    2, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    
    -- channel=106
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 4, 11, 11, 11, 7, 1, 1, 0, 0, 0, 0, 
    0, 0, 0, 48, 10, 4, 21, 13, 11, 16, 12, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 43, 51, 35, 25, 23, 34, 36, 34, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 5, 5, 4, 4, 9, 12, 
    13, 7, 6, 5, 9, 12, 12, 12, 12, 14, 8, 9, 12, 0, 0, 
    
    -- channel=107
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=108
    38, 6, 0, 3, 16, 2, 1, 6, 5, 6, 6, 3, 14, 15, 9, 
    36, 12, 0, 0, 21, 4, 0, 6, 0, 3, 0, 6, 21, 1, 6, 
    32, 13, 0, 0, 0, 8, 0, 11, 0, 0, 1, 12, 18, 5, 6, 
    29, 13, 0, 0, 4, 0, 0, 0, 1, 0, 5, 0, 36, 6, 7, 
    19, 14, 0, 0, 0, 0, 0, 1, 0, 0, 1, 17, 3, 5, 5, 
    19, 4, 0, 2, 8, 8, 12, 5, 2, 7, 10, 17, 0, 2, 8, 
    25, 0, 0, 6, 8, 7, 5, 2, 1, 0, 4, 0, 2, 1, 3, 
    33, 4, 0, 0, 5, 33, 17, 3, 0, 0, 3, 1, 3, 1, 5, 
    34, 10, 3, 0, 0, 22, 32, 11, 0, 0, 6, 2, 1, 1, 4, 
    33, 9, 4, 0, 0, 4, 16, 15, 19, 0, 8, 0, 0, 3, 7, 
    34, 2, 5, 0, 0, 0, 32, 72, 30, 0, 43, 24, 85, 36, 17, 
    11, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 0, 5, 2, 7, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 4, 6, 9, 6, 6, 12, 11, 12, 15, 49, 
    0, 8, 8, 15, 9, 21, 15, 22, 16, 19, 16, 17, 31, 53, 3, 
    
    -- channel=109
    29, 45, 51, 32, 35, 39, 39, 38, 37, 38, 37, 41, 34, 28, 33, 
    32, 51, 49, 23, 0, 0, 0, 0, 0, 0, 4, 9, 22, 37, 36, 
    35, 51, 41, 10, 0, 0, 0, 0, 0, 0, 0, 0, 18, 37, 36, 
    35, 50, 51, 0, 3, 9, 8, 0, 3, 11, 1, 3, 5, 39, 44, 
    35, 47, 51, 49, 40, 43, 43, 39, 40, 47, 37, 37, 30, 43, 43, 
    34, 45, 52, 39, 36, 32, 30, 32, 31, 33, 32, 31, 44, 43, 41, 
    31, 57, 45, 49, 37, 36, 40, 40, 39, 39, 38, 41, 42, 43, 44, 
    30, 44, 41, 13, 26, 28, 28, 36, 42, 43, 38, 40, 41, 43, 44, 
    26, 37, 38, 43, 48, 8, 21, 40, 31, 31, 37, 40, 42, 43, 43, 
    25, 36, 38, 37, 74, 23, 9, 3, 16, 48, 50, 42, 31, 32, 36, 
    27, 38, 38, 55, 16, 6, 15, 0, 0, 21, 0, 17, 0, 17, 34, 
    33, 47, 49, 50, 50, 55, 29, 29, 62, 46, 48, 45, 50, 63, 59, 
    16, 23, 21, 18, 12, 13, 12, 17, 26, 25, 28, 28, 30, 30, 34, 
    28, 29, 29, 24, 24, 23, 19, 16, 17, 16, 13, 12, 14, 19, 7, 
    12, 13, 14, 11, 12, 6, 7, 5, 9, 8, 8, 8, 12, 5, 40, 
    
    -- channel=110
    0, 0, 21, 11, 0, 6, 16, 4, 10, 9, 11, 11, 0, 0, 0, 
    0, 0, 0, 68, 31, 19, 35, 17, 27, 21, 21, 0, 0, 0, 0, 
    0, 0, 5, 16, 19, 4, 19, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 30, 48, 27, 24, 32, 25, 34, 57, 35, 34, 0, 0, 0, 
    0, 0, 0, 23, 1, 0, 0, 0, 2, 10, 3, 0, 0, 0, 0, 
    0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 30, 69, 31, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 5, 50, 49, 0, 0, 0, 7, 5, 0, 0, 0, 0, 0, 
    0, 0, 2, 14, 130, 6, 7, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 2, 2, 43, 134, 16, 1, 5, 20, 50, 1, 0, 0, 0, 0, 
    0, 1, 1, 43, 16, 67, 18, 0, 7, 31, 0, 30, 0, 0, 0, 
    0, 4, 8, 7, 2, 14, 0, 0, 9, 0, 0, 0, 0, 2, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 5, 5, 
    36, 28, 30, 21, 32, 25, 20, 17, 23, 22, 16, 15, 15, 5, 0, 
    28, 15, 16, 14, 17, 6, 18, 8, 19, 18, 19, 17, 0, 0, 25, 
    
    -- channel=111
    24, 45, 26, 18, 17, 26, 24, 19, 16, 16, 20, 19, 20, 31, 29, 
    23, 29, 44, 7, 0, 0, 1, 0, 4, 5, 11, 2, 27, 27, 27, 
    20, 30, 27, 21, 36, 18, 18, 16, 34, 34, 22, 11, 28, 30, 27, 
    20, 33, 46, 0, 5, 1, 8, 0, 0, 6, 3, 19, 0, 26, 24, 
    31, 29, 38, 38, 21, 19, 17, 16, 22, 25, 17, 21, 30, 31, 27, 
    41, 31, 23, 59, 41, 42, 40, 43, 45, 43, 40, 24, 30, 28, 25, 
    35, 43, 1, 0, 19, 40, 28, 31, 33, 33, 29, 33, 30, 28, 26, 
    33, 36, 70, 83, 0, 0, 33, 34, 26, 32, 28, 32, 33, 31, 27, 
    30, 33, 31, 52, 43, 0, 0, 0, 19, 36, 32, 31, 29, 28, 28, 
    31, 28, 30, 25, 57, 0, 1, 8, 0, 0, 0, 0, 27, 39, 32, 
    27, 30, 27, 71, 60, 39, 0, 1, 58, 12, 40, 0, 0, 3, 10, 
    15, 19, 16, 14, 9, 47, 38, 13, 18, 37, 24, 43, 19, 12, 19, 
    11, 23, 24, 29, 24, 27, 23, 6, 16, 9, 9, 2, 3, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 5, 0, 
    0, 0, 4, 0, 3, 1, 2, 0, 4, 2, 1, 3, 9, 2, 11, 
    
    -- channel=112
    12, 10, 13, 23, 19, 20, 24, 20, 21, 21, 23, 23, 18, 25, 24, 
    5, 1, 10, 66, 77, 70, 72, 69, 74, 72, 66, 54, 29, 27, 26, 
    1, 2, 20, 70, 68, 73, 79, 77, 69, 71, 67, 64, 33, 22, 24, 
    3, 2, 25, 81, 64, 54, 63, 67, 63, 72, 67, 63, 48, 21, 20, 
    8, 3, 6, 29, 21, 21, 15, 23, 24, 23, 24, 14, 27, 15, 16, 
    13, 18, 16, 4, 7, 8, 11, 16, 15, 10, 11, 15, 16, 18, 15, 
    17, 11, 18, 38, 22, 12, 17, 20, 19, 21, 19, 20, 19, 20, 20, 
    17, 16, 15, 20, 33, 22, 20, 22, 27, 25, 22, 21, 18, 17, 15, 
    18, 24, 24, 28, 51, 16, 26, 39, 37, 30, 18, 22, 21, 18, 17, 
    23, 30, 28, 44, 57, 19, 17, 20, 23, 35, 30, 40, 32, 21, 20, 
    26, 26, 26, 32, 7, 12, 0, 0, 8, 0, 0, 0, 0, 15, 23, 
    43, 43, 45, 45, 44, 42, 28, 25, 35, 25, 24, 22, 23, 27, 24, 
    21, 15, 14, 13, 12, 12, 12, 14, 20, 18, 19, 19, 20, 24, 20, 
    29, 24, 22, 16, 20, 19, 15, 14, 15, 13, 11, 12, 11, 2, 0, 
    23, 13, 12, 12, 12, 7, 10, 7, 10, 7, 11, 9, 0, 0, 2, 
    
    -- channel=113
    56, 64, 48, 49, 57, 54, 48, 49, 46, 49, 49, 50, 50, 51, 54, 
    63, 71, 54, 46, 65, 79, 72, 75, 72, 72, 75, 71, 65, 63, 63, 
    64, 68, 63, 59, 32, 34, 33, 39, 34, 29, 34, 45, 68, 60, 64, 
    59, 67, 46, 42, 49, 50, 38, 49, 56, 50, 51, 48, 65, 65, 68, 
    54, 66, 59, 54, 60, 63, 59, 59, 63, 58, 58, 59, 61, 60, 66, 
    52, 62, 78, 57, 41, 43, 47, 48, 46, 44, 44, 58, 63, 60, 61, 
    54, 43, 24, 87, 106, 77, 65, 64, 60, 59, 63, 62, 64, 66, 69, 
    58, 61, 30, 0, 32, 100, 96, 69, 62, 61, 60, 60, 60, 60, 65, 
    58, 60, 57, 45, 0, 31, 69, 103, 102, 83, 74, 62, 62, 63, 65, 
    55, 59, 59, 55, 22, 32, 28, 23, 36, 67, 111, 111, 100, 80, 67, 
    59, 62, 62, 38, 0, 0, 0, 0, 0, 0, 0, 0, 14, 37, 62, 
    90, 99, 100, 102, 107, 82, 72, 91, 95, 78, 83, 73, 85, 95, 95, 
    34, 42, 37, 37, 35, 32, 39, 58, 62, 66, 70, 75, 79, 78, 82, 
    35, 46, 42, 35, 25, 26, 27, 25, 18, 15, 15, 15, 15, 13, 0, 
    11, 16, 14, 13, 10, 7, 4, 4, 1, 0, 3, 3, 8, 0, 26, 
    
    -- channel=114
    33, 2, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 11, 0, 0, 17, 28, 9, 26, 13, 18, 19, 26, 10, 0, 0, 
    32, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 
    13, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 
    0, 0, 8, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 52, 120, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 0, 0, 0, 0, 128, 103, 5, 0, 0, 0, 0, 0, 0, 0, 
    22, 0, 0, 0, 0, 20, 63, 122, 109, 46, 23, 0, 0, 0, 0, 
    23, 0, 0, 0, 0, 22, 33, 10, 9, 35, 129, 132, 108, 46, 0, 
    30, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 21, 0, 0, 
    87, 64, 68, 77, 85, 47, 51, 74, 49, 30, 43, 29, 31, 41, 46, 
    0, 0, 0, 0, 0, 0, 4, 27, 17, 33, 34, 45, 48, 39, 47, 
    0, 25, 18, 19, 7, 11, 12, 12, 5, 0, 6, 2, 4, 7, 8, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 
    
    -- channel=115
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 20, 30, 28, 25, 23, 24, 23, 20, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 9, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 74, 83, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 86, 53, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 57, 112, 83, 30, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 27, 18, 0, 15, 73, 131, 123, 77, 21, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    64, 69, 79, 85, 91, 68, 32, 43, 63, 34, 34, 22, 25, 51, 49, 
    0, 0, 0, 0, 0, 0, 0, 9, 23, 32, 37, 45, 50, 50, 59, 
    30, 44, 40, 32, 25, 24, 21, 18, 13, 6, 7, 3, 4, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    
    -- channel=116
    75, 72, 51, 49, 62, 57, 55, 57, 54, 57, 59, 57, 63, 68, 68, 
    76, 84, 69, 7, 36, 31, 25, 30, 28, 34, 31, 42, 70, 70, 71, 
    75, 82, 67, 10, 10, 16, 0, 14, 16, 19, 21, 31, 60, 75, 73, 
    72, 80, 51, 11, 30, 29, 23, 25, 32, 23, 30, 29, 58, 75, 77, 
    68, 78, 72, 51, 53, 55, 55, 57, 59, 50, 52, 72, 62, 75, 76, 
    71, 77, 67, 64, 66, 65, 67, 65, 63, 64, 66, 71, 73, 70, 76, 
    75, 43, 33, 63, 76, 67, 73, 73, 71, 70, 72, 72, 73, 74, 76, 
    80, 74, 60, 8, 24, 69, 72, 68, 71, 69, 70, 70, 72, 71, 76, 
    79, 75, 73, 59, 0, 12, 33, 66, 66, 61, 67, 70, 71, 72, 76, 
    77, 72, 74, 69, 0, 6, 8, 4, 10, 23, 56, 67, 65, 64, 70, 
    79, 69, 72, 37, 22, 0, 6, 43, 22, 1, 14, 7, 65, 57, 71, 
    73, 64, 62, 61, 61, 49, 50, 59, 63, 62, 61, 62, 61, 69, 69, 
    30, 27, 25, 21, 21, 20, 22, 29, 25, 28, 26, 30, 31, 26, 27, 
    7, 10, 8, 6, 3, 3, 4, 4, 3, 0, 0, 0, 0, 0, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 41, 16, 
    
    -- channel=117
    0, 0, 29, 2, 0, 0, 9, 0, 3, 0, 2, 2, 0, 0, 0, 
    0, 0, 4, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 16, 15, 0, 11, 0, 2, 11, 2, 0, 0, 0, 0, 
    0, 0, 20, 19, 0, 0, 16, 0, 0, 20, 0, 6, 0, 0, 0, 
    0, 0, 0, 29, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 1, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 
    0, 41, 64, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 24, 94, 30, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 17, 174, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 33, 172, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 54, 50, 103, 8, 0, 29, 50, 10, 30, 0, 0, 0, 
    0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 0, 4, 0, 8, 3, 0, 0, 5, 7, 0, 1, 0, 0, 0, 
    23, 4, 3, 0, 5, 0, 7, 0, 9, 7, 7, 3, 0, 0, 11, 
    
    -- channel=118
    0, 0, 7, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 6, 8, 7, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 20, 17, 14, 9, 9, 9, 9, 0, 0, 0, 0, 
    0, 8, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 65, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 74, 127, 92, 80, 88, 90, 102, 97, 61, 26, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 
    0, 2, 2, 3, 0, 15, 18, 15, 17, 20, 11, 2, 9, 44, 0, 
    
    -- channel=119
    0, 0, 23, 2, 0, 6, 10, 6, 15, 9, 9, 7, 9, 13, 2, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 30, 45, 34, 33, 48, 50, 43, 33, 0, 0, 0, 
    0, 0, 6, 52, 17, 14, 41, 24, 13, 12, 3, 17, 0, 0, 0, 
    3, 0, 2, 13, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 
    0, 0, 0, 0, 36, 34, 31, 30, 31, 28, 26, 10, 0, 0, 0, 
    0, 27, 44, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 30, 124, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 77, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 16, 118, 181, 98, 83, 133, 124, 132, 117, 59, 40, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 
    1, 0, 0, 0, 0, 12, 20, 15, 19, 21, 12, 2, 9, 41, 0, 
    
    -- channel=120
    83, 120, 128, 105, 94, 109, 110, 100, 106, 102, 109, 107, 103, 122, 122, 
    86, 114, 138, 119, 89, 96, 100, 92, 105, 105, 101, 87, 118, 126, 125, 
    85, 113, 137, 110, 112, 91, 98, 81, 102, 115, 103, 100, 105, 129, 126, 
    93, 112, 143, 86, 87, 86, 92, 84, 87, 100, 84, 100, 66, 123, 121, 
    112, 112, 127, 132, 99, 97, 97, 100, 108, 105, 93, 93, 124, 128, 125, 
    117, 129, 114, 122, 131, 130, 128, 134, 136, 131, 126, 120, 125, 124, 124, 
    112, 131, 109, 39, 65, 111, 125, 132, 134, 136, 127, 131, 127, 127, 122, 
    108, 132, 152, 167, 60, 23, 79, 123, 130, 130, 124, 128, 128, 128, 124, 
    109, 129, 135, 141, 172, 26, 3, 27, 74, 109, 110, 131, 129, 126, 125, 
    108, 125, 131, 150, 153, 13, 19, 33, 21, 12, 0, 48, 77, 106, 122, 
    101, 127, 128, 149, 126, 125, 35, 27, 118, 82, 79, 59, 40, 91, 103, 
    78, 103, 98, 92, 84, 110, 94, 76, 97, 110, 96, 111, 97, 97, 98, 
    61, 75, 79, 74, 70, 69, 66, 56, 70, 60, 59, 53, 56, 61, 46, 
    22, 18, 24, 16, 20, 14, 17, 16, 23, 19, 14, 20, 17, 11, 7, 
    28, 21, 22, 18, 20, 17, 28, 19, 27, 25, 25, 21, 4, 38, 48, 
    
    -- channel=121
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 1, 15, 20, 14, 16, 12, 19, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 68, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 60, 31, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 41, 89, 67, 23, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 41, 22, 5, 0, 9, 66, 102, 103, 60, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    59, 73, 81, 86, 91, 74, 37, 38, 62, 32, 36, 21, 29, 46, 45, 
    0, 0, 0, 0, 0, 0, 0, 10, 27, 32, 37, 43, 46, 48, 53, 
    23, 33, 30, 21, 19, 16, 12, 9, 5, 3, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 
    
    -- channel=122
    0, 5, 26, 19, 1, 14, 20, 14, 19, 16, 18, 17, 11, 18, 21, 
    0, 1, 12, 30, 10, 0, 10, 3, 9, 8, 8, 1, 4, 14, 17, 
    0, 5, 14, 19, 16, 17, 24, 11, 18, 27, 26, 20, 5, 13, 16, 
    1, 3, 3, 14, 4, 7, 12, 4, 4, 8, 0, 9, 3, 12, 11, 
    13, 5, 10, 24, 9, 7, 7, 6, 10, 10, 10, 0, 21, 13, 14, 
    15, 21, 7, 0, 22, 19, 16, 18, 22, 21, 17, 15, 13, 16, 16, 
    11, 31, 46, 0, 0, 0, 11, 15, 18, 21, 14, 16, 14, 12, 10, 
    6, 19, 32, 71, 39, 0, 0, 7, 18, 17, 15, 17, 15, 15, 13, 
    8, 19, 22, 29, 96, 0, 0, 0, 0, 0, 0, 16, 17, 15, 13, 
    8, 19, 19, 38, 74, 0, 0, 2, 3, 0, 0, 0, 0, 0, 8, 
    3, 17, 19, 36, 45, 78, 19, 0, 48, 50, 32, 38, 0, 14, 12, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 4, 9, 9, 10, 8, 3, 0, 1, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 8, 3, 2, 3, 8, 10, 6, 7, 6, 1, 8, 
    20, 8, 7, 7, 10, 6, 16, 11, 18, 17, 17, 13, 0, 25, 25, 
    
    -- channel=123
    0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 48, 0, 3, 9, 7, 9, 0, 3, 19, 0, 0, 0, 
    0, 0, 5, 61, 5, 0, 24, 1, 8, 0, 0, 12, 0, 0, 1, 
    0, 0, 10, 41, 5, 13, 25, 9, 16, 14, 0, 0, 0, 0, 0, 
    0, 0, 2, 0, 0, 3, 2, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 12, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 35, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 77, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 74, 8, 0, 0, 0, 0, 12, 9, 1, 0, 0, 
    0, 0, 0, 0, 14, 6, 0, 0, 0, 27, 0, 0, 0, 0, 0, 
    0, 19, 19, 19, 22, 24, 14, 1, 10, 26, 4, 14, 1, 10, 11, 
    0, 3, 5, 4, 4, 6, 6, 2, 9, 8, 9, 9, 10, 11, 12, 
    21, 6, 4, 8, 6, 3, 5, 3, 0, 6, 3, 1, 1, 1, 0, 
    25, 5, 0, 0, 4, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    
    -- channel=124
    78, 110, 111, 93, 82, 98, 97, 88, 91, 89, 95, 94, 91, 111, 114, 
    81, 108, 126, 98, 71, 89, 91, 83, 96, 97, 95, 79, 108, 116, 116, 
    82, 105, 129, 86, 95, 69, 78, 61, 81, 93, 86, 82, 101, 120, 118, 
    86, 104, 124, 50, 59, 63, 66, 56, 58, 71, 58, 77, 44, 115, 111, 
    101, 102, 114, 117, 89, 87, 86, 87, 97, 96, 87, 85, 110, 117, 114, 
    112, 121, 115, 115, 113, 111, 110, 116, 117, 117, 113, 107, 115, 113, 111, 
    107, 113, 82, 43, 81, 111, 112, 118, 120, 122, 116, 121, 118, 118, 114, 
    107, 122, 138, 133, 42, 41, 96, 118, 119, 118, 113, 116, 117, 116, 111, 
    111, 123, 127, 133, 135, 27, 15, 49, 96, 117, 106, 116, 116, 116, 113, 
    111, 120, 124, 142, 137, 15, 22, 31, 24, 19, 12, 77, 103, 114, 112, 
    101, 119, 120, 136, 83, 73, 3, 1, 85, 47, 44, 26, 20, 75, 91, 
    99, 121, 119, 115, 108, 126, 108, 90, 103, 106, 101, 107, 97, 92, 96, 
    53, 63, 67, 67, 65, 65, 60, 55, 68, 62, 62, 57, 61, 65, 50, 
    21, 21, 26, 21, 26, 17, 18, 19, 26, 22, 18, 22, 19, 14, 9, 
    22, 20, 22, 19, 21, 13, 22, 17, 24, 21, 24, 23, 8, 40, 75, 
    
    -- channel=125
    46, 57, 47, 37, 41, 39, 36, 36, 34, 36, 36, 36, 37, 37, 43, 
    57, 71, 61, 5, 6, 23, 19, 18, 19, 22, 23, 26, 47, 48, 46, 
    59, 69, 64, 4, 0, 0, 0, 0, 0, 0, 0, 0, 39, 49, 49, 
    56, 70, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 53, 55, 
    54, 66, 62, 44, 44, 45, 48, 44, 45, 45, 40, 46, 42, 56, 57, 
    54, 61, 67, 64, 48, 46, 46, 45, 45, 47, 47, 48, 58, 53, 55, 
    50, 48, 28, 48, 74, 66, 56, 55, 54, 53, 54, 55, 56, 56, 57, 
    51, 58, 46, 4, 7, 61, 68, 55, 50, 50, 50, 52, 54, 54, 57, 
    51, 52, 50, 44, 4, 17, 29, 59, 67, 61, 58, 51, 53, 56, 58, 
    46, 46, 48, 46, 23, 15, 15, 9, 12, 32, 60, 71, 70, 62, 56, 
    46, 48, 49, 39, 4, 0, 0, 3, 0, 0, 0, 0, 14, 26, 45, 
    58, 67, 66, 67, 68, 67, 56, 57, 67, 60, 62, 60, 60, 67, 68, 
    23, 32, 30, 30, 28, 30, 32, 41, 47, 50, 51, 54, 58, 56, 54, 
    16, 26, 26, 22, 16, 17, 18, 17, 15, 12, 11, 10, 10, 10, 20, 
    0, 9, 10, 8, 7, 8, 5, 5, 4, 4, 5, 8, 12, 26, 39, 
    
    -- channel=126
    35, 29, 7, 25, 32, 28, 29, 28, 23, 29, 30, 30, 28, 29, 35, 
    36, 38, 26, 16, 49, 64, 62, 61, 62, 63, 62, 55, 42, 43, 40, 
    36, 36, 43, 8, 7, 0, 0, 2, 0, 0, 0, 3, 52, 39, 40, 
    26, 33, 29, 0, 10, 10, 0, 10, 13, 21, 26, 24, 26, 44, 43, 
    23, 33, 24, 20, 28, 32, 31, 31, 32, 31, 33, 39, 21, 38, 37, 
    38, 32, 44, 31, 0, 0, 2, 5, 0, 3, 7, 20, 39, 36, 36, 
    46, 11, 0, 82, 96, 52, 36, 35, 32, 30, 35, 34, 38, 43, 44, 
    53, 40, 9, 0, 0, 90, 87, 51, 40, 38, 35, 34, 33, 32, 34, 
    58, 49, 43, 35, 0, 2, 57, 115, 102, 67, 48, 32, 36, 38, 37, 
    60, 49, 46, 47, 0, 0, 0, 0, 12, 65, 112, 122, 97, 62, 39, 
    63, 44, 48, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 39, 
    92, 84, 91, 96, 100, 69, 34, 54, 71, 34, 44, 27, 39, 57, 55, 
    0, 0, 0, 0, 0, 0, 0, 6, 19, 25, 29, 38, 43, 44, 45, 
    18, 28, 24, 15, 10, 6, 1, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
    
    -- channel=127
    0, 0, 0, 0, 0, 0, 3, 1, 3, 5, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 19, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 0, 0, 11, 22, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 28, 59, 75, 29, 17, 48, 43, 70, 15, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 7, 5, 7, 10, 11, 7, 6, 4, 8, 7, 2, 4, 18, 28, 
    6, 6, 4, 5, 8, 13, 11, 13, 17, 15, 5, 3, 24, 3, 0, 
    
    -- channel=128
    29, 11, 30, 31, 0, 33, 31, 35, 49, 54, 38, 69, 24, 32, 39, 
    38, 34, 32, 35, 0, 20, 22, 43, 39, 46, 33, 75, 35, 44, 39, 
    42, 49, 45, 24, 0, 31, 43, 37, 45, 17, 54, 77, 61, 58, 64, 
    12, 53, 34, 28, 20, 57, 59, 16, 59, 29, 53, 92, 75, 68, 30, 
    25, 78, 41, 18, 63, 65, 22, 52, 48, 67, 74, 83, 81, 68, 5, 
    18, 75, 76, 30, 61, 73, 53, 70, 71, 76, 60, 96, 76, 70, 3, 
    24, 56, 73, 77, 64, 62, 63, 62, 67, 65, 63, 76, 68, 77, 21, 
    39, 60, 71, 75, 63, 35, 70, 77, 64, 65, 69, 75, 66, 75, 5, 
    53, 65, 55, 62, 74, 75, 60, 66, 71, 77, 72, 77, 64, 53, 32, 
    63, 49, 44, 67, 51, 58, 78, 76, 76, 72, 70, 68, 36, 37, 60, 
    33, 67, 43, 49, 63, 59, 86, 83, 74, 66, 70, 67, 56, 53, 62, 
    72, 81, 62, 72, 51, 68, 82, 88, 79, 63, 75, 66, 60, 71, 68, 
    73, 110, 102, 90, 71, 75, 71, 51, 79, 75, 67, 59, 46, 54, 73, 
    31, 53, 113, 114, 90, 80, 75, 55, 63, 74, 79, 61, 14, 71, 73, 
    28, 26, 55, 119, 114, 99, 88, 84, 67, 67, 57, 50, 37, 37, 95, 
    
    -- channel=129
    33, 44, 42, 38, 29, 45, 38, 44, 37, 37, 30, 49, 25, 29, 36, 
    37, 51, 39, 35, 33, 34, 26, 40, 39, 44, 31, 46, 32, 52, 37, 
    18, 31, 32, 28, 35, 46, 57, 42, 36, 26, 31, 50, 29, 41, 34, 
    33, 43, 33, 29, 48, 59, 44, 31, 30, 46, 45, 53, 24, 36, 8, 
    40, 34, 36, 31, 51, 51, 31, 55, 54, 55, 46, 54, 31, 26, 8, 
    32, 26, 31, 49, 53, 33, 40, 52, 51, 44, 38, 63, 32, 29, 21, 
    45, 33, 34, 36, 34, 28, 39, 24, 22, 25, 32, 32, 36, 38, 31, 
    32, 32, 33, 24, 36, 28, 21, 28, 35, 34, 22, 25, 25, 30, 21, 
    44, 41, 30, 28, 11, 30, 26, 24, 19, 13, 25, 22, 3, 24, 38, 
    32, 24, 28, 25, 28, 13, 20, 21, 19, 14, 23, 19, 16, 28, 38, 
    21, 40, 39, 36, 34, 34, 20, 14, 15, 8, 15, 20, 26, 37, 43, 
    51, 62, 62, 47, 37, 24, 22, 12, 11, 19, 16, 20, 29, 40, 42, 
    14, 22, 56, 63, 45, 43, 18, 2, 10, 19, 16, 16, 24, 39, 40, 
    27, 18, 23, 55, 61, 56, 42, 42, 36, 12, 21, 16, 13, 40, 45, 
    32, 42, 33, 32, 52, 63, 64, 45, 32, 6, 8, 19, 44, 43, 54, 
    
    -- channel=130
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 12, 0, 0, 0, 0, 0, 11, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 6, 0, 0, 18, 8, 11, 3, 18, 17, 14, 3, 0, 0, 
    0, 0, 0, 0, 10, 14, 23, 24, 27, 18, 12, 47, 0, 0, 0, 
    0, 0, 0, 0, 20, 0, 42, 35, 26, 28, 27, 27, 8, 3, 0, 
    0, 0, 0, 0, 0, 45, 13, 30, 37, 28, 22, 18, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 45, 32, 28, 25, 22, 20, 1, 0, 0, 
    0, 8, 0, 0, 0, 0, 26, 38, 34, 12, 24, 27, 5, 11, 0, 
    0, 36, 0, 0, 0, 5, 15, 23, 39, 23, 46, 11, 3, 2, 0, 
    0, 0, 23, 4, 0, 0, 0, 0, 3, 35, 28, 14, 0, 0, 0, 
    0, 0, 10, 27, 12, 0, 0, 0, 0, 16, 32, 1, 0, 0, 21, 
    
    -- channel=131
    18, 13, 12, 14, 28, 0, 18, 9, 28, 23, 34, 0, 54, 13, 15, 
    13, 16, 24, 13, 25, 11, 19, 8, 23, 16, 32, 0, 46, 1, 22, 
    27, 20, 17, 17, 20, 0, 15, 27, 12, 35, 18, 0, 41, 20, 23, 
    31, 4, 24, 15, 5, 20, 44, 31, 8, 13, 17, 19, 40, 18, 45, 
    21, 0, 30, 27, 0, 23, 40, 0, 25, 20, 39, 22, 35, 21, 52, 
    24, 5, 19, 19, 25, 14, 14, 0, 22, 24, 32, 6, 42, 19, 50, 
    21, 9, 16, 20, 19, 14, 16, 20, 24, 12, 6, 14, 35, 19, 39, 
    24, 13, 13, 25, 10, 28, 15, 19, 10, 13, 20, 10, 21, 26, 43, 
    11, 13, 24, 24, 15, 5, 10, 14, 18, 26, 27, 12, 31, 23, 23, 
    18, 25, 29, 18, 24, 24, 2, 9, 17, 20, 18, 24, 33, 25, 10, 
    36, 13, 27, 11, 18, 12, 8, 15, 18, 26, 16, 25, 26, 12, 19, 
    2, 8, 40, 24, 28, 11, 9, 21, 17, 20, 11, 23, 33, 18, 33, 
    29, 29, 38, 40, 35, 20, 13, 40, 11, 12, 19, 23, 34, 24, 35, 
    37, 33, 31, 35, 45, 38, 43, 34, 5, 18, 16, 30, 46, 17, 11, 
    40, 20, 23, 28, 37, 36, 46, 40, 37, 19, 25, 27, 25, 21, 17, 
    
    -- channel=132
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=133
    0, 0, 0, 0, 10, 0, 0, 0, 16, 18, 7, 0, 8, 10, 0, 
    0, 0, 0, 0, 7, 12, 12, 0, 0, 0, 5, 0, 0, 0, 0, 
    40, 24, 0, 10, 7, 0, 0, 9, 13, 31, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 21, 37, 0, 0, 0, 0, 5, 0, 31, 
    0, 0, 0, 3, 0, 0, 4, 0, 0, 0, 1, 24, 0, 0, 31, 
    17, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 1, 9, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 39, 
    0, 0, 25, 15, 29, 0, 0, 0, 0, 0, 0, 1, 25, 44, 0, 
    0, 32, 20, 7, 11, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 0, 0, 0, 0, 0, 0, 0, 0, 8, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 8, 0, 6, 
    60, 51, 0, 0, 0, 0, 16, 62, 42, 0, 0, 0, 0, 20, 17, 
    8, 78, 49, 0, 0, 0, 0, 0, 0, 8, 0, 10, 49, 0, 0, 
    14, 0, 40, 39, 0, 0, 0, 0, 20, 32, 57, 11, 0, 0, 0, 
    
    -- channel=134
    42, 15, 27, 26, 33, 0, 33, 5, 35, 17, 49, 1, 86, 0, 18, 
    44, 31, 40, 34, 24, 0, 4, 2, 45, 33, 47, 6, 93, 36, 62, 
    34, 10, 29, 23, 11, 0, 36, 43, 14, 31, 16, 20, 103, 57, 72, 
    31, 28, 55, 30, 0, 39, 55, 0, 4, 33, 36, 44, 86, 71, 91, 
    40, 36, 96, 30, 13, 59, 54, 1, 57, 51, 65, 22, 76, 73, 83, 
    31, 20, 70, 82, 50, 44, 35, 66, 66, 52, 44, 34, 81, 62, 84, 
    47, 34, 38, 87, 57, 43, 44, 49, 36, 44, 50, 57, 55, 63, 76, 
    37, 34, 56, 75, 87, 34, 42, 57, 66, 65, 56, 54, 92, 52, 47, 
    43, 62, 44, 47, 47, 92, 52, 63, 71, 59, 54, 64, 52, 36, 51, 
    65, 36, 39, 34, 51, 24, 71, 82, 70, 87, 58, 67, 61, 37, 21, 
    61, 24, 49, 38, 47, 66, 45, 90, 88, 68, 57, 58, 51, 34, 76, 
    58, 112, 90, 44, 64, 43, 73, 72, 71, 75, 74, 64, 50, 31, 54, 
    39, 27, 98, 88, 67, 50, 71, 54, 18, 70, 73, 65, 59, 0, 57, 
    53, 0, 5, 84, 97, 66, 52, 59, 51, 64, 67, 61, 33, 9, 31, 
    55, 25, 0, 25, 88, 108, 88, 70, 45, 40, 42, 31, 51, 42, 51, 
    
    -- channel=135
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=136
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 21, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 31, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 
    0, 4, 0, 0, 0, 0, 0, 0, 15, 0, 0, 10, 0, 0, 0, 
    0, 20, 0, 0, 8, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 
    0, 8, 12, 0, 0, 9, 3, 11, 11, 14, 14, 17, 0, 0, 0, 
    0, 5, 10, 0, 1, 6, 22, 16, 6, 14, 22, 28, 0, 2, 0, 
    0, 0, 0, 0, 25, 5, 24, 18, 23, 27, 14, 24, 10, 0, 0, 
    0, 0, 0, 4, 0, 25, 24, 28, 26, 18, 21, 11, 0, 0, 5, 
    0, 5, 0, 0, 1, 0, 41, 24, 22, 18, 23, 13, 0, 0, 0, 
    2, 0, 0, 0, 0, 12, 25, 27, 27, 11, 24, 15, 0, 7, 0, 
    12, 24, 0, 0, 0, 2, 9, 6, 36, 22, 21, 10, 0, 7, 0, 
    0, 11, 24, 0, 0, 0, 0, 0, 19, 25, 24, 8, 0, 7, 0, 
    0, 0, 16, 19, 0, 0, 0, 0, 0, 18, 15, 3, 0, 0, 19, 
    
    -- channel=137
    0, 0, 0, 0, 0, 0, 0, 0, 7, 6, 6, 0, 38, 0, 0, 
    0, 0, 2, 0, 0, 0, 0, 0, 5, 0, 12, 0, 38, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 36, 0, 3, 
    0, 0, 0, 0, 0, 0, 9, 7, 0, 0, 0, 0, 39, 4, 28, 
    0, 0, 6, 0, 0, 14, 23, 0, 11, 0, 14, 15, 28, 5, 28, 
    3, 0, 9, 0, 0, 6, 28, 20, 19, 23, 36, 0, 30, 4, 27, 
    0, 0, 3, 8, 34, 38, 27, 22, 25, 32, 27, 20, 42, 0, 22, 
    0, 0, 0, 8, 30, 23, 26, 37, 46, 24, 15, 38, 25, 17, 13, 
    0, 0, 9, 10, 14, 15, 33, 44, 30, 34, 44, 26, 46, 36, 0, 
    0, 12, 0, 0, 12, 32, 23, 25, 39, 44, 29, 39, 40, 0, 0, 
    15, 0, 1, 1, 0, 0, 16, 39, 36, 41, 34, 39, 33, 2, 0, 
    0, 12, 16, 0, 12, 0, 22, 47, 40, 34, 32, 43, 47, 16, 0, 
    9, 39, 43, 20, 0, 7, 28, 59, 33, 36, 49, 39, 42, 9, 0, 
    8, 1, 28, 38, 32, 5, 5, 9, 0, 39, 35, 42, 48, 0, 0, 
    20, 0, 0, 29, 45, 26, 19, 10, 14, 35, 49, 34, 0, 0, 0, 
    
    -- channel=138
    3, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 14, 
    0, 14, 0, 0, 10, 0, 0, 4, 0, 0, 0, 0, 25, 2, 0, 
    0, 0, 0, 0, 17, 18, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 9, 25, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 
    0, 0, 7, 0, 9, 0, 6, 26, 0, 2, 0, 0, 0, 0, 0, 
    1, 0, 0, 31, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 14, 
    20, 0, 0, 0, 0, 11, 32, 4, 8, 6, 15, 4, 0, 0, 11, 
    1, 0, 0, 0, 21, 13, 12, 16, 20, 30, 17, 0, 17, 0, 0, 
    0, 0, 0, 0, 0, 43, 0, 8, 14, 11, 14, 0, 0, 0, 26, 
    0, 0, 0, 0, 0, 0, 17, 9, 3, 5, 13, 8, 18, 9, 0, 
    0, 0, 1, 0, 0, 12, 0, 0, 6, 0, 8, 13, 13, 0, 0, 
    18, 4, 20, 0, 0, 0, 0, 0, 0, 10, 10, 11, 13, 0, 0, 
    0, 0, 0, 1, 1, 0, 0, 0, 0, 12, 0, 20, 16, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 23, 0, 0, 10, 8, 11, 0, 0, 
    0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 39, 2, 0, 
    
    -- channel=139
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=140
    22, 4, 54, 31, 0, 70, 27, 36, 36, 31, 0, 78, 0, 49, 29, 
    18, 19, 19, 33, 0, 54, 16, 55, 21, 43, 0, 97, 0, 72, 23, 
    11, 15, 25, 11, 0, 64, 57, 27, 32, 0, 45, 93, 0, 36, 24, 
    0, 83, 16, 4, 19, 85, 26, 0, 84, 0, 83, 88, 1, 30, 0, 
    0, 99, 0, 0, 70, 39, 0, 75, 44, 62, 37, 46, 26, 27, 0, 
    0, 95, 24, 0, 81, 28, 5, 64, 37, 34, 18, 92, 11, 27, 0, 
    0, 73, 49, 13, 6, 26, 18, 35, 15, 24, 19, 46, 13, 52, 0, 
    0, 56, 47, 21, 15, 0, 34, 23, 14, 29, 28, 29, 3, 41, 0, 
    33, 51, 14, 16, 29, 0, 33, 10, 26, 18, 4, 32, 0, 3, 0, 
    33, 1, 3, 47, 19, 21, 15, 29, 11, 11, 9, 9, 0, 21, 50, 
    0, 57, 5, 46, 45, 16, 64, 14, 8, 0, 12, 6, 5, 24, 56, 
    31, 77, 15, 61, 2, 45, 45, 18, 10, 0, 29, 10, 0, 55, 19, 
    35, 41, 15, 37, 24, 49, 17, 0, 19, 8, 14, 0, 0, 36, 35, 
    0, 52, 69, 33, 29, 42, 33, 0, 56, 22, 16, 0, 0, 72, 36, 
    0, 20, 87, 80, 26, 38, 40, 44, 13, 17, 2, 0, 0, 42, 125, 
    
    -- channel=141
    12, 19, 0, 27, 44, 0, 14, 13, 17, 26, 32, 0, 37, 13, 14, 
    27, 16, 29, 26, 43, 3, 28, 5, 21, 11, 32, 0, 38, 0, 17, 
    25, 19, 25, 34, 36, 0, 0, 18, 28, 42, 11, 0, 29, 22, 21, 
    41, 0, 22, 16, 17, 0, 27, 54, 0, 21, 0, 0, 38, 22, 45, 
    33, 0, 36, 29, 0, 15, 49, 0, 14, 1, 13, 27, 26, 31, 64, 
    37, 3, 36, 32, 0, 9, 0, 0, 10, 16, 25, 0, 31, 32, 55, 
    23, 7, 30, 25, 7, 0, 0, 0, 1, 0, 0, 0, 26, 22, 54, 
    33, 16, 16, 29, 0, 16, 0, 0, 0, 0, 0, 0, 0, 19, 67, 
    18, 14, 41, 40, 20, 0, 0, 0, 0, 0, 1, 0, 25, 18, 28, 
    19, 43, 32, 13, 24, 27, 0, 0, 0, 0, 0, 0, 15, 16, 22, 
    48, 0, 27, 22, 21, 9, 0, 0, 0, 9, 0, 0, 2, 20, 11, 
    12, 0, 14, 15, 38, 22, 0, 0, 5, 8, 0, 0, 0, 0, 47, 
    29, 25, 15, 13, 22, 11, 12, 16, 2, 0, 0, 1, 1, 21, 35, 
    30, 23, 18, 13, 20, 16, 22, 21, 0, 0, 0, 5, 34, 0, 35, 
    36, 2, 7, 9, 15, 16, 25, 22, 18, 1, 6, 21, 14, 22, 0, 
    
    -- channel=142
    18, 18, 0, 0, 63, 0, 17, 0, 19, 0, 54, 0, 130, 0, 8, 
    3, 13, 20, 1, 61, 0, 9, 0, 15, 0, 50, 0, 102, 0, 26, 
    39, 1, 9, 18, 44, 0, 0, 28, 0, 63, 0, 0, 74, 7, 31, 
    43, 0, 43, 31, 0, 0, 51, 43, 0, 16, 0, 0, 44, 8, 102, 
    33, 0, 56, 46, 0, 7, 91, 0, 2, 0, 31, 0, 35, 13, 133, 
    53, 0, 0, 50, 0, 13, 29, 0, 23, 23, 43, 0, 53, 0, 134, 
    36, 0, 0, 19, 43, 21, 23, 37, 41, 15, 7, 23, 38, 0, 94, 
    33, 0, 0, 16, 6, 56, 9, 29, 18, 29, 45, 0, 70, 13, 98, 
    0, 0, 11, 3, 0, 30, 8, 17, 37, 38, 37, 21, 64, 25, 46, 
    13, 21, 36, 0, 1, 0, 8, 13, 27, 43, 29, 46, 69, 30, 0, 
    69, 0, 41, 0, 16, 9, 0, 30, 32, 53, 29, 41, 52, 0, 0, 
    0, 0, 64, 0, 20, 0, 0, 31, 27, 48, 24, 45, 56, 0, 8, 
    17, 0, 29, 48, 39, 0, 9, 74, 0, 21, 26, 56, 70, 0, 21, 
    64, 10, 0, 3, 61, 26, 22, 27, 0, 22, 17, 67, 91, 0, 0, 
    69, 24, 0, 0, 4, 39, 44, 32, 43, 20, 24, 25, 45, 10, 0, 
    
    -- channel=143
    29, 7, 7, 10, 32, 0, 15, 0, 0, 4, 27, 0, 60, 0, 0, 
    16, 0, 18, 15, 20, 0, 18, 0, 35, 0, 40, 0, 91, 0, 23, 
    0, 11, 10, 0, 12, 0, 2, 0, 18, 0, 39, 0, 67, 6, 32, 
    33, 13, 0, 13, 0, 2, 6, 15, 0, 41, 11, 0, 63, 22, 51, 
    9, 12, 66, 0, 0, 18, 38, 0, 33, 0, 6, 0, 29, 20, 68, 
    5, 0, 46, 40, 0, 0, 14, 31, 15, 10, 28, 0, 21, 32, 73, 
    19, 0, 0, 30, 10, 4, 12, 0, 0, 6, 11, 0, 35, 2, 67, 
    7, 4, 0, 21, 63, 0, 2, 5, 30, 0, 0, 23, 13, 14, 21, 
    17, 0, 0, 15, 0, 51, 0, 19, 0, 0, 12, 0, 8, 2, 44, 
    0, 5, 0, 0, 38, 0, 11, 11, 2, 18, 0, 10, 39, 1, 0, 
    25, 14, 14, 29, 0, 16, 0, 11, 22, 3, 2, 14, 14, 8, 20, 
    27, 39, 35, 0, 45, 0, 4, 16, 6, 15, 14, 6, 9, 0, 17, 
    0, 12, 58, 18, 4, 16, 6, 0, 0, 24, 14, 6, 19, 0, 5, 
    28, 0, 7, 50, 30, 4, 0, 38, 0, 6, 17, 0, 21, 0, 37, 
    39, 26, 0, 0, 53, 31, 24, 9, 0, 2, 3, 27, 13, 19, 0, 
    
    -- channel=144
    3, 0, 0, 0, 3, 0, 0, 0, 1, 0, 9, 0, 45, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 8, 0, 34, 0, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 30, 0, 1, 
    0, 0, 8, 2, 0, 0, 1, 1, 0, 0, 0, 0, 24, 0, 37, 
    0, 0, 6, 13, 0, 0, 20, 0, 0, 0, 2, 0, 18, 3, 39, 
    11, 0, 0, 0, 0, 16, 34, 0, 2, 10, 19, 0, 24, 0, 40, 
    1, 0, 0, 3, 34, 46, 41, 39, 42, 45, 36, 28, 28, 0, 26, 
    0, 0, 0, 7, 35, 50, 40, 54, 49, 44, 49, 41, 47, 7, 24, 
    0, 0, 1, 0, 29, 38, 46, 53, 53, 57, 57, 49, 59, 27, 1, 
    1, 3, 6, 0, 7, 37, 40, 45, 56, 60, 48, 57, 53, 8, 0, 
    17, 0, 2, 0, 0, 1, 24, 53, 55, 63, 51, 56, 46, 0, 0, 
    0, 0, 10, 0, 0, 0, 31, 61, 56, 52, 49, 63, 52, 12, 0, 
    14, 11, 14, 6, 1, 0, 31, 78, 39, 49, 60, 58, 60, 0, 0, 
    13, 8, 0, 9, 8, 0, 5, 13, 4, 56, 50, 67, 59, 0, 0, 
    19, 0, 0, 0, 14, 0, 0, 1, 32, 49, 57, 35, 9, 0, 0, 
    
    -- channel=145
    0, 0, 0, 0, 0, 4, 0, 7, 0, 11, 0, 19, 0, 14, 0, 
    0, 0, 0, 1, 0, 12, 9, 3, 0, 0, 0, 22, 0, 0, 0, 
    18, 16, 0, 12, 0, 0, 0, 0, 15, 3, 0, 19, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 4, 0, 0, 0, 3, 0, 0, 
    0, 18, 0, 0, 2, 0, 0, 0, 0, 0, 0, 13, 0, 10, 0, 
    0, 33, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 
    0, 12, 29, 0, 0, 7, 0, 6, 13, 15, 8, 6, 2, 4, 0, 
    0, 12, 12, 9, 0, 10, 16, 3, 0, 0, 5, 28, 0, 10, 0, 
    0, 0, 23, 19, 36, 0, 19, 17, 11, 21, 11, 20, 26, 29, 0, 
    8, 24, 7, 15, 15, 51, 15, 15, 20, 14, 18, 10, 4, 0, 0, 
    7, 8, 0, 5, 0, 0, 31, 21, 20, 25, 24, 12, 4, 3, 3, 
    0, 0, 0, 0, 2, 10, 23, 25, 28, 13, 11, 13, 0, 17, 4, 
    41, 54, 0, 0, 0, 15, 22, 36, 56, 18, 26, 9, 0, 29, 0, 
    0, 42, 47, 0, 0, 0, 0, 0, 2, 30, 21, 14, 13, 7, 0, 
    0, 0, 31, 34, 0, 0, 0, 0, 4, 33, 46, 20, 0, 0, 0, 
    
    -- channel=146
    0, 0, 0, 0, 0, 62, 0, 26, 11, 35, 0, 78, 0, 63, 0, 
    0, 0, 0, 1, 0, 54, 25, 28, 0, 3, 0, 94, 0, 8, 0, 
    5, 31, 0, 0, 0, 31, 0, 0, 44, 0, 58, 73, 0, 0, 0, 
    0, 50, 0, 0, 0, 24, 0, 0, 58, 0, 31, 32, 0, 0, 0, 
    0, 104, 0, 0, 44, 0, 0, 24, 0, 0, 0, 52, 0, 0, 0, 
    0, 122, 11, 0, 6, 0, 0, 12, 0, 0, 0, 33, 0, 20, 0, 
    0, 51, 49, 0, 0, 3, 0, 0, 0, 9, 0, 0, 0, 9, 0, 
    0, 43, 3, 7, 0, 0, 29, 0, 0, 0, 0, 34, 0, 6, 0, 
    0, 0, 2, 20, 51, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 47, 19, 85, 0, 0, 0, 0, 0, 0, 0, 0, 35, 
    0, 47, 0, 37, 0, 0, 82, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 29, 26, 8, 0, 0, 0, 0, 0, 19, 0, 
    55, 129, 0, 0, 0, 41, 21, 0, 85, 0, 0, 0, 0, 31, 2, 
    0, 86, 168, 3, 0, 0, 0, 0, 2, 17, 0, 0, 0, 52, 23, 
    0, 0, 115, 143, 4, 0, 0, 0, 0, 47, 43, 0, 0, 0, 72, 
    
    -- channel=147
    0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 3, 0, 22, 0, 
    0, 0, 0, 0, 0, 15, 14, 0, 0, 0, 0, 3, 0, 0, 0, 
    20, 25, 0, 0, 0, 0, 0, 0, 11, 2, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 13, 2, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 
    0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 5, 10, 26, 0, 0, 0, 0, 4, 0, 0, 25, 13, 0, 
    0, 13, 1, 16, 5, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 14, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    44, 74, 0, 0, 0, 0, 0, 34, 57, 0, 0, 0, 0, 23, 0, 
    0, 72, 88, 0, 0, 0, 0, 0, 0, 7, 0, 0, 16, 13, 0, 
    0, 0, 51, 60, 0, 0, 0, 0, 8, 32, 44, 17, 0, 0, 0, 
    
    -- channel=148
    7, 0, 17, 19, 0, 12, 9, 10, 24, 21, 10, 32, 0, 11, 12, 
    11, 8, 14, 23, 0, 9, 3, 20, 16, 21, 4, 42, 0, 26, 14, 
    25, 11, 20, 15, 0, 1, 16, 22, 18, 8, 19, 45, 21, 29, 35, 
    0, 30, 19, 0, 0, 34, 29, 0, 38, 0, 29, 53, 36, 37, 16, 
    5, 58, 11, 7, 19, 25, 0, 20, 16, 32, 31, 34, 38, 43, 0, 
    0, 59, 43, 0, 37, 17, 3, 25, 23, 23, 11, 47, 31, 41, 0, 
    0, 39, 51, 39, 8, 0, 0, 8, 11, 11, 4, 16, 25, 51, 0, 
    9, 39, 43, 45, 3, 0, 10, 16, 0, 0, 10, 29, 4, 44, 0, 
    23, 37, 35, 33, 43, 0, 18, 8, 11, 15, 12, 17, 16, 10, 0, 
    42, 17, 20, 41, 21, 45, 5, 22, 20, 14, 10, 12, 0, 15, 31, 
    5, 32, 10, 27, 35, 9, 49, 21, 22, 17, 7, 6, 0, 17, 48, 
    19, 32, 5, 40, 27, 37, 29, 25, 23, 9, 12, 11, 0, 33, 38, 
    47, 57, 27, 28, 19, 52, 27, 10, 22, 12, 20, 0, 1, 16, 49, 
    6, 36, 56, 40, 23, 26, 30, 2, 31, 20, 17, 5, 0, 40, 10, 
    3, 0, 41, 59, 43, 30, 33, 29, 30, 21, 18, 0, 0, 5, 72, 
    
    -- channel=149
    14, 22, 0, 0, 74, 0, 13, 0, 0, 0, 53, 0, 143, 0, 0, 
    0, 12, 18, 0, 75, 0, 0, 0, 12, 0, 51, 0, 128, 0, 25, 
    18, 0, 6, 8, 57, 0, 0, 20, 0, 50, 0, 0, 77, 0, 25, 
    45, 0, 33, 30, 0, 0, 38, 43, 0, 36, 0, 0, 39, 0, 100, 
    39, 0, 80, 32, 0, 0, 96, 0, 0, 0, 11, 0, 22, 5, 153, 
    59, 0, 0, 82, 0, 0, 28, 0, 11, 0, 24, 0, 48, 0, 165, 
    53, 0, 0, 15, 19, 0, 9, 0, 8, 0, 0, 0, 29, 0, 127, 
    31, 0, 0, 0, 4, 29, 0, 0, 4, 5, 10, 0, 58, 0, 109, 
    0, 0, 0, 0, 0, 46, 0, 0, 3, 0, 14, 0, 38, 10, 71, 
    0, 8, 31, 0, 0, 0, 0, 0, 0, 21, 4, 22, 65, 19, 0, 
    67, 0, 44, 0, 0, 13, 0, 6, 15, 23, 0, 16, 37, 0, 0, 
    0, 0, 74, 0, 23, 0, 0, 0, 4, 34, 0, 16, 37, 0, 2, 
    0, 0, 27, 43, 36, 0, 0, 41, 0, 4, 0, 37, 51, 0, 7, 
    55, 0, 0, 0, 56, 16, 0, 40, 0, 0, 0, 43, 89, 0, 0, 
    74, 26, 0, 0, 0, 37, 36, 10, 17, 0, 0, 17, 56, 0, 0, 
    
    -- channel=150
    10, 17, 26, 8, 4, 11, 6, 0, 0, 0, 0, 0, 0, 0, 12, 
    4, 22, 0, 6, 5, 0, 0, 12, 0, 2, 0, 0, 1, 38, 8, 
    0, 0, 0, 0, 1, 28, 34, 3, 0, 0, 0, 0, 0, 6, 2, 
    0, 30, 14, 2, 18, 16, 0, 0, 17, 0, 15, 0, 0, 0, 0, 
    8, 0, 11, 0, 1, 0, 0, 40, 1, 15, 0, 0, 0, 0, 0, 
    0, 0, 0, 42, 27, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 11, 4, 0, 3, 0, 0, 
    4, 12, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 3, 
    0, 0, 1, 0, 14, 4, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    23, 47, 21, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 
    0, 15, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 34, 26, 4, 
    
    -- channel=151
    18, 26, 22, 0, 10, 0, 9, 0, 0, 0, 0, 0, 31, 0, 8, 
    10, 33, 2, 0, 14, 0, 0, 0, 2, 2, 0, 0, 47, 41, 22, 
    0, 0, 0, 0, 6, 18, 42, 6, 0, 0, 0, 0, 27, 11, 11, 
    0, 18, 24, 7, 16, 16, 0, 0, 0, 20, 16, 0, 0, 2, 0, 
    15, 0, 43, 8, 0, 2, 16, 30, 19, 28, 0, 0, 0, 0, 7, 
    0, 0, 0, 81, 24, 0, 12, 15, 13, 0, 0, 5, 0, 0, 36, 
    37, 0, 0, 1, 0, 0, 22, 11, 0, 0, 11, 14, 0, 0, 30, 
    0, 0, 2, 0, 34, 22, 0, 7, 24, 52, 31, 0, 44, 0, 0, 
    11, 16, 0, 0, 0, 49, 7, 3, 22, 0, 0, 6, 0, 0, 24, 
    2, 0, 0, 0, 0, 0, 15, 24, 4, 15, 3, 5, 8, 11, 0, 
    0, 0, 15, 0, 14, 21, 0, 9, 10, 0, 0, 0, 10, 2, 12, 
    42, 89, 69, 11, 0, 0, 0, 0, 0, 12, 17, 5, 0, 0, 0, 
    0, 0, 3, 37, 21, 0, 0, 0, 0, 4, 0, 13, 9, 0, 0, 
    0, 0, 0, 0, 40, 17, 0, 30, 33, 0, 0, 1, 0, 0, 0, 
    1, 21, 0, 0, 0, 46, 31, 2, 0, 0, 0, 0, 63, 34, 0, 
    
    -- channel=152
    38, 19, 13, 18, 51, 0, 29, 0, 24, 9, 56, 0, 114, 0, 15, 
    34, 28, 33, 26, 47, 0, 4, 0, 41, 15, 55, 0, 117, 7, 53, 
    38, 18, 28, 26, 32, 0, 12, 36, 5, 40, 11, 0, 111, 39, 71, 
    40, 0, 50, 39, 0, 5, 46, 12, 0, 46, 6, 1, 90, 60, 108, 
    45, 0, 104, 33, 0, 42, 69, 0, 34, 21, 49, 0, 68, 62, 121, 
    50, 0, 64, 84, 13, 35, 60, 49, 58, 45, 49, 3, 77, 51, 128, 
    57, 3, 19, 84, 67, 39, 49, 40, 47, 47, 52, 44, 66, 43, 107, 
    43, 11, 34, 69, 81, 33, 30, 60, 65, 53, 49, 53, 99, 53, 73, 
    34, 38, 41, 40, 25, 109, 42, 65, 62, 55, 65, 53, 78, 45, 71, 
    53, 38, 43, 26, 44, 12, 68, 74, 70, 88, 60, 72, 80, 37, 3, 
    75, 15, 55, 16, 24, 55, 19, 86, 93, 76, 60, 65, 65, 31, 56, 
    44, 78, 85, 16, 67, 20, 53, 76, 74, 89, 66, 71, 61, 26, 45, 
    26, 15, 95, 74, 54, 39, 55, 71, 17, 78, 70, 75, 77, 0, 45, 
    62, 0, 0, 71, 85, 41, 32, 55, 11, 60, 71, 76, 65, 0, 10, 
    71, 24, 0, 0, 80, 86, 68, 39, 49, 43, 50, 41, 50, 17, 0, 
    
    -- channel=153
    0, 0, 0, 0, 12, 0, 0, 0, 8, 15, 8, 0, 11, 8, 0, 
    0, 0, 0, 0, 8, 7, 16, 0, 0, 0, 6, 0, 0, 0, 0, 
    28, 17, 0, 11, 4, 0, 0, 0, 8, 27, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 10, 32, 0, 0, 0, 0, 14, 0, 26, 
    0, 0, 0, 7, 0, 0, 5, 0, 0, 0, 0, 9, 0, 0, 36, 
    9, 2, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 3, 2, 12, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 
    0, 0, 19, 16, 19, 0, 0, 0, 0, 0, 0, 0, 29, 25, 0, 
    0, 28, 12, 5, 5, 46, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    24, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 1, 0, 6, 
    46, 49, 0, 0, 0, 0, 5, 49, 30, 0, 0, 0, 0, 18, 12, 
    13, 63, 54, 0, 0, 0, 0, 0, 0, 2, 0, 5, 42, 0, 0, 
    14, 0, 35, 33, 0, 0, 0, 0, 11, 22, 44, 11, 0, 0, 0, 
    
    -- channel=154
    26, 28, 23, 19, 41, 0, 28, 7, 30, 12, 45, 0, 92, 0, 19, 
    24, 39, 34, 19, 42, 0, 4, 5, 28, 24, 42, 0, 82, 14, 42, 
    26, 8, 20, 22, 31, 0, 32, 44, 0, 41, 1, 0, 72, 35, 43, 
    33, 0, 46, 29, 11, 29, 58, 23, 0, 29, 19, 20, 49, 33, 62, 
    41, 0, 60, 37, 1, 38, 62, 6, 39, 32, 57, 8, 49, 30, 78, 
    43, 0, 25, 67, 37, 20, 41, 23, 52, 37, 43, 14, 63, 18, 87, 
    48, 3, 9, 39, 41, 19, 36, 31, 30, 18, 20, 35, 46, 28, 73, 
    35, 4, 23, 25, 25, 45, 8, 31, 31, 39, 42, 4, 66, 31, 59, 
    22, 33, 27, 19, 4, 41, 19, 23, 34, 25, 35, 31, 35, 32, 46, 
    35, 25, 35, 10, 9, 0, 21, 25, 30, 38, 30, 37, 47, 29, 7, 
    49, 6, 50, 6, 37, 25, 0, 36, 32, 36, 22, 33, 48, 23, 38, 
    22, 56, 91, 36, 36, 10, 13, 26, 26, 41, 24, 36, 49, 23, 39, 
    13, 0, 64, 83, 59, 15, 17, 38, 0, 25, 26, 42, 47, 16, 42, 
    46, 0, 0, 46, 91, 61, 39, 46, 15, 18, 22, 48, 50, 14, 8, 
    56, 30, 0, 0, 47, 81, 77, 53, 38, 8, 10, 18, 56, 30, 14, 
    
    -- channel=155
    0, 27, 0, 0, 9, 0, 0, 14, 0, 1, 0, 9, 0, 0, 3, 
    0, 41, 0, 0, 41, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 
    9, 11, 0, 10, 52, 0, 0, 0, 0, 23, 0, 3, 0, 0, 0, 
    0, 0, 0, 6, 46, 0, 0, 36, 0, 29, 0, 3, 0, 0, 0, 
    26, 0, 0, 20, 0, 0, 0, 1, 0, 0, 0, 27, 0, 0, 0, 
    49, 0, 0, 36, 0, 1, 24, 0, 0, 0, 0, 12, 0, 0, 2, 
    40, 0, 0, 1, 16, 4, 8, 0, 2, 3, 12, 0, 0, 0, 22, 
    25, 0, 5, 0, 0, 62, 0, 0, 1, 0, 9, 0, 4, 0, 55, 
    0, 0, 17, 0, 7, 16, 3, 4, 0, 0, 11, 10, 6, 15, 26, 
    0, 20, 27, 0, 0, 0, 15, 0, 8, 0, 21, 0, 0, 0, 0, 
    13, 0, 10, 0, 7, 20, 0, 0, 0, 4, 5, 0, 0, 4, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 2, 10, 0, 0, 
    3, 0, 0, 0, 3, 0, 0, 13, 12, 0, 0, 16, 0, 30, 0, 
    0, 14, 0, 0, 0, 0, 0, 0, 14, 0, 2, 21, 26, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 6, 16, 18, 0, 0, 
    
    -- channel=156
    47, 22, 26, 36, 57, 0, 45, 19, 56, 44, 72, 1, 120, 3, 21, 
    48, 34, 53, 43, 49, 0, 25, 3, 61, 39, 74, 0, 118, 16, 68, 
    58, 46, 40, 41, 35, 0, 26, 58, 38, 53, 38, 3, 122, 60, 86, 
    53, 10, 55, 45, 0, 40, 83, 35, 0, 52, 33, 32, 119, 78, 119, 
    55, 33, 108, 42, 17, 75, 79, 0, 65, 45, 87, 48, 93, 81, 124, 
    57, 28, 91, 80, 40, 52, 57, 73, 84, 72, 74, 29, 101, 79, 122, 
    56, 30, 52, 104, 82, 53, 48, 47, 53, 54, 57, 54, 83, 69, 109, 
    57, 35, 51, 90, 86, 31, 43, 63, 71, 48, 43, 62, 94, 72, 81, 
    48, 57, 67, 71, 52, 96, 48, 69, 63, 60, 69, 57, 88, 71, 73, 
    70, 67, 57, 53, 67, 41, 71, 72, 73, 89, 63, 75, 79, 39, 24, 
    91, 37, 66, 46, 44, 65, 37, 91, 89, 79, 66, 68, 66, 43, 79, 
    50, 88, 94, 39, 90, 42, 71, 84, 77, 86, 70, 72, 77, 44, 84, 
    66, 75, 131, 98, 75, 65, 82, 87, 43, 78, 77, 74, 76, 13, 83, 
    78, 6, 53, 113, 113, 73, 65, 66, 21, 71, 74, 76, 74, 20, 52, 
    90, 37, 0, 60, 122, 117, 102, 75, 63, 63, 75, 58, 44, 36, 31, 
    
    -- channel=157
    12, 6, 14, 33, 20, 20, 15, 22, 22, 27, 21, 26, 3, 19, 14, 
    21, 8, 22, 33, 16, 16, 24, 18, 18, 19, 21, 24, 2, 7, 17, 
    28, 29, 27, 30, 13, 11, 10, 20, 37, 18, 30, 20, 12, 24, 28, 
    20, 18, 12, 16, 8, 16, 26, 20, 21, 12, 11, 17, 32, 27, 24, 
    20, 40, 19, 9, 15, 19, 7, 9, 14, 12, 20, 27, 24, 32, 22, 
    16, 43, 45, 7, 12, 11, 0, 13, 15, 14, 11, 12, 18, 43, 9, 
    7, 27, 41, 33, 1, 0, 0, 0, 0, 0, 0, 0, 12, 34, 16, 
    23, 31, 29, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 18, 
    22, 23, 35, 38, 21, 0, 0, 0, 0, 0, 0, 0, 10, 17, 16, 
    28, 34, 25, 35, 21, 19, 0, 0, 0, 0, 0, 0, 0, 8, 28, 
    26, 23, 17, 31, 24, 13, 11, 0, 0, 0, 0, 0, 0, 18, 30, 
    17, 0, 0, 21, 32, 27, 5, 0, 0, 0, 0, 0, 0, 11, 47, 
    37, 45, 12, 6, 15, 27, 15, 0, 14, 0, 0, 0, 0, 17, 44, 
    17, 25, 48, 19, 5, 13, 14, 2, 0, 0, 0, 0, 0, 25, 43, 
    19, 5, 22, 39, 20, 8, 12, 17, 5, 7, 5, 1, 0, 11, 16, 
    
    -- channel=158
    0, 0, 0, 0, 0, 0, 0, 0, 17, 25, 3, 7, 0, 13, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 3, 14, 0, 0, 0, 
    20, 18, 0, 0, 0, 0, 0, 0, 18, 0, 22, 14, 16, 2, 7, 
    0, 0, 0, 0, 0, 0, 22, 2, 7, 0, 7, 25, 55, 13, 21, 
    0, 37, 0, 0, 0, 10, 0, 0, 0, 0, 26, 46, 43, 23, 1, 
    0, 52, 31, 0, 6, 28, 0, 0, 2, 28, 24, 5, 36, 38, 0, 
    0, 17, 42, 21, 12, 16, 0, 17, 27, 17, 0, 7, 30, 23, 0, 
    0, 22, 10, 39, 3, 0, 32, 18, 0, 0, 7, 35, 0, 31, 0, 
    0, 1, 28, 39, 56, 0, 14, 19, 18, 43, 28, 20, 46, 23, 0, 
    7, 29, 7, 31, 31, 72, 6, 14, 28, 25, 18, 25, 6, 0, 2, 
    15, 16, 0, 14, 0, 0, 56, 34, 26, 38, 29, 28, 7, 0, 5, 
    0, 0, 0, 11, 20, 25, 39, 54, 38, 12, 22, 22, 19, 15, 32, 
    69, 117, 36, 6, 10, 33, 43, 52, 69, 23, 37, 13, 7, 17, 33, 
    6, 61, 126, 55, 10, 18, 43, 1, 0, 45, 30, 22, 11, 7, 25, 
    1, 0, 49, 112, 60, 9, 16, 41, 34, 49, 56, 26, 0, 0, 38, 
    
    -- channel=159
    14, 27, 15, 21, 23, 7, 8, 9, 5, 12, 19, 9, 19, 17, 27, 
    23, 28, 19, 16, 23, 2, 18, 22, 13, 13, 17, 9, 34, 14, 16, 
    0, 5, 19, 10, 26, 32, 33, 6, 11, 24, 13, 13, 13, 26, 3, 
    33, 34, 20, 18, 35, 20, 20, 40, 20, 27, 21, 29, 3, 10, 3, 
    21, 0, 32, 12, 0, 11, 43, 29, 21, 27, 10, 15, 13, 9, 19, 
    13, 0, 4, 56, 31, 14, 0, 0, 8, 13, 14, 11, 15, 6, 23, 
    28, 9, 6, 2, 0, 0, 5, 11, 0, 0, 0, 5, 8, 13, 21, 
    25, 17, 22, 1, 0, 17, 1, 0, 0, 17, 10, 0, 2, 2, 39, 
    17, 15, 4, 9, 0, 0, 0, 0, 3, 7, 0, 0, 0, 0, 30, 
    0, 11, 24, 0, 17, 0, 0, 0, 0, 0, 0, 0, 10, 28, 21, 
    20, 8, 20, 13, 19, 27, 0, 0, 0, 0, 0, 0, 0, 12, 6, 
    32, 14, 49, 33, 13, 10, 0, 0, 0, 0, 0, 0, 0, 0, 27, 
    0, 0, 13, 35, 41, 0, 0, 0, 0, 0, 0, 0, 0, 16, 16, 
    20, 2, 0, 11, 36, 48, 37, 40, 19, 0, 0, 0, 6, 1, 46, 
    6, 29, 0, 0, 0, 37, 46, 52, 9, 0, 0, 10, 50, 57, 20, 
    
    -- channel=160
    50, 63, 56, 61, 60, 58, 54, 55, 36, 24, 25, 24, 29, 36, 26, 
    79, 70, 66, 66, 67, 67, 58, 59, 40, 19, 27, 30, 39, 32, 32, 
    56, 76, 70, 72, 74, 70, 65, 65, 65, 48, 45, 31, 31, 36, 37, 
    66, 66, 73, 77, 80, 76, 68, 62, 64, 67, 55, 36, 25, 35, 38, 
    52, 75, 76, 77, 80, 67, 55, 60, 44, 62, 66, 32, 36, 33, 36, 
    73, 58, 79, 75, 63, 93, 55, 56, 46, 51, 39, 16, 23, 30, 37, 
    56, 87, 77, 72, 78, 87, 74, 53, 54, 61, 29, 10, 18, 30, 28, 
    34, 79, 75, 70, 93, 82, 76, 91, 80, 73, 41, 14, 23, 42, 14, 
    47, 75, 75, 56, 90, 87, 64, 73, 74, 54, 17, 8, 32, 64, 15, 
    38, 79, 82, 20, 57, 73, 45, 69, 28, 15, 12, 6, 29, 78, 17, 
    49, 71, 73, 4, 19, 25, 26, 44, 16, 6, 7, 12, 26, 74, 40, 
    47, 59, 61, 57, 25, 36, 35, 5, 0, 0, 0, 0, 25, 42, 62, 
    57, 54, 61, 64, 55, 35, 45, 30, 17, 5, 0, 7, 14, 19, 44, 
    44, 59, 49, 56, 40, 48, 54, 41, 42, 34, 34, 41, 34, 40, 24, 
    52, 57, 51, 55, 53, 51, 52, 44, 44, 42, 46, 52, 47, 37, 47, 
    
    -- channel=161
    45, 53, 32, 33, 32, 32, 35, 34, 25, 25, 22, 24, 24, 24, 24, 
    35, 32, 37, 33, 35, 37, 37, 37, 33, 27, 19, 22, 23, 21, 25, 
    27, 29, 35, 34, 34, 36, 34, 35, 41, 47, 41, 31, 16, 21, 25, 
    26, 30, 32, 35, 33, 33, 29, 34, 30, 31, 32, 26, 20, 20, 19, 
    30, 30, 33, 32, 34, 29, 23, 27, 25, 20, 29, 23, 23, 21, 20, 
    27, 25, 28, 31, 29, 39, 28, 11, 18, 22, 15, 13, 21, 23, 19, 
    27, 24, 23, 24, 37, 24, 24, 32, 35, 26, 19, 21, 24, 23, 17, 
    19, 24, 21, 25, 31, 32, 36, 22, 21, 22, 22, 22, 28, 32, 24, 
    22, 26, 22, 25, 4, 14, 13, 1, 5, 0, 0, 13, 28, 19, 19, 
    14, 21, 17, 6, 8, 17, 13, 38, 17, 17, 25, 27, 29, 25, 15, 
    16, 17, 6, 13, 13, 0, 0, 0, 5, 19, 11, 20, 29, 20, 11, 
    17, 15, 20, 39, 41, 45, 37, 14, 18, 21, 20, 13, 17, 15, 13, 
    23, 15, 16, 23, 38, 20, 18, 32, 37, 35, 33, 34, 25, 20, 0, 
    8, 13, 17, 20, 21, 19, 17, 18, 29, 35, 38, 41, 41, 36, 24, 
    18, 21, 19, 26, 30, 20, 17, 17, 20, 18, 24, 24, 25, 24, 31, 
    
    -- channel=162
    16, 29, 43, 47, 40, 42, 35, 33, 0, 4, 8, 0, 0, 20, 0, 
    38, 36, 42, 45, 53, 46, 44, 48, 18, 0, 9, 19, 26, 17, 13, 
    33, 36, 44, 55, 55, 55, 46, 55, 49, 0, 24, 17, 27, 27, 21, 
    14, 46, 48, 57, 54, 61, 58, 50, 59, 52, 39, 13, 18, 21, 24, 
    40, 39, 47, 51, 54, 61, 43, 40, 30, 59, 50, 4, 14, 24, 24, 
    36, 39, 45, 55, 51, 58, 25, 42, 14, 43, 31, 0, 12, 12, 21, 
    40, 57, 50, 40, 41, 53, 26, 5, 23, 23, 3, 0, 0, 5, 16, 
    15, 71, 43, 51, 53, 45, 51, 57, 42, 36, 0, 0, 0, 21, 1, 
    35, 68, 44, 28, 41, 47, 34, 47, 41, 40, 0, 0, 2, 37, 0, 
    38, 73, 42, 0, 70, 54, 19, 62, 20, 0, 0, 0, 15, 60, 0, 
    42, 66, 36, 0, 0, 6, 8, 47, 10, 0, 0, 0, 9, 77, 0, 
    50, 47, 45, 0, 17, 7, 19, 8, 0, 0, 0, 0, 2, 37, 31, 
    50, 56, 33, 61, 18, 31, 36, 13, 0, 0, 0, 0, 0, 0, 20, 
    42, 59, 40, 34, 24, 22, 54, 31, 21, 13, 4, 14, 3, 15, 23, 
    41, 50, 42, 49, 32, 46, 49, 47, 39, 29, 42, 48, 39, 27, 30, 
    
    -- channel=163
    28, 10, 24, 21, 27, 26, 26, 16, 27, 11, 10, 13, 9, 5, 12, 
    24, 33, 23, 26, 28, 27, 27, 21, 33, 20, 8, 10, 3, 13, 11, 
    40, 28, 25, 29, 29, 33, 33, 28, 25, 14, 1, 9, 11, 13, 9, 
    25, 25, 29, 27, 30, 28, 32, 29, 24, 23, 23, 32, 18, 12, 13, 
    21, 22, 26, 30, 32, 34, 28, 22, 31, 21, 23, 40, 10, 14, 12, 
    0, 28, 30, 31, 37, 21, 25, 30, 22, 14, 29, 35, 10, 14, 10, 
    0, 11, 29, 30, 19, 26, 26, 15, 8, 11, 28, 20, 8, 12, 13, 
    16, 0, 27, 25, 12, 24, 18, 15, 17, 18, 30, 17, 0, 4, 22, 
    14, 0, 22, 29, 25, 21, 39, 29, 26, 34, 46, 19, 0, 2, 33, 
    23, 6, 19, 52, 11, 9, 34, 0, 29, 23, 5, 6, 0, 0, 39, 
    20, 6, 26, 48, 7, 35, 24, 24, 40, 17, 16, 7, 1, 0, 39, 
    17, 10, 20, 11, 11, 0, 0, 24, 25, 14, 11, 10, 3, 10, 19, 
    9, 16, 18, 22, 20, 14, 7, 14, 3, 1, 5, 0, 4, 9, 18, 
    23, 7, 23, 10, 29, 9, 7, 19, 8, 2, 0, 0, 0, 0, 15, 
    14, 5, 14, 7, 6, 12, 19, 18, 16, 12, 9, 11, 14, 19, 5, 
    
    -- channel=164
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=165
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 2, 0, 
    0, 0, 0, 0, 3, 0, 0, 36, 19, 0, 4, 22, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 
    0, 0, 0, 14, 19, 6, 12, 55, 44, 75, 84, 17, 0, 0, 0, 
    0, 0, 0, 29, 43, 22, 22, 0, 0, 17, 0, 0, 0, 0, 0, 
    0, 1, 19, 21, 0, 63, 41, 46, 50, 21, 28, 1, 0, 7, 0, 
    2, 0, 0, 0, 0, 0, 0, 7, 9, 4, 3, 21, 1, 32, 2, 
    0, 0, 0, 9, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 1, 2, 5, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=166
    37, 43, 25, 29, 26, 20, 12, 7, 16, 0, 6, 10, 2, 11, 16, 
    43, 47, 22, 30, 30, 29, 25, 19, 16, 0, 0, 4, 15, 20, 5, 
    56, 37, 34, 30, 35, 31, 32, 12, 23, 39, 21, 20, 11, 6, 18, 
    33, 41, 35, 31, 39, 29, 30, 23, 22, 26, 18, 25, 6, 4, 13, 
    26, 37, 41, 32, 36, 37, 45, 51, 38, 13, 22, 44, 4, 10, 14, 
    0, 45, 43, 48, 32, 40, 91, 39, 36, 27, 34, 10, 0, 5, 9, 
    7, 21, 64, 59, 35, 69, 40, 67, 64, 63, 48, 12, 0, 6, 9, 
    24, 10, 64, 38, 62, 79, 62, 63, 71, 74, 76, 19, 0, 30, 27, 
    29, 27, 69, 44, 63, 24, 69, 21, 26, 21, 8, 0, 0, 23, 58, 
    31, 13, 76, 78, 0, 50, 46, 51, 51, 0, 3, 14, 0, 19, 99, 
    44, 12, 58, 41, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 85, 
    21, 34, 31, 60, 30, 19, 24, 17, 0, 0, 0, 0, 0, 0, 23, 
    28, 27, 32, 19, 55, 37, 20, 30, 18, 7, 0, 0, 0, 0, 5, 
    35, 9, 38, 15, 29, 23, 25, 33, 19, 29, 18, 26, 26, 20, 19, 
    19, 39, 32, 30, 37, 40, 24, 19, 21, 11, 20, 25, 30, 29, 14, 
    
    -- channel=167
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=168
    0, 8, 8, 14, 7, 9, 3, 12, 0, 5, 9, 5, 11, 19, 1, 
    15, 1, 12, 12, 11, 10, 4, 11, 0, 0, 15, 12, 16, 9, 11, 
    0, 13, 13, 15, 15, 10, 5, 17, 4, 0, 11, 5, 18, 14, 13, 
    7, 12, 13, 19, 14, 16, 13, 11, 17, 13, 14, 0, 8, 20, 18, 
    11, 20, 14, 17, 15, 14, 15, 18, 8, 29, 22, 0, 13, 11, 15, 
    54, 14, 25, 15, 11, 25, 0, 14, 0, 24, 12, 0, 10, 9, 17, 
    46, 37, 15, 11, 24, 21, 11, 0, 17, 19, 0, 0, 9, 8, 12, 
    8, 54, 15, 20, 33, 11, 17, 29, 21, 14, 0, 0, 12, 12, 0, 
    15, 50, 21, 11, 27, 41, 9, 25, 25, 19, 0, 0, 26, 34, 0, 
    15, 57, 25, 0, 38, 32, 0, 21, 0, 1, 0, 0, 22, 47, 0, 
    17, 48, 22, 0, 22, 25, 17, 46, 0, 0, 3, 3, 18, 55, 0, 
    21, 34, 22, 0, 0, 5, 12, 0, 0, 0, 0, 5, 21, 34, 14, 
    31, 28, 29, 26, 0, 6, 26, 0, 0, 0, 0, 0, 10, 12, 31, 
    23, 43, 13, 30, 1, 20, 34, 12, 13, 4, 2, 7, 0, 12, 0, 
    24, 34, 22, 27, 18, 21, 25, 19, 18, 22, 23, 23, 17, 7, 21, 
    
    -- channel=169
    63, 34, 67, 64, 71, 67, 68, 50, 46, 24, 27, 21, 15, 23, 30, 
    55, 72, 62, 67, 75, 71, 74, 69, 66, 19, 20, 36, 40, 41, 31, 
    67, 57, 62, 74, 73, 80, 78, 69, 81, 40, 30, 39, 42, 46, 36, 
    49, 63, 69, 71, 76, 85, 86, 76, 74, 77, 60, 48, 40, 28, 38, 
    54, 51, 67, 69, 74, 81, 60, 53, 52, 65, 64, 66, 29, 42, 40, 
    4, 56, 52, 73, 76, 56, 47, 61, 61, 45, 52, 45, 23, 32, 34, 
    0, 55, 71, 64, 43, 57, 60, 38, 18, 24, 44, 20, 5, 24, 33, 
    43, 33, 67, 63, 45, 66, 64, 62, 54, 55, 43, 23, 7, 28, 31, 
    59, 38, 57, 50, 55, 44, 68, 72, 65, 67, 70, 14, 0, 27, 33, 
    63, 36, 50, 58, 55, 52, 77, 65, 63, 30, 1, 16, 7, 32, 46, 
    66, 48, 56, 70, 0, 15, 31, 44, 64, 15, 7, 22, 9, 36, 68, 
    70, 49, 55, 29, 51, 25, 30, 50, 0, 0, 0, 0, 5, 24, 63, 
    52, 68, 39, 67, 49, 58, 43, 47, 17, 0, 0, 0, 1, 7, 19, 
    59, 49, 72, 37, 61, 37, 50, 63, 39, 35, 30, 28, 28, 24, 56, 
    56, 45, 61, 54, 46, 59, 62, 67, 56, 45, 51, 57, 56, 55, 34, 
    
    -- channel=170
    62, 46, 49, 53, 56, 53, 57, 44, 41, 30, 36, 42, 42, 30, 40, 
    41, 44, 56, 51, 55, 63, 66, 61, 67, 41, 28, 30, 33, 40, 39, 
    33, 38, 52, 52, 54, 57, 67, 59, 62, 66, 44, 49, 36, 38, 41, 
    39, 23, 46, 50, 45, 61, 56, 60, 46, 53, 58, 59, 43, 44, 38, 
    20, 39, 46, 50, 55, 56, 53, 59, 49, 46, 49, 45, 33, 31, 36, 
    30, 42, 50, 45, 45, 42, 19, 0, 35, 37, 37, 38, 22, 35, 33, 
    4, 26, 24, 36, 47, 5, 25, 55, 38, 28, 35, 38, 26, 38, 32, 
    38, 12, 27, 20, 22, 27, 42, 13, 4, 13, 40, 28, 20, 38, 37, 
    53, 20, 29, 26, 0, 24, 32, 3, 6, 0, 8, 31, 20, 19, 49, 
    55, 19, 11, 41, 0, 5, 36, 37, 39, 34, 44, 34, 17, 11, 42, 
    48, 18, 1, 43, 28, 0, 27, 13, 39, 33, 15, 27, 32, 0, 23, 
    43, 38, 18, 64, 39, 52, 43, 35, 37, 25, 20, 12, 25, 7, 15, 
    54, 42, 33, 11, 53, 38, 54, 58, 48, 41, 35, 32, 17, 41, 11, 
    43, 33, 37, 36, 33, 46, 33, 57, 50, 41, 49, 43, 51, 41, 24, 
    51, 46, 54, 47, 52, 41, 45, 42, 43, 52, 50, 46, 49, 49, 48, 
    
    -- channel=171
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=172
    0, 57, 11, 21, 12, 18, 9, 28, 0, 11, 10, 11, 16, 31, 0, 
    19, 5, 14, 18, 21, 18, 10, 22, 0, 7, 20, 9, 19, 7, 8, 
    0, 25, 20, 19, 21, 12, 9, 21, 13, 7, 42, 6, 13, 6, 15, 
    0, 24, 16, 26, 16, 14, 5, 12, 19, 11, 12, 0, 2, 22, 13, 
    5, 27, 19, 22, 17, 16, 1, 20, 0, 22, 16, 0, 18, 10, 11, 
    58, 8, 33, 19, 5, 48, 0, 0, 0, 28, 0, 0, 23, 11, 18, 
    98, 29, 8, 7, 26, 39, 0, 3, 47, 33, 0, 0, 19, 19, 13, 
    5, 77, 1, 10, 46, 0, 17, 35, 11, 7, 0, 0, 20, 37, 0, 
    3, 69, 9, 0, 41, 12, 0, 6, 5, 0, 0, 0, 50, 54, 0, 
    0, 73, 11, 0, 45, 29, 0, 47, 0, 0, 0, 13, 45, 80, 0, 
    0, 45, 5, 0, 50, 3, 0, 26, 0, 0, 2, 2, 36, 78, 0, 
    0, 29, 13, 0, 0, 26, 35, 0, 0, 4, 4, 20, 24, 35, 4, 
    17, 6, 22, 11, 0, 0, 11, 0, 6, 15, 12, 30, 42, 2, 40, 
    2, 18, 0, 23, 0, 20, 30, 0, 12, 12, 16, 40, 21, 37, 0, 
    4, 35, 0, 21, 9, 14, 12, 0, 5, 0, 18, 19, 8, 0, 25, 
    
    -- channel=173
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 5, 0, 0, 2, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 15, 
    0, 0, 0, 30, 0, 21, 0, 0, 6, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 7, 8, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=174
    67, 26, 51, 46, 60, 59, 59, 37, 73, 24, 27, 40, 31, 18, 46, 
    44, 63, 46, 54, 54, 58, 67, 50, 83, 50, 16, 27, 21, 47, 31, 
    80, 39, 50, 51, 52, 62, 74, 51, 52, 60, 19, 46, 40, 32, 31, 
    56, 39, 52, 42, 59, 59, 70, 59, 44, 52, 58, 81, 42, 31, 35, 
    25, 37, 50, 53, 57, 59, 51, 48, 76, 34, 43, 100, 19, 32, 31, 
    0, 58, 49, 55, 64, 1, 63, 50, 51, 17, 66, 85, 13, 31, 26, 
    0, 0, 57, 58, 21, 45, 50, 49, 19, 32, 80, 56, 15, 30, 35, 
    60, 0, 58, 35, 4, 49, 51, 24, 34, 36, 98, 56, 0, 5, 71, 
    56, 0, 46, 68, 31, 17, 101, 53, 43, 61, 96, 46, 0, 0, 113, 
    71, 0, 33, 158, 0, 12, 90, 0, 108, 47, 27, 40, 0, 0, 138, 
    70, 1, 51, 130, 25, 42, 36, 41, 78, 42, 29, 9, 7, 0, 110, 
    48, 42, 21, 60, 54, 16, 23, 74, 52, 26, 24, 12, 0, 11, 20, 
    36, 45, 55, 9, 61, 45, 28, 65, 43, 28, 34, 8, 7, 18, 37, 
    67, 10, 69, 32, 59, 39, 25, 72, 35, 38, 29, 18, 34, 25, 38, 
    41, 35, 53, 34, 36, 52, 54, 46, 49, 46, 35, 33, 50, 60, 20, 
    
    -- channel=175
    19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 5, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 
    0, 5, 0, 0, 0, 0, 0, 0, 4, 12, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 16, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 13, 0, 24, 0, 0, 1, 0, 0, 0, 
    0, 0, 1, 8, 0, 0, 10, 41, 9, 0, 5, 0, 0, 0, 0, 
    0, 0, 9, 0, 0, 21, 0, 9, 8, 27, 23, 0, 0, 18, 0, 
    1, 0, 7, 0, 16, 0, 0, 0, 0, 0, 23, 0, 0, 0, 17, 
    0, 0, 15, 18, 9, 0, 26, 50, 0, 0, 0, 6, 0, 0, 63, 
    0, 0, 3, 62, 0, 0, 0, 0, 15, 0, 0, 17, 0, 0, 81, 
    0, 0, 11, 22, 3, 10, 0, 2, 0, 0, 2, 0, 0, 0, 50, 
    0, 0, 0, 8, 0, 3, 0, 8, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 27, 0, 0, 7, 0, 5, 9, 5, 3, 0, 28, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    
    -- channel=176
    79, 59, 93, 94, 96, 97, 95, 76, 72, 51, 55, 53, 47, 55, 60, 
    81, 91, 90, 92, 100, 100, 106, 100, 93, 56, 49, 64, 65, 71, 60, 
    91, 76, 90, 98, 100, 105, 109, 101, 102, 68, 57, 73, 76, 73, 67, 
    69, 76, 94, 94, 103, 111, 116, 103, 101, 100, 89, 91, 71, 66, 71, 
    68, 76, 90, 95, 101, 110, 92, 86, 93, 98, 92, 95, 58, 69, 69, 
    24, 80, 83, 98, 97, 70, 73, 83, 76, 72, 88, 73, 47, 60, 65, 
    30, 68, 88, 87, 64, 82, 72, 60, 43, 53, 75, 53, 32, 53, 65, 
    73, 51, 88, 76, 61, 80, 90, 77, 66, 65, 78, 53, 23, 47, 68, 
    95, 54, 81, 80, 72, 66, 111, 93, 86, 91, 87, 41, 16, 46, 74, 
    101, 60, 70, 102, 45, 72, 101, 73, 100, 57, 34, 44, 28, 40, 77, 
    106, 73, 75, 90, 25, 54, 68, 88, 95, 49, 38, 41, 40, 48, 78, 
    100, 88, 66, 62, 71, 49, 58, 75, 37, 22, 18, 18, 31, 60, 63, 
    94, 97, 79, 72, 86, 87, 80, 79, 43, 24, 16, 6, 30, 39, 59, 
    102, 83, 101, 72, 83, 71, 85, 100, 69, 62, 51, 50, 51, 56, 68, 
    89, 88, 97, 87, 77, 93, 100, 99, 90, 85, 85, 87, 88, 86, 68, 
    
    -- channel=177
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 8, 0, 0, 10, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 12, 9, 4, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 11, 4, 
    2, 2, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 7, 7, 10, 
    18, 0, 0, 0, 0, 0, 0, 0, 0, 13, 5, 0, 9, 11, 11, 
    38, 0, 0, 0, 0, 0, 0, 29, 7, 10, 10, 3, 13, 8, 11, 
    19, 26, 5, 0, 0, 12, 13, 0, 0, 0, 0, 3, 9, 1, 10, 
    0, 33, 8, 16, 10, 0, 0, 14, 17, 9, 0, 3, 16, 0, 0, 
    0, 24, 5, 11, 27, 32, 8, 37, 37, 46, 34, 11, 18, 17, 0, 
    5, 31, 18, 0, 61, 30, 8, 0, 0, 15, 0, 0, 18, 23, 0, 
    5, 35, 27, 0, 12, 50, 36, 49, 25, 12, 21, 14, 7, 48, 0, 
    17, 15, 21, 0, 0, 0, 0, 3, 4, 6, 6, 19, 23, 38, 22, 
    8, 16, 13, 29, 0, 6, 7, 0, 0, 0, 0, 0, 10, 12, 26, 
    12, 32, 11, 19, 10, 0, 16, 2, 0, 0, 0, 0, 0, 0, 6, 
    9, 6, 7, 5, 0, 4, 10, 17, 9, 9, 4, 5, 0, 0, 1, 
    
    -- channel=178
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 7, 6, 0, 0, 
    0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 3, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 3, 0, 
    3, 2, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 20, 4, 2, 
    129, 0, 0, 0, 0, 13, 0, 17, 0, 20, 0, 0, 35, 1, 12, 
    78, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 3, 5, 
    0, 98, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 31, 6, 0, 
    0, 55, 0, 0, 55, 29, 0, 39, 39, 30, 0, 0, 57, 53, 0, 
    0, 71, 0, 0, 183, 30, 0, 24, 0, 0, 0, 0, 50, 87, 0, 
    0, 47, 0, 0, 3, 68, 48, 80, 0, 0, 24, 33, 9, 117, 0, 
    0, 0, 13, 0, 0, 0, 0, 0, 0, 6, 4, 39, 64, 46, 43, 
    0, 0, 0, 52, 0, 0, 0, 0, 0, 0, 0, 0, 24, 2, 45, 
    0, 40, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=179
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 7, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 4, 1, 1, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 22, 2, 0, 9, 6, 3, 
    53, 0, 0, 0, 6, 0, 0, 32, 11, 1, 4, 14, 15, 5, 7, 
    4, 25, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 3, 0, 7, 
    0, 22, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 
    0, 0, 0, 0, 27, 32, 0, 51, 47, 62, 63, 23, 13, 3, 0, 
    0, 16, 0, 0, 94, 12, 9, 0, 0, 19, 0, 0, 7, 3, 0, 
    0, 19, 16, 0, 0, 87, 65, 72, 54, 12, 33, 19, 0, 36, 0, 
    7, 0, 11, 0, 0, 0, 0, 0, 13, 17, 8, 29, 33, 35, 27, 
    0, 0, 0, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 32, 
    5, 26, 0, 3, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 11, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=180
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 10, 0, 0, 0, 0, 0, 0, 0, 
    21, 0, 0, 0, 0, 13, 0, 0, 3, 0, 0, 0, 0, 0, 0, 
    0, 15, 0, 0, 11, 0, 0, 8, 9, 1, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 17, 0, 0, 0, 0, 2, 0, 0, 0, 4, 0, 
    0, 16, 13, 0, 29, 5, 0, 0, 0, 0, 0, 0, 0, 16, 0, 
    0, 0, 7, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 23, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=181
    60, 0, 10, 1, 17, 10, 21, 0, 51, 0, 0, 13, 0, 0, 32, 
    6, 26, 6, 6, 6, 12, 25, 3, 58, 27, 0, 0, 0, 17, 4, 
    48, 0, 4, 1, 5, 13, 31, 0, 19, 54, 0, 22, 0, 0, 2, 
    33, 0, 6, 0, 8, 8, 21, 16, 0, 8, 16, 57, 9, 0, 0, 
    0, 0, 3, 3, 5, 18, 18, 14, 36, 0, 2, 90, 0, 0, 0, 
    0, 17, 0, 11, 15, 0, 49, 9, 33, 0, 29, 73, 0, 0, 0, 
    0, 0, 18, 24, 0, 0, 24, 51, 0, 1, 69, 50, 0, 0, 0, 
    28, 0, 25, 0, 0, 22, 16, 0, 5, 14, 96, 51, 0, 0, 51, 
    27, 0, 15, 39, 0, 0, 67, 0, 0, 13, 80, 31, 0, 0, 121, 
    40, 0, 7, 161, 0, 0, 76, 0, 80, 32, 16, 22, 0, 0, 159, 
    38, 0, 13, 147, 0, 0, 0, 0, 65, 25, 0, 0, 0, 0, 120, 
    16, 0, 0, 52, 38, 1, 0, 52, 38, 10, 12, 0, 0, 0, 0, 
    0, 3, 7, 0, 53, 21, 0, 51, 38, 21, 25, 0, 0, 0, 0, 
    27, 0, 38, 0, 38, 0, 0, 44, 11, 18, 10, 0, 16, 0, 16, 
    5, 0, 21, 0, 11, 6, 8, 9, 10, 9, 0, 0, 15, 30, 0, 
    
    -- channel=182
    0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 13, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 11, 37, 16, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 16, 0, 0, 11, 
    0, 0, 0, 0, 31, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 0, 0, 17, 0, 23, 24, 0, 2, 2, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 23, 35, 38, 34, 12, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 10, 21, 21, 14, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=183
    44, 64, 18, 22, 20, 18, 12, 10, 11, 1, 6, 21, 18, 13, 16, 
    14, 12, 20, 21, 20, 31, 34, 23, 31, 21, 0, 0, 8, 18, 9, 
    17, 0, 24, 12, 20, 18, 31, 16, 24, 70, 49, 40, 9, 0, 18, 
    3, 4, 9, 11, 11, 12, 12, 16, 3, 9, 29, 34, 7, 14, 8, 
    0, 10, 16, 14, 15, 21, 25, 48, 33, 0, 5, 20, 0, 0, 4, 
    0, 27, 26, 20, 3, 16, 49, 0, 0, 11, 10, 0, 0, 1, 1, 
    9, 0, 10, 14, 24, 5, 0, 65, 74, 54, 27, 15, 6, 11, 3, 
    25, 0, 6, 0, 14, 24, 40, 2, 3, 11, 52, 12, 0, 32, 39, 
    28, 3, 22, 9, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 52, 
    25, 0, 6, 35, 0, 0, 0, 28, 49, 0, 26, 34, 0, 0, 72, 
    27, 0, 0, 5, 21, 0, 0, 0, 0, 0, 0, 0, 20, 0, 16, 
    0, 21, 0, 75, 49, 58, 58, 20, 2, 0, 0, 0, 0, 0, 0, 
    22, 7, 14, 0, 50, 19, 23, 52, 53, 50, 42, 31, 11, 1, 0, 
    15, 0, 5, 1, 0, 25, 9, 25, 31, 42, 44, 55, 59, 44, 0, 
    10, 39, 21, 30, 41, 30, 10, 0, 9, 13, 22, 19, 29, 28, 27, 
    
    -- channel=184
    56, 32, 33, 33, 35, 26, 32, 14, 45, 9, 15, 20, 10, 14, 40, 
    50, 56, 26, 34, 35, 36, 35, 26, 42, 10, 1, 18, 26, 35, 19, 
    65, 35, 33, 33, 36, 36, 42, 14, 36, 59, 25, 36, 20, 21, 28, 
    48, 35, 38, 33, 43, 38, 42, 35, 23, 38, 25, 44, 18, 8, 22, 
    31, 39, 42, 31, 41, 39, 43, 46, 43, 15, 31, 73, 8, 20, 23, 
    0, 41, 37, 47, 34, 27, 92, 54, 57, 19, 43, 40, 0, 14, 14, 
    0, 19, 68, 63, 30, 58, 66, 80, 48, 50, 68, 35, 0, 10, 16, 
    39, 0, 75, 42, 46, 87, 65, 63, 77, 80, 104, 45, 0, 25, 42, 
    52, 8, 73, 58, 55, 24, 92, 34, 48, 45, 57, 9, 0, 9, 94, 
    48, 0, 80, 124, 0, 40, 85, 54, 69, 15, 16, 28, 0, 0, 139, 
    64, 9, 69, 99, 0, 0, 8, 0, 43, 7, 0, 4, 0, 0, 130, 
    44, 39, 40, 78, 49, 38, 32, 35, 0, 0, 0, 0, 0, 0, 46, 
    37, 40, 38, 30, 73, 45, 27, 56, 41, 18, 11, 0, 0, 0, 0, 
    50, 11, 66, 20, 60, 27, 26, 61, 35, 48, 37, 34, 40, 25, 40, 
    36, 43, 53, 40, 50, 48, 39, 37, 36, 29, 30, 32, 44, 46, 21, 
    
    -- channel=185
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 33, 7, 0, 1, 20, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 2, 9, 40, 32, 58, 76, 16, 0, 0, 0, 
    0, 0, 0, 20, 58, 0, 18, 0, 0, 13, 0, 0, 0, 0, 0, 
    0, 0, 11, 29, 0, 66, 42, 43, 50, 7, 21, 4, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 1, 8, 8, 6, 14, 3, 14, 11, 
    0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=186
    60, 40, 31, 30, 37, 35, 37, 26, 44, 8, 9, 19, 12, 8, 26, 
    38, 44, 34, 36, 36, 39, 45, 32, 54, 27, 0, 9, 9, 23, 15, 
    54, 24, 36, 34, 36, 43, 46, 30, 44, 58, 23, 31, 13, 12, 17, 
    40, 28, 35, 32, 41, 37, 41, 38, 24, 32, 38, 49, 13, 9, 14, 
    18, 25, 36, 38, 38, 41, 28, 34, 43, 9, 29, 60, 4, 12, 11, 
    0, 38, 32, 41, 39, 24, 56, 26, 24, 6, 34, 38, 0, 12, 6, 
    0, 0, 43, 40, 28, 42, 35, 46, 30, 35, 50, 29, 1, 12, 9, 
    32, 0, 41, 28, 21, 46, 49, 30, 36, 35, 69, 33, 0, 9, 42, 
    34, 0, 37, 51, 11, 5, 59, 18, 12, 17, 29, 10, 0, 0, 69, 
    34, 0, 29, 92, 0, 10, 45, 8, 66, 17, 10, 23, 0, 0, 90, 
    39, 0, 28, 70, 2, 0, 0, 0, 22, 16, 0, 0, 1, 0, 70, 
    21, 24, 14, 54, 48, 25, 23, 35, 17, 2, 1, 0, 0, 0, 4, 
    18, 21, 33, 1, 55, 25, 9, 49, 36, 24, 24, 5, 0, 0, 4, 
    27, 0, 38, 16, 27, 16, 7, 38, 25, 32, 27, 25, 33, 24, 19, 
    17, 20, 26, 24, 29, 28, 25, 18, 23, 17, 17, 18, 30, 33, 16, 
    
    -- channel=187
    34, 0, 14, 3, 1, 5, 8, 8, 7, 20, 4, 6, 5, 2, 22, 
    22, 8, 27, 2, 0, 8, 17, 5, 0, 28, 0, 11, 0, 5, 15, 
    12, 0, 18, 11, 6, 14, 7, 22, 5, 12, 0, 25, 4, 9, 9, 
    47, 0, 11, 9, 12, 19, 14, 23, 12, 6, 24, 24, 6, 5, 7, 
    30, 0, 8, 11, 10, 9, 17, 0, 31, 7, 24, 18, 5, 7, 4, 
    24, 10, 0, 9, 26, 0, 10, 7, 25, 0, 15, 32, 0, 11, 2, 
    0, 15, 0, 1, 25, 0, 30, 0, 0, 0, 29, 31, 8, 0, 3, 
    6, 0, 6, 17, 0, 11, 29, 0, 0, 0, 14, 32, 20, 0, 30, 
    7, 0, 3, 54, 0, 31, 26, 0, 0, 22, 30, 16, 11, 0, 34, 
    7, 0, 0, 30, 0, 15, 39, 0, 12, 31, 20, 0, 5, 0, 0, 
    9, 3, 0, 26, 0, 12, 23, 0, 45, 36, 12, 0, 11, 0, 0, 
    30, 0, 0, 17, 17, 4, 1, 0, 27, 9, 2, 6, 5, 27, 0, 
    23, 0, 15, 7, 57, 16, 0, 11, 12, 4, 0, 0, 0, 32, 0, 
    2, 19, 15, 32, 9, 0, 0, 12, 7, 8, 5, 0, 5, 3, 0, 
    0, 0, 18, 8, 20, 0, 9, 15, 12, 23, 5, 1, 14, 7, 17, 
    
    -- channel=188
    50, 28, 34, 33, 37, 27, 29, 13, 37, 7, 11, 11, 1, 7, 28, 
    53, 65, 27, 37, 37, 35, 32, 24, 30, 0, 2, 14, 22, 26, 11, 
    68, 47, 37, 39, 39, 41, 40, 17, 36, 38, 13, 20, 15, 18, 19, 
    53, 51, 44, 39, 50, 42, 43, 35, 30, 39, 20, 28, 13, 0, 16, 
    43, 43, 49, 38, 46, 41, 42, 37, 36, 20, 32, 66, 10, 20, 20, 
    0, 42, 38, 51, 46, 32, 86, 66, 66, 21, 39, 34, 6, 13, 12, 
    0, 35, 75, 67, 31, 66, 72, 60, 35, 43, 57, 21, 0, 8, 13, 
    29, 1, 77, 51, 55, 88, 61, 65, 82, 83, 84, 35, 0, 21, 27, 
    34, 15, 70, 56, 77, 34, 84, 54, 62, 61, 69, 6, 0, 16, 71, 
    33, 0, 81, 105, 16, 56, 82, 51, 54, 9, 1, 15, 0, 8, 114, 
    48, 13, 76, 86, 0, 0, 13, 0, 42, 3, 2, 8, 0, 0, 122, 
    36, 29, 45, 57, 35, 16, 15, 28, 0, 0, 0, 0, 0, 0, 59, 
    24, 33, 30, 46, 59, 44, 14, 33, 19, 1, 0, 0, 0, 0, 0, 
    37, 11, 58, 16, 55, 18, 20, 43, 19, 31, 22, 19, 23, 12, 39, 
    23, 26, 37, 27, 34, 39, 29, 33, 28, 16, 21, 25, 32, 35, 8, 
    
    -- channel=189
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=190
    0, 0, 8, 5, 9, 9, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 22, 6, 15, 16, 6, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    18, 35, 12, 22, 20, 21, 10, 13, 0, 0, 0, 0, 0, 0, 0, 
    11, 30, 25, 24, 28, 23, 21, 6, 20, 16, 0, 0, 0, 0, 0, 
    21, 23, 21, 26, 29, 18, 9, 0, 0, 28, 10, 0, 0, 0, 0, 
    34, 15, 26, 22, 28, 21, 0, 43, 13, 9, 6, 0, 0, 0, 0, 
    5, 43, 33, 26, 8, 41, 37, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 38, 30, 31, 28, 23, 0, 35, 30, 25, 0, 0, 0, 0, 0, 
    0, 16, 20, 3, 75, 57, 26, 69, 63, 62, 42, 0, 0, 21, 0, 
    0, 34, 33, 0, 89, 32, 18, 1, 0, 0, 0, 0, 0, 29, 0, 
    0, 29, 50, 0, 0, 56, 37, 61, 18, 0, 0, 0, 0, 49, 9, 
    11, 4, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 17, 47, 
    0, 15, 7, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 
    8, 25, 9, 2, 16, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 2, 8, 11, 2, 0, 0, 0, 0, 0, 0, 
    
    -- channel=191
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 13, 1, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 12, 8, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 5, 0, 0, 0, 8, 
    0, 0, 0, 7, 29, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 27, 11, 4, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 18, 14, 0, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=192
    83, 77, 78, 78, 69, 60, 58, 50, 45, 40, 38, 22, 0, 11, 16, 
    63, 61, 46, 43, 37, 33, 33, 32, 29, 28, 27, 7, 6, 18, 16, 
    40, 30, 28, 23, 27, 28, 27, 33, 31, 29, 33, 0, 7, 27, 22, 
    23, 24, 25, 25, 28, 30, 32, 34, 37, 33, 2, 21, 34, 28, 21, 
    21, 23, 25, 25, 28, 34, 38, 32, 37, 26, 6, 0, 3, 14, 20, 
    25, 23, 24, 24, 24, 39, 53, 47, 59, 47, 75, 0, 13, 6, 12, 
    25, 25, 20, 19, 36, 26, 28, 5, 10, 56, 88, 7, 0, 0, 0, 
    26, 21, 23, 12, 13, 23, 6, 22, 45, 86, 91, 18, 9, 0, 26, 
    23, 20, 8, 22, 0, 9, 48, 99, 92, 99, 71, 0, 9, 42, 49, 
    16, 78, 0, 8, 0, 11, 65, 81, 87, 63, 84, 48, 44, 52, 49, 
    51, 37, 22, 0, 0, 11, 66, 75, 49, 6, 24, 90, 55, 48, 0, 
    19, 26, 27, 0, 0, 27, 88, 78, 0, 4, 0, 36, 63, 0, 2, 
    9, 18, 26, 0, 28, 36, 71, 78, 0, 16, 0, 0, 46, 0, 0, 
    10, 20, 20, 13, 28, 39, 45, 45, 5, 27, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    
    -- channel=193
    54, 45, 40, 40, 35, 31, 30, 31, 24, 11, 25, 19, 9, 20, 26, 
    30, 34, 27, 21, 19, 21, 21, 23, 23, 28, 21, 23, 24, 28, 21, 
    18, 9, 14, 16, 21, 21, 22, 27, 28, 29, 15, 21, 35, 32, 26, 
    18, 21, 22, 23, 24, 22, 21, 27, 32, 26, 6, 23, 28, 20, 21, 
    20, 20, 20, 20, 20, 22, 22, 16, 19, 12, 27, 34, 13, 23, 22, 
    20, 19, 20, 19, 17, 18, 36, 37, 11, 3, 28, 22, 16, 11, 20, 
    20, 19, 16, 18, 16, 0, 0, 0, 0, 17, 0, 12, 29, 1, 13, 
    19, 16, 20, 14, 0, 20, 17, 33, 54, 50, 0, 0, 19, 28, 27, 
    16, 16, 6, 2, 7, 9, 30, 19, 0, 0, 0, 0, 6, 41, 16, 
    20, 23, 16, 9, 15, 19, 27, 0, 0, 0, 0, 24, 26, 2, 0, 
    15, 0, 0, 9, 19, 26, 25, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 12, 0, 14, 27, 13, 10, 0, 0, 15, 17, 6, 0, 0, 24, 
    12, 8, 0, 21, 30, 22, 6, 0, 0, 20, 15, 16, 0, 4, 17, 
    16, 13, 0, 6, 0, 0, 0, 0, 0, 3, 0, 18, 0, 16, 22, 
    16, 11, 14, 25, 26, 24, 23, 20, 21, 7, 8, 19, 26, 27, 28, 
    
    -- channel=194
    119, 123, 133, 134, 125, 113, 110, 95, 93, 65, 51, 45, 12, 0, 23, 
    130, 114, 112, 110, 101, 88, 85, 75, 67, 55, 53, 29, 0, 0, 36, 
    92, 82, 79, 79, 73, 67, 67, 63, 60, 61, 53, 0, 0, 26, 44, 
    54, 62, 65, 63, 66, 68, 67, 65, 63, 62, 0, 0, 16, 44, 44, 
    56, 66, 67, 67, 71, 72, 65, 66, 53, 15, 0, 0, 27, 43, 44, 
    64, 68, 65, 64, 71, 59, 61, 65, 70, 49, 0, 0, 3, 0, 37, 
    70, 68, 63, 63, 61, 44, 0, 0, 0, 9, 60, 0, 0, 0, 6, 
    69, 67, 67, 38, 0, 0, 0, 0, 0, 45, 28, 0, 0, 0, 0, 
    67, 70, 22, 0, 0, 0, 9, 62, 50, 33, 3, 0, 1, 0, 32, 
    81, 66, 0, 0, 0, 0, 34, 34, 15, 26, 49, 0, 25, 6, 0, 
    88, 76, 0, 0, 0, 0, 26, 18, 0, 0, 0, 57, 0, 0, 0, 
    61, 0, 0, 0, 0, 0, 23, 19, 0, 0, 0, 22, 0, 0, 0, 
    31, 0, 0, 0, 0, 0, 30, 5, 0, 0, 0, 0, 11, 0, 0, 
    10, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=195
    25, 43, 50, 55, 56, 49, 46, 46, 35, 42, 30, 20, 32, 10, 12, 
    51, 48, 45, 42, 39, 35, 32, 33, 26, 24, 16, 31, 11, 0, 12, 
    39, 37, 30, 28, 25, 20, 20, 22, 19, 16, 22, 14, 5, 0, 18, 
    18, 15, 14, 16, 14, 14, 13, 20, 21, 19, 39, 0, 0, 17, 21, 
    9, 11, 13, 14, 12, 17, 18, 17, 14, 29, 18, 0, 17, 23, 17, 
    10, 12, 15, 17, 11, 7, 4, 0, 5, 10, 0, 28, 9, 8, 16, 
    13, 13, 17, 12, 13, 17, 33, 33, 21, 0, 0, 26, 10, 16, 11, 
    12, 15, 9, 12, 20, 0, 10, 0, 0, 0, 0, 47, 0, 0, 0, 
    12, 9, 30, 12, 21, 8, 0, 0, 0, 1, 21, 36, 0, 0, 0, 
    6, 0, 26, 0, 14, 0, 0, 0, 0, 22, 0, 0, 0, 0, 16, 
    0, 20, 18, 5, 7, 0, 0, 0, 34, 26, 15, 0, 6, 16, 36, 
    10, 0, 2, 15, 0, 0, 0, 0, 50, 0, 8, 0, 0, 34, 1, 
    7, 0, 0, 5, 0, 0, 0, 2, 42, 0, 3, 0, 1, 24, 1, 
    0, 0, 5, 3, 2, 19, 23, 25, 31, 0, 16, 16, 12, 10, 1, 
    2, 6, 3, 2, 0, 0, 0, 0, 4, 0, 5, 9, 2, 2, 0, 
    
    -- channel=196
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=197
    0, 0, 0, 4, 5, 4, 3, 3, 10, 25, 6, 0, 26, 15, 0, 
    0, 0, 4, 4, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 26, 4, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 67, 75, 0, 0, 18, 0, 0, 
    0, 0, 0, 0, 0, 70, 74, 83, 44, 0, 0, 0, 0, 24, 5, 
    0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 62, 0, 0, 0, 
    0, 0, 11, 18, 38, 25, 0, 0, 18, 9, 21, 12, 0, 0, 0, 
    0, 0, 0, 2, 21, 7, 0, 3, 0, 86, 69, 0, 0, 0, 34, 
    0, 116, 17, 9, 5, 0, 0, 0, 66, 84, 76, 61, 38, 54, 103, 
    10, 0, 0, 6, 0, 0, 0, 0, 41, 0, 0, 41, 5, 50, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 9, 50, 46, 6, 
    0, 7, 58, 64, 107, 151, 163, 167, 94, 10, 19, 8, 52, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 36, 13, 0, 0, 0, 
    
    -- channel=198
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 22, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 3, 24, 66, 48, 23, 10, 0, 0, 
    0, 0, 0, 0, 0, 7, 82, 104, 87, 62, 132, 85, 0, 29, 0, 
    0, 0, 0, 0, 10, 16, 17, 0, 0, 0, 117, 164, 14, 0, 0, 
    0, 0, 0, 33, 29, 15, 33, 47, 87, 147, 143, 134, 39, 0, 49, 
    0, 0, 14, 5, 34, 0, 0, 133, 143, 130, 154, 51, 12, 60, 99, 
    0, 65, 110, 7, 6, 0, 0, 115, 119, 112, 64, 147, 128, 109, 91, 
    0, 33, 80, 28, 0, 0, 28, 115, 135, 0, 0, 0, 108, 82, 20, 
    0, 6, 66, 31, 0, 32, 47, 129, 129, 10, 10, 0, 59, 74, 0, 
    0, 11, 56, 37, 36, 97, 100, 112, 122, 14, 56, 1, 12, 21, 0, 
    0, 0, 22, 0, 0, 0, 0, 0, 6, 5, 21, 2, 0, 0, 0, 
    1, 5, 11, 34, 9, 12, 10, 2, 0, 0, 14, 0, 0, 0, 0, 
    
    -- channel=199
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=200
    26, 21, 24, 21, 17, 19, 22, 13, 23, 19, 9, 15, 1, 5, 7, 
    29, 22, 21, 27, 26, 23, 24, 17, 18, 14, 20, 3, 0, 18, 13, 
    22, 24, 27, 25, 23, 23, 24, 18, 17, 20, 24, 0, 0, 14, 8, 
    22, 25, 24, 23, 24, 27, 28, 24, 18, 21, 0, 13, 16, 18, 12, 
    24, 28, 28, 27, 31, 28, 22, 30, 38, 20, 0, 5, 12, 13, 14, 
    28, 29, 27, 25, 34, 43, 29, 12, 20, 7, 10, 0, 16, 2, 15, 
    29, 28, 25, 29, 37, 26, 19, 10, 13, 72, 63, 0, 0, 7, 7, 
    29, 29, 34, 24, 6, 17, 0, 13, 28, 54, 48, 0, 0, 7, 19, 
    30, 37, 19, 18, 0, 12, 47, 58, 47, 53, 26, 0, 32, 39, 31, 
    42, 65, 0, 18, 0, 15, 73, 52, 49, 28, 43, 6, 28, 28, 19, 
    70, 33, 0, 0, 0, 16, 77, 44, 8, 0, 39, 82, 25, 17, 0, 
    37, 23, 5, 0, 2, 29, 77, 41, 0, 6, 0, 57, 38, 0, 0, 
    25, 17, 17, 0, 30, 25, 62, 46, 0, 19, 0, 11, 37, 0, 1, 
    16, 18, 9, 1, 29, 35, 37, 36, 0, 29, 0, 0, 3, 0, 0, 
    12, 5, 1, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 
    
    -- channel=201
    146, 158, 167, 173, 170, 150, 143, 135, 115, 102, 87, 71, 39, 10, 54, 
    157, 145, 144, 138, 128, 114, 109, 104, 91, 84, 69, 55, 13, 0, 63, 
    116, 111, 101, 101, 93, 87, 88, 86, 84, 79, 55, 20, 15, 37, 74, 
    75, 79, 82, 82, 83, 85, 82, 83, 82, 75, 47, 0, 40, 72, 76, 
    72, 82, 83, 85, 83, 86, 78, 74, 43, 24, 0, 0, 46, 67, 68, 
    80, 83, 82, 83, 74, 44, 35, 56, 68, 78, 1, 0, 2, 33, 58, 
    84, 83, 85, 74, 50, 43, 17, 0, 0, 0, 4, 15, 0, 11, 25, 
    83, 84, 64, 34, 16, 0, 10, 0, 0, 0, 1, 61, 0, 0, 0, 
    82, 69, 21, 2, 14, 0, 0, 3, 25, 19, 20, 7, 0, 0, 9, 
    75, 10, 11, 0, 0, 0, 0, 6, 0, 32, 48, 3, 0, 0, 8, 
    47, 68, 3, 0, 0, 0, 0, 0, 17, 0, 0, 1, 12, 5, 32, 
    58, 0, 0, 0, 0, 0, 0, 0, 44, 0, 0, 0, 0, 17, 0, 
    34, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 2, 0, 
    20, 7, 5, 0, 0, 11, 16, 18, 28, 0, 0, 0, 0, 0, 0, 
    23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=202
    133, 138, 137, 140, 137, 129, 122, 122, 105, 67, 84, 85, 37, 31, 72, 
    142, 135, 126, 128, 121, 112, 106, 106, 98, 93, 91, 62, 31, 39, 83, 
    92, 98, 109, 106, 100, 98, 98, 96, 94, 94, 44, 27, 45, 58, 77, 
    90, 94, 94, 97, 97, 98, 103, 102, 95, 85, 12, 11, 57, 75, 85, 
    88, 96, 95, 96, 96, 92, 72, 87, 106, 96, 45, 28, 74, 82, 81, 
    95, 97, 97, 95, 92, 84, 38, 0, 0, 0, 1, 35, 10, 60, 75, 
    97, 96, 95, 91, 58, 0, 0, 0, 5, 4, 0, 56, 17, 3, 52, 
    94, 98, 89, 62, 20, 19, 7, 61, 59, 0, 0, 0, 31, 18, 46, 
    94, 94, 35, 0, 0, 0, 0, 0, 0, 0, 0, 44, 43, 38, 0, 
    100, 63, 18, 0, 11, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 
    62, 0, 0, 0, 25, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    47, 14, 0, 6, 21, 0, 0, 0, 0, 11, 12, 0, 0, 0, 32, 
    43, 0, 0, 27, 9, 0, 0, 0, 10, 0, 19, 3, 0, 9, 16, 
    42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 23, 16, 
    39, 26, 21, 26, 13, 14, 13, 15, 19, 0, 0, 22, 18, 18, 16, 
    
    -- channel=203
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=204
    38, 17, 16, 10, 4, 3, 8, 0, 10, 0, 0, 8, 0, 0, 1, 
    5, 3, 0, 0, 0, 0, 0, 0, 1, 3, 17, 3, 0, 33, 2, 
    0, 0, 0, 0, 0, 0, 2, 6, 9, 11, 45, 0, 2, 29, 1, 
    0, 2, 3, 1, 6, 6, 9, 14, 13, 21, 0, 12, 14, 8, 0, 
    4, 3, 1, 1, 6, 16, 13, 9, 26, 17, 0, 17, 0, 0, 2, 
    5, 1, 0, 0, 15, 37, 51, 14, 5, 0, 32, 0, 7, 0, 0, 
    3, 0, 0, 7, 42, 0, 0, 0, 0, 80, 80, 0, 4, 0, 0, 
    0, 0, 18, 15, 0, 18, 0, 38, 92, 138, 18, 0, 0, 26, 49, 
    0, 16, 10, 0, 0, 17, 51, 109, 16, 0, 0, 0, 32, 74, 44, 
    15, 107, 0, 20, 0, 37, 103, 33, 3, 0, 0, 0, 41, 4, 0, 
    66, 1, 0, 0, 0, 56, 123, 17, 0, 0, 32, 62, 0, 0, 0, 
    35, 13, 14, 0, 28, 72, 92, 10, 0, 17, 0, 81, 11, 0, 0, 
    19, 23, 28, 0, 76, 48, 87, 2, 0, 38, 0, 20, 52, 0, 15, 
    18, 30, 9, 0, 22, 0, 0, 0, 0, 51, 0, 0, 18, 0, 16, 
    10, 6, 5, 12, 15, 17, 14, 9, 6, 41, 0, 0, 14, 16, 24, 
    
    -- channel=205
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 41, 9, 0, 0, 
    0, 0, 0, 0, 0, 1, 47, 62, 28, 2, 21, 56, 16, 19, 0, 
    0, 0, 0, 0, 10, 0, 17, 3, 0, 0, 41, 80, 9, 4, 0, 
    0, 0, 0, 28, 41, 26, 14, 0, 34, 51, 52, 75, 0, 0, 5, 
    0, 0, 43, 18, 36, 2, 0, 42, 49, 58, 52, 16, 0, 33, 33, 
    0, 40, 58, 23, 23, 0, 0, 46, 59, 86, 33, 35, 59, 54, 76, 
    0, 10, 31, 44, 6, 3, 4, 43, 98, 11, 23, 4, 35, 73, 6, 
    0, 11, 33, 47, 0, 17, 13, 53, 84, 10, 22, 7, 20, 65, 0, 
    0, 0, 29, 35, 35, 64, 69, 74, 78, 2, 47, 28, 26, 24, 3, 
    0, 3, 32, 16, 18, 16, 15, 14, 13, 12, 18, 24, 5, 5, 2, 
    
    -- channel=206
    93, 112, 113, 121, 126, 113, 103, 108, 85, 92, 80, 59, 65, 9, 57, 
    110, 111, 113, 107, 98, 90, 84, 85, 75, 71, 47, 79, 44, 0, 63, 
    83, 93, 83, 84, 73, 71, 73, 70, 67, 55, 34, 31, 31, 27, 68, 
    65, 64, 64, 68, 64, 67, 64, 71, 65, 55, 86, 0, 41, 68, 71, 
    58, 64, 65, 69, 58, 60, 48, 51, 39, 98, 58, 0, 60, 67, 60, 
    62, 66, 68, 69, 42, 14, 0, 0, 0, 0, 0, 145, 0, 60, 58, 
    65, 68, 77, 45, 27, 19, 64, 71, 39, 0, 0, 153, 43, 10, 37, 
    64, 70, 23, 43, 55, 0, 23, 0, 0, 0, 0, 138, 53, 0, 0, 
    67, 32, 60, 0, 52, 0, 0, 0, 0, 0, 75, 148, 0, 0, 0, 
    23, 0, 120, 0, 54, 0, 0, 0, 0, 51, 0, 5, 0, 5, 56, 
    0, 0, 73, 36, 25, 0, 0, 0, 110, 73, 20, 0, 28, 55, 96, 
    27, 0, 7, 66, 0, 0, 0, 0, 174, 0, 31, 0, 0, 118, 12, 
    19, 0, 0, 40, 0, 0, 0, 2, 160, 0, 49, 11, 0, 88, 6, 
    24, 0, 8, 8, 0, 7, 11, 21, 67, 0, 38, 51, 14, 25, 3, 
    23, 25, 10, 27, 0, 1, 10, 15, 20, 0, 19, 33, 10, 7, 0, 
    
    -- channel=207
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 21, 30, 17, 78, 118, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 130, 0, 14, 0, 
    0, 0, 0, 0, 0, 0, 29, 37, 17, 0, 29, 83, 45, 0, 25, 
    0, 0, 0, 7, 26, 0, 0, 47, 27, 42, 47, 19, 16, 0, 32, 
    0, 3, 29, 0, 4, 0, 0, 30, 26, 3, 69, 96, 24, 24, 3, 
    0, 4, 88, 3, 0, 5, 0, 35, 30, 5, 0, 11, 41, 15, 26, 
    0, 0, 71, 17, 3, 0, 0, 33, 99, 7, 8, 0, 44, 43, 2, 
    0, 4, 49, 17, 6, 33, 0, 20, 81, 14, 21, 0, 9, 32, 0, 
    0, 0, 10, 0, 0, 0, 0, 0, 70, 0, 29, 1, 0, 5, 0, 
    0, 0, 8, 13, 6, 9, 3, 1, 0, 0, 21, 9, 0, 0, 0, 
    
    -- channel=208
    194, 213, 219, 226, 223, 206, 195, 190, 173, 139, 133, 114, 80, 45, 96, 
    217, 206, 205, 203, 191, 174, 166, 159, 146, 131, 112, 103, 37, 33, 111, 
    171, 171, 165, 163, 151, 145, 143, 138, 133, 125, 95, 41, 47, 74, 119, 
    132, 136, 138, 138, 139, 141, 139, 135, 131, 122, 73, 8, 77, 117, 124, 
    128, 140, 142, 142, 140, 137, 121, 119, 94, 93, 29, 16, 99, 119, 118, 
    138, 142, 141, 140, 126, 85, 64, 68, 71, 51, 0, 43, 24, 80, 109, 
    143, 144, 143, 122, 103, 68, 48, 31, 26, 0, 6, 46, 13, 35, 70, 
    142, 142, 107, 89, 49, 23, 21, 0, 0, 0, 12, 75, 23, 0, 1, 
    143, 115, 75, 24, 26, 1, 0, 0, 30, 24, 47, 55, 22, 0, 13, 
    118, 55, 48, 0, 15, 0, 0, 11, 10, 52, 22, 15, 11, 13, 40, 
    99, 60, 21, 8, 3, 0, 0, 5, 55, 19, 11, 0, 23, 29, 45, 
    100, 5, 1, 12, 0, 0, 0, 7, 58, 0, 7, 0, 0, 40, 6, 
    74, 9, 0, 0, 0, 0, 0, 6, 46, 0, 8, 4, 6, 25, 13, 
    61, 28, 14, 7, 6, 24, 29, 34, 34, 0, 17, 14, 8, 4, 4, 
    58, 26, 0, 0, 0, 0, 0, 0, 0, 3, 19, 6, 0, 0, 0, 
    
    -- channel=209
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 14, 17, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 
    2, 8, 0, 0, 0, 0, 0, 0, 0, 0, 6, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 25, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 15, 57, 71, 0, 0, 30, 0, 0, 
    0, 0, 0, 1, 10, 61, 62, 59, 43, 54, 58, 0, 1, 31, 10, 
    1, 0, 0, 2, 16, 19, 14, 0, 0, 0, 53, 36, 0, 12, 0, 
    3, 7, 18, 41, 26, 35, 40, 36, 67, 71, 52, 9, 7, 0, 25, 
    8, 0, 0, 36, 15, 30, 68, 68, 63, 84, 96, 0, 14, 39, 46, 
    38, 102, 19, 19, 10, 5, 50, 59, 56, 60, 71, 120, 65, 57, 52, 
    36, 29, 23, 6, 4, 35, 64, 54, 7, 17, 5, 75, 58, 24, 8, 
    27, 30, 36, 0, 5, 1, 48, 57, 0, 25, 0, 25, 71, 20, 15, 
    13, 35, 56, 54, 89, 116, 122, 124, 59, 44, 32, 10, 41, 14, 10, 
    10, 13, 4, 0, 0, 0, 1, 4, 2, 38, 34, 9, 1, 1, 3, 
    
    -- channel=210
    0, 0, 0, 0, 0, 0, 3, 0, 0, 10, 0, 0, 0, 40, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 29, 0, 
    7, 4, 3, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 4, 0, 0, 46, 55, 0, 0, 79, 0, 0, 
    0, 0, 0, 4, 16, 35, 26, 12, 43, 114, 78, 0, 0, 67, 10, 
    0, 0, 8, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 8, 5, 
    0, 3, 0, 46, 0, 47, 83, 73, 2, 6, 0, 0, 9, 0, 6, 
    8, 30, 0, 27, 0, 54, 136, 43, 1, 0, 119, 0, 0, 0, 0, 
    65, 99, 0, 0, 0, 32, 89, 10, 0, 0, 66, 238, 0, 0, 0, 
    28, 0, 24, 0, 10, 61, 112, 0, 0, 5, 0, 121, 54, 0, 0, 
    19, 21, 47, 0, 22, 0, 31, 0, 0, 44, 0, 0, 134, 0, 31, 
    0, 30, 52, 24, 110, 134, 136, 126, 11, 76, 0, 0, 59, 1, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 72, 13, 0, 0, 2, 13, 
    
    -- channel=211
    0, 1, 22, 29, 29, 29, 32, 23, 27, 50, 19, 12, 16, 37, 0, 
    30, 14, 24, 32, 33, 27, 26, 20, 16, 8, 3, 0, 0, 0, 0, 
    41, 47, 36, 25, 20, 11, 9, 5, 0, 0, 3, 4, 0, 0, 0, 
    19, 10, 7, 5, 3, 3, 0, 0, 0, 0, 16, 26, 0, 10, 11, 
    4, 6, 8, 8, 8, 1, 6, 1, 0, 0, 0, 0, 3, 9, 8, 
    5, 5, 7, 9, 10, 0, 0, 0, 23, 50, 0, 0, 53, 0, 8, 
    5, 6, 8, 12, 1, 48, 74, 84, 66, 27, 0, 0, 0, 50, 20, 
    9, 7, 1, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 5, 8, 43, 11, 36, 15, 0, 0, 4, 0, 0, 0, 0, 0, 
    6, 0, 0, 10, 3, 21, 15, 4, 0, 38, 75, 0, 0, 0, 7, 
    23, 87, 0, 0, 9, 0, 0, 0, 13, 70, 76, 128, 8, 29, 58, 
    25, 3, 0, 0, 0, 0, 3, 0, 0, 0, 0, 49, 26, 0, 7, 
    19, 6, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 68, 16, 17, 
    0, 12, 40, 44, 87, 140, 151, 153, 85, 22, 20, 0, 50, 25, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 23, 8, 0, 0, 0, 
    
    -- channel=212
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 25, 22, 38, 22, 32, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 14, 0, 0, 36, 103, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 25, 93, 79, 22, 0, 0, 1, 
    0, 0, 0, 12, 0, 5, 34, 101, 82, 76, 55, 0, 0, 25, 43, 
    0, 29, 0, 13, 0, 10, 61, 84, 79, 80, 66, 12, 45, 49, 42, 
    0, 45, 2, 0, 0, 2, 79, 76, 60, 0, 35, 99, 54, 47, 0, 
    0, 9, 34, 0, 0, 45, 82, 76, 0, 0, 0, 44, 52, 0, 0, 
    0, 13, 40, 0, 32, 39, 87, 74, 0, 15, 0, 1, 54, 0, 0, 
    0, 9, 30, 9, 40, 48, 52, 48, 0, 21, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 
    
    -- channel=213
    0, 18, 7, 19, 32, 26, 13, 35, 12, 17, 21, 16, 45, 0, 13, 
    17, 31, 29, 26, 23, 22, 12, 23, 15, 15, 0, 51, 40, 0, 14, 
    15, 25, 17, 20, 11, 12, 11, 12, 10, 1, 7, 38, 12, 0, 25, 
    7, 5, 6, 12, 4, 5, 3, 12, 11, 11, 80, 0, 0, 9, 20, 
    0, 4, 5, 10, 0, 4, 0, 0, 0, 73, 75, 0, 16, 17, 11, 
    3, 7, 10, 11, 0, 0, 0, 0, 0, 0, 0, 161, 0, 29, 12, 
    6, 9, 20, 0, 0, 0, 33, 41, 8, 0, 0, 234, 33, 0, 3, 
    5, 14, 0, 19, 40, 0, 27, 0, 0, 0, 0, 168, 81, 0, 0, 
    10, 0, 33, 0, 51, 0, 0, 0, 0, 0, 68, 169, 0, 0, 0, 
    0, 0, 166, 0, 61, 0, 0, 0, 0, 34, 0, 66, 0, 4, 42, 
    0, 0, 114, 29, 29, 0, 0, 0, 100, 81, 0, 0, 36, 45, 97, 
    0, 0, 4, 77, 0, 0, 0, 0, 216, 0, 30, 0, 0, 133, 7, 
    0, 0, 0, 67, 0, 0, 0, 0, 212, 0, 61, 0, 0, 115, 0, 
    0, 0, 0, 9, 0, 0, 0, 0, 84, 0, 37, 53, 0, 25, 0, 
    0, 19, 10, 35, 2, 3, 7, 10, 13, 0, 16, 39, 1, 0, 0, 
    
    -- channel=214
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 18, 66, 46, 32, 0, 0, 0, 
    0, 0, 0, 0, 0, 12, 38, 0, 0, 0, 37, 72, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 54, 51, 0, 0, 
    0, 0, 0, 22, 0, 0, 0, 102, 164, 126, 0, 0, 7, 20, 75, 
    0, 0, 8, 0, 0, 0, 4, 21, 0, 0, 0, 0, 37, 100, 20, 
    0, 69, 41, 7, 0, 0, 3, 0, 0, 0, 0, 48, 68, 9, 0, 
    0, 0, 0, 15, 5, 52, 58, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 1, 15, 36, 28, 10, 0, 0, 20, 20, 0, 0, 0, 3, 
    0, 2, 0, 42, 77, 87, 43, 0, 6, 18, 53, 24, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 16, 
    0, 15, 41, 69, 45, 47, 41, 33, 27, 0, 0, 0, 21, 22, 22, 
    
    -- channel=215
    53, 38, 21, 16, 14, 15, 11, 18, 10, 0, 0, 16, 11, 0, 20, 
    25, 37, 28, 20, 17, 19, 18, 20, 20, 19, 32, 34, 0, 22, 31, 
    0, 0, 12, 20, 19, 26, 27, 27, 29, 30, 23, 5, 39, 36, 30, 
    15, 25, 28, 30, 31, 31, 42, 50, 46, 39, 0, 0, 6, 11, 15, 
    29, 29, 27, 27, 28, 34, 24, 33, 83, 128, 74, 49, 43, 24, 22, 
    30, 31, 31, 27, 26, 57, 89, 50, 0, 0, 68, 119, 0, 46, 22, 
    31, 30, 27, 23, 34, 0, 0, 0, 0, 0, 0, 129, 51, 0, 10, 
    27, 30, 37, 70, 12, 5, 12, 109, 186, 145, 12, 0, 23, 7, 86, 
    27, 30, 26, 0, 0, 0, 0, 28, 0, 0, 0, 14, 46, 113, 38, 
    26, 103, 92, 0, 0, 0, 0, 0, 0, 0, 0, 106, 97, 22, 0, 
    0, 0, 0, 7, 0, 29, 17, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 23, 19, 0, 0, 2, 19, 5, 12, 0, 0, 0, 0, 
    0, 0, 0, 50, 59, 92, 29, 0, 50, 1, 63, 7, 0, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 2, 
    18, 16, 29, 68, 33, 36, 30, 21, 15, 0, 0, 0, 8, 8, 8, 
    
    -- channel=216
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 3, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 20, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 37, 9, 6, 16, 
    0, 0, 0, 0, 0, 1, 3, 7, 5, 3, 39, 0, 16, 3, 0, 
    0, 0, 0, 3, 0, 8, 13, 7, 5, 55, 63, 13, 9, 1, 0, 
    0, 0, 3, 1, 0, 0, 63, 93, 86, 90, 127, 109, 0, 32, 0, 
    0, 4, 7, 0, 12, 13, 41, 15, 4, 0, 77, 227, 14, 2, 0, 
    1, 4, 0, 25, 33, 16, 44, 22, 34, 81, 131, 203, 87, 0, 24, 
    4, 0, 11, 14, 57, 0, 0, 91, 132, 133, 167, 123, 8, 34, 78, 
    0, 26, 139, 8, 40, 0, 0, 97, 120, 139, 90, 161, 97, 103, 109, 
    0, 37, 136, 41, 9, 0, 0, 108, 166, 53, 0, 0, 132, 111, 74, 
    0, 20, 74, 59, 0, 5, 11, 126, 197, 15, 28, 0, 72, 121, 9, 
    0, 19, 51, 58, 0, 69, 55, 112, 189, 3, 69, 3, 8, 82, 0, 
    0, 18, 41, 36, 0, 17, 25, 31, 84, 0, 48, 31, 0, 6, 0, 
    11, 15, 10, 35, 8, 10, 11, 8, 3, 0, 41, 17, 0, 0, 0, 
    
    -- channel=217
    0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 15, 14, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    12, 19, 1, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 37, 67, 0, 0, 22, 0, 0, 
    0, 0, 0, 0, 0, 46, 72, 81, 48, 0, 0, 0, 0, 34, 5, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 67, 0, 0, 0, 
    0, 0, 0, 27, 37, 21, 0, 0, 0, 3, 9, 22, 0, 0, 0, 
    0, 0, 0, 1, 19, 2, 0, 2, 0, 71, 60, 0, 0, 0, 23, 
    0, 97, 16, 5, 5, 0, 0, 0, 54, 76, 58, 69, 26, 45, 92, 
    4, 0, 0, 8, 0, 0, 0, 0, 48, 0, 0, 17, 5, 49, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 46, 44, 3, 
    0, 1, 48, 48, 81, 132, 142, 147, 100, 0, 27, 12, 47, 16, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 26, 10, 0, 0, 0, 
    
    -- channel=218
    49, 51, 42, 46, 45, 37, 31, 38, 24, 18, 28, 13, 23, 0, 17, 
    34, 43, 35, 26, 23, 22, 18, 23, 19, 24, 5, 41, 22, 0, 15, 
    19, 14, 10, 17, 15, 16, 17, 22, 21, 15, 19, 14, 19, 5, 25, 
    8, 11, 12, 16, 14, 14, 14, 25, 29, 26, 44, 0, 5, 14, 19, 
    7, 11, 11, 14, 8, 18, 12, 9, 10, 60, 48, 0, 8, 17, 13, 
    9, 12, 14, 15, 0, 2, 20, 31, 12, 0, 15, 100, 0, 13, 10, 
    12, 13, 18, 1, 12, 0, 5, 0, 0, 0, 0, 111, 29, 0, 0, 
    11, 14, 0, 24, 22, 0, 18, 0, 24, 27, 22, 89, 31, 0, 0, 
    11, 0, 28, 0, 23, 0, 0, 0, 20, 12, 47, 65, 0, 11, 4, 
    0, 0, 93, 0, 22, 0, 0, 0, 11, 36, 0, 41, 32, 21, 34, 
    0, 0, 35, 14, 4, 0, 0, 8, 59, 9, 0, 0, 22, 25, 26, 
    3, 0, 0, 35, 0, 0, 0, 20, 97, 0, 13, 0, 0, 58, 0, 
    1, 0, 0, 29, 0, 12, 0, 15, 98, 0, 34, 4, 0, 35, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 5, 0, 6, 22, 0, 0, 0, 
    2, 9, 0, 21, 1, 1, 6, 4, 4, 0, 0, 8, 0, 0, 0, 
    
    -- channel=219
    17, 32, 23, 34, 28, 32, 25, 32, 24, 7, 13, 10, 9, 32, 17, 
    34, 33, 39, 35, 29, 31, 23, 25, 23, 20, 5, 13, 9, 13, 15, 
    32, 35, 38, 30, 24, 22, 19, 16, 15, 19, 0, 43, 22, 0, 9, 
    22, 24, 23, 24, 22, 18, 13, 9, 13, 14, 0, 36, 18, 14, 17, 
    20, 25, 27, 23, 23, 7, 5, 10, 2, 0, 11, 43, 21, 23, 17, 
    22, 26, 25, 22, 15, 0, 0, 18, 14, 10, 0, 105, 23, 16, 22, 
    24, 26, 19, 17, 0, 9, 0, 43, 0, 16, 0, 35, 56, 0, 35, 
    29, 25, 8, 13, 0, 18, 0, 0, 0, 0, 0, 23, 43, 13, 0, 
    27, 10, 15, 2, 4, 6, 39, 0, 0, 0, 0, 109, 0, 0, 0, 
    24, 0, 60, 4, 52, 7, 22, 0, 0, 29, 7, 29, 0, 0, 9, 
    17, 0, 9, 4, 41, 0, 0, 0, 0, 80, 8, 0, 13, 9, 52, 
    0, 35, 0, 35, 0, 0, 0, 0, 15, 0, 4, 10, 0, 28, 36, 
    0, 0, 0, 58, 0, 0, 0, 0, 45, 0, 2, 37, 0, 76, 6, 
    0, 0, 0, 45, 0, 6, 15, 24, 33, 0, 2, 30, 0, 32, 3, 
    1, 0, 0, 0, 4, 0, 0, 1, 3, 0, 9, 37, 1, 2, 0, 
    
    -- channel=220
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 37, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 8, 30, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 42, 95, 108, 122, 116, 71, 0, 24, 0, 
    0, 0, 0, 0, 0, 26, 45, 18, 5, 0, 85, 177, 0, 9, 0, 
    0, 0, 0, 0, 28, 9, 37, 0, 0, 49, 123, 192, 70, 0, 6, 
    0, 0, 0, 16, 60, 0, 0, 95, 138, 135, 156, 85, 0, 0, 73, 
    0, 0, 103, 4, 30, 0, 0, 105, 114, 146, 122, 130, 74, 94, 103, 
    0, 70, 122, 33, 1, 0, 0, 108, 159, 56, 0, 24, 129, 112, 85, 
    0, 1, 73, 47, 0, 6, 16, 120, 180, 6, 16, 0, 74, 111, 0, 
    0, 11, 55, 34, 0, 43, 47, 103, 157, 2, 45, 0, 31, 72, 0, 
    0, 8, 54, 42, 26, 52, 62, 66, 94, 2, 41, 18, 0, 0, 0, 
    0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 41, 13, 0, 0, 0, 
    
    -- channel=221
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 43, 32, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 29, 34, 22, 31, 53, 7, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 2, 55, 42, 11, 0, 0, 
    0, 0, 0, 21, 21, 22, 31, 40, 51, 62, 45, 6, 0, 0, 19, 
    0, 0, 0, 27, 14, 20, 42, 63, 64, 62, 80, 15, 9, 38, 34, 
    0, 40, 49, 21, 12, 15, 37, 63, 56, 53, 38, 88, 63, 58, 36, 
    0, 16, 48, 16, 11, 34, 62, 59, 37, 16, 14, 37, 64, 31, 6, 
    0, 20, 50, 17, 21, 29, 44, 60, 29, 25, 9, 10, 57, 29, 0, 
    0, 8, 49, 48, 64, 82, 84, 85, 61, 34, 29, 9, 27, 17, 1, 
    0, 0, 17, 7, 14, 14, 13, 12, 8, 24, 25, 13, 4, 4, 5, 
    
    -- channel=222
    2, 16, 35, 35, 31, 22, 24, 10, 10, 36, 4, 0, 0, 0, 0, 
    24, 10, 12, 10, 7, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 18, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 32, 56, 0, 0, 5, 0, 0, 
    0, 0, 0, 0, 0, 35, 65, 43, 30, 0, 63, 0, 0, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 26, 0, 0, 0, 
    0, 0, 0, 13, 0, 1, 0, 20, 52, 69, 55, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 65, 44, 66, 96, 0, 0, 4, 25, 
    0, 92, 0, 0, 0, 0, 0, 43, 55, 29, 45, 133, 36, 41, 31, 
    0, 0, 10, 0, 0, 0, 20, 25, 0, 0, 0, 19, 41, 0, 0, 
    0, 0, 16, 0, 0, 0, 13, 38, 0, 0, 0, 0, 69, 0, 0, 
    0, 0, 27, 0, 60, 114, 125, 127, 46, 4, 0, 0, 14, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=223
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 39, 50, 27, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 39, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 24, 14, 29, 0, 30, 29, 0, 0, 
    0, 0, 0, 0, 3, 0, 7, 84, 79, 0, 0, 0, 0, 12, 22, 
    0, 0, 14, 0, 0, 14, 8, 0, 0, 0, 0, 45, 20, 8, 0, 
    0, 0, 17, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 12, 30, 8, 0, 0, 21, 16, 0, 0, 0, 0, 
    0, 6, 0, 11, 16, 0, 0, 0, 2, 13, 9, 0, 0, 1, 3, 
    0, 0, 0, 40, 34, 34, 6, 0, 15, 0, 16, 4, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 13, 1, 9, 3, 
    0, 12, 44, 31, 20, 22, 21, 18, 17, 0, 0, 7, 8, 9, 8, 
    
    -- channel=224
    34, 31, 37, 33, 45, 53, 40, 32, 23, 23, 19, 12, 8, 7, 4, 
    33, 30, 33, 32, 44, 61, 59, 49, 30, 22, 23, 23, 23, 22, 19, 
    32, 30, 22, 33, 43, 54, 59, 70, 64, 45, 39, 40, 34, 27, 23, 
    31, 31, 17, 19, 47, 55, 59, 65, 70, 69, 60, 46, 37, 28, 27, 
    49, 57, 40, 21, 47, 66, 65, 57, 70, 73, 77, 67, 50, 42, 41, 
    70, 73, 40, 17, 44, 66, 66, 65, 68, 66, 71, 72, 64, 51, 42, 
    66, 66, 61, 22, 38, 64, 67, 71, 70, 60, 63, 76, 62, 47, 28, 
    67, 71, 68, 58, 23, 46, 55, 70, 80, 66, 62, 67, 62, 44, 38, 
    75, 83, 85, 73, 82, 58, 65, 59, 79, 69, 67, 64, 66, 53, 29, 
    102, 110, 100, 83, 81, 61, 65, 66, 79, 75, 74, 66, 65, 37, 19, 
    117, 105, 48, 67, 75, 65, 68, 61, 76, 76, 66, 66, 61, 41, 17, 
    84, 72, 60, 42, 34, 51, 68, 29, 54, 68, 67, 61, 47, 49, 29, 
    55, 48, 48, 50, 42, 40, 49, 50, 52, 74, 71, 64, 51, 42, 43, 
    43, 48, 47, 40, 39, 41, 37, 48, 55, 63, 68, 64, 53, 38, 41, 
    36, 32, 34, 27, 31, 42, 44, 35, 32, 37, 44, 48, 40, 30, 26, 
    
    -- channel=225
    23, 23, 20, 21, 29, 37, 30, 25, 25, 25, 24, 24, 25, 26, 27, 
    22, 23, 21, 28, 41, 46, 49, 44, 29, 28, 32, 35, 39, 35, 32, 
    22, 22, 19, 35, 47, 59, 61, 62, 55, 38, 36, 31, 26, 20, 19, 
    26, 25, 24, 45, 60, 61, 66, 68, 56, 41, 40, 29, 22, 25, 30, 
    38, 42, 28, 51, 60, 60, 65, 69, 69, 67, 61, 51, 33, 32, 35, 
    22, 16, 12, 47, 55, 58, 54, 64, 65, 71, 69, 60, 39, 26, 24, 
    9, 9, 16, 32, 34, 46, 60, 65, 59, 63, 67, 68, 41, 21, 15, 
    19, 20, 18, 36, 45, 51, 53, 64, 62, 62, 69, 68, 50, 34, 30, 
    24, 22, 30, 40, 35, 30, 41, 62, 58, 59, 68, 71, 61, 45, 20, 
    33, 23, 7, 14, 23, 24, 39, 61, 63, 62, 66, 71, 62, 33, 24, 
    0, 0, 0, 2, 34, 34, 46, 51, 60, 59, 56, 65, 59, 39, 31, 
    0, 0, 17, 32, 37, 58, 51, 39, 45, 56, 58, 59, 50, 34, 31, 
    10, 12, 12, 25, 40, 50, 41, 47, 60, 64, 54, 56, 53, 35, 31, 
    22, 28, 26, 19, 21, 30, 44, 45, 53, 44, 39, 55, 47, 36, 29, 
    22, 18, 24, 30, 32, 29, 36, 33, 37, 38, 41, 37, 35, 31, 26, 
    
    -- channel=226
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    16, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 15, 9, 
    10, 7, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 11, 0, 
    1, 7, 7, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 22, 13, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 55, 59, 0, 22, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    51, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 7, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 15, 
    0, 0, 0, 0, 10, 11, 0, 0, 0, 0, 0, 0, 0, 4, 8, 
    
    -- channel=227
    10, 11, 6, 11, 19, 23, 21, 13, 11, 11, 10, 10, 8, 4, 5, 
    10, 12, 11, 13, 28, 33, 33, 28, 17, 11, 10, 6, 2, 0, 2, 
    12, 12, 18, 14, 39, 42, 48, 44, 19, 7, 9, 12, 10, 11, 14, 
    11, 9, 13, 25, 42, 44, 45, 46, 44, 35, 24, 26, 12, 11, 11, 
    0, 0, 19, 25, 37, 28, 36, 49, 53, 49, 46, 36, 14, 11, 11, 
    4, 11, 34, 24, 27, 28, 48, 51, 48, 52, 56, 45, 24, 17, 19, 
    14, 14, 14, 21, 29, 27, 46, 45, 42, 48, 55, 44, 35, 24, 24, 
    10, 8, 16, 12, 18, 14, 36, 41, 41, 47, 53, 51, 43, 26, 14, 
    6, 2, 4, 16, 18, 28, 25, 44, 45, 48, 50, 55, 42, 27, 22, 
    0, 0, 17, 37, 33, 47, 30, 50, 46, 44, 47, 55, 44, 31, 16, 
    9, 22, 48, 57, 46, 55, 46, 42, 43, 44, 47, 54, 39, 18, 17, 
    33, 38, 24, 22, 41, 46, 27, 32, 46, 43, 39, 44, 36, 17, 22, 
    23, 16, 16, 13, 18, 13, 25, 36, 34, 29, 37, 45, 37, 25, 21, 
    15, 12, 19, 24, 20, 19, 23, 32, 31, 32, 42, 44, 43, 25, 20, 
    17, 22, 22, 19, 12, 18, 22, 23, 22, 23, 24, 27, 27, 20, 21, 
    
    -- channel=228
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=229
    0, 0, 0, 6, 6, 0, 0, 1, 0, 0, 4, 3, 0, 0, 0, 
    0, 0, 0, 6, 2, 18, 4, 0, 2, 0, 0, 0, 0, 0, 0, 
    4, 1, 20, 10, 7, 2, 10, 0, 0, 0, 0, 0, 0, 4, 9, 
    0, 0, 0, 0, 1, 0, 0, 0, 9, 16, 0, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 5, 0, 0, 0, 
    12, 8, 0, 0, 0, 27, 10, 0, 0, 0, 0, 0, 8, 13, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 8, 30, 
    0, 0, 29, 17, 29, 10, 3, 0, 0, 0, 0, 0, 7, 10, 0, 
    0, 14, 70, 52, 44, 50, 30, 21, 1, 7, 9, 0, 0, 0, 0, 
    111, 93, 6, 1, 2, 12, 0, 0, 7, 0, 0, 0, 0, 0, 0, 
    29, 29, 8, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 20, 40, 20, 0, 0, 0, 7, 27, 32, 7, 10, 6, 6, 
    26, 36, 11, 0, 0, 0, 0, 3, 0, 0, 10, 18, 6, 0, 3, 
    
    -- channel=230
    37, 35, 31, 34, 24, 29, 30, 23, 26, 22, 14, 9, 4, 1, 3, 
    36, 37, 32, 8, 24, 8, 20, 18, 13, 17, 18, 20, 25, 30, 28, 
    29, 30, 24, 1, 3, 1, 0, 0, 14, 43, 43, 40, 32, 29, 18, 
    26, 30, 37, 0, 0, 4, 4, 6, 4, 5, 26, 31, 25, 25, 18, 
    58, 78, 106, 11, 2, 14, 38, 24, 7, 3, 0, 22, 29, 29, 29, 
    84, 82, 98, 17, 18, 15, 26, 23, 19, 12, 8, 6, 20, 31, 33, 
    71, 69, 74, 73, 6, 5, 26, 14, 23, 27, 14, 1, 26, 22, 26, 
    66, 73, 84, 59, 85, 19, 38, 14, 30, 39, 17, 8, 16, 14, 21, 
    80, 90, 119, 109, 106, 93, 45, 28, 22, 34, 25, 18, 10, 23, 11, 
    144, 158, 131, 134, 62, 86, 25, 31, 22, 30, 30, 23, 12, 15, 0, 
    149, 150, 81, 26, 22, 9, 16, 5, 21, 26, 22, 17, 14, 21, 10, 
    94, 58, 59, 60, 31, 0, 18, 25, 0, 8, 29, 37, 14, 3, 25, 
    37, 38, 33, 39, 44, 37, 11, 20, 8, 18, 53, 35, 32, 3, 8, 
    27, 32, 30, 11, 0, 12, 8, 13, 0, 1, 5, 21, 23, 0, 0, 
    22, 0, 0, 0, 0, 7, 15, 2, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=231
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=232
    0, 0, 8, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    9, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    21, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 5, 
    21, 20, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    18, 22, 13, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 33, 24, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    40, 44, 36, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    52, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 24, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    9, 8, 10, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 4, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=233
    0, 0, 0, 3, 5, 11, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 15, 22, 25, 12, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 0, 14, 19, 29, 28, 16, 3, 8, 12, 12, 12, 11, 
    0, 0, 0, 0, 12, 14, 19, 36, 34, 27, 16, 20, 10, 7, 10, 
    0, 0, 19, 8, 14, 21, 25, 30, 41, 36, 33, 31, 19, 20, 24, 
    12, 17, 39, 0, 9, 7, 24, 26, 33, 40, 43, 33, 27, 36, 33, 
    15, 15, 19, 0, 10, 31, 39, 32, 29, 26, 40, 29, 30, 32, 26, 
    5, 7, 18, 34, 21, 0, 26, 33, 33, 29, 34, 30, 30, 17, 10, 
    11, 7, 6, 0, 34, 22, 31, 35, 29, 26, 28, 33, 27, 23, 39, 
    5, 25, 49, 60, 42, 64, 26, 38, 27, 23, 30, 35, 26, 23, 25, 
    31, 42, 32, 30, 24, 44, 27, 40, 36, 32, 38, 32, 25, 28, 26, 
    54, 34, 13, 32, 15, 20, 17, 6, 15, 18, 22, 30, 32, 36, 31, 
    10, 12, 5, 8, 29, 17, 33, 21, 14, 14, 22, 26, 32, 32, 41, 
    3, 8, 24, 32, 26, 24, 17, 31, 32, 25, 35, 25, 35, 40, 37, 
    24, 30, 27, 26, 25, 35, 26, 35, 36, 30, 28, 37, 39, 34, 38, 
    
    -- channel=234
    0, 0, 0, 0, 0, 6, 2, 0, 0, 0, 1, 3, 8, 11, 18, 
    0, 0, 0, 0, 2, 0, 9, 11, 7, 9, 18, 24, 22, 18, 18, 
    0, 0, 0, 3, 12, 18, 14, 24, 21, 11, 10, 10, 8, 5, 9, 
    0, 1, 28, 14, 18, 26, 32, 26, 22, 2, 3, 9, 12, 13, 21, 
    15, 8, 4, 26, 14, 8, 19, 28, 29, 24, 14, 18, 15, 28, 30, 
    0, 0, 0, 24, 26, 7, 4, 23, 25, 30, 29, 16, 17, 26, 25, 
    0, 0, 0, 46, 1, 0, 8, 16, 15, 25, 27, 18, 20, 12, 11, 
    0, 0, 0, 0, 40, 26, 24, 20, 7, 14, 25, 24, 15, 14, 23, 
    0, 0, 15, 18, 8, 23, 17, 23, 3, 9, 23, 24, 12, 11, 15, 
    0, 0, 0, 0, 0, 0, 0, 27, 6, 5, 14, 21, 14, 28, 42, 
    0, 0, 0, 0, 0, 0, 7, 8, 7, 4, 11, 25, 23, 36, 40, 
    0, 0, 4, 0, 13, 14, 13, 22, 10, 14, 16, 20, 30, 22, 49, 
    0, 0, 0, 1, 10, 13, 0, 23, 10, 6, 2, 8, 39, 33, 31, 
    2, 0, 0, 0, 17, 28, 24, 11, 14, 0, 0, 10, 20, 37, 28, 
    0, 6, 26, 38, 34, 21, 28, 35, 39, 32, 16, 13, 30, 42, 40, 
    
    -- channel=235
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=236
    14, 11, 22, 9, 19, 23, 15, 10, 10, 14, 9, 5, 8, 16, 11, 
    14, 10, 22, 6, 23, 38, 22, 26, 12, 14, 19, 23, 27, 28, 19, 
    14, 11, 3, 22, 20, 39, 43, 45, 45, 33, 23, 21, 15, 6, 0, 
    17, 20, 0, 31, 37, 47, 50, 51, 50, 37, 26, 8, 12, 6, 10, 
    43, 48, 7, 0, 46, 60, 49, 31, 47, 50, 50, 31, 24, 16, 22, 
    31, 20, 0, 0, 38, 76, 34, 26, 47, 43, 51, 52, 34, 16, 9, 
    10, 6, 0, 0, 39, 46, 25, 44, 53, 32, 36, 61, 32, 17, 0, 
    21, 24, 16, 0, 0, 59, 31, 54, 57, 28, 33, 51, 40, 24, 12, 
    33, 38, 30, 22, 19, 9, 29, 31, 54, 31, 37, 40, 52, 26, 0, 
    55, 47, 0, 0, 15, 0, 34, 13, 56, 42, 41, 34, 46, 3, 5, 
    11, 0, 0, 0, 22, 0, 31, 22, 50, 42, 32, 33, 38, 22, 4, 
    0, 0, 0, 1, 2, 39, 54, 11, 45, 46, 45, 30, 19, 36, 0, 
    0, 5, 4, 15, 0, 26, 45, 15, 48, 64, 44, 25, 11, 28, 17, 
    12, 23, 13, 0, 5, 20, 27, 27, 38, 51, 32, 26, 20, 11, 29, 
    6, 0, 6, 10, 26, 28, 19, 5, 20, 26, 37, 28, 12, 18, 14, 
    
    -- channel=237
    20, 20, 13, 18, 12, 5, 9, 14, 16, 13, 14, 15, 12, 7, 9, 
    21, 20, 13, 20, 3, 0, 0, 0, 9, 10, 4, 0, 0, 0, 0, 
    21, 20, 20, 4, 8, 0, 0, 0, 0, 0, 0, 0, 1, 5, 6, 
    16, 15, 16, 3, 2, 0, 0, 0, 0, 0, 0, 4, 0, 2, 0, 
    0, 0, 3, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 18, 43, 18, 0, 0, 11, 3, 0, 0, 0, 0, 0, 0, 0, 
    25, 25, 26, 14, 5, 0, 2, 0, 0, 0, 0, 0, 0, 0, 8, 
    17, 12, 11, 13, 1, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    9, 9, 9, 3, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 
    0, 0, 29, 33, 25, 22, 0, 0, 0, 7, 0, 0, 0, 0, 0, 
    32, 38, 70, 51, 17, 24, 2, 7, 0, 0, 2, 1, 0, 0, 0, 
    60, 73, 33, 20, 26, 9, 0, 8, 9, 4, 0, 0, 0, 0, 0, 
    32, 25, 23, 5, 3, 0, 0, 2, 0, 0, 3, 7, 0, 0, 0, 
    13, 0, 0, 4, 0, 0, 0, 0, 0, 0, 16, 12, 0, 0, 0, 
    2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=238
    10, 14, 0, 13, 18, 16, 29, 15, 18, 18, 18, 20, 16, 9, 17, 
    10, 18, 10, 12, 29, 17, 25, 27, 21, 15, 18, 14, 8, 7, 16, 
    12, 13, 36, 2, 35, 29, 34, 31, 0, 8, 12, 21, 21, 26, 31, 
    11, 8, 44, 27, 24, 33, 33, 33, 37, 16, 13, 38, 22, 27, 25, 
    0, 0, 66, 44, 24, 0, 22, 50, 43, 38, 27, 25, 17, 30, 29, 
    0, 11, 78, 46, 20, 0, 44, 45, 36, 46, 51, 20, 16, 32, 40, 
    12, 17, 23, 87, 33, 0, 41, 31, 24, 45, 52, 17, 33, 25, 43, 
    5, 5, 30, 5, 66, 8, 52, 26, 17, 45, 49, 39, 30, 22, 28, 
    0, 0, 7, 56, 26, 76, 22, 51, 21, 38, 43, 48, 17, 27, 52, 
    0, 0, 23, 79, 21, 78, 15, 59, 23, 27, 37, 53, 27, 55, 40, 
    10, 47, 116, 72, 35, 51, 34, 28, 28, 30, 43, 52, 35, 29, 48, 
    44, 53, 40, 32, 76, 29, 2, 58, 26, 18, 24, 46, 49, 14, 61, 
    29, 16, 21, 17, 31, 29, 15, 41, 15, 0, 30, 40, 49, 37, 26, 
    17, 15, 31, 43, 32, 30, 28, 40, 32, 22, 21, 37, 51, 41, 32, 
    33, 41, 40, 41, 18, 26, 41, 47, 43, 39, 30, 38, 50, 39, 42, 
    
    -- channel=239
    10, 7, 3, 8, 0, 12, 0, 8, 8, 8, 4, 5, 4, 0, 3, 
    10, 12, 7, 0, 6, 0, 17, 0, 0, 8, 3, 5, 8, 8, 8, 
    5, 13, 0, 0, 0, 0, 0, 0, 4, 9, 13, 9, 3, 6, 2, 
    7, 9, 20, 0, 0, 0, 0, 0, 0, 0, 3, 0, 4, 4, 4, 
    15, 23, 46, 0, 0, 14, 12, 0, 0, 0, 0, 8, 2, 2, 1, 
    14, 13, 76, 0, 15, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    11, 13, 37, 13, 0, 0, 18, 1, 3, 0, 0, 0, 0, 0, 2, 
    12, 12, 13, 46, 48, 0, 2, 0, 5, 11, 0, 0, 8, 0, 2, 
    15, 18, 44, 0, 62, 18, 33, 0, 0, 10, 2, 0, 0, 0, 0, 
    30, 30, 12, 90, 5, 76, 0, 0, 0, 2, 6, 2, 0, 0, 0, 
    28, 35, 0, 0, 0, 5, 0, 1, 1, 0, 2, 0, 0, 18, 0, 
    18, 11, 30, 38, 0, 0, 14, 0, 0, 0, 2, 8, 0, 0, 5, 
    6, 7, 4, 4, 35, 6, 0, 15, 0, 0, 16, 2, 9, 0, 11, 
    2, 0, 0, 0, 0, 10, 0, 0, 0, 0, 6, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=240
    5, 6, 8, 13, 8, 14, 18, 10, 8, 8, 8, 6, 5, 3, 3, 
    4, 6, 10, 3, 13, 16, 17, 18, 16, 6, 9, 7, 7, 10, 14, 
    5, 6, 20, 2, 8, 11, 15, 21, 19, 11, 18, 24, 28, 30, 30, 
    4, 3, 10, 3, 0, 5, 11, 25, 34, 30, 17, 33, 30, 25, 27, 
    0, 0, 33, 9, 5, 0, 10, 20, 28, 27, 24, 31, 35, 39, 42, 
    19, 25, 39, 12, 1, 0, 14, 13, 19, 24, 29, 23, 42, 55, 55, 
    25, 26, 22, 25, 19, 11, 18, 12, 15, 17, 26, 16, 42, 51, 49, 
    14, 18, 32, 28, 28, 0, 22, 18, 15, 14, 17, 20, 26, 30, 31, 
    17, 14, 14, 26, 32, 46, 26, 26, 12, 9, 11, 17, 14, 35, 59, 
    16, 33, 54, 54, 30, 58, 21, 28, 9, 5, 11, 15, 17, 44, 54, 
    40, 55, 54, 33, 26, 29, 24, 25, 15, 17, 21, 17, 26, 43, 58, 
    56, 43, 29, 22, 14, 7, 12, 18, 6, 7, 12, 19, 43, 49, 59, 
    24, 20, 19, 21, 26, 15, 21, 22, 0, 0, 10, 16, 43, 56, 54, 
    17, 21, 34, 46, 41, 38, 24, 30, 22, 20, 14, 9, 39, 59, 57, 
    37, 44, 44, 49, 49, 47, 43, 53, 52, 42, 32, 39, 48, 60, 64, 
    
    -- channel=241
    15, 14, 20, 23, 13, 0, 3, 11, 8, 8, 10, 9, 6, 6, 0, 
    15, 10, 16, 17, 0, 0, 0, 0, 3, 4, 0, 0, 0, 0, 0, 
    16, 13, 14, 14, 0, 0, 0, 0, 0, 0, 0, 0, 6, 14, 14, 
    9, 8, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 10, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 
    37, 35, 18, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 13, 17, 
    23, 20, 18, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    3, 24, 61, 18, 25, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    55, 53, 39, 29, 13, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    88, 77, 23, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    35, 34, 26, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 11, 13, 20, 16, 0, 0, 0, 0, 0, 4, 0, 0, 0, 4, 
    16, 20, 6, 0, 4, 3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    
    -- channel=242
    0, 0, 11, 1, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 24, 3, 5, 11, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 8, 0, 0, 8, 0, 25, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 41, 0, 0, 0, 0, 16, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 29, 0, 0, 0, 0, 0, 19, 11, 0, 0, 
    6, 0, 0, 0, 21, 63, 0, 1, 5, 0, 0, 19, 0, 18, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 9, 0, 0, 0, 11, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 0, 14, 0, 0, 0, 14, 0, 0, 
    0, 0, 0, 0, 24, 0, 22, 0, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 26, 30, 22, 14, 24, 12, 4, 0, 0, 0, 0, 0, 
    25, 27, 0, 0, 0, 19, 26, 0, 40, 21, 0, 0, 0, 27, 0, 
    11, 13, 5, 0, 0, 0, 32, 0, 6, 28, 0, 0, 0, 0, 11, 
    2, 0, 0, 5, 14, 2, 0, 0, 3, 34, 48, 0, 0, 0, 15, 
    2, 11, 8, 0, 13, 14, 0, 0, 0, 0, 15, 19, 0, 3, 0, 
    
    -- channel=243
    0, 0, 0, 1, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 12, 7, 0, 3, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    5, 4, 0, 0, 13, 26, 0, 0, 0, 0, 0, 0, 0, 15, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 0, 0, 0, 17, 0, 4, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 16, 63, 39, 41, 19, 22, 0, 0, 0, 0, 0, 0, 0, 
    67, 80, 12, 0, 0, 14, 0, 0, 25, 4, 0, 0, 0, 5, 0, 
    30, 18, 12, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 3, 
    2, 0, 5, 25, 25, 0, 0, 0, 0, 18, 34, 0, 0, 4, 11, 
    10, 28, 19, 2, 4, 3, 0, 1, 0, 0, 8, 16, 7, 5, 9, 
    
    -- channel=244
    16, 13, 16, 13, 7, 4, 5, 5, 4, 2, 0, 0, 0, 0, 0, 
    15, 11, 14, 0, 1, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 11, 5, 0, 0, 0, 0, 0, 0, 5, 2, 1, 2, 0, 0, 
    9, 8, 0, 0, 0, 0, 0, 0, 0, 6, 4, 0, 0, 0, 0, 
    18, 27, 13, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 41, 8, 0, 0, 14, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 34, 24, 0, 14, 10, 0, 0, 3, 0, 0, 0, 0, 0, 0, 
    32, 33, 33, 11, 0, 6, 0, 0, 11, 0, 0, 0, 0, 0, 0, 
    36, 38, 36, 29, 19, 4, 3, 0, 12, 3, 0, 0, 1, 0, 0, 
    66, 73, 71, 25, 32, 4, 7, 0, 10, 9, 1, 0, 0, 0, 0, 
    79, 72, 1, 24, 23, 0, 9, 0, 5, 8, 0, 0, 0, 0, 0, 
    57, 38, 25, 8, 0, 0, 8, 0, 3, 6, 7, 0, 0, 0, 0, 
    28, 19, 13, 13, 0, 0, 0, 0, 0, 14, 14, 1, 0, 0, 0, 
    7, 9, 4, 0, 0, 0, 0, 0, 0, 9, 12, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=245
    1, 5, 0, 0, 0, 2, 16, 6, 10, 6, 9, 12, 8, 0, 10, 
    1, 10, 0, 0, 4, 0, 8, 10, 10, 2, 6, 5, 2, 0, 9, 
    1, 3, 19, 0, 6, 0, 0, 0, 0, 0, 1, 6, 6, 10, 15, 
    0, 0, 42, 0, 0, 0, 0, 0, 0, 0, 0, 20, 7, 13, 8, 
    0, 0, 67, 37, 0, 0, 0, 20, 5, 0, 0, 5, 0, 8, 7, 
    0, 0, 88, 39, 3, 0, 12, 21, 3, 8, 12, 0, 0, 4, 17, 
    0, 1, 16, 103, 0, 0, 19, 0, 0, 17, 19, 0, 6, 0, 26, 
    0, 0, 12, 8, 85, 0, 23, 0, 0, 24, 20, 5, 2, 0, 11, 
    0, 0, 6, 45, 24, 68, 0, 21, 0, 15, 17, 21, 0, 4, 23, 
    0, 0, 3, 95, 0, 74, 0, 40, 0, 1, 10, 28, 0, 34, 14, 
    0, 33, 113, 27, 0, 17, 2, 0, 0, 0, 10, 25, 9, 10, 25, 
    23, 30, 45, 25, 53, 0, 0, 38, 0, 0, 0, 21, 23, 0, 47, 
    12, 0, 1, 0, 30, 15, 0, 28, 0, 0, 10, 14, 34, 0, 0, 
    0, 0, 5, 13, 0, 4, 1, 7, 0, 0, 0, 12, 23, 9, 0, 
    8, 9, 6, 12, 0, 0, 12, 17, 8, 5, 0, 0, 17, 1, 7, 
    
    -- channel=246
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 11, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 25, 30, 30, 22, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 3, 0, 0, 0, 0, 
    0, 3, 26, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    42, 45, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 37, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 36, 53, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    42, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=247
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 20, 33, 40, 40, 34, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 31, 22, 17, 7, 0, 0, 
    0, 2, 40, 7, 0, 1, 6, 0, 0, 0, 0, 0, 1, 8, 11, 
    55, 67, 66, 15, 0, 0, 20, 16, 0, 0, 0, 0, 8, 23, 27, 
    13, 0, 11, 26, 15, 3, 0, 0, 1, 2, 0, 0, 0, 7, 11, 
    0, 0, 0, 80, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 
    0, 8, 8, 0, 91, 47, 25, 0, 0, 5, 0, 0, 0, 0, 11, 
    11, 26, 77, 96, 34, 59, 3, 15, 0, 0, 5, 2, 0, 0, 0, 
    83, 54, 0, 0, 0, 0, 0, 3, 0, 0, 0, 1, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 30, 
    0, 0, 0, 0, 8, 0, 0, 23, 0, 0, 5, 11, 5, 0, 32, 
    0, 0, 0, 0, 10, 28, 0, 0, 0, 0, 10, 0, 20, 3, 0, 
    0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 3, 0, 0, 0, 0, 0, 0, 1, 0, 
    
    -- channel=248
    39, 38, 29, 41, 26, 27, 34, 32, 33, 27, 23, 21, 14, 6, 11, 
    38, 41, 31, 13, 26, 1, 22, 16, 20, 21, 18, 22, 25, 29, 33, 
    32, 35, 35, 7, 3, 0, 0, 0, 8, 40, 40, 41, 37, 38, 30, 
    28, 28, 43, 0, 0, 0, 0, 0, 0, 3, 26, 33, 31, 36, 27, 
    43, 61, 112, 24, 0, 0, 17, 7, 0, 0, 0, 16, 26, 38, 35, 
    73, 79, 121, 27, 7, 0, 12, 14, 0, 0, 0, 0, 9, 36, 41, 
    70, 72, 82, 92, 4, 0, 26, 1, 3, 11, 0, 0, 12, 21, 37, 
    61, 67, 85, 75, 92, 0, 29, 0, 9, 28, 4, 0, 2, 4, 29, 
    67, 69, 102, 96, 104, 98, 44, 19, 0, 21, 10, 1, 0, 17, 29, 
    117, 135, 136, 172, 52, 107, 12, 33, 2, 13, 16, 11, 0, 19, 9, 
    142, 159, 113, 38, 24, 17, 7, 3, 6, 12, 12, 6, 1, 22, 19, 
    116, 83, 92, 67, 32, 0, 0, 20, 0, 0, 11, 22, 11, 0, 41, 
    55, 46, 41, 46, 65, 38, 0, 25, 0, 0, 36, 23, 28, 1, 17, 
    31, 37, 39, 29, 8, 24, 5, 15, 1, 0, 5, 14, 16, 4, 0, 
    35, 18, 9, 10, 0, 13, 23, 14, 2, 3, 0, 4, 13, 0, 3, 
    
    -- channel=249
    0, 0, 0, 5, 5, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 4, 3, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 16, 7, 11, 0, 8, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 4, 0, 0, 11, 22, 9, 0, 0, 0, 2, 0, 0, 7, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    0, 0, 17, 15, 25, 17, 4, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 8, 51, 64, 36, 52, 14, 22, 0, 1, 8, 0, 0, 0, 0, 
    86, 83, 12, 2, 7, 13, 0, 0, 19, 0, 0, 0, 0, 0, 0, 
    28, 19, 8, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 29, 16, 0, 0, 5, 1, 18, 36, 6, 4, 1, 0, 
    16, 28, 10, 0, 0, 0, 0, 0, 0, 0, 3, 15, 5, 0, 0, 
    
    -- channel=250
    15, 16, 6, 14, 20, 26, 31, 17, 17, 15, 14, 13, 9, 4, 11, 
    15, 18, 11, 14, 33, 27, 37, 37, 21, 13, 18, 20, 20, 18, 21, 
    14, 13, 22, 7, 34, 39, 42, 42, 28, 28, 25, 26, 20, 16, 16, 
    14, 12, 30, 29, 35, 40, 42, 43, 45, 26, 27, 33, 16, 21, 20, 
    21, 28, 64, 45, 37, 21, 47, 59, 53, 52, 42, 37, 21, 28, 28, 
    23, 26, 55, 45, 32, 26, 53, 53, 47, 54, 58, 35, 21, 23, 27, 
    17, 20, 26, 70, 23, 11, 51, 46, 41, 53, 59, 39, 33, 14, 22, 
    19, 22, 36, 27, 71, 27, 53, 43, 44, 58, 58, 52, 34, 22, 23, 
    21, 19, 40, 77, 47, 68, 28, 63, 42, 51, 57, 60, 37, 31, 21, 
    38, 40, 43, 70, 29, 60, 27, 67, 47, 48, 55, 66, 43, 31, 13, 
    33, 48, 72, 32, 30, 40, 37, 29, 45, 45, 48, 57, 41, 22, 30, 
    24, 13, 31, 34, 55, 33, 20, 47, 24, 31, 41, 53, 41, 11, 39, 
    17, 11, 13, 21, 39, 39, 20, 42, 37, 26, 50, 50, 47, 24, 16, 
    15, 20, 26, 20, 10, 19, 30, 36, 36, 24, 24, 43, 40, 23, 16, 
    19, 13, 13, 18, 8, 17, 31, 24, 25, 25, 22, 21, 23, 15, 17, 
    
    -- channel=251
    0, 5, 0, 5, 3, 0, 2, 0, 2, 0, 3, 5, 4, 1, 3, 
    0, 0, 0, 34, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 15, 2, 0, 0, 0, 0, 0, 0, 0, 6, 5, 9, 
    0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 3, 0, 5, 5, 
    0, 0, 0, 57, 0, 0, 0, 16, 0, 0, 0, 0, 0, 3, 2, 
    0, 0, 0, 69, 0, 0, 0, 7, 0, 1, 0, 0, 2, 0, 6, 
    1, 2, 0, 44, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 12, 
    0, 0, 0, 19, 5, 1, 0, 0, 0, 0, 1, 0, 0, 0, 3, 
    0, 0, 0, 44, 0, 0, 0, 15, 0, 0, 0, 0, 0, 13, 13, 
    0, 0, 21, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 16, 9, 
    0, 0, 95, 0, 11, 1, 4, 15, 0, 0, 0, 0, 2, 0, 17, 
    23, 20, 39, 0, 14, 2, 0, 23, 0, 0, 0, 0, 19, 0, 16, 
    13, 5, 3, 4, 2, 9, 0, 0, 0, 0, 0, 5, 15, 5, 0, 
    3, 0, 3, 14, 13, 0, 11, 0, 1, 0, 0, 2, 2, 15, 0, 
    9, 13, 7, 12, 13, 0, 7, 17, 8, 0, 0, 0, 5, 13, 4, 
    
    -- channel=252
    46, 45, 35, 48, 47, 45, 40, 39, 37, 33, 27, 24, 16, 6, 7, 
    45, 46, 39, 25, 52, 39, 54, 35, 26, 27, 17, 17, 19, 22, 26, 
    40, 43, 44, 28, 36, 30, 31, 27, 22, 44, 45, 45, 39, 40, 33, 
    36, 34, 35, 6, 27, 24, 23, 30, 25, 32, 49, 47, 31, 34, 28, 
    36, 54, 106, 39, 26, 36, 53, 47, 37, 31, 34, 44, 33, 35, 33, 
    78, 86, 125, 32, 31, 19, 52, 57, 42, 40, 37, 27, 27, 40, 41, 
    80, 79, 86, 72, 23, 42, 70, 47, 42, 49, 46, 24, 37, 33, 41, 
    68, 70, 88, 83, 82, 3, 54, 37, 52, 68, 51, 33, 37, 20, 28, 
    73, 70, 89, 80, 113, 93, 65, 52, 46, 64, 54, 47, 30, 36, 38, 
    102, 129, 146, 184, 90, 125, 46, 67, 46, 59, 60, 57, 33, 30, 5, 
    143, 161, 119, 74, 62, 68, 50, 46, 52, 57, 58, 49, 30, 27, 12, 
    146, 108, 92, 85, 56, 25, 27, 35, 20, 29, 46, 58, 30, 14, 34, 
    66, 60, 49, 51, 72, 53, 34, 47, 32, 31, 69, 62, 47, 11, 26, 
    38, 44, 54, 46, 19, 30, 20, 40, 33, 28, 52, 57, 45, 17, 8, 
    47, 33, 18, 11, 0, 23, 32, 24, 10, 15, 15, 28, 27, 2, 5, 
    
    -- channel=253
    22, 20, 19, 20, 15, 5, 7, 16, 14, 14, 14, 14, 11, 8, 4, 
    22, 20, 17, 15, 4, 2, 0, 0, 4, 8, 0, 0, 0, 0, 0, 
    22, 21, 15, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    17, 15, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 22, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 25, 23, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 17, 14, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 13, 4, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 16, 32, 26, 20, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    39, 38, 21, 31, 12, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    57, 56, 24, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 26, 21, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 6, 4, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=254
    0, 0, 0, 0, 11, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 8, 29, 18, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 14, 28, 26, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 9, 6, 18, 28, 41, 20, 12, 0, 0, 0, 
    0, 0, 0, 0, 0, 16, 1, 2, 23, 27, 39, 24, 2, 0, 0, 
    11, 27, 16, 0, 0, 14, 26, 19, 18, 15, 22, 35, 23, 4, 0, 
    35, 33, 20, 0, 6, 36, 26, 25, 22, 8, 19, 26, 22, 22, 5, 
    22, 16, 19, 4, 0, 0, 0, 17, 27, 14, 15, 20, 30, 12, 0, 
    17, 17, 0, 0, 12, 0, 14, 1, 36, 25, 13, 15, 24, 7, 8, 
    0, 16, 64, 45, 70, 44, 34, 11, 31, 29, 21, 15, 21, 1, 0, 
    69, 73, 40, 92, 61, 70, 40, 30, 30, 32, 30, 20, 10, 0, 0, 
    113, 109, 17, 4, 0, 19, 16, 0, 35, 30, 12, 11, 2, 11, 0, 
    38, 30, 23, 5, 0, 0, 20, 4, 3, 18, 15, 22, 0, 1, 6, 
    7, 1, 16, 26, 18, 0, 0, 12, 7, 32, 56, 25, 19, 0, 5, 
    9, 19, 9, 0, 0, 4, 0, 0, 0, 0, 6, 18, 5, 0, 0, 
    
    -- channel=255
    1, 2, 0, 0, 1, 14, 9, 0, 2, 1, 1, 2, 5, 8, 15, 
    2, 4, 0, 9, 4, 2, 7, 17, 8, 11, 20, 17, 9, 1, 0, 
    3, 2, 0, 0, 24, 28, 31, 30, 10, 0, 0, 0, 0, 0, 0, 
    6, 12, 34, 25, 38, 48, 44, 27, 27, 6, 0, 8, 0, 0, 0, 
    21, 6, 0, 19, 23, 13, 25, 37, 32, 31, 20, 13, 1, 0, 0, 
    0, 0, 4, 25, 34, 31, 32, 35, 34, 36, 35, 33, 5, 0, 0, 
    0, 0, 0, 40, 2, 0, 14, 30, 30, 36, 34, 28, 14, 0, 0, 
    2, 0, 0, 0, 30, 36, 25, 23, 20, 29, 37, 38, 25, 20, 4, 
    0, 16, 29, 22, 0, 7, 0, 26, 28, 33, 39, 41, 29, 1, 0, 
    0, 0, 0, 0, 0, 0, 3, 27, 32, 32, 31, 38, 32, 19, 0, 
    0, 0, 26, 24, 8, 11, 17, 11, 18, 19, 25, 43, 29, 5, 0, 
    0, 0, 0, 0, 35, 39, 21, 35, 39, 40, 27, 33, 20, 0, 3, 
    0, 0, 5, 0, 0, 0, 0, 20, 22, 25, 21, 24, 21, 1, 0, 
    6, 0, 0, 0, 0, 0, 15, 5, 6, 7, 5, 29, 19, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    
    -- channel=256
    0, 44, 86, 71, 63, 75, 75, 79, 60, 23, 74, 83, 90, 93, 90, 
    0, 23, 78, 78, 67, 60, 77, 89, 84, 34, 95, 93, 92, 95, 92, 
    0, 4, 65, 78, 91, 48, 44, 69, 63, 65, 89, 102, 99, 98, 94, 
    10, 39, 78, 69, 93, 70, 52, 36, 45, 79, 91, 118, 105, 96, 111, 
    81, 90, 95, 55, 87, 83, 71, 40, 51, 69, 93, 123, 115, 93, 111, 
    100, 99, 97, 79, 86, 78, 61, 48, 55, 70, 84, 128, 119, 101, 102, 
    102, 100, 79, 97, 71, 76, 57, 64, 59, 69, 87, 126, 127, 117, 96, 
    100, 99, 61, 98, 80, 77, 66, 64, 80, 79, 84, 100, 136, 117, 123, 
    92, 86, 73, 86, 95, 85, 73, 45, 70, 74, 79, 60, 90, 101, 127, 
    102, 93, 92, 88, 94, 97, 97, 72, 60, 84, 59, 71, 75, 69, 84, 
    110, 91, 101, 95, 99, 72, 93, 95, 79, 61, 69, 71, 74, 61, 64, 
    110, 91, 106, 99, 94, 76, 93, 90, 82, 51, 76, 70, 78, 67, 55, 
    105, 97, 108, 99, 70, 66, 95, 87, 72, 57, 72, 65, 64, 65, 59, 
    101, 93, 106, 103, 73, 75, 70, 74, 63, 51, 62, 62, 50, 63, 70, 
    91, 91, 93, 104, 88, 78, 60, 63, 44, 61, 57, 62, 53, 60, 63, 
    
    -- channel=257
    20, 28, 21, 21, 17, 27, 28, 29, 28, 20, 28, 26, 29, 31, 29, 
    21, 24, 9, 19, 15, 18, 20, 25, 15, 22, 33, 22, 22, 23, 22, 
    22, 21, 16, 21, 3, 7, 4, 0, 0, 24, 19, 14, 16, 20, 24, 
    43, 53, 46, 19, 0, 10, 27, 17, 14, 17, 7, 19, 15, 11, 17, 
    40, 45, 23, 24, 4, 0, 7, 9, 11, 13, 15, 17, 14, 22, 24, 
    25, 23, 20, 27, 13, 4, 0, 12, 12, 14, 12, 12, 17, 30, 35, 
    26, 25, 16, 12, 3, 4, 2, 23, 10, 13, 14, 14, 17, 25, 40, 
    26, 21, 10, 10, 14, 6, 9, 7, 13, 21, 7, 10, 9, 9, 29, 
    25, 19, 12, 10, 13, 17, 13, 4, 20, 18, 15, 24, 1, 0, 23, 
    30, 32, 10, 15, 4, 0, 2, 15, 23, 19, 8, 16, 28, 20, 9, 
    25, 21, 12, 13, 18, 8, 4, 3, 10, 8, 18, 20, 14, 13, 17, 
    22, 22, 14, 7, 5, 16, 15, 13, 8, 14, 24, 14, 12, 18, 18, 
    25, 27, 22, 4, 0, 3, 5, 9, 6, 17, 15, 16, 5, 12, 17, 
    26, 31, 27, 7, 11, 27, 9, 9, 10, 20, 17, 16, 15, 17, 19, 
    22, 31, 30, 2, 11, 7, 14, 13, 12, 22, 17, 17, 22, 22, 13, 
    
    -- channel=258
    0, 33, 43, 40, 26, 46, 41, 44, 18, 0, 35, 48, 52, 52, 49, 
    0, 0, 48, 47, 21, 20, 40, 43, 35, 0, 53, 41, 45, 49, 51, 
    0, 0, 48, 39, 44, 0, 15, 32, 24, 20, 42, 41, 42, 45, 43, 
    0, 0, 48, 21, 55, 11, 0, 1, 10, 45, 31, 52, 47, 35, 45, 
    8, 37, 26, 2, 46, 32, 18, 0, 10, 35, 42, 58, 40, 10, 38, 
    28, 34, 28, 6, 47, 33, 7, 0, 4, 23, 36, 64, 40, 6, 22, 
    29, 32, 25, 29, 16, 18, 4, 33, 14, 25, 27, 60, 46, 28, 21, 
    23, 35, 3, 79, 26, 24, 16, 4, 30, 32, 19, 73, 60, 38, 31, 
    6, 27, 29, 65, 28, 32, 16, 0, 49, 15, 25, 0, 59, 28, 59, 
    16, 27, 38, 38, 37, 38, 32, 15, 0, 29, 24, 27, 23, 27, 39, 
    30, 12, 40, 34, 37, 12, 42, 38, 21, 21, 17, 34, 33, 18, 23, 
    31, 6, 49, 42, 37, 36, 40, 36, 25, 1, 35, 28, 33, 16, 8, 
    25, 14, 45, 33, 13, 35, 48, 36, 24, 9, 30, 22, 28, 21, 16, 
    22, 7, 40, 37, 17, 29, 38, 26, 15, 12, 25, 15, 5, 25, 23, 
    17, 7, 32, 40, 24, 20, 18, 26, 3, 9, 17, 16, 7, 22, 24, 
    
    -- channel=259
    1, 0, 16, 25, 23, 25, 27, 25, 22, 28, 0, 14, 22, 25, 27, 
    1, 0, 14, 12, 4, 18, 15, 12, 19, 26, 0, 20, 26, 26, 26, 
    0, 0, 0, 12, 0, 21, 20, 24, 27, 5, 5, 21, 22, 20, 21, 
    8, 0, 0, 26, 0, 9, 3, 16, 10, 0, 14, 1, 7, 24, 17, 
    20, 0, 20, 32, 0, 8, 15, 21, 7, 0, 9, 8, 22, 42, 25, 
    24, 18, 28, 19, 1, 8, 20, 13, 2, 0, 8, 13, 26, 42, 36, 
    31, 23, 35, 13, 18, 10, 21, 0, 9, 2, 6, 8, 23, 26, 29, 
    35, 19, 26, 1, 13, 6, 11, 2, 7, 8, 15, 24, 12, 34, 21, 
    41, 22, 11, 3, 6, 1, 6, 23, 6, 13, 18, 19, 27, 38, 16, 
    34, 16, 10, 15, 16, 19, 6, 6, 12, 10, 26, 17, 5, 19, 21, 
    28, 29, 9, 12, 11, 24, 10, 11, 17, 27, 14, 11, 12, 23, 19, 
    28, 35, 6, 11, 16, 14, 5, 10, 17, 29, 6, 16, 11, 17, 17, 
    31, 39, 12, 13, 32, 8, 16, 19, 27, 23, 12, 16, 20, 16, 17, 
    33, 41, 18, 13, 21, 0, 24, 23, 27, 18, 15, 15, 20, 8, 13, 
    35, 38, 23, 6, 17, 25, 28, 18, 28, 8, 14, 14, 13, 11, 15, 
    
    -- channel=260
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=261
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 23, 37, 44, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 6, 0, 0, 0, 0, 0, 0, 0, 0, 8, 1, 
    0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 1, 8, 
    0, 0, 0, 0, 0, 6, 14, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 5, 0, 0, 0, 0, 0, 0, 0, 0, 16, 70, 24, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 47, 52, 13, 
    0, 0, 0, 0, 5, 26, 0, 0, 0, 0, 19, 0, 0, 0, 31, 
    0, 0, 0, 0, 0, 4, 4, 6, 0, 18, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 1, 2, 0, 0, 0, 4, 0, 2, 0, 0, 0, 
    0, 4, 0, 0, 21, 19, 0, 13, 18, 7, 0, 3, 24, 10, 0, 
    2, 5, 6, 0, 0, 0, 16, 15, 16, 10, 0, 0, 2, 0, 0, 
    24, 0, 16, 2, 0, 3, 28, 14, 15, 0, 2, 0, 0, 0, 8, 
    
    -- channel=262
    0, 0, 55, 65, 69, 57, 68, 65, 90, 64, 5, 90, 83, 80, 78, 
    0, 0, 31, 43, 95, 83, 69, 80, 88, 73, 46, 108, 100, 91, 88, 
    0, 0, 5, 56, 88, 116, 46, 36, 50, 49, 97, 93, 111, 115, 115, 
    73, 14, 90, 84, 70, 114, 103, 75, 47, 44, 101, 99, 134, 128, 92, 
    107, 99, 103, 83, 63, 96, 105, 81, 49, 47, 81, 115, 129, 114, 78, 
    101, 92, 102, 83, 86, 97, 93, 56, 77, 64, 79, 102, 133, 130, 88, 
    100, 89, 82, 79, 86, 68, 100, 62, 98, 80, 77, 104, 126, 140, 118, 
    101, 87, 96, 62, 115, 101, 88, 95, 63, 68, 88, 46, 90, 130, 103, 
    114, 72, 96, 83, 112, 131, 118, 107, 37, 66, 88, 68, 21, 60, 67, 
    117, 97, 107, 103, 94, 97, 104, 112, 110, 72, 78, 56, 63, 80, 53, 
    113, 109, 90, 111, 112, 110, 75, 87, 105, 91, 42, 71, 80, 68, 60, 
    106, 112, 84, 117, 120, 90, 97, 95, 100, 72, 53, 69, 78, 77, 61, 
    105, 95, 79, 112, 119, 23, 80, 81, 77, 59, 51, 58, 58, 49, 63, 
    101, 87, 63, 110, 118, 94, 83, 62, 55, 32, 50, 52, 51, 38, 63, 
    75, 80, 56, 93, 109, 101, 64, 48, 48, 28, 44, 53, 52, 53, 50, 
    
    -- channel=263
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=264
    0, 56, 28, 15, 20, 19, 14, 19, 0, 0, 54, 25, 23, 21, 18, 
    0, 34, 35, 31, 27, 19, 24, 25, 21, 0, 66, 26, 24, 25, 24, 
    0, 9, 45, 34, 53, 3, 22, 36, 21, 24, 41, 34, 29, 29, 24, 
    0, 22, 34, 5, 57, 19, 10, 5, 20, 56, 30, 50, 37, 21, 35, 
    0, 25, 19, 0, 57, 41, 21, 1, 25, 47, 39, 46, 35, 1, 30, 
    16, 26, 14, 8, 40, 35, 18, 16, 23, 44, 42, 52, 30, 0, 6, 
    13, 21, 8, 29, 29, 43, 15, 34, 17, 32, 43, 50, 34, 15, 3, 
    8, 24, 3, 57, 21, 31, 22, 29, 30, 31, 25, 42, 45, 23, 27, 
    0, 24, 24, 55, 31, 30, 30, 2, 43, 22, 17, 8, 53, 24, 43, 
    1, 18, 34, 30, 40, 43, 39, 22, 14, 33, 10, 21, 27, 15, 36, 
    17, 9, 39, 34, 33, 12, 46, 45, 18, 9, 23, 26, 28, 15, 18, 
    21, 0, 47, 39, 32, 21, 36, 34, 25, 0, 32, 22, 29, 16, 10, 
    15, 0, 34, 38, 13, 51, 41, 29, 17, 8, 28, 20, 24, 21, 16, 
    10, 0, 28, 38, 12, 37, 21, 22, 14, 13, 22, 20, 9, 29, 22, 
    9, 0, 19, 45, 26, 19, 8, 18, 2, 23, 18, 19, 11, 21, 22, 
    
    -- channel=265
    0, 0, 50, 55, 35, 52, 54, 49, 44, 11, 0, 45, 59, 60, 62, 
    0, 0, 45, 43, 19, 23, 44, 44, 47, 41, 0, 41, 49, 53, 60, 
    0, 0, 18, 23, 18, 25, 20, 32, 47, 22, 11, 34, 42, 41, 42, 
    0, 0, 2, 42, 25, 28, 7, 19, 12, 1, 35, 23, 37, 46, 38, 
    41, 15, 33, 42, 7, 23, 33, 32, 10, 4, 30, 31, 37, 46, 30, 
    40, 32, 45, 28, 26, 28, 32, 14, 4, 0, 18, 34, 42, 46, 36, 
    43, 37, 54, 39, 16, 2, 23, 14, 25, 11, 7, 32, 43, 47, 37, 
    43, 38, 47, 46, 33, 22, 26, 2, 34, 20, 31, 58, 55, 53, 32, 
    44, 26, 39, 28, 28, 24, 9, 31, 18, 26, 40, 19, 29, 54, 42, 
    45, 25, 30, 35, 25, 31, 31, 24, 2, 21, 50, 40, 20, 41, 33, 
    41, 31, 28, 28, 32, 36, 23, 26, 42, 47, 29, 30, 31, 37, 33, 
    38, 42, 20, 34, 40, 51, 30, 33, 36, 44, 20, 35, 35, 33, 31, 
    38, 46, 27, 28, 43, 20, 42, 42, 48, 36, 28, 31, 37, 36, 29, 
    42, 45, 26, 29, 41, 11, 51, 41, 40, 29, 28, 24, 28, 20, 29, 
    42, 41, 23, 26, 31, 37, 47, 42, 38, 10, 27, 26, 25, 22, 33, 
    
    -- channel=266
    12, 0, 15, 19, 16, 20, 25, 22, 34, 30, 3, 8, 24, 23, 26, 
    12, 1, 0, 8, 0, 1, 0, 0, 0, 33, 0, 2, 12, 16, 18, 
    13, 7, 0, 16, 0, 3, 0, 0, 0, 14, 0, 0, 0, 0, 3, 
    59, 46, 0, 0, 0, 0, 23, 11, 4, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 15, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 18, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 17, 0, 0, 0, 0, 1, 0, 8, 0, 29, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 25, 4, 0, 10, 19, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 1, 0, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 1, 0, 0, 6, 12, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 10, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 27, 0, 0, 4, 10, 0, 6, 9, 1, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 15, 2, 5, 15, 2, 0, 
    
    -- channel=267
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=268
    7, 86, 38, 12, 11, 20, 15, 25, 0, 0, 69, 33, 21, 23, 15, 
    10, 56, 57, 23, 15, 7, 17, 28, 12, 0, 119, 17, 12, 16, 13, 
    9, 27, 83, 39, 40, 0, 0, 20, 0, 9, 74, 22, 15, 18, 13, 
    10, 68, 110, 0, 47, 0, 0, 0, 18, 64, 20, 52, 14, 0, 22, 
    0, 68, 23, 0, 67, 6, 0, 0, 18, 41, 32, 61, 11, 0, 43, 
    15, 26, 10, 0, 46, 5, 0, 0, 26, 42, 32, 63, 14, 0, 30, 
    17, 19, 0, 33, 12, 14, 0, 19, 6, 28, 30, 63, 23, 6, 10, 
    8, 17, 0, 75, 1, 12, 0, 14, 14, 22, 10, 29, 35, 7, 21, 
    0, 20, 0, 55, 5, 20, 6, 0, 43, 0, 17, 2, 59, 0, 55, 
    3, 26, 20, 10, 22, 6, 0, 0, 5, 35, 0, 13, 29, 17, 37, 
    16, 1, 32, 15, 20, 0, 34, 14, 0, 0, 3, 29, 21, 0, 11, 
    20, 0, 54, 9, 2, 0, 35, 14, 1, 0, 49, 10, 20, 0, 0, 
    15, 2, 48, 11, 0, 0, 32, 4, 0, 0, 34, 5, 7, 0, 9, 
    7, 5, 50, 24, 0, 23, 0, 2, 0, 0, 27, 11, 0, 32, 18, 
    0, 13, 40, 35, 0, 0, 0, 7, 0, 31, 14, 17, 3, 30, 13, 
    
    -- channel=269
    9, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 9, 9, 0, 0, 0, 18, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 3, 31, 19, 9, 19, 5, 0, 17, 14, 7, 4, 
    0, 0, 0, 6, 3, 24, 2, 10, 5, 0, 14, 0, 10, 19, 14, 
    5, 0, 7, 23, 0, 22, 20, 24, 5, 0, 11, 0, 18, 30, 5, 
    9, 7, 13, 8, 0, 19, 30, 23, 2, 0, 12, 5, 25, 28, 10, 
    11, 8, 18, 0, 19, 23, 27, 3, 16, 8, 11, 0, 20, 24, 21, 
    17, 5, 8, 0, 16, 14, 29, 0, 6, 9, 10, 15, 8, 26, 14, 
    23, 13, 3, 0, 16, 9, 17, 33, 0, 5, 0, 0, 10, 30, 2, 
    23, 6, 7, 6, 21, 27, 21, 25, 0, 0, 16, 0, 0, 0, 1, 
    20, 20, 12, 12, 8, 26, 8, 15, 24, 10, 4, 0, 0, 12, 0, 
    19, 24, 4, 18, 15, 19, 0, 5, 11, 23, 0, 4, 0, 2, 5, 
    20, 23, 4, 21, 29, 13, 0, 8, 16, 8, 0, 5, 9, 8, 0, 
    21, 20, 5, 19, 28, 0, 5, 5, 9, 8, 0, 0, 7, 0, 0, 
    25, 14, 7, 16, 23, 16, 14, 0, 9, 0, 0, 0, 1, 0, 2, 
    
    -- channel=270
    11, 0, 13, 39, 41, 23, 40, 25, 45, 92, 0, 22, 39, 37, 45, 
    9, 0, 0, 1, 10, 41, 9, 9, 39, 85, 0, 26, 41, 41, 45, 
    10, 0, 0, 13, 0, 80, 37, 24, 41, 0, 0, 9, 26, 21, 26, 
    70, 0, 0, 54, 0, 34, 39, 50, 15, 0, 18, 0, 14, 45, 0, 
    38, 0, 27, 71, 0, 12, 42, 64, 7, 0, 0, 0, 27, 76, 6, 
    27, 14, 35, 43, 0, 14, 58, 33, 14, 0, 0, 0, 27, 74, 33, 
    36, 22, 70, 13, 38, 7, 60, 0, 32, 0, 0, 0, 17, 36, 39, 
    48, 14, 90, 0, 34, 16, 19, 39, 0, 6, 31, 0, 0, 49, 3, 
    69, 15, 27, 0, 3, 7, 30, 74, 0, 28, 31, 56, 2, 41, 0, 
    46, 11, 11, 18, 16, 24, 2, 23, 58, 6, 58, 24, 9, 40, 20, 
    25, 51, 0, 22, 14, 64, 0, 13, 37, 70, 12, 12, 19, 47, 33, 
    25, 59, 0, 13, 36, 30, 6, 18, 41, 72, 0, 26, 13, 42, 40, 
    34, 51, 0, 18, 84, 17, 14, 30, 54, 49, 6, 25, 35, 20, 34, 
    41, 57, 0, 5, 51, 9, 48, 39, 53, 26, 16, 26, 45, 0, 18, 
    38, 43, 0, 0, 31, 56, 55, 26, 61, 4, 20, 23, 29, 16, 19, 
    
    -- channel=271
    2, 0, 18, 8, 0, 6, 5, 4, 44, 0, 0, 13, 8, 3, 4, 
    0, 0, 15, 0, 33, 0, 17, 16, 15, 49, 0, 18, 9, 5, 9, 
    0, 0, 2, 0, 22, 35, 0, 0, 13, 32, 0, 9, 23, 24, 23, 
    0, 0, 0, 0, 16, 58, 21, 15, 6, 0, 34, 14, 28, 26, 17, 
    56, 3, 17, 23, 0, 19, 34, 28, 8, 0, 20, 14, 24, 22, 0, 
    24, 4, 25, 12, 13, 15, 26, 11, 19, 0, 0, 15, 27, 40, 2, 
    13, 6, 0, 38, 0, 0, 25, 18, 30, 15, 0, 11, 21, 52, 18, 
    9, 6, 24, 26, 25, 17, 42, 0, 41, 0, 8, 0, 32, 27, 20, 
    30, 0, 48, 0, 46, 46, 11, 53, 0, 0, 41, 0, 0, 13, 0, 
    41, 4, 17, 26, 0, 5, 42, 44, 0, 9, 14, 17, 0, 13, 0, 
    29, 10, 24, 11, 26, 21, 0, 1, 51, 10, 10, 5, 9, 12, 1, 
    14, 40, 0, 26, 23, 36, 12, 13, 16, 26, 0, 5, 24, 10, 14, 
    16, 25, 0, 21, 31, 0, 17, 6, 17, 11, 0, 3, 0, 16, 9, 
    16, 18, 0, 29, 50, 0, 5, 3, 4, 0, 1, 0, 6, 0, 14, 
    9, 29, 0, 25, 26, 13, 11, 11, 10, 0, 0, 6, 11, 0, 3, 
    
    -- channel=272
    5, 0, 59, 73, 56, 66, 71, 63, 60, 56, 1, 56, 77, 75, 79, 
    5, 0, 49, 60, 29, 48, 52, 50, 64, 60, 0, 51, 67, 71, 77, 
    8, 3, 14, 59, 30, 50, 46, 53, 64, 28, 22, 39, 50, 51, 53, 
    12, 0, 9, 65, 31, 39, 32, 43, 33, 19, 36, 28, 45, 53, 35, 
    40, 21, 36, 59, 26, 38, 50, 54, 30, 22, 26, 33, 44, 52, 35, 
    44, 38, 46, 48, 36, 42, 51, 36, 26, 18, 25, 31, 39, 46, 36, 
    46, 43, 67, 48, 41, 26, 48, 25, 36, 24, 21, 28, 40, 39, 32, 
    47, 48, 79, 42, 48, 37, 37, 41, 30, 35, 42, 53, 38, 54, 28, 
    48, 40, 60, 46, 34, 31, 34, 49, 33, 46, 49, 45, 45, 55, 29, 
    40, 35, 46, 46, 40, 49, 39, 31, 40, 42, 61, 54, 40, 54, 47, 
    37, 45, 31, 41, 41, 53, 37, 44, 49, 67, 41, 47, 50, 56, 53, 
    37, 46, 28, 45, 54, 58, 40, 48, 53, 60, 37, 51, 47, 53, 47, 
    37, 43, 30, 41, 70, 54, 53, 57, 63, 56, 42, 49, 55, 47, 48, 
    40, 42, 28, 36, 53, 49, 63, 59, 61, 44, 44, 45, 49, 36, 45, 
    41, 36, 34, 28, 43, 58, 64, 57, 59, 33, 42, 44, 42, 43, 46, 
    
    -- channel=273
    9, 49, 15, 8, 11, 10, 2, 4, 0, 0, 37, 7, 3, 2, 1, 
    10, 35, 34, 27, 17, 15, 26, 18, 19, 0, 27, 14, 10, 10, 9, 
    10, 20, 35, 19, 47, 14, 38, 48, 43, 22, 24, 31, 21, 16, 11, 
    0, 0, 0, 12, 63, 20, 0, 6, 20, 46, 38, 35, 34, 36, 40, 
    0, 2, 14, 2, 48, 47, 29, 20, 29, 46, 41, 33, 32, 10, 29, 
    16, 26, 19, 3, 36, 46, 34, 22, 15, 34, 44, 43, 30, 0, 5, 
    12, 20, 22, 19, 29, 38, 21, 37, 22, 36, 39, 42, 33, 10, 0, 
    12, 26, 5, 44, 23, 38, 32, 27, 41, 33, 36, 73, 55, 34, 25, 
    0, 23, 14, 43, 30, 19, 21, 13, 44, 24, 18, 2, 63, 49, 46, 
    0, 10, 30, 33, 44, 59, 49, 19, 0, 20, 26, 18, 10, 13, 42, 
    18, 13, 38, 27, 26, 23, 48, 51, 27, 23, 24, 17, 25, 22, 21, 
    24, 6, 41, 40, 38, 34, 26, 33, 29, 12, 21, 27, 28, 16, 12, 
    20, 9, 34, 42, 30, 56, 38, 37, 31, 19, 27, 26, 38, 31, 16, 
    17, 4, 26, 39, 14, 13, 31, 30, 24, 23, 22, 21, 17, 27, 18, 
    25, 4, 22, 51, 30, 24, 27, 28, 16, 18, 22, 18, 10, 17, 29, 
    
    -- channel=274
    0, 129, 44, 0, 0, 9, 0, 0, 0, 0, 101, 0, 0, 0, 0, 
    1, 70, 113, 9, 0, 0, 19, 1, 0, 0, 89, 0, 0, 0, 0, 
    0, 24, 150, 0, 35, 0, 0, 57, 25, 9, 19, 12, 0, 0, 0, 
    0, 0, 24, 0, 77, 0, 0, 0, 0, 59, 8, 34, 0, 0, 21, 
    0, 0, 0, 0, 61, 0, 0, 0, 11, 40, 37, 26, 0, 0, 19, 
    0, 0, 0, 0, 22, 0, 0, 0, 0, 14, 21, 62, 0, 0, 0, 
    0, 0, 0, 14, 0, 0, 0, 13, 0, 6, 10, 50, 0, 0, 0, 
    0, 0, 0, 92, 0, 0, 0, 0, 35, 0, 0, 95, 72, 0, 0, 
    0, 0, 0, 10, 0, 0, 0, 0, 44, 0, 0, 0, 94, 43, 79, 
    0, 0, 0, 0, 1, 13, 4, 0, 0, 7, 0, 6, 0, 0, 31, 
    0, 0, 31, 0, 0, 0, 37, 3, 0, 0, 8, 0, 0, 0, 0, 
    0, 0, 43, 0, 0, 0, 0, 0, 0, 0, 24, 0, 10, 0, 0, 
    0, 0, 31, 0, 0, 6, 31, 0, 0, 0, 27, 0, 10, 10, 0, 
    0, 0, 34, 10, 0, 0, 0, 0, 0, 0, 13, 0, 0, 25, 0, 
    0, 0, 10, 49, 0, 0, 0, 11, 0, 17, 2, 0, 0, 0, 10, 
    
    -- channel=275
    0, 37, 6, 0, 0, 1, 0, 0, 0, 0, 16, 0, 0, 0, 0, 
    0, 24, 41, 2, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 8, 38, 0, 0, 0, 19, 51, 42, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 21, 0, 0, 0, 0, 4, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 4, 0, 0, 0, 1, 6, 2, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 0, 0, 0, 0, 11, 0, 0, 68, 28, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 65, 57, 28, 
    0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 1, 0, 0, 24, 
    0, 0, 0, 0, 0, 0, 14, 6, 0, 0, 9, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 31, 11, 3, 7, 0, 6, 1, 18, 14, 0, 
    0, 0, 6, 0, 0, 0, 0, 11, 11, 8, 1, 0, 0, 5, 0, 
    11, 0, 4, 10, 0, 0, 11, 13, 4, 3, 2, 0, 0, 0, 8, 
    
    -- channel=276
    0, 21, 9, 8, 10, 7, 1, 10, 0, 0, 26, 18, 7, 7, 2, 
    0, 8, 18, 17, 30, 23, 24, 22, 24, 0, 53, 29, 21, 19, 14, 
    0, 0, 21, 22, 57, 12, 14, 33, 16, 12, 56, 52, 45, 43, 33, 
    0, 0, 51, 18, 56, 29, 8, 2, 15, 47, 45, 66, 54, 47, 52, 
    19, 39, 39, 0, 57, 48, 33, 4, 22, 37, 49, 68, 57, 27, 52, 
    38, 43, 38, 14, 50, 46, 19, 10, 26, 39, 46, 78, 62, 32, 39, 
    38, 37, 20, 31, 29, 42, 29, 33, 27, 38, 48, 69, 68, 52, 35, 
    39, 38, 0, 52, 42, 39, 34, 30, 29, 40, 34, 63, 59, 59, 53, 
    29, 35, 17, 46, 46, 46, 41, 11, 35, 14, 29, 0, 55, 41, 64, 
    38, 41, 43, 37, 54, 61, 51, 26, 12, 35, 10, 12, 14, 20, 32, 
    50, 39, 52, 45, 49, 24, 52, 51, 30, 15, 8, 23, 25, 9, 18, 
    52, 31, 63, 55, 47, 24, 40, 37, 33, 0, 27, 21, 29, 14, 0, 
    46, 33, 55, 52, 27, 10, 44, 30, 19, 4, 23, 16, 23, 11, 10, 
    40, 26, 53, 59, 25, 19, 17, 17, 10, 0, 17, 12, 2, 16, 19, 
    31, 24, 47, 60, 40, 31, 8, 9, 0, 10, 9, 14, 0, 18, 13, 
    
    -- channel=277
    3, 0, 0, 18, 8, 0, 9, 0, 46, 88, 0, 0, 5, 3, 12, 
    1, 0, 0, 0, 0, 18, 0, 0, 14, 104, 0, 1, 13, 7, 12, 
    2, 0, 0, 0, 0, 88, 5, 0, 12, 0, 0, 0, 6, 2, 11, 
    79, 0, 0, 42, 0, 42, 45, 41, 0, 0, 0, 0, 2, 29, 0, 
    45, 0, 2, 76, 0, 0, 34, 66, 0, 0, 0, 0, 6, 65, 0, 
    11, 0, 12, 42, 0, 0, 47, 30, 0, 0, 0, 0, 5, 69, 5, 
    13, 0, 41, 0, 14, 0, 51, 0, 21, 0, 0, 0, 0, 29, 32, 
    27, 0, 85, 0, 28, 2, 19, 19, 0, 0, 6, 0, 0, 24, 0, 
    60, 0, 20, 0, 2, 4, 26, 74, 0, 16, 7, 39, 0, 1, 0, 
    38, 0, 0, 5, 0, 0, 0, 28, 51, 0, 31, 0, 0, 12, 0, 
    9, 41, 0, 2, 0, 53, 0, 0, 32, 45, 0, 0, 0, 29, 7, 
    1, 55, 0, 0, 17, 24, 0, 0, 20, 68, 0, 2, 0, 27, 26, 
    11, 33, 0, 0, 68, 0, 0, 3, 32, 36, 0, 4, 0, 0, 12, 
    20, 36, 0, 0, 52, 0, 17, 10, 29, 7, 0, 2, 27, 0, 0, 
    15, 20, 0, 0, 20, 35, 37, 0, 43, 0, 0, 0, 14, 0, 0, 
    
    -- channel=278
    14, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 0, 0, 
    14, 5, 0, 0, 1, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 
    13, 10, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    105, 78, 47, 0, 0, 0, 35, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 13, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 37, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=279
    3, 0, 0, 10, 16, 0, 18, 18, 54, 61, 0, 31, 28, 23, 22, 
    3, 0, 0, 0, 30, 29, 0, 0, 3, 33, 21, 24, 25, 18, 15, 
    4, 0, 0, 16, 0, 39, 0, 0, 0, 0, 23, 0, 8, 21, 32, 
    148, 86, 71, 9, 0, 24, 79, 41, 6, 0, 0, 0, 19, 0, 0, 
    45, 53, 11, 20, 0, 0, 6, 11, 0, 0, 0, 0, 1, 6, 0, 
    1, 0, 0, 24, 0, 0, 0, 4, 29, 9, 0, 0, 0, 23, 0, 
    0, 0, 0, 0, 8, 0, 19, 0, 21, 0, 0, 0, 0, 16, 35, 
    0, 0, 29, 0, 20, 0, 0, 31, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 28, 10, 3, 43, 48, 29, 0, 0, 0, 33, 0, 0, 0, 
    10, 21, 7, 2, 0, 0, 0, 33, 81, 7, 0, 0, 27, 11, 0, 
    0, 9, 0, 14, 11, 11, 0, 0, 0, 1, 0, 15, 5, 0, 0, 
    0, 3, 0, 0, 0, 0, 10, 1, 0, 5, 1, 0, 0, 12, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 22, 65, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 1, 4, 0, 0, 0, 0, 0, 0, 11, 6, 0, 
    
    -- channel=280
    5, 0, 48, 66, 61, 48, 61, 55, 88, 76, 0, 75, 77, 73, 75, 
    3, 0, 14, 43, 92, 75, 67, 72, 91, 114, 0, 95, 90, 85, 85, 
    5, 0, 0, 42, 82, 138, 49, 38, 63, 52, 59, 80, 103, 102, 103, 
    65, 0, 39, 88, 56, 133, 106, 79, 45, 21, 100, 79, 130, 133, 85, 
    116, 69, 94, 101, 37, 98, 120, 104, 51, 32, 72, 85, 124, 125, 59, 
    99, 82, 100, 93, 72, 101, 109, 71, 72, 49, 67, 74, 124, 135, 73, 
    92, 81, 94, 80, 77, 65, 113, 62, 101, 70, 68, 76, 119, 138, 106, 
    99, 80, 121, 42, 119, 99, 103, 95, 72, 66, 93, 46, 82, 129, 98, 
    117, 60, 102, 60, 116, 122, 115, 127, 20, 76, 95, 71, 0, 75, 51, 
    116, 83, 95, 103, 84, 101, 115, 120, 104, 68, 87, 61, 58, 81, 39, 
    106, 108, 78, 103, 109, 119, 66, 91, 123, 100, 51, 61, 75, 79, 66, 
    97, 120, 60, 116, 123, 111, 88, 95, 107, 97, 39, 71, 78, 87, 70, 
    99, 98, 57, 109, 135, 35, 81, 86, 94, 77, 44, 64, 63, 60, 66, 
    100, 89, 39, 100, 131, 89, 87, 70, 72, 43, 45, 56, 64, 31, 65, 
    78, 79, 37, 82, 114, 107, 85, 56, 66, 26, 44, 56, 59, 49, 51, 
    
    -- channel=281
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 19, 34, 39, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 61, 9, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 52, 6, 
    0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 13, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 13, 13, 0, 3, 13, 2, 0, 0, 18, 6, 0, 
    0, 3, 0, 0, 0, 0, 5, 8, 12, 3, 0, 0, 0, 0, 0, 
    17, 0, 0, 0, 0, 0, 20, 7, 11, 0, 0, 0, 0, 0, 1, 
    
    -- channel=282
    0, 0, 12, 35, 28, 23, 38, 32, 48, 66, 0, 32, 43, 44, 46, 
    0, 0, 0, 14, 22, 40, 17, 26, 39, 63, 0, 39, 45, 42, 42, 
    0, 0, 0, 26, 1, 60, 16, 2, 13, 6, 19, 24, 37, 38, 44, 
    73, 1, 15, 53, 0, 39, 51, 41, 12, 0, 25, 9, 42, 54, 21, 
    60, 32, 42, 61, 0, 18, 39, 45, 7, 0, 11, 20, 47, 74, 29, 
    45, 36, 44, 50, 12, 23, 37, 26, 19, 2, 13, 9, 48, 79, 52, 
    50, 38, 53, 18, 32, 11, 44, 1, 37, 11, 16, 13, 44, 59, 66, 
    57, 28, 58, 0, 46, 26, 25, 37, 4, 26, 31, 2, 4, 55, 38, 
    69, 23, 26, 20, 27, 36, 44, 51, 1, 31, 30, 46, 0, 22, 5, 
    61, 41, 25, 36, 25, 23, 17, 38, 59, 19, 39, 19, 25, 38, 15, 
    47, 58, 9, 37, 37, 55, 6, 21, 36, 51, 12, 22, 24, 35, 28, 
    44, 62, 6, 28, 41, 34, 25, 32, 39, 50, 10, 26, 18, 39, 33, 
    50, 57, 15, 29, 52, 3, 16, 30, 37, 36, 10, 23, 21, 14, 29, 
    53, 59, 15, 21, 46, 33, 40, 27, 33, 20, 16, 22, 31, 5, 22, 
    41, 48, 26, 3, 37, 46, 37, 17, 36, 8, 17, 21, 27, 21, 15, 
    
    -- channel=283
    2, 26, 0, 2, 9, 4, 5, 0, 0, 38, 3, 0, 0, 2, 5, 
    4, 36, 0, 10, 0, 25, 1, 0, 0, 36, 0, 0, 3, 4, 5, 
    5, 16, 0, 12, 0, 26, 20, 0, 2, 9, 0, 0, 0, 0, 3, 
    2, 0, 0, 26, 0, 2, 22, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 40, 0, 0, 3, 23, 0, 10, 0, 0, 0, 21, 0, 
    0, 1, 0, 38, 0, 6, 8, 28, 0, 4, 0, 0, 0, 10, 0, 
    0, 9, 25, 0, 0, 7, 0, 21, 0, 0, 5, 0, 0, 0, 24, 
    10, 13, 33, 0, 6, 0, 4, 18, 0, 25, 0, 11, 0, 0, 15, 
    2, 12, 0, 0, 0, 0, 13, 0, 15, 41, 0, 31, 0, 0, 0, 
    0, 19, 0, 0, 0, 0, 0, 10, 30, 0, 1, 0, 13, 0, 1, 
    0, 19, 0, 0, 0, 10, 0, 7, 2, 0, 17, 0, 0, 14, 4, 
    0, 0, 0, 0, 0, 30, 0, 2, 1, 31, 0, 6, 0, 15, 11, 
    2, 0, 0, 0, 0, 72, 0, 10, 8, 26, 0, 14, 0, 6, 0, 
    7, 4, 3, 0, 9, 34, 0, 7, 13, 33, 0, 9, 13, 0, 0, 
    19, 0, 25, 0, 11, 2, 32, 0, 11, 9, 4, 0, 11, 0, 0, 
    
    -- channel=284
    0, 0, 67, 67, 67, 60, 69, 62, 81, 53, 0, 82, 80, 79, 80, 
    0, 0, 47, 42, 87, 74, 79, 83, 93, 96, 6, 102, 94, 89, 90, 
    0, 0, 3, 33, 81, 121, 52, 53, 77, 53, 69, 96, 109, 107, 106, 
    30, 0, 47, 88, 69, 120, 84, 68, 42, 26, 113, 87, 129, 142, 105, 
    115, 73, 106, 96, 42, 98, 114, 95, 49, 36, 90, 101, 132, 136, 83, 
    110, 96, 118, 88, 75, 102, 107, 61, 63, 44, 80, 97, 141, 147, 96, 
    109, 96, 105, 85, 73, 59, 102, 58, 97, 71, 73, 100, 135, 151, 119, 
    116, 94, 108, 56, 113, 99, 97, 82, 85, 69, 104, 85, 119, 148, 117, 
    129, 70, 91, 61, 114, 114, 97, 116, 33, 74, 100, 66, 28, 105, 87, 
    131, 89, 99, 104, 91, 109, 117, 111, 84, 65, 96, 67, 53, 85, 59, 
    124, 114, 91, 104, 109, 117, 75, 93, 124, 104, 57, 63, 77, 79, 68, 
    117, 130, 74, 117, 126, 110, 90, 95, 108, 95, 44, 75, 83, 84, 69, 
    119, 119, 77, 112, 132, 30, 89, 94, 99, 77, 54, 66, 72, 68, 66, 
    120, 113, 63, 110, 124, 68, 96, 77, 75, 48, 52, 57, 63, 38, 67, 
    103, 105, 54, 99, 115, 109, 91, 65, 68, 29, 50, 59, 58, 51, 60, 
    
    -- channel=285
    7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    7, 3, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 4, 2, 0, 24, 7, 2, 7, 7, 4, 8, 16, 4, 0, 0, 
    0, 0, 0, 0, 31, 18, 0, 0, 1, 11, 24, 19, 15, 17, 22, 
    0, 0, 9, 0, 18, 26, 14, 2, 9, 14, 24, 17, 19, 8, 11, 
    6, 10, 11, 0, 13, 23, 16, 7, 8, 13, 20, 27, 24, 6, 2, 
    4, 5, 0, 3, 7, 20, 12, 12, 15, 18, 22, 25, 25, 18, 1, 
    6, 6, 0, 6, 12, 20, 23, 8, 23, 12, 19, 27, 34, 23, 22, 
    4, 3, 0, 0, 24, 15, 11, 10, 3, 0, 5, 0, 12, 28, 25, 
    10, 2, 10, 9, 22, 32, 33, 16, 0, 0, 0, 0, 0, 0, 2, 
    17, 9, 23, 11, 13, 10, 22, 22, 17, 0, 0, 0, 0, 0, 0, 
    18, 11, 21, 21, 17, 8, 6, 8, 9, 0, 0, 0, 4, 0, 0, 
    15, 11, 17, 24, 11, 0, 8, 6, 3, 0, 0, 0, 5, 3, 0, 
    13, 6, 13, 27, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 6, 6, 36, 17, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=286
    0, 5, 47, 22, 17, 32, 23, 23, 0, 0, 21, 26, 27, 31, 32, 
    0, 0, 76, 30, 5, 4, 35, 33, 37, 0, 10, 36, 37, 39, 37, 
    0, 0, 58, 14, 42, 0, 29, 65, 61, 10, 32, 65, 47, 38, 31, 
    0, 0, 0, 21, 68, 11, 0, 0, 6, 25, 55, 55, 37, 54, 72, 
    0, 0, 40, 7, 49, 46, 26, 1, 12, 23, 55, 68, 62, 48, 70, 
    46, 47, 57, 7, 36, 39, 34, 2, 0, 8, 43, 90, 70, 41, 52, 
    53, 49, 51, 46, 33, 35, 16, 4, 10, 25, 35, 81, 76, 52, 21, 
    52, 53, 8, 64, 20, 30, 24, 0, 49, 25, 45, 107, 106, 84, 61, 
    44, 48, 19, 30, 36, 13, 0, 9, 35, 17, 39, 0, 99, 106, 93, 
    46, 21, 43, 37, 61, 76, 54, 7, 0, 25, 38, 33, 0, 22, 61, 
    59, 36, 61, 36, 35, 31, 65, 54, 39, 32, 28, 19, 27, 24, 23, 
    64, 45, 62, 50, 50, 33, 32, 36, 39, 14, 21, 29, 38, 13, 9, 
    59, 58, 63, 56, 53, 33, 63, 52, 47, 17, 35, 26, 45, 37, 16, 
    56, 51, 63, 61, 26, 0, 42, 46, 34, 16, 27, 19, 13, 23, 22, 
    62, 51, 47, 74, 40, 39, 33, 35, 16, 9, 20, 19, 2, 11, 33, 
    
    -- channel=287
    1, 0, 0, 0, 0, 0, 0, 0, 10, 20, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    64, 44, 0, 0, 0, 0, 4, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 
    0, 0, 0, 1, 0, 0, 0, 4, 0, 0, 0, 0, 0, 14, 12, 
    0, 0, 0, 0, 17, 11, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 7, 0, 0, 0, 0, 1, 0, 0, 0, 0, 20, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=288
    103, 103, 97, 71, 80, 76, 84, 100, 109, 110, 109, 113, 99, 102, 94, 
    111, 111, 101, 43, 41, 44, 47, 55, 76, 93, 106, 114, 111, 99, 121, 
    113, 114, 91, 20, 23, 18, 15, 7, 6, 29, 93, 107, 98, 89, 114, 
    112, 107, 93, 13, 52, 53, 34, 30, 29, 32, 43, 112, 98, 86, 85, 
    114, 105, 57, 15, 30, 35, 27, 23, 32, 39, 35, 76, 108, 88, 90, 
    115, 95, 69, 0, 16, 17, 11, 15, 14, 31, 37, 57, 115, 113, 113, 
    94, 65, 60, 36, 11, 12, 5, 0, 15, 14, 13, 42, 73, 99, 120, 
    75, 32, 73, 29, 16, 1, 1, 3, 4, 2, 6, 13, 28, 40, 108, 
    68, 21, 61, 3, 32, 33, 31, 0, 24, 35, 9, 14, 41, 30, 86, 
    76, 11, 30, 9, 9, 3, 8, 47, 24, 34, 26, 28, 35, 12, 83, 
    80, 8, 16, 4, 0, 8, 18, 0, 34, 13, 16, 36, 0, 40, 59, 
    63, 0, 23, 25, 0, 0, 25, 0, 38, 38, 32, 44, 6, 10, 76, 
    55, 17, 15, 26, 0, 0, 0, 0, 7, 80, 55, 16, 0, 10, 58, 
    55, 42, 24, 15, 12, 0, 0, 1, 14, 32, 53, 8, 0, 17, 54, 
    42, 36, 20, 0, 10, 0, 0, 0, 4, 13, 25, 6, 0, 13, 69, 
    
    -- channel=289
    14, 14, 3, 8, 8, 14, 29, 34, 19, 13, 12, 10, 22, 27, 27, 
    4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 8, 3, 6, 17, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 5, 3, 11, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 22, 21, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 10, 27, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 15, 0, 0, 0, 2, 2, 15, 33, 40, 36, 40, 19, 0, 0, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 2, 2, 11, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 14, 0, 3, 13, 13, 11, 10, 25, 21, 1, 8, 7, 2, 
    0, 0, 0, 0, 0, 8, 19, 16, 16, 0, 0, 0, 13, 5, 0, 
    0, 0, 0, 0, 0, 6, 13, 9, 4, 0, 0, 0, 15, 4, 0, 
    
    -- channel=290
    33, 36, 28, 17, 25, 30, 34, 35, 46, 41, 36, 42, 19, 31, 9, 
    46, 46, 34, 4, 17, 23, 26, 34, 43, 42, 34, 44, 44, 22, 40, 
    48, 47, 36, 0, 0, 0, 0, 0, 0, 0, 50, 48, 33, 12, 49, 
    47, 41, 31, 0, 28, 40, 3, 0, 0, 5, 9, 53, 31, 17, 29, 
    50, 37, 29, 0, 18, 6, 0, 0, 3, 5, 0, 56, 56, 24, 26, 
    60, 35, 0, 0, 4, 0, 0, 0, 0, 0, 6, 18, 55, 47, 48, 
    50, 25, 24, 0, 3, 0, 0, 0, 0, 6, 0, 22, 51, 62, 48, 
    46, 1, 33, 9, 0, 0, 0, 0, 0, 0, 0, 0, 8, 16, 71, 
    31, 0, 31, 0, 0, 13, 0, 0, 0, 0, 0, 0, 8, 12, 82, 
    25, 0, 22, 0, 4, 0, 0, 17, 0, 5, 0, 0, 15, 0, 58, 
    35, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 55, 
    29, 0, 11, 0, 0, 0, 0, 0, 31, 0, 4, 23, 0, 1, 40, 
    21, 0, 2, 0, 0, 0, 0, 0, 0, 40, 24, 0, 0, 0, 49, 
    22, 13, 0, 0, 0, 0, 0, 0, 0, 31, 15, 0, 0, 0, 39, 
    12, 3, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 36, 
    
    -- channel=291
    11, 7, 13, 21, 6, 0, 0, 0, 0, 12, 16, 11, 11, 13, 15, 
    5, 5, 15, 22, 3, 0, 3, 11, 10, 12, 23, 9, 16, 33, 15, 
    8, 7, 15, 19, 0, 0, 0, 0, 0, 0, 0, 8, 21, 35, 20, 
    8, 13, 7, 22, 0, 0, 0, 0, 0, 0, 0, 9, 12, 22, 17, 
    6, 13, 20, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 
    2, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 
    1, 23, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 0, 
    8, 26, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 6, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 24, 3, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 
    4, 18, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 6, 0, 0, 
    0, 29, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 3, 4, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 24, 2, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    
    -- channel=292
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=293
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 46, 53, 50, 66, 90, 80, 48, 21, 0, 0, 6, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 6, 0, 0, 2, 19, 13, 
    0, 0, 0, 20, 0, 0, 10, 5, 0, 0, 10, 12, 0, 0, 17, 
    0, 0, 58, 30, 0, 25, 25, 6, 7, 8, 0, 0, 0, 0, 0, 
    4, 17, 0, 12, 34, 0, 5, 27, 32, 15, 35, 25, 0, 0, 0, 
    7, 38, 32, 0, 0, 3, 5, 0, 0, 16, 25, 34, 69, 56, 0, 
    17, 60, 0, 3, 24, 3, 0, 23, 61, 53, 38, 69, 57, 25, 0, 
    0, 0, 0, 79, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
    0, 23, 37, 0, 29, 16, 37, 19, 54, 37, 53, 44, 34, 39, 0, 
    0, 0, 0, 0, 8, 9, 0, 9, 7, 0, 0, 0, 12, 0, 0, 
    6, 45, 0, 0, 0, 17, 73, 39, 25, 26, 0, 35, 48, 60, 0, 
    1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 19, 0, 0, 
    0, 17, 0, 10, 0, 0, 0, 0, 0, 62, 38, 26, 1, 0, 0, 
    12, 0, 0, 22, 5, 0, 0, 0, 0, 2, 25, 12, 0, 0, 0, 
    
    -- channel=294
    134, 135, 138, 103, 100, 104, 119, 138, 145, 135, 130, 122, 136, 123, 114, 
    148, 148, 153, 106, 82, 75, 64, 66, 80, 82, 98, 119, 123, 115, 103, 
    145, 144, 143, 127, 64, 101, 100, 111, 94, 75, 73, 130, 129, 100, 70, 
    144, 149, 119, 130, 76, 114, 133, 103, 111, 107, 113, 84, 118, 131, 87, 
    138, 149, 115, 88, 77, 82, 91, 91, 96, 95, 119, 102, 135, 154, 140, 
    111, 144, 110, 101, 21, 67, 80, 66, 63, 66, 64, 65, 101, 145, 144, 
    104, 102, 68, 71, 93, 85, 89, 71, 72, 90, 66, 51, 66, 78, 132, 
    107, 58, 40, 119, 52, 43, 31, 36, 5, 0, 15, 3, 7, 52, 87, 
    122, 87, 67, 28, 42, 56, 74, 84, 97, 101, 136, 106, 103, 96, 64, 
    123, 89, 34, 34, 19, 37, 19, 18, 78, 52, 59, 52, 71, 47, 26, 
    115, 100, 48, 38, 14, 0, 46, 64, 4, 56, 44, 54, 44, 63, 42, 
    120, 84, 12, 80, 53, 6, 0, 9, 2, 53, 79, 77, 37, 13, 0, 
    101, 125, 87, 83, 56, 31, 0, 0, 0, 67, 141, 141, 24, 5, 33, 
    110, 106, 90, 76, 49, 42, 7, 10, 26, 32, 44, 100, 9, 9, 31, 
    100, 99, 104, 49, 39, 30, 22, 23, 22, 27, 32, 55, 23, 9, 41, 
    
    -- channel=295
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=296
    36, 38, 37, 23, 29, 35, 26, 32, 39, 35, 33, 40, 22, 26, 12, 
    47, 47, 34, 9, 39, 54, 59, 54, 55, 46, 30, 48, 40, 16, 33, 
    52, 53, 33, 0, 59, 56, 57, 48, 53, 62, 61, 44, 34, 11, 39, 
    52, 46, 48, 0, 78, 61, 45, 63, 58, 60, 55, 63, 35, 10, 21, 
    54, 42, 32, 17, 67, 74, 51, 65, 67, 70, 51, 69, 53, 23, 34, 
    66, 35, 30, 9, 62, 59, 55, 56, 56, 67, 60, 70, 80, 52, 53, 
    63, 30, 45, 21, 45, 57, 44, 44, 53, 41, 33, 58, 70, 68, 61, 
    40, 21, 59, 10, 50, 44, 48, 34, 33, 35, 31, 35, 62, 76, 91, 
    35, 1, 56, 5, 51, 39, 33, 11, 22, 32, 0, 9, 46, 45, 94, 
    37, 0, 33, 7, 40, 26, 46, 71, 41, 65, 51, 54, 50, 34, 108, 
    49, 0, 24, 11, 17, 32, 43, 15, 60, 35, 42, 56, 27, 47, 89, 
    53, 0, 31, 25, 0, 17, 49, 0, 60, 26, 29, 44, 2, 35, 104, 
    59, 5, 33, 29, 6, 0, 2, 10, 27, 62, 22, 0, 0, 26, 94, 
    61, 45, 27, 18, 26, 0, 2, 11, 23, 57, 63, 0, 0, 38, 89, 
    55, 50, 26, 16, 24, 5, 7, 13, 22, 35, 51, 10, 0, 32, 98, 
    
    -- channel=297
    25, 18, 24, 27, 24, 20, 26, 16, 25, 34, 31, 33, 26, 24, 25, 
    28, 28, 38, 33, 17, 7, 5, 24, 34, 36, 36, 27, 36, 40, 30, 
    28, 27, 40, 6, 0, 0, 0, 0, 0, 0, 6, 30, 35, 43, 32, 
    27, 31, 18, 27, 0, 2, 0, 0, 0, 0, 0, 23, 34, 37, 31, 
    29, 33, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 33, 6, 
    30, 43, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 27, 
    21, 43, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 33, 28, 
    44, 29, 1, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    26, 13, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    27, 7, 20, 0, 0, 0, 0, 0, 4, 0, 0, 0, 1, 0, 0, 
    23, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 8, 1, 0, 0, 0, 0, 0, 0, 11, 0, 5, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 15, 23, 0, 0, 0, 
    0, 7, 0, 11, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 
    
    -- channel=298
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 11, 0, 0, 0, 0, 0, 4, 34, 18, 21, 33, 0, 0, 0, 
    0, 8, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 18, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 0, 1, 11, 0, 0, 4, 0, 0, 0, 0, 9, 0, 0, 
    0, 37, 0, 0, 11, 12, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 13, 12, 4, 0, 0, 0, 0, 19, 0, 0, 
    0, 0, 0, 0, 0, 3, 7, 3, 0, 0, 0, 0, 13, 0, 0, 
    
    -- channel=299
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=300
    13, 23, 7, 0, 7, 14, 26, 52, 46, 14, 13, 17, 0, 34, 2, 
    10, 12, 0, 0, 0, 0, 0, 0, 0, 6, 5, 32, 12, 0, 39, 
    7, 8, 0, 0, 10, 4, 0, 0, 0, 7, 50, 26, 1, 0, 50, 
    6, 0, 0, 0, 55, 4, 0, 0, 0, 0, 9, 39, 0, 0, 21, 
    9, 0, 0, 0, 29, 0, 0, 0, 0, 0, 0, 44, 28, 0, 26, 
    22, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 6, 52, 6, 8, 
    18, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 26, 25, 5, 17, 
    0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 10, 62, 
    0, 0, 56, 0, 19, 7, 0, 0, 40, 52, 0, 35, 71, 3, 64, 
    0, 0, 9, 0, 16, 0, 5, 24, 0, 0, 0, 0, 0, 0, 85, 
    0, 0, 12, 0, 0, 6, 24, 0, 22, 0, 0, 29, 0, 17, 66, 
    0, 0, 14, 15, 0, 15, 22, 0, 73, 0, 5, 22, 0, 4, 75, 
    0, 0, 37, 0, 0, 0, 5, 11, 21, 103, 13, 0, 0, 18, 99, 
    4, 0, 0, 0, 0, 0, 11, 20, 32, 39, 0, 0, 0, 48, 68, 
    0, 0, 0, 0, 0, 0, 5, 11, 13, 13, 14, 0, 0, 36, 96, 
    
    -- channel=301
    24, 18, 24, 35, 16, 10, 6, 0, 5, 24, 21, 23, 23, 11, 23, 
    28, 28, 35, 60, 50, 52, 59, 68, 53, 38, 34, 17, 25, 30, 8, 
    33, 32, 46, 58, 44, 44, 45, 52, 63, 58, 18, 19, 25, 33, 15, 
    33, 35, 42, 77, 11, 29, 51, 66, 54, 51, 42, 24, 32, 17, 11, 
    31, 38, 61, 79, 34, 55, 72, 59, 56, 55, 64, 22, 17, 36, 5, 
    22, 40, 29, 61, 46, 52, 57, 56, 61, 51, 58, 47, 19, 33, 32, 
    19, 50, 30, 42, 22, 44, 55, 48, 36, 41, 43, 31, 44, 47, 27, 
    13, 51, 1, 17, 50, 54, 51, 40, 36, 42, 36, 30, 41, 45, 21, 
    18, 32, 0, 73, 16, 15, 19, 33, 0, 0, 2, 0, 0, 19, 16, 
    30, 52, 23, 25, 31, 41, 41, 23, 61, 58, 69, 64, 51, 64, 5, 
    29, 56, 14, 25, 21, 25, 12, 32, 28, 42, 38, 19, 53, 10, 7, 
    43, 71, 18, 9, 30, 10, 25, 53, 0, 28, 20, 20, 51, 42, 3, 
    45, 40, 3, 31, 36, 22, 12, 11, 12, 0, 3, 28, 31, 13, 0, 
    33, 52, 46, 35, 30, 33, 8, 5, 0, 33, 53, 69, 27, 0, 8, 
    54, 50, 49, 50, 27, 30, 14, 14, 16, 20, 25, 54, 23, 7, 0, 
    
    -- channel=302
    14, 8, 30, 51, 4, 0, 0, 0, 0, 9, 20, 2, 24, 15, 24, 
    6, 6, 40, 73, 15, 0, 0, 12, 0, 0, 11, 2, 14, 52, 0, 
    10, 10, 36, 119, 0, 0, 0, 0, 2, 7, 0, 1, 46, 61, 0, 
    10, 26, 20, 111, 0, 0, 15, 0, 0, 0, 7, 0, 18, 54, 22, 
    5, 33, 52, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 5, 
    0, 49, 19, 86, 0, 0, 1, 0, 0, 0, 0, 0, 0, 10, 9, 
    5, 63, 29, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 84, 0, 62, 0, 18, 18, 34, 0, 0, 18, 0, 0, 0, 0, 
    33, 60, 0, 74, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    34, 111, 0, 37, 0, 19, 0, 0, 25, 5, 24, 12, 4, 35, 0, 
    18, 99, 20, 20, 18, 0, 0, 65, 0, 37, 14, 0, 49, 0, 0, 
    16, 132, 0, 1, 52, 3, 0, 41, 0, 0, 0, 7, 53, 9, 0, 
    0, 50, 0, 24, 31, 44, 4, 0, 0, 0, 0, 80, 39, 0, 0, 
    0, 21, 41, 27, 3, 51, 3, 0, 0, 0, 0, 113, 28, 0, 0, 
    1, 0, 41, 36, 4, 21, 5, 0, 0, 0, 0, 44, 33, 0, 0, 
    
    -- channel=303
    32, 22, 35, 7, 38, 33, 52, 41, 28, 36, 19, 31, 45, 13, 31, 
    35, 33, 43, 14, 28, 22, 0, 3, 26, 29, 19, 19, 27, 20, 25, 
    29, 27, 50, 32, 37, 32, 32, 32, 14, 0, 27, 31, 14, 22, 0, 
    29, 34, 14, 73, 22, 61, 30, 41, 53, 43, 0, 19, 40, 37, 0, 
    28, 39, 7, 58, 34, 0, 50, 31, 25, 16, 57, 14, 35, 68, 34, 
    19, 43, 44, 24, 0, 27, 14, 17, 19, 7, 15, 0, 11, 29, 28, 
    0, 30, 0, 49, 23, 15, 59, 26, 30, 52, 16, 0, 0, 12, 40, 
    29, 0, 17, 44, 13, 3, 0, 0, 0, 0, 0, 0, 0, 0, 28, 
    28, 20, 0, 0, 19, 9, 48, 64, 41, 23, 94, 49, 7, 13, 0, 
    40, 0, 29, 0, 0, 11, 0, 0, 23, 0, 5, 3, 34, 0, 0, 
    26, 53, 0, 23, 0, 1, 26, 0, 9, 0, 3, 20, 0, 38, 0, 
    31, 17, 41, 36, 12, 0, 0, 44, 0, 46, 45, 0, 15, 0, 0, 
    32, 86, 0, 47, 41, 4, 3, 0, 0, 50, 63, 94, 0, 8, 0, 
    21, 39, 31, 57, 21, 31, 3, 0, 5, 0, 4, 75, 6, 0, 0, 
    28, 34, 47, 13, 18, 24, 5, 6, 0, 0, 0, 67, 0, 0, 0, 
    
    -- channel=304
    31, 31, 41, 45, 37, 26, 18, 12, 23, 33, 38, 35, 29, 27, 25, 
    36, 35, 49, 58, 38, 30, 30, 39, 42, 26, 36, 35, 41, 42, 30, 
    38, 39, 48, 59, 0, 0, 0, 0, 0, 0, 4, 36, 51, 47, 27, 
    38, 45, 38, 67, 0, 5, 23, 0, 0, 0, 0, 30, 36, 47, 38, 
    38, 46, 60, 41, 0, 0, 15, 0, 0, 0, 0, 5, 29, 38, 24, 
    39, 58, 35, 37, 0, 0, 5, 1, 0, 0, 5, 0, 12, 38, 38, 
    45, 64, 50, 22, 0, 4, 3, 0, 0, 6, 8, 9, 28, 37, 31, 
    64, 67, 19, 62, 11, 0, 6, 16, 14, 5, 13, 12, 0, 5, 5, 
    54, 45, 29, 59, 0, 18, 1, 0, 0, 0, 0, 0, 0, 14, 0, 
    48, 57, 32, 22, 9, 12, 9, 4, 29, 20, 25, 21, 30, 22, 0, 
    45, 52, 15, 17, 12, 1, 0, 26, 0, 16, 5, 0, 28, 0, 0, 
    40, 57, 10, 8, 16, 10, 15, 21, 4, 20, 14, 34, 28, 22, 0, 
    23, 12, 9, 28, 10, 14, 6, 2, 0, 0, 20, 45, 18, 0, 0, 
    22, 33, 24, 32, 11, 14, 2, 1, 3, 17, 20, 50, 12, 0, 0, 
    22, 14, 25, 24, 11, 9, 5, 4, 5, 9, 14, 27, 11, 0, 0, 
    
    -- channel=305
    29, 29, 33, 34, 31, 33, 20, 10, 29, 39, 36, 42, 15, 18, 9, 
    47, 46, 41, 48, 74, 87, 94, 104, 98, 77, 44, 46, 46, 28, 30, 
    56, 56, 48, 12, 69, 59, 60, 53, 66, 76, 63, 43, 39, 27, 43, 
    55, 54, 57, 34, 79, 81, 72, 94, 80, 74, 70, 71, 37, 5, 29, 
    58, 48, 71, 62, 88, 102, 92, 96, 95, 97, 74, 70, 52, 20, 0, 
    70, 52, 39, 45, 94, 83, 83, 96, 98, 96, 106, 100, 76, 55, 56, 
    66, 61, 66, 34, 51, 83, 84, 72, 77, 81, 62, 77, 98, 98, 66, 
    56, 56, 56, 28, 87, 65, 61, 63, 83, 82, 68, 87, 101, 100, 93, 
    34, 20, 53, 63, 60, 59, 54, 20, 0, 0, 0, 0, 13, 57, 107, 
    43, 25, 65, 24, 72, 53, 74, 89, 82, 92, 92, 89, 85, 71, 105, 
    55, 13, 28, 30, 36, 54, 40, 38, 81, 50, 55, 50, 53, 46, 91, 
    69, 34, 53, 17, 12, 38, 87, 45, 72, 59, 45, 68, 47, 77, 98, 
    80, 0, 21, 50, 23, 9, 22, 28, 37, 35, 22, 7, 30, 36, 83, 
    67, 74, 50, 47, 47, 15, 11, 19, 33, 91, 91, 38, 21, 44, 90, 
    81, 70, 44, 51, 46, 28, 17, 22, 34, 50, 75, 48, 16, 41, 78, 
    
    -- channel=306
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 38, 66, 60, 75, 97, 76, 9, 15, 0, 0, 16, 
    0, 0, 0, 0, 31, 0, 0, 0, 0, 26, 105, 0, 0, 0, 60, 
    0, 0, 0, 0, 91, 26, 0, 5, 0, 0, 0, 92, 0, 0, 0, 
    0, 0, 0, 0, 68, 27, 0, 13, 18, 10, 0, 73, 6, 0, 0, 
    35, 0, 0, 0, 71, 16, 0, 17, 22, 30, 43, 58, 84, 0, 0, 
    17, 0, 0, 0, 0, 0, 0, 0, 25, 23, 0, 71, 109, 91, 27, 
    0, 0, 74, 0, 0, 0, 0, 0, 39, 43, 17, 63, 105, 66, 146, 
    0, 0, 53, 0, 46, 14, 0, 0, 0, 0, 0, 0, 0, 0, 136, 
    0, 0, 81, 0, 57, 0, 42, 93, 2, 44, 23, 36, 54, 0, 151, 
    0, 0, 0, 0, 0, 45, 7, 0, 91, 0, 0, 14, 0, 17, 85, 
    0, 0, 80, 0, 0, 8, 93, 0, 125, 23, 0, 41, 0, 66, 147, 
    0, 0, 0, 0, 0, 0, 5, 15, 28, 114, 0, 0, 0, 37, 111, 
    0, 0, 0, 0, 0, 0, 0, 7, 28, 98, 74, 0, 0, 56, 105, 
    0, 0, 0, 0, 5, 0, 0, 0, 6, 21, 47, 0, 0, 43, 114, 
    
    -- channel=307
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 41, 58, 69, 87, 83, 54, 14, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 29, 0, 0, 2, 23, 
    0, 0, 0, 0, 4, 0, 0, 5, 0, 0, 0, 45, 0, 0, 0, 
    0, 0, 14, 10, 11, 24, 21, 4, 7, 4, 0, 4, 0, 0, 0, 
    14, 0, 0, 0, 46, 12, 3, 21, 29, 23, 38, 34, 20, 0, 0, 
    9, 17, 23, 0, 0, 0, 0, 0, 0, 2, 7, 40, 76, 70, 3, 
    2, 28, 20, 0, 18, 8, 16, 19, 51, 53, 37, 59, 72, 48, 46, 
    0, 0, 3, 44, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 
    0, 0, 50, 0, 34, 16, 43, 56, 30, 56, 56, 56, 50, 28, 44, 
    0, 0, 0, 0, 2, 26, 0, 0, 44, 0, 4, 0, 0, 0, 6, 
    0, 0, 34, 0, 0, 9, 78, 40, 44, 18, 0, 23, 15, 60, 53, 
    2, 0, 0, 0, 0, 0, 2, 4, 4, 0, 0, 0, 0, 6, 4, 
    0, 1, 0, 4, 0, 0, 0, 0, 0, 57, 66, 5, 0, 5, 17, 
    5, 0, 0, 4, 6, 0, 0, 0, 0, 9, 31, 17, 0, 5, 4, 
    
    -- channel=308
    61, 61, 60, 38, 49, 43, 50, 64, 72, 65, 63, 65, 47, 57, 38, 
    74, 74, 67, 33, 54, 67, 66, 67, 79, 63, 60, 69, 64, 45, 64, 
    77, 78, 60, 8, 50, 52, 54, 46, 52, 61, 74, 67, 55, 36, 63, 
    76, 74, 59, 18, 89, 69, 60, 72, 65, 68, 56, 81, 47, 40, 38, 
    76, 70, 58, 22, 71, 74, 57, 68, 73, 72, 64, 81, 71, 45, 50, 
    77, 65, 32, 11, 48, 54, 54, 53, 49, 59, 64, 58, 94, 76, 77, 
    62, 35, 35, 13, 50, 55, 45, 39, 57, 53, 32, 64, 81, 83, 76, 
    42, 8, 39, 31, 32, 15, 33, 25, 20, 15, 21, 23, 43, 62, 97, 
    38, 0, 44, 0, 37, 46, 23, 0, 21, 29, 3, 10, 46, 53, 81, 
    42, 0, 30, 0, 30, 13, 32, 66, 30, 61, 46, 47, 63, 17, 83, 
    55, 0, 11, 1, 1, 16, 22, 12, 26, 24, 24, 31, 24, 39, 65, 
    59, 0, 26, 21, 0, 5, 36, 0, 59, 19, 31, 64, 0, 26, 74, 
    56, 3, 34, 35, 0, 0, 0, 0, 6, 75, 43, 12, 0, 11, 75, 
    68, 47, 24, 30, 21, 0, 0, 2, 21, 49, 59, 9, 0, 27, 68, 
    57, 51, 32, 10, 18, 0, 0, 3, 10, 22, 37, 7, 0, 18, 82, 
    
    -- channel=309
    7, 0, 19, 42, 0, 0, 0, 0, 0, 0, 5, 0, 29, 0, 27, 
    0, 0, 33, 93, 3, 0, 0, 0, 0, 0, 0, 0, 0, 34, 0, 
    0, 0, 37, 168, 0, 0, 0, 20, 5, 0, 0, 0, 25, 45, 0, 
    0, 15, 13, 166, 0, 0, 43, 0, 0, 0, 0, 0, 11, 50, 0, 
    0, 25, 56, 105, 0, 0, 23, 0, 0, 0, 9, 0, 0, 46, 8, 
    0, 42, 51, 118, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 54, 9, 63, 0, 0, 15, 2, 0, 0, 5, 0, 0, 0, 0, 
    10, 78, 0, 77, 3, 17, 5, 25, 0, 0, 6, 0, 0, 0, 0, 
    34, 92, 0, 88, 0, 0, 0, 30, 0, 0, 52, 15, 0, 0, 0, 
    35, 139, 0, 62, 0, 21, 0, 0, 20, 0, 10, 0, 0, 39, 0, 
    9, 153, 5, 29, 10, 0, 0, 61, 0, 32, 6, 0, 43, 0, 0, 
    12, 165, 0, 11, 70, 0, 0, 61, 0, 0, 0, 0, 86, 0, 0, 
    0, 109, 0, 17, 54, 48, 0, 0, 0, 0, 7, 115, 46, 0, 0, 
    0, 25, 58, 26, 7, 68, 0, 0, 0, 0, 0, 124, 40, 0, 0, 
    5, 9, 55, 39, 1, 28, 4, 0, 0, 0, 0, 52, 40, 0, 0, 
    
    -- channel=310
    0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 22, 26, 59, 62, 70, 48, 16, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 0, 13, 2, 18, 27, 16, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 6, 1, 0, 5, 0, 0, 0, 40, 
    0, 0, 0, 22, 0, 6, 18, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 66, 23, 5, 22, 17, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 13, 18, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 5, 0, 1, 44, 120, 116, 97, 124, 104, 20, 0, 
    0, 1, 0, 15, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 31, 10, 14, 0, 43, 38, 0, 24, 17, 33, 9, 27, 0, 
    0, 0, 0, 55, 39, 10, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 64, 79, 0, 23, 36, 11, 12, 16, 24, 26, 21, 6, 11, 26, 
    2, 0, 5, 0, 5, 19, 28, 28, 18, 0, 0, 0, 8, 19, 6, 
    0, 0, 14, 0, 1, 8, 30, 28, 21, 8, 0, 0, 28, 15, 32, 
    
    -- channel=311
    20, 26, 19, 3, 0, 17, 30, 56, 24, 0, 0, 0, 34, 26, 23, 
    6, 7, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 60, 0, 44, 52, 65, 28, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 29, 0, 0, 23, 0, 5, 20, 14, 0, 0, 38, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 41, 87, 
    0, 0, 19, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 60, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    37, 42, 0, 0, 0, 0, 6, 67, 140, 139, 146, 155, 112, 25, 0, 
    10, 36, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 47, 26, 6, 0, 0, 32, 39, 0, 15, 0, 17, 6, 15, 0, 
    0, 15, 0, 61, 52, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 
    0, 102, 85, 0, 29, 37, 0, 0, 0, 13, 66, 66, 7, 0, 0, 
    2, 0, 14, 0, 0, 27, 19, 15, 5, 0, 0, 0, 5, 0, 0, 
    0, 0, 22, 0, 0, 6, 22, 17, 5, 0, 0, 0, 29, 0, 0, 
    
    -- channel=312
    128, 120, 136, 115, 104, 104, 115, 122, 122, 130, 124, 117, 139, 108, 113, 
    143, 141, 158, 143, 90, 84, 71, 79, 92, 84, 96, 106, 121, 122, 90, 
    142, 140, 156, 171, 68, 100, 105, 116, 92, 65, 51, 116, 129, 115, 48, 
    141, 149, 126, 189, 69, 125, 156, 124, 129, 121, 96, 73, 123, 136, 78, 
    136, 154, 138, 143, 75, 91, 125, 109, 113, 108, 140, 76, 121, 157, 123, 
    110, 160, 142, 146, 28, 85, 102, 92, 87, 83, 89, 64, 81, 142, 140, 
    99, 133, 86, 118, 93, 97, 127, 92, 91, 112, 85, 48, 56, 85, 127, 
    122, 97, 41, 144, 78, 65, 49, 71, 42, 33, 49, 33, 16, 52, 63, 
    132, 125, 49, 77, 53, 78, 94, 102, 86, 80, 140, 90, 72, 109, 34, 
    138, 138, 42, 70, 24, 59, 22, 29, 93, 62, 81, 67, 88, 78, 0, 
    124, 160, 49, 60, 28, 14, 45, 84, 5, 75, 60, 49, 70, 79, 9, 
    130, 146, 24, 84, 79, 12, 0, 67, 0, 80, 87, 81, 90, 18, 0, 
    117, 167, 69, 98, 89, 51, 13, 9, 0, 44, 142, 178, 53, 12, 0, 
    114, 128, 124, 99, 69, 76, 15, 14, 28, 13, 57, 150, 41, 0, 4, 
    117, 116, 128, 76, 57, 57, 29, 29, 26, 32, 38, 99, 44, 4, 4, 
    
    -- channel=313
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 28, 42, 44, 59, 83, 71, 44, 10, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 1, 0, 0, 12, 9, 
    0, 0, 0, 11, 0, 0, 0, 1, 0, 0, 0, 20, 0, 0, 0, 
    0, 0, 36, 29, 0, 12, 23, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 0, 0, 25, 0, 1, 18, 25, 9, 35, 16, 0, 0, 0, 
    0, 32, 21, 0, 0, 0, 1, 0, 0, 10, 8, 17, 53, 49, 0, 
    6, 41, 0, 0, 14, 0, 0, 16, 44, 40, 31, 51, 38, 23, 7, 
    0, 0, 0, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 8, 40, 0, 27, 12, 29, 19, 34, 37, 51, 44, 43, 30, 0, 
    0, 0, 0, 0, 1, 5, 0, 0, 6, 0, 0, 0, 12, 0, 0, 
    2, 35, 10, 0, 0, 2, 56, 39, 12, 11, 0, 25, 26, 55, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    0, 9, 0, 14, 0, 0, 0, 0, 0, 43, 41, 38, 0, 0, 0, 
    4, 0, 0, 20, 1, 0, 0, 0, 0, 0, 15, 27, 0, 0, 0, 
    
    -- channel=314
    41, 37, 41, 48, 19, 22, 26, 35, 33, 39, 43, 28, 51, 48, 50, 
    35, 34, 48, 53, 0, 0, 0, 0, 0, 0, 25, 21, 33, 58, 25, 
    32, 31, 42, 80, 0, 0, 0, 0, 0, 0, 0, 25, 49, 52, 10, 
    31, 37, 29, 68, 0, 0, 21, 0, 0, 0, 5, 0, 32, 66, 36, 
    27, 41, 36, 22, 0, 0, 0, 0, 0, 0, 0, 0, 16, 50, 43, 
    6, 44, 34, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 31, 
    9, 34, 11, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    23, 37, 0, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 53, 0, 28, 0, 0, 0, 12, 21, 16, 45, 32, 7, 6, 0, 
    34, 70, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 73, 7, 4, 0, 0, 0, 35, 0, 13, 0, 0, 24, 0, 0, 
    10, 70, 0, 8, 34, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 
    0, 47, 14, 4, 14, 24, 0, 0, 0, 0, 32, 63, 20, 0, 0, 
    0, 9, 21, 6, 0, 24, 0, 0, 0, 0, 0, 42, 9, 0, 0, 
    0, 0, 19, 12, 0, 5, 0, 0, 0, 0, 0, 7, 18, 0, 0, 
    
    -- channel=315
    0, 0, 0, 38, 0, 0, 0, 0, 0, 0, 3, 0, 7, 0, 15, 
    0, 0, 0, 76, 0, 0, 30, 15, 0, 2, 4, 0, 0, 16, 0, 
    0, 0, 5, 69, 0, 0, 5, 4, 0, 1, 0, 0, 3, 12, 0, 
    0, 0, 30, 42, 0, 0, 17, 0, 0, 6, 14, 0, 4, 0, 17, 
    0, 0, 53, 54, 0, 22, 19, 0, 1, 23, 0, 0, 0, 0, 1, 
    0, 0, 50, 43, 0, 0, 9, 7, 7, 0, 2, 14, 0, 0, 0, 
    0, 22, 24, 35, 4, 11, 0, 16, 2, 0, 33, 7, 0, 14, 0, 
    0, 73, 0, 0, 18, 15, 5, 9, 11, 15, 12, 10, 0, 13, 0, 
    13, 89, 0, 81, 0, 15, 20, 21, 0, 3, 0, 0, 0, 13, 0, 
    8, 94, 0, 79, 0, 19, 7, 34, 0, 7, 16, 5, 0, 58, 6, 
    3, 92, 0, 10, 30, 5, 0, 38, 0, 9, 0, 0, 55, 0, 42, 
    6, 108, 0, 0, 45, 17, 8, 42, 0, 17, 0, 0, 107, 0, 40, 
    3, 34, 5, 0, 28, 24, 5, 2, 17, 0, 0, 0, 56, 0, 0, 
    0, 3, 24, 0, 3, 31, 3, 1, 0, 0, 3, 0, 51, 0, 8, 
    7, 10, 0, 31, 0, 20, 8, 0, 1, 0, 0, 0, 47, 0, 0, 
    
    -- channel=316
    127, 116, 128, 112, 100, 99, 113, 119, 128, 138, 132, 126, 135, 115, 118, 
    141, 139, 155, 127, 90, 84, 73, 94, 112, 117, 114, 115, 129, 136, 105, 
    140, 139, 151, 121, 35, 56, 56, 66, 54, 54, 67, 122, 133, 130, 79, 
    139, 146, 117, 143, 51, 110, 117, 91, 91, 86, 95, 89, 126, 134, 93, 
    136, 149, 126, 104, 55, 66, 92, 77, 85, 79, 113, 82, 124, 147, 100, 
    114, 157, 109, 99, 15, 51, 62, 63, 62, 55, 71, 65, 87, 141, 139, 
    96, 125, 75, 78, 49, 60, 90, 58, 58, 95, 73, 49, 78, 102, 135, 
    116, 82, 37, 112, 46, 33, 13, 40, 31, 22, 30, 31, 16, 37, 81, 
    110, 93, 48, 62, 35, 59, 73, 70, 37, 36, 97, 45, 27, 79, 58, 
    121, 100, 52, 37, 16, 38, 10, 15, 85, 43, 67, 54, 77, 55, 0, 
    111, 118, 34, 38, 7, 2, 15, 48, 0, 38, 30, 20, 35, 49, 8, 
    113, 110, 23, 53, 50, 0, 0, 56, 0, 77, 73, 78, 69, 22, 0, 
    94, 112, 33, 81, 60, 27, 3, 0, 0, 39, 122, 147, 35, 0, 0, 
    89, 107, 92, 84, 48, 54, 2, 1, 15, 26, 52, 130, 21, 0, 0, 
    92, 89, 97, 56, 40, 40, 12, 12, 9, 16, 26, 85, 22, 0, 0, 
    
    -- channel=317
    27, 21, 25, 17, 23, 24, 24, 22, 30, 34, 27, 32, 21, 17, 18, 
    36, 35, 34, 27, 49, 58, 58, 66, 65, 55, 35, 32, 31, 22, 24, 
    40, 41, 37, 15, 61, 57, 54, 51, 55, 56, 44, 29, 22, 19, 26, 
    40, 39, 37, 31, 75, 71, 62, 89, 80, 75, 53, 47, 29, 10, 11, 
    41, 39, 36, 54, 72, 77, 79, 85, 84, 81, 74, 49, 34, 21, 1, 
    41, 39, 32, 37, 68, 71, 69, 78, 79, 77, 82, 69, 53, 40, 40, 
    30, 29, 26, 38, 39, 66, 75, 63, 65, 71, 54, 54, 63, 61, 51, 
    18, 13, 27, 11, 62, 55, 50, 50, 58, 59, 51, 57, 66, 60, 65, 
    9, 4, 19, 28, 52, 42, 48, 24, 2, 5, 4, 0, 13, 43, 62, 
    25, 8, 35, 12, 43, 39, 44, 55, 55, 57, 61, 58, 59, 48, 58, 
    30, 11, 19, 22, 21, 38, 32, 20, 55, 35, 43, 40, 28, 45, 45, 
    44, 18, 35, 23, 11, 18, 47, 40, 37, 45, 36, 43, 32, 47, 54, 
    55, 23, 8, 42, 26, 9, 15, 18, 23, 40, 27, 22, 18, 28, 41, 
    49, 53, 42, 39, 38, 19, 10, 14, 20, 48, 60, 42, 15, 25, 54, 
    61, 56, 43, 35, 37, 25, 13, 17, 22, 32, 44, 46, 9, 25, 52, 
    
    -- channel=318
    37, 34, 42, 26, 30, 7, 0, 0, 31, 55, 54, 63, 20, 29, 21, 
    52, 52, 53, 7, 44, 52, 57, 86, 100, 93, 78, 69, 69, 58, 67, 
    64, 65, 53, 0, 0, 0, 0, 0, 0, 13, 64, 61, 54, 56, 85, 
    64, 66, 48, 0, 6, 0, 0, 3, 0, 0, 4, 100, 50, 17, 37, 
    67, 62, 41, 0, 12, 12, 12, 0, 4, 0, 1, 38, 49, 25, 0, 
    79, 65, 0, 0, 21, 0, 0, 1, 11, 14, 37, 48, 84, 64, 65, 
    62, 57, 42, 0, 0, 0, 0, 0, 0, 0, 0, 24, 92, 100, 79, 
    50, 20, 28, 0, 0, 0, 0, 0, 14, 14, 0, 22, 44, 31, 101, 
    6, 0, 24, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 67, 
    27, 0, 48, 0, 10, 0, 11, 20, 32, 40, 42, 42, 50, 0, 44, 
    38, 0, 0, 0, 0, 0, 0, 0, 34, 0, 0, 0, 0, 0, 5, 
    31, 0, 15, 0, 0, 0, 41, 0, 14, 6, 0, 31, 0, 44, 26, 
    26, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 21, 0, 8, 0, 0, 0, 0, 0, 56, 60, 12, 0, 0, 5, 
    17, 1, 0, 0, 0, 0, 0, 0, 0, 0, 15, 8, 0, 0, 3, 
    
    -- channel=319
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 0, 0, 0, 6, 7, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 19, 16, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 17, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 12, 22, 6, 0, 0, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    
    
    others => 0);
end gold_package;
