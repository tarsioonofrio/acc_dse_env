library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    -11, 313, -277, -14, 5, 234, 184, -488, 251, -170, 663, 806, -343, 233, 92, 293, -118, -663, -225, -760, 911, 382, -307, 159, -85, -306, -572, -462, 777, -455, 779, -175, -433, 303, -128, 1178, -748, -308, 86, -576, -293, -225, -214, 165, 925, 374, 537, -108, -49, -1201, -1428, 690, -226, 75, -154, 569, 1354, -237, -765, 135, -1192, 765, -228, 473, -448, 1488, 815, -463, -761, -581, -559, -658, -208, -165, 494, 605, 541, 677, -216, -522, 72, -215, -315, 369, 812, 1069, 163, -101, -761, -1149, 1339, 42, -336, 464, -301, -534, -1128, 308, -241, 344, 
    
    
    others => 0);
end gold_package;
