library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package inmem_package is
  type mem is array(0 to 4000000) of integer;

  constant input_mem : mem := (
    -- bias
    -1951, -2797, -14671, 3654, 3015, 1817, 2111, -762, 5167, -2454, -1388, -1390, 2736, -2045, 2488, 1138, -4497, -2030, -1124, 3216, -3699, 2732, 4299, 1974, -6667, 3268, -4680, -5118, 482, 3638, 4848, 1600,

    -- weights
    -- filter=0 channel=0
    -14, 2, 5, 13, 12, 4, -12, -20, -5,
    -- filter=0 channel=1
    -18, -8, 0, 3, -11, 7, 12, -17, 2,
    -- filter=0 channel=2
    17, -7, 15, 16, 12, -13, 5, -19, 18,
    -- filter=0 channel=3
    9, 18, -18, 17, 19, 5, 11, -14, 3,
    -- filter=0 channel=4
    14, -19, -15, -7, -2, -10, -5, -8, -13,
    -- filter=0 channel=5
    -10, -17, 0, 2, 1, 4, 15, 7, 6,
    -- filter=0 channel=6
    -2, -4, 7, 12, 0, 6, 2, 17, -5,
    -- filter=0 channel=7
    -1, 3, 15, -21, -8, 13, 12, -18, 6,
    -- filter=0 channel=8
    -11, 14, 9, -15, 17, 0, -4, 16, 7,
    -- filter=0 channel=9
    -3, 7, 1, -11, -14, -13, 4, -11, -1,
    -- filter=0 channel=10
    -12, -3, 1, -4, -16, 20, -11, 8, -10,
    -- filter=0 channel=11
    6, 8, -5, 19, -8, 11, -19, 5, -10,
    -- filter=0 channel=12
    11, -13, 17, -20, 0, 7, -1, -3, 19,
    -- filter=0 channel=13
    -16, 16, 14, 10, 3, 0, -1, -14, 6,
    -- filter=0 channel=14
    9, 6, -16, 14, -20, 20, -14, 0, -10,
    -- filter=0 channel=15
    -13, 16, 13, -3, 16, -14, -8, -3, 9,
    -- filter=1 channel=0
    -9, 12, 0, 4, -20, -9, -18, -8, -17,
    -- filter=1 channel=1
    18, -11, 19, 6, 7, -5, 0, -19, 11,
    -- filter=1 channel=2
    -6, -5, 12, 0, 20, -16, -19, 13, 0,
    -- filter=1 channel=3
    1, 9, 18, -7, -16, 14, -15, 15, -13,
    -- filter=1 channel=4
    18, -17, -20, 4, 0, 19, -10, 12, 8,
    -- filter=1 channel=5
    13, -2, 8, 7, 13, -18, -6, 13, 12,
    -- filter=1 channel=6
    -1, -6, -7, 8, 2, -19, -16, 11, 0,
    -- filter=1 channel=7
    17, 10, -10, 7, 17, -12, 0, -14, 17,
    -- filter=1 channel=8
    -1, -14, -4, 10, 3, -19, -21, 7, -14,
    -- filter=1 channel=9
    -9, 7, -1, 20, -12, 14, 0, -15, 13,
    -- filter=1 channel=10
    -4, 13, 5, 10, 11, -12, -18, 0, -16,
    -- filter=1 channel=11
    0, 6, -13, 17, -19, -6, 17, 11, 16,
    -- filter=1 channel=12
    20, -9, -3, 9, 3, 1, -19, 0, 4,
    -- filter=1 channel=13
    -16, 3, -1, -19, -20, 10, 4, 0, -2,
    -- filter=1 channel=14
    -17, -6, -13, 18, -16, -11, 9, 11, -6,
    -- filter=1 channel=15
    -16, -9, 18, 10, -2, 1, -19, -2, -11,
    -- filter=2 channel=0
    -53, -50, -8, -39, -53, -51, -39, -26, -41,
    -- filter=2 channel=1
    -6, 0, 18, 23, 15, 27, 17, 34, 28,
    -- filter=2 channel=2
    -22, -20, -1, -29, -16, 1, -10, -18, -9,
    -- filter=2 channel=3
    -8, -38, -27, -47, -43, -43, -21, -33, -23,
    -- filter=2 channel=4
    20, 35, 12, 23, 20, 12, 24, 1, 23,
    -- filter=2 channel=5
    12, 6, 19, 25, 2, 18, 15, 13, 0,
    -- filter=2 channel=6
    -4, -7, -5, -13, -10, -27, 3, -28, -12,
    -- filter=2 channel=7
    3, 2, -36, 0, -11, -12, 14, -31, -32,
    -- filter=2 channel=8
    4, 6, 17, 6, 17, 13, -7, 8, -17,
    -- filter=2 channel=9
    11, 13, 32, 52, 53, 15, 53, 26, 38,
    -- filter=2 channel=10
    32, 23, -11, 35, 30, 23, 27, 24, 16,
    -- filter=2 channel=11
    -17, -29, -38, -35, 0, -14, -12, -25, -18,
    -- filter=2 channel=12
    14, 18, 0, 1, -16, 3, -17, -12, 6,
    -- filter=2 channel=13
    12, 54, 25, 66, 54, 40, 55, 67, 46,
    -- filter=2 channel=14
    -25, 14, 18, 4, 16, -15, -25, -1, 19,
    -- filter=2 channel=15
    2, -29, -5, -4, -28, -13, 0, -30, -24,
    -- filter=3 channel=0
    22, 16, 16, -7, -1, 10, -14, 18, 11,
    -- filter=3 channel=1
    13, -15, -4, -19, 10, 6, -9, -18, 14,
    -- filter=3 channel=2
    1, 17, -12, 21, 11, 15, 16, 16, 12,
    -- filter=3 channel=3
    -8, -18, 4, -6, 12, -5, 0, -10, -2,
    -- filter=3 channel=4
    15, 15, 25, 15, -18, -7, -22, 21, 11,
    -- filter=3 channel=5
    -15, -8, -9, 16, 8, -1, -3, 23, 10,
    -- filter=3 channel=6
    16, 12, -5, 3, 10, 4, 19, -9, -13,
    -- filter=3 channel=7
    2, 9, 7, -11, 7, 12, -2, 16, -2,
    -- filter=3 channel=8
    6, 2, 2, -10, 2, -9, 8, -7, 5,
    -- filter=3 channel=9
    18, 14, 17, -17, 0, -10, -1, -17, 23,
    -- filter=3 channel=10
    -24, 7, 3, -24, 16, 13, 20, -8, -14,
    -- filter=3 channel=11
    1, 1, -18, 20, -9, 20, -13, -18, 14,
    -- filter=3 channel=12
    -19, 8, -15, 12, 8, -12, -20, 7, 15,
    -- filter=3 channel=13
    -14, -4, 17, -14, -18, 8, 0, 0, 13,
    -- filter=3 channel=14
    12, -14, -12, 18, -12, -7, 4, 9, -15,
    -- filter=3 channel=15
    11, -13, 20, 13, 1, 16, 2, 1, -11,
    -- filter=4 channel=0
    8, -9, -13, -15, -3, 29, -5, 14, 9,
    -- filter=4 channel=1
    6, 33, 23, 0, 14, 27, 24, -5, 25,
    -- filter=4 channel=2
    -20, 8, -12, 5, -22, -17, -19, 6, 12,
    -- filter=4 channel=3
    10, 16, 24, 8, 15, 39, 0, 29, 28,
    -- filter=4 channel=4
    -9, -6, 0, -12, -30, -18, -32, -14, -19,
    -- filter=4 channel=5
    29, 23, 42, 26, 19, 14, -5, 20, 33,
    -- filter=4 channel=6
    -10, -4, 31, 7, 18, 15, -9, 15, 5,
    -- filter=4 channel=7
    2, -12, -19, 5, -27, -28, -24, 0, -25,
    -- filter=4 channel=8
    8, -10, 0, 6, 10, 1, 1, -4, 5,
    -- filter=4 channel=9
    -36, -13, -7, -32, -21, -32, -13, -37, -12,
    -- filter=4 channel=10
    30, 25, 24, -7, -9, 11, -20, 16, 17,
    -- filter=4 channel=11
    2, -6, 12, -22, 2, -6, 14, 14, 4,
    -- filter=4 channel=12
    8, 14, 3, 19, -10, 10, 2, -10, 1,
    -- filter=4 channel=13
    34, 28, 40, -10, -2, 5, 8, -8, 9,
    -- filter=4 channel=14
    34, 8, 45, 29, 13, 36, 10, 12, 13,
    -- filter=4 channel=15
    -21, 8, -9, -19, -1, -6, -32, -32, 2,
    -- filter=5 channel=0
    18, 6, -17, -7, -8, 0, 14, -15, -8,
    -- filter=5 channel=1
    6, -17, 18, -2, 21, -13, -24, 13, -1,
    -- filter=5 channel=2
    -8, -8, -17, 28, 0, -2, 14, 4, -7,
    -- filter=5 channel=3
    6, -5, -15, -11, 0, 8, -8, 0, -18,
    -- filter=5 channel=4
    -2, 1, 0, -9, -1, 1, -14, 0, -10,
    -- filter=5 channel=5
    12, 15, 1, -15, 15, 25, -24, 21, 6,
    -- filter=5 channel=6
    16, -7, -4, -17, -19, 4, 9, 2, 11,
    -- filter=5 channel=7
    0, -9, 2, -4, -3, -1, 24, 7, 15,
    -- filter=5 channel=8
    17, -7, -10, -16, 14, 1, 15, 2, -5,
    -- filter=5 channel=9
    17, 0, 8, 20, 0, 10, 0, -12, 18,
    -- filter=5 channel=10
    -15, 1, 12, -10, 11, 26, 19, 7, -15,
    -- filter=5 channel=11
    9, 2, 6, 5, 4, -10, 8, -18, -12,
    -- filter=5 channel=12
    -9, 7, -19, 17, 0, -6, -17, -7, 14,
    -- filter=5 channel=13
    -24, 22, 27, -32, -10, 26, -28, 23, -1,
    -- filter=5 channel=14
    -13, -1, 2, -5, -11, -14, -4, -18, -6,
    -- filter=5 channel=15
    24, 0, -13, 23, -6, -2, 12, 9, -19,
    -- filter=6 channel=0
    -2, 23, -9, 10, 5, -13, 13, 23, -13,
    -- filter=6 channel=1
    20, 12, -11, 14, 8, -15, -3, 20, -25,
    -- filter=6 channel=2
    -4, 8, 23, 1, -13, 25, -10, -17, 1,
    -- filter=6 channel=3
    -2, -7, 0, -17, -8, -17, -10, -17, -19,
    -- filter=6 channel=4
    16, 20, 11, 13, 27, -20, 22, 20, -19,
    -- filter=6 channel=5
    -3, -14, -27, -14, -21, -5, -5, 15, -16,
    -- filter=6 channel=6
    -6, -4, 10, -11, 4, 14, 5, -10, -2,
    -- filter=6 channel=7
    -8, 0, -4, -10, 17, 9, 4, 17, 13,
    -- filter=6 channel=8
    -13, -12, -15, 16, -6, 0, 0, 14, 0,
    -- filter=6 channel=9
    26, 11, 24, 13, 10, -15, 8, 1, -15,
    -- filter=6 channel=10
    5, -12, 5, 28, -17, 4, 29, -7, -9,
    -- filter=6 channel=11
    0, 11, -15, -8, 22, -3, 10, -8, -17,
    -- filter=6 channel=12
    -8, 17, -4, 19, -12, -13, 6, -12, 21,
    -- filter=6 channel=13
    23, -7, -5, 24, 19, -9, 39, 10, -35,
    -- filter=6 channel=14
    -5, -8, -26, 11, 15, -4, -7, 18, 13,
    -- filter=6 channel=15
    22, 14, 10, 6, 8, -3, 20, -11, 0,
    -- filter=7 channel=0
    -13, -16, -14, -31, -28, -27, -25, -5, 14,
    -- filter=7 channel=1
    -6, 20, -3, 14, 28, 15, -16, 15, 18,
    -- filter=7 channel=2
    6, -9, -23, -1, -14, 15, 5, 0, -20,
    -- filter=7 channel=3
    -11, -29, -9, -9, -27, -11, -10, -2, -1,
    -- filter=7 channel=4
    5, 28, 30, 7, 30, 13, 21, 17, 15,
    -- filter=7 channel=5
    -9, -4, -11, -7, 0, -19, 10, -1, -12,
    -- filter=7 channel=6
    10, 0, -10, -17, 13, 8, 3, 6, 15,
    -- filter=7 channel=7
    29, 14, -5, 0, 13, 10, -10, 11, 17,
    -- filter=7 channel=8
    13, -2, 2, 7, 7, 17, -11, 17, 15,
    -- filter=7 channel=9
    46, 36, 41, 25, 50, 42, 44, 45, 37,
    -- filter=7 channel=10
    -2, 20, 9, 15, -6, 4, 17, 31, -7,
    -- filter=7 channel=11
    -24, 12, -12, -3, 3, 8, -1, 1, -10,
    -- filter=7 channel=12
    -1, 10, 7, -11, 20, 1, 11, -14, -2,
    -- filter=7 channel=13
    28, 10, 29, 32, 16, 23, 33, 44, -5,
    -- filter=7 channel=14
    -18, -6, -3, 2, -21, -5, -25, -1, -14,
    -- filter=7 channel=15
    15, 9, 0, 0, 9, 6, 14, 14, -15,
    -- filter=8 channel=0
    -4, -20, 9, 0, 11, 0, -16, -19, 11,
    -- filter=8 channel=1
    24, 20, 11, 20, 25, 3, 29, 10, 19,
    -- filter=8 channel=2
    -5, 3, 5, 0, -11, -19, -20, -15, -12,
    -- filter=8 channel=3
    12, -2, 29, -1, 21, 15, 3, 21, 22,
    -- filter=8 channel=4
    7, -3, -18, -3, -7, -26, -24, 8, 16,
    -- filter=8 channel=5
    21, -6, 20, 6, 28, 18, 14, 4, 17,
    -- filter=8 channel=6
    19, 9, -12, 10, 0, 16, -2, 23, -5,
    -- filter=8 channel=7
    -16, -1, 2, -26, -2, -6, -15, -18, 3,
    -- filter=8 channel=8
    -13, 5, 17, 11, 20, -1, 17, 15, 7,
    -- filter=8 channel=9
    -18, -23, -31, -1, -24, -26, -7, -14, 2,
    -- filter=8 channel=10
    10, 12, 29, 9, -15, 24, -5, 12, 14,
    -- filter=8 channel=11
    -3, 17, -4, -17, 6, -18, -3, 18, 20,
    -- filter=8 channel=12
    -2, 2, -4, -5, 0, -21, 4, -5, -10,
    -- filter=8 channel=13
    17, 14, 16, -11, 6, -3, 21, 6, 2,
    -- filter=8 channel=14
    -3, 21, 33, 13, 2, -4, -1, 28, 13,
    -- filter=8 channel=15
    -28, -19, 2, -29, 0, 4, -20, 9, -13,
    -- filter=9 channel=0
    -28, -30, -13, -21, -25, -31, -22, -35, -37,
    -- filter=9 channel=1
    -10, 3, 8, -5, -1, 11, -10, 25, -7,
    -- filter=9 channel=2
    17, -13, 12, -1, -1, -28, 3, 11, -5,
    -- filter=9 channel=3
    -1, -5, -24, -2, -8, -21, -19, 6, -28,
    -- filter=9 channel=4
    7, 4, -3, -12, 6, 17, -12, 26, 25,
    -- filter=9 channel=5
    0, 2, 6, 2, 3, -8, 22, 9, 0,
    -- filter=9 channel=6
    -14, -19, 6, -3, -14, -10, -11, 0, 3,
    -- filter=9 channel=7
    18, -11, 0, 22, -17, -4, -9, -19, -19,
    -- filter=9 channel=8
    4, -20, -10, 15, -12, 7, 11, -18, -14,
    -- filter=9 channel=9
    19, 29, 0, 15, 30, 4, 12, 25, 13,
    -- filter=9 channel=10
    11, 29, 10, 4, 18, 1, 20, 17, 11,
    -- filter=9 channel=11
    -17, 11, 4, 1, 5, -3, 9, 11, 0,
    -- filter=9 channel=12
    -4, 5, 1, -14, 6, -18, 18, 16, -9,
    -- filter=9 channel=13
    27, 37, 26, 41, 14, 22, 14, 21, 11,
    -- filter=9 channel=14
    -23, -3, -9, -8, -16, -20, -4, 16, -18,
    -- filter=9 channel=15
    -9, 12, 6, -14, -7, 8, 11, 10, -20,
    -- filter=10 channel=0
    1, -22, 11, 0, -17, 12, 13, 3, -12,
    -- filter=10 channel=1
    -8, -15, 7, 17, -5, 8, -3, -15, -21,
    -- filter=10 channel=2
    0, 11, 14, -2, -16, 5, 17, 6, 11,
    -- filter=10 channel=3
    -30, -1, -2, 5, -29, -23, -9, -23, -10,
    -- filter=10 channel=4
    30, 17, 0, 24, 12, 4, -6, -9, -13,
    -- filter=10 channel=5
    8, 15, -20, 8, 12, -6, -13, 7, 12,
    -- filter=10 channel=6
    12, 6, 0, -3, -12, 19, -21, -15, 12,
    -- filter=10 channel=7
    0, 5, -18, 2, -18, -17, 20, 16, -14,
    -- filter=10 channel=8
    -6, -16, -7, 13, 2, -21, -15, -18, -13,
    -- filter=10 channel=9
    27, 36, 4, 30, 4, -8, 5, 14, 23,
    -- filter=10 channel=10
    30, 0, 4, 25, 0, 6, 26, -9, -5,
    -- filter=10 channel=11
    18, -21, 0, 18, -17, 12, 16, -1, 13,
    -- filter=10 channel=12
    0, -10, -18, 3, -20, -17, 17, 4, -18,
    -- filter=10 channel=13
    29, 26, 0, 35, -4, 0, 13, -6, -21,
    -- filter=10 channel=14
    -20, -15, -24, -16, -24, -1, -3, -4, -24,
    -- filter=10 channel=15
    23, 4, 11, 18, -7, 20, -11, -5, 5,
    -- filter=11 channel=0
    -2, -20, -4, 18, 3, -6, -7, 1, -18,
    -- filter=11 channel=1
    19, -12, 7, -4, -4, -14, -14, 5, 13,
    -- filter=11 channel=2
    8, 14, 15, 0, 14, 1, 16, 11, 9,
    -- filter=11 channel=3
    -7, 12, 2, 13, 9, 13, -12, -8, -15,
    -- filter=11 channel=4
    -17, 6, -16, 10, 1, 3, -12, 6, -13,
    -- filter=11 channel=5
    -18, 1, -9, 14, 4, 17, 5, 14, 0,
    -- filter=11 channel=6
    12, -16, 1, -12, -7, 20, -8, -20, -12,
    -- filter=11 channel=7
    5, 0, -17, -19, 6, -5, 3, -6, 20,
    -- filter=11 channel=8
    -18, -20, 7, -4, 9, 4, 9, 10, 1,
    -- filter=11 channel=9
    11, -4, -13, -20, 14, 6, 10, 16, 14,
    -- filter=11 channel=10
    -1, -18, -5, 2, 17, 18, 9, -5, 18,
    -- filter=11 channel=11
    -8, 1, 13, 15, 11, 14, -16, 19, -10,
    -- filter=11 channel=12
    -6, -4, -20, 1, -4, 7, 3, -14, 15,
    -- filter=11 channel=13
    2, -13, -12, 17, 15, 8, -13, -20, -16,
    -- filter=11 channel=14
    -2, -16, -4, -3, 0, 14, 8, 15, 20,
    -- filter=11 channel=15
    -12, 14, -7, -11, -2, 8, 7, -8, -3,
    -- filter=12 channel=0
    -10, 11, 7, -20, 20, 7, -9, 21, -2,
    -- filter=12 channel=1
    25, 11, 14, 11, -1, 5, 22, 31, 24,
    -- filter=12 channel=2
    -8, -2, -20, 5, -18, 13, 0, -2, -20,
    -- filter=12 channel=3
    1, 3, 22, 26, 26, 0, 21, 17, -8,
    -- filter=12 channel=4
    5, 10, -5, 1, -8, -18, 15, -4, 8,
    -- filter=12 channel=5
    -4, 10, -6, -2, 3, 10, 26, 23, 2,
    -- filter=12 channel=6
    -18, 6, 8, -15, 12, 12, 21, -9, -15,
    -- filter=12 channel=7
    0, -28, -26, 8, -26, 1, -25, -18, 2,
    -- filter=12 channel=8
    18, -17, 16, 11, 12, 2, -15, 4, 3,
    -- filter=12 channel=9
    1, -27, -3, -12, -17, -29, -27, 4, -12,
    -- filter=12 channel=10
    -14, 23, -12, 20, 18, 12, 16, 14, -1,
    -- filter=12 channel=11
    2, -12, 0, 12, -15, -8, 8, -10, -11,
    -- filter=12 channel=12
    12, 13, 0, -20, -10, 2, 14, -18, -9,
    -- filter=12 channel=13
    -11, 17, 5, 18, 22, 11, 1, 8, 0,
    -- filter=12 channel=14
    26, 26, 28, 11, 13, 0, 0, 25, 24,
    -- filter=12 channel=15
    13, -9, 0, -24, -26, -5, -6, 11, 9,
    -- filter=13 channel=0
    7, 7, -6, -20, -4, -18, -24, -3, 13,
    -- filter=13 channel=1
    3, 4, -11, -13, -12, 0, 7, 1, 12,
    -- filter=13 channel=2
    -9, 9, -16, -4, -11, 6, -13, 14, 6,
    -- filter=13 channel=3
    -20, -19, -13, -14, 4, 6, 0, -18, -9,
    -- filter=13 channel=4
    -12, 23, 20, 17, -1, -9, 1, 28, 0,
    -- filter=13 channel=5
    14, 7, -13, 2, 16, -24, -8, 16, 2,
    -- filter=13 channel=6
    0, 0, 1, -9, -13, 6, -23, 8, 9,
    -- filter=13 channel=7
    6, -4, -16, 23, -2, 4, 2, -12, -6,
    -- filter=13 channel=8
    -19, -15, -18, 8, -1, 17, 0, 14, 4,
    -- filter=13 channel=9
    29, 14, 10, 36, 22, 24, 20, 35, 20,
    -- filter=13 channel=10
    11, -17, 4, -6, 15, -8, 6, 13, -9,
    -- filter=13 channel=11
    5, 3, 15, 8, -21, -6, -19, -20, 15,
    -- filter=13 channel=12
    19, 5, 6, -15, 7, -16, -18, 16, -7,
    -- filter=13 channel=13
    22, -7, 0, 22, 20, 27, 29, 24, 29,
    -- filter=13 channel=14
    -1, -3, -22, -16, -5, -10, -5, 10, -11,
    -- filter=13 channel=15
    -7, -11, -12, -10, -3, 21, 3, 2, 16,
    -- filter=14 channel=0
    5, 1, 26, 11, 8, 2, 10, 13, 28,
    -- filter=14 channel=1
    2, 25, 1, 9, -2, 20, 10, 3, 34,
    -- filter=14 channel=2
    11, -12, 16, 4, -12, 8, 11, 11, -9,
    -- filter=14 channel=3
    35, 18, 24, 30, 24, -2, 12, 28, 26,
    -- filter=14 channel=4
    -29, -29, 17, -20, 0, -3, -11, -25, 22,
    -- filter=14 channel=5
    5, 27, 3, 0, 23, 30, 22, 38, 4,
    -- filter=14 channel=6
    22, 9, 4, -9, 12, 26, 15, 12, 32,
    -- filter=14 channel=7
    -22, -25, 1, -4, -12, 4, 0, -26, -17,
    -- filter=14 channel=8
    -3, -5, -14, 7, 5, -21, -18, 20, 15,
    -- filter=14 channel=9
    -22, -38, -24, -32, -13, -27, -25, -24, -18,
    -- filter=14 channel=10
    8, 5, 21, 9, 24, 9, 7, 5, -1,
    -- filter=14 channel=11
    -18, -9, 16, -11, -20, -17, 0, -11, -6,
    -- filter=14 channel=12
    4, 18, 11, 5, -7, -15, -8, 17, 2,
    -- filter=14 channel=13
    14, -4, 35, -10, 14, 38, 19, 24, 6,
    -- filter=14 channel=14
    8, 0, 35, 29, 31, 1, 17, 35, 22,
    -- filter=14 channel=15
    8, -26, -12, -13, -23, 0, 1, -19, -11,
    -- filter=15 channel=0
    -4, -10, 20, -19, 18, -4, 4, 2, 17,
    -- filter=15 channel=1
    -15, -11, 13, -3, 0, 9, 18, 0, -15,
    -- filter=15 channel=2
    -20, 14, -13, 5, -21, -20, -6, 16, -18,
    -- filter=15 channel=3
    12, 11, 0, -5, -14, -18, -20, -12, 2,
    -- filter=15 channel=4
    10, -3, 9, 3, 10, 0, -15, 1, 20,
    -- filter=15 channel=5
    -13, 9, 19, -7, 0, -10, -13, 17, 1,
    -- filter=15 channel=6
    3, -9, 3, 17, -16, -11, -13, -20, -19,
    -- filter=15 channel=7
    7, 11, -16, 2, -14, 7, -9, 11, 7,
    -- filter=15 channel=8
    14, 18, 16, 5, -14, -12, 9, 5, 16,
    -- filter=15 channel=9
    6, -2, -3, -7, 9, -3, -15, 13, -10,
    -- filter=15 channel=10
    -6, 0, -2, -19, 12, -4, -14, -12, -17,
    -- filter=15 channel=11
    -10, 11, -21, -3, -19, 12, 20, 0, -9,
    -- filter=15 channel=12
    -18, -13, -3, -21, -20, 6, 1, 12, 6,
    -- filter=15 channel=13
    2, -3, 2, 22, -14, 15, -20, -13, -7,
    -- filter=15 channel=14
    -6, 0, -12, -14, 5, -9, 3, -1, 14,
    -- filter=15 channel=15
    19, -9, 2, 13, 15, 18, 5, -18, -7,
    -- filter=16 channel=0
    -3, -6, 13, -14, -20, -15, 16, 18, -3,
    -- filter=16 channel=1
    -7, -10, -4, -2, 8, -2, -13, 10, 26,
    -- filter=16 channel=2
    13, 4, 15, 19, 22, -9, 4, 9, 1,
    -- filter=16 channel=3
    -8, 8, 15, -8, -7, 19, 14, -4, 13,
    -- filter=16 channel=4
    -11, -18, 26, -13, -2, -3, 13, 24, 31,
    -- filter=16 channel=5
    -17, 14, 25, -7, 8, 20, -15, 20, 13,
    -- filter=16 channel=6
    14, 12, 7, 10, -12, 4, -11, 18, 7,
    -- filter=16 channel=7
    0, 15, 10, -13, 2, 8, -8, 14, -1,
    -- filter=16 channel=8
    -1, 8, -19, -7, 9, -3, -2, 14, -14,
    -- filter=16 channel=9
    -16, 1, -1, 6, -19, 21, -11, 15, 11,
    -- filter=16 channel=10
    12, 24, 8, -4, 0, 24, 21, 19, 20,
    -- filter=16 channel=11
    7, -21, 1, -1, -20, -3, -16, -5, 17,
    -- filter=16 channel=12
    13, 18, -19, 19, -19, -17, -1, -21, -8,
    -- filter=16 channel=13
    -25, 18, 13, -13, 27, 3, -7, 22, 12,
    -- filter=16 channel=14
    8, -10, 0, -10, -13, 4, -8, 4, -5,
    -- filter=16 channel=15
    -2, 19, 10, -5, -16, -11, -5, 1, 12,
    -- filter=17 channel=0
    -5, 8, 0, 17, 5, -3, 16, 16, -6,
    -- filter=17 channel=1
    22, 3, -18, 17, 36, -15, 15, 19, -5,
    -- filter=17 channel=2
    0, -11, 16, 32, 13, 22, 21, 12, 6,
    -- filter=17 channel=3
    3, -11, -18, -23, -3, -10, -11, -6, -15,
    -- filter=17 channel=4
    31, 20, -10, 8, 17, -5, 34, 47, 6,
    -- filter=17 channel=5
    15, -11, -37, 6, 19, -16, 25, -13, -10,
    -- filter=17 channel=6
    15, -12, 15, 25, 19, -9, 19, 27, 17,
    -- filter=17 channel=7
    -3, 11, -9, 18, 6, 7, 31, -12, 19,
    -- filter=17 channel=8
    16, 2, 18, 14, -18, 10, 10, -4, 20,
    -- filter=17 channel=9
    31, 28, 9, 15, 31, -7, 28, 18, 3,
    -- filter=17 channel=10
    36, 2, -27, 24, -3, -3, 17, 7, -22,
    -- filter=17 channel=11
    16, 15, 1, 0, 7, 4, 3, -2, 12,
    -- filter=17 channel=12
    18, -5, -14, 19, -14, -1, 2, 8, 3,
    -- filter=17 channel=13
    33, 24, -48, 41, 29, -26, 52, 39, -4,
    -- filter=17 channel=14
    -18, 1, 4, 11, 10, 1, -9, 9, -21,
    -- filter=17 channel=15
    19, 19, 32, -14, -5, 27, 5, 8, 30,
    -- filter=18 channel=0
    13, 0, 9, 1, 13, -4, 7, 3, 10,
    -- filter=18 channel=1
    3, -15, 9, 14, 19, -9, -15, 0, -2,
    -- filter=18 channel=2
    14, 14, -16, -7, 11, -8, -11, 9, -4,
    -- filter=18 channel=3
    -8, 8, -1, -14, -1, 6, -6, 11, 7,
    -- filter=18 channel=4
    -15, 16, -18, -5, 4, -16, -4, -16, 0,
    -- filter=18 channel=5
    -15, 3, -12, -16, -14, 5, 17, -4, 13,
    -- filter=18 channel=6
    21, 14, 8, 18, 13, -17, 9, 22, 23,
    -- filter=18 channel=7
    -3, 9, -7, -5, -4, -2, 22, -6, -6,
    -- filter=18 channel=8
    15, 0, -2, 11, 0, -16, -8, -4, -2,
    -- filter=18 channel=9
    -11, 16, 21, 16, 2, -16, -19, 9, -15,
    -- filter=18 channel=10
    11, -3, 9, 24, -3, 11, 23, -18, -10,
    -- filter=18 channel=11
    11, -17, 14, 7, -4, 13, 18, 11, -7,
    -- filter=18 channel=12
    -19, 20, 16, -19, 11, -2, -4, -16, -2,
    -- filter=18 channel=13
    -11, 12, -17, -17, 20, 10, -5, 22, -13,
    -- filter=18 channel=14
    0, -14, 8, -7, 8, 20, 5, 1, 17,
    -- filter=18 channel=15
    -13, 0, 0, -13, -6, 16, -18, 19, 23,
    -- filter=19 channel=0
    12, 18, -5, 29, 15, 27, 36, 6, 25,
    -- filter=19 channel=1
    3, -15, -6, -38, -21, 24, -28, 8, 6,
    -- filter=19 channel=2
    17, 17, 4, 0, 19, 36, 25, 32, 35,
    -- filter=19 channel=3
    -9, 16, 15, 16, 4, -6, -16, 18, -11,
    -- filter=19 channel=4
    7, 18, 7, -3, -17, -1, -3, -16, 38,
    -- filter=19 channel=5
    5, 6, -11, -2, -12, 12, -27, 13, 38,
    -- filter=19 channel=6
    6, 4, 18, 5, -9, 2, 16, 19, -10,
    -- filter=19 channel=7
    25, 37, 0, 8, 27, -7, 18, -1, 31,
    -- filter=19 channel=8
    9, -8, -10, -12, 11, 11, 0, 12, -10,
    -- filter=19 channel=9
    -27, -17, 9, -13, -1, 1, -34, -8, 0,
    -- filter=19 channel=10
    10, 19, 4, 0, 10, 26, -12, 32, 36,
    -- filter=19 channel=11
    27, -7, 6, 24, -12, -6, 30, -13, 14,
    -- filter=19 channel=12
    16, 10, 13, 9, 10, -18, -17, 4, -8,
    -- filter=19 channel=13
    -26, 7, 30, -60, -19, 43, -59, -21, 60,
    -- filter=19 channel=14
    -4, -17, 14, -20, 6, 29, 11, 21, 25,
    -- filter=19 channel=15
    -1, 32, 16, 22, 7, 11, 10, 2, 26,
    -- filter=20 channel=0
    1, 16, -12, -17, 7, -17, 16, -4, -6,
    -- filter=20 channel=1
    -17, -18, -2, -26, 6, -9, -16, -2, -11,
    -- filter=20 channel=2
    -1, -10, 11, 12, -12, -8, 30, -5, 10,
    -- filter=20 channel=3
    0, -12, 1, 12, 3, -7, -7, 0, 12,
    -- filter=20 channel=4
    -6, -1, -1, 17, 33, 29, -16, 33, 24,
    -- filter=20 channel=5
    -2, 4, -22, 16, 4, -14, 13, -9, 17,
    -- filter=20 channel=6
    1, 0, 19, 10, 14, 2, 16, -15, -2,
    -- filter=20 channel=7
    16, 2, 3, 0, -6, 22, 21, 2, -18,
    -- filter=20 channel=8
    8, -19, -16, 5, 4, 14, 19, -16, -4,
    -- filter=20 channel=9
    15, 10, 15, 14, 23, 32, 27, 32, 9,
    -- filter=20 channel=10
    20, 22, 6, 8, 24, 0, 22, 13, 2,
    -- filter=20 channel=11
    -6, 6, 11, -16, 14, -9, 10, -4, 7,
    -- filter=20 channel=12
    19, -14, 5, -6, -16, 0, -1, -5, -15,
    -- filter=20 channel=13
    12, -6, 7, 6, 10, 28, -9, 28, -1,
    -- filter=20 channel=14
    -23, -16, 14, -26, 6, 0, -14, -14, 4,
    -- filter=20 channel=15
    2, 12, 14, -8, 17, 2, -16, -13, 8,
    -- filter=21 channel=0
    -16, 3, -3, -29, -4, 7, -30, -23, -7,
    -- filter=21 channel=1
    -4, 9, -10, 8, -6, 8, -9, -5, 21,
    -- filter=21 channel=2
    -5, 5, 2, 23, -8, -19, 3, -3, -5,
    -- filter=21 channel=3
    -12, -22, -30, -17, -28, -16, 4, -9, -27,
    -- filter=21 channel=4
    0, 13, -5, -6, 19, 25, 31, 24, 2,
    -- filter=21 channel=5
    -24, -28, -8, -2, -21, -20, 10, -12, -7,
    -- filter=21 channel=6
    -6, -6, -9, -5, 5, -5, 14, -21, 13,
    -- filter=21 channel=7
    -8, -8, -8, 9, -5, -4, 3, 5, -1,
    -- filter=21 channel=8
    -9, 10, -9, 14, -16, 20, 17, -19, -6,
    -- filter=21 channel=9
    34, 40, 40, 12, 28, 37, 19, 32, 15,
    -- filter=21 channel=10
    9, 20, 9, 4, 19, 14, 2, -4, -21,
    -- filter=21 channel=11
    -20, -10, 4, -7, -14, 16, 0, 3, 11,
    -- filter=21 channel=12
    -3, 9, -15, -12, -4, -20, 20, -8, -15,
    -- filter=21 channel=13
    18, 3, -2, 23, 33, 17, 7, 41, 24,
    -- filter=21 channel=14
    -22, -1, -9, -32, -31, -28, -34, -14, -21,
    -- filter=21 channel=15
    -5, -10, 7, 2, -9, 22, -2, 11, -3,
    -- filter=22 channel=0
    -8, 1, -19, -12, 7, 4, 2, -10, 10,
    -- filter=22 channel=1
    6, 7, -2, -12, 24, -6, 13, -12, -12,
    -- filter=22 channel=2
    -14, -18, -8, -13, 17, -11, 14, -8, -19,
    -- filter=22 channel=3
    0, 2, -10, 26, 17, 19, -13, 13, 5,
    -- filter=22 channel=4
    -16, 16, -18, -15, 2, -2, 8, -10, 6,
    -- filter=22 channel=5
    16, -4, -10, -2, -8, -6, -3, 4, -16,
    -- filter=22 channel=6
    1, -15, 0, 11, 8, 10, -3, 15, 6,
    -- filter=22 channel=7
    -15, -2, -1, -1, 5, 0, 6, 9, 19,
    -- filter=22 channel=8
    -12, -15, 20, -18, 16, 6, 3, -16, -4,
    -- filter=22 channel=9
    -18, -23, -10, -1, 9, -8, 7, -25, -19,
    -- filter=22 channel=10
    0, 26, 17, 8, 4, -8, 2, -16, -20,
    -- filter=22 channel=11
    -18, 20, -17, 18, -15, 15, 21, 0, -15,
    -- filter=22 channel=12
    15, 0, -15, -20, 11, -18, -6, -12, -17,
    -- filter=22 channel=13
    26, 10, -9, -5, 20, 3, 24, -6, -3,
    -- filter=22 channel=14
    -7, 28, 14, 16, 12, -2, 20, -2, -3,
    -- filter=22 channel=15
    -12, -3, 0, 9, -14, 8, -16, 5, -19,
    -- filter=23 channel=0
    -33, -15, -12, -28, -39, -8, -1, -6, -13,
    -- filter=23 channel=1
    49, 27, 36, 20, 7, 35, -11, 9, 22,
    -- filter=23 channel=2
    -45, -37, -11, -47, -22, -28, -26, -24, -27,
    -- filter=23 channel=3
    -2, 17, 26, 30, 24, 6, 44, 34, 32,
    -- filter=23 channel=4
    0, -31, -14, -31, -10, -32, -8, -35, -35,
    -- filter=23 channel=5
    40, 46, 52, 11, 26, 20, 8, 35, 22,
    -- filter=23 channel=6
    0, 8, 14, -15, -8, 13, -16, -17, 19,
    -- filter=23 channel=7
    -20, -25, -43, -28, -45, -45, -8, -19, -12,
    -- filter=23 channel=8
    8, 16, -5, -7, 2, -2, -17, 18, -14,
    -- filter=23 channel=9
    -37, -48, -18, -13, -36, -46, -36, -47, -19,
    -- filter=23 channel=10
    20, 17, 43, 6, 21, 42, 19, -4, 16,
    -- filter=23 channel=11
    -2, -14, -25, -14, -7, 2, 10, 11, -10,
    -- filter=23 channel=12
    -3, -15, -10, -11, 7, -11, 17, -19, -16,
    -- filter=23 channel=13
    46, 39, 42, 6, 39, 34, -11, -8, 28,
    -- filter=23 channel=14
    40, 12, 45, 43, 31, 23, 3, 11, 44,
    -- filter=23 channel=15
    -14, -14, -9, -12, -12, -37, -40, -16, -35,
    -- filter=24 channel=0
    -19, -7, -27, -1, -15, -17, -34, -33, 6,
    -- filter=24 channel=1
    -12, 4, 13, 12, 28, 15, 22, 29, 29,
    -- filter=24 channel=2
    6, 5, -12, 18, 5, -2, 19, -19, -12,
    -- filter=24 channel=3
    -3, -29, -35, -18, -2, -34, -16, -20, -16,
    -- filter=24 channel=4
    17, 13, 1, 9, 26, 17, 28, 43, 4,
    -- filter=24 channel=5
    -23, -11, -31, -5, -21, 7, -18, -7, -23,
    -- filter=24 channel=6
    -10, 6, 6, -9, -13, -11, -21, -25, 0,
    -- filter=24 channel=7
    -1, -14, -22, 26, 9, -15, -4, -15, 13,
    -- filter=24 channel=8
    11, -7, 6, 18, 17, -4, 0, 10, 3,
    -- filter=24 channel=9
    17, 41, 27, 47, 18, 20, 40, 11, 39,
    -- filter=24 channel=10
    10, 14, -13, 25, 12, 10, -5, 21, 19,
    -- filter=24 channel=11
    -8, 11, -15, 6, -7, -6, 8, -20, -24,
    -- filter=24 channel=12
    -2, 4, 15, 13, 12, -13, 14, -11, 10,
    -- filter=24 channel=13
    29, 27, 11, 46, 41, 20, 15, 52, 18,
    -- filter=24 channel=14
    -9, -27, -19, -2, 0, -20, -27, 10, 15,
    -- filter=24 channel=15
    12, 1, 5, 12, -6, 23, 3, -3, 5,
    -- filter=25 channel=0
    20, -2, 10, 12, -4, -11, 13, 18, -19,
    -- filter=25 channel=1
    11, 16, 12, 0, 9, 7, 11, 11, -12,
    -- filter=25 channel=2
    -19, 2, -5, 6, -19, -3, 11, -19, 14,
    -- filter=25 channel=3
    -15, -11, 3, 5, 10, 19, -11, -13, 11,
    -- filter=25 channel=4
    11, 14, 13, -8, 11, -16, -19, -3, -7,
    -- filter=25 channel=5
    17, 12, -13, -20, -15, 16, -3, -16, 7,
    -- filter=25 channel=6
    8, -10, -8, -13, 11, -11, 19, 17, 20,
    -- filter=25 channel=7
    5, 13, 7, -3, -14, -18, 4, 0, -9,
    -- filter=25 channel=8
    20, -12, -18, 1, 3, -17, -20, -16, -17,
    -- filter=25 channel=9
    2, -5, -20, -20, 5, -2, -10, 19, -11,
    -- filter=25 channel=10
    -4, -20, -15, 9, -2, 18, -10, -12, -3,
    -- filter=25 channel=11
    -6, -17, -1, 0, 3, 3, 13, 3, -5,
    -- filter=25 channel=12
    2, 13, -17, 19, 9, 9, -20, 19, -15,
    -- filter=25 channel=13
    -8, 2, -4, -13, -10, -1, 5, -4, -21,
    -- filter=25 channel=14
    -9, -9, -17, -4, -7, 9, -6, 15, -11,
    -- filter=25 channel=15
    18, 14, 6, -4, -12, -4, -15, -4, 10,
    -- filter=26 channel=0
    -8, -21, 19, 7, 18, 6, 9, 13, -14,
    -- filter=26 channel=1
    -12, 16, 10, 7, 21, -27, 3, 2, -10,
    -- filter=26 channel=2
    10, 1, -2, 27, 10, -7, 17, 12, 12,
    -- filter=26 channel=3
    -37, 3, -30, -28, -21, -3, 4, -12, 5,
    -- filter=26 channel=4
    38, 37, 33, 43, 18, 8, 34, 33, 27,
    -- filter=26 channel=5
    8, -19, 0, -5, -9, -10, 10, -24, -6,
    -- filter=26 channel=6
    -1, -17, 9, 5, 20, -2, 12, -5, -2,
    -- filter=26 channel=7
    -6, 7, -2, 12, 24, 22, 2, 4, -10,
    -- filter=26 channel=8
    11, 12, 2, 8, -16, 2, -11, 16, 15,
    -- filter=26 channel=9
    31, 39, 18, 41, 22, -5, 39, 33, -3,
    -- filter=26 channel=10
    -5, -2, 15, 7, 11, -6, 0, 18, -24,
    -- filter=26 channel=11
    15, 1, 14, 8, -5, -14, 19, -14, 13,
    -- filter=26 channel=12
    -10, -7, -12, -3, -11, 16, 14, -12, 3,
    -- filter=26 channel=13
    18, 11, 23, 37, 28, -13, 44, 6, -4,
    -- filter=26 channel=14
    -19, -8, -26, -29, 5, -18, -8, -7, -18,
    -- filter=26 channel=15
    -1, 7, -2, 0, 31, 26, 15, -1, 12,
    -- filter=27 channel=0
    1, 0, -8, 21, -2, 15, 7, 5, 20,
    -- filter=27 channel=1
    -2, 2, 18, 9, 12, 21, -15, 0, 14,
    -- filter=27 channel=2
    12, -17, -5, 12, 19, -5, 19, 10, 21,
    -- filter=27 channel=3
    -3, -7, -8, -5, 8, -18, 19, 18, -5,
    -- filter=27 channel=4
    2, 0, -9, 15, -11, 20, -3, -7, -4,
    -- filter=27 channel=5
    8, -9, -4, 0, 10, 13, 20, -10, 3,
    -- filter=27 channel=6
    -16, 0, -5, -11, 14, -3, 13, -15, -18,
    -- filter=27 channel=7
    -3, -13, -16, -4, 18, -15, -10, -3, 16,
    -- filter=27 channel=8
    10, 12, 15, 3, -15, 10, 16, 11, -10,
    -- filter=27 channel=9
    -14, -2, 15, -15, 0, -10, -14, 8, -11,
    -- filter=27 channel=10
    6, 2, 12, 11, -13, 19, 9, -5, 15,
    -- filter=27 channel=11
    -16, 18, -3, 13, 8, 2, -14, -2, -7,
    -- filter=27 channel=12
    -14, -9, 19, 2, -11, -19, -10, 4, 0,
    -- filter=27 channel=13
    -3, 10, 8, -3, -17, -18, -11, -20, -6,
    -- filter=27 channel=14
    5, 16, 14, -14, -19, 14, -11, -15, 10,
    -- filter=27 channel=15
    -20, -2, -4, 4, 7, 21, 8, 20, -8,
    -- filter=28 channel=0
    -17, 20, 21, -11, -5, -16, 0, 9, 20,
    -- filter=28 channel=1
    -13, 21, -3, 4, 8, 15, 24, 12, -22,
    -- filter=28 channel=2
    -12, -19, 5, -2, -19, -3, -6, 6, -17,
    -- filter=28 channel=3
    -21, 16, 19, 1, 6, 5, 20, 2, 8,
    -- filter=28 channel=4
    0, 5, -8, -3, -3, 7, 15, -4, 9,
    -- filter=28 channel=5
    22, -16, -8, -3, 0, -20, 0, 14, -20,
    -- filter=28 channel=6
    -3, -8, -15, -5, -5, -16, 19, 5, 17,
    -- filter=28 channel=7
    -13, -9, -3, 13, -12, -11, 8, 22, 7,
    -- filter=28 channel=8
    -13, -12, -16, -9, 16, -9, -16, 10, -6,
    -- filter=28 channel=9
    -16, -8, 11, 12, -5, -19, 0, 21, 0,
    -- filter=28 channel=10
    12, -6, 10, 9, -9, -4, 14, 10, -14,
    -- filter=28 channel=11
    8, 6, -11, 0, 20, 0, -4, -15, 8,
    -- filter=28 channel=12
    -7, 10, 19, -6, 17, -3, 7, -12, -15,
    -- filter=28 channel=13
    -3, -3, -20, 29, -2, -34, 7, 15, -21,
    -- filter=28 channel=14
    18, -14, -14, -2, 13, 11, -15, -13, -5,
    -- filter=28 channel=15
    -6, -4, 24, -15, -8, -3, -8, 7, 4,
    -- filter=29 channel=0
    21, -12, -10, -17, 9, -11, -20, -2, -12,
    -- filter=29 channel=1
    -11, -15, -18, 3, -17, -6, -5, -10, -4,
    -- filter=29 channel=2
    19, -10, -16, 8, 2, 8, -21, 20, -11,
    -- filter=29 channel=3
    -17, 12, -2, 20, 2, 1, 11, -11, -4,
    -- filter=29 channel=4
    -16, 19, 5, -10, 9, 6, -15, 13, -20,
    -- filter=29 channel=5
    8, 15, 0, 4, -18, 8, 5, 11, -2,
    -- filter=29 channel=6
    -7, 20, -7, 9, -9, 0, 18, 6, 16,
    -- filter=29 channel=7
    2, -5, 4, 19, 4, 17, -21, 10, 9,
    -- filter=29 channel=8
    -7, 1, 3, 0, -3, 15, -14, -4, -17,
    -- filter=29 channel=9
    4, -6, 15, -20, -7, -7, -21, 6, -16,
    -- filter=29 channel=10
    -20, -16, 9, -15, -4, -13, -6, 13, -12,
    -- filter=29 channel=11
    13, -3, -8, -18, 5, -13, 6, -2, -21,
    -- filter=29 channel=12
    19, 6, -1, -5, -3, -2, -15, -17, -10,
    -- filter=29 channel=13
    2, 3, -9, 7, -10, 4, 16, 13, -9,
    -- filter=29 channel=14
    5, -2, 0, 12, -12, -8, -1, 0, -2,
    -- filter=29 channel=15
    -2, 15, -12, -20, 19, -19, 3, 10, -7,
    -- filter=30 channel=0
    -7, 5, 25, 13, 29, 5, -10, 9, 0,
    -- filter=30 channel=1
    2, 6, -21, 6, -27, 4, 2, 3, -12,
    -- filter=30 channel=2
    18, 5, 10, 1, 21, -6, -7, 2, -4,
    -- filter=30 channel=3
    -1, -18, 8, 9, 2, -8, 8, -17, -2,
    -- filter=30 channel=4
    4, -11, -3, 20, 4, -17, 12, -3, 3,
    -- filter=30 channel=5
    13, -26, -19, 3, -26, -7, -13, 5, 12,
    -- filter=30 channel=6
    25, -2, 6, 5, 16, -15, 10, -3, -3,
    -- filter=30 channel=7
    -13, 11, 3, -17, -8, 0, -1, 23, 25,
    -- filter=30 channel=8
    16, -19, 15, -17, 1, -19, 18, -10, 12,
    -- filter=30 channel=9
    -7, 9, 6, 11, 7, 18, -9, 15, 1,
    -- filter=30 channel=10
    21, 3, 20, 19, -11, 17, 6, 18, -6,
    -- filter=30 channel=11
    8, -8, 8, 1, 17, 6, -5, 10, 0,
    -- filter=30 channel=12
    -13, -20, 10, -5, 7, 13, -3, -8, 17,
    -- filter=30 channel=13
    20, -10, 3, -5, -29, -8, 22, -23, 11,
    -- filter=30 channel=14
    9, 8, 5, 5, -16, 9, -2, -15, -13,
    -- filter=30 channel=15
    -6, -11, 14, 25, -11, 9, 18, 19, 0,
    -- filter=31 channel=0
    10, 12, -17, -6, -14, 5, -9, -16, 20,
    -- filter=31 channel=1
    2, -14, 18, -17, 0, -12, -1, 2, 16,
    -- filter=31 channel=2
    3, -5, 19, 12, -15, 7, 8, 8, 1,
    -- filter=31 channel=3
    15, -6, -13, -16, -18, -17, -9, -12, 22,
    -- filter=31 channel=4
    16, -19, 9, -11, -8, 10, 3, 8, 0,
    -- filter=31 channel=5
    -3, -9, 12, -14, -9, -13, 12, -4, -17,
    -- filter=31 channel=6
    -10, 11, 0, -10, 17, -7, 11, -10, -10,
    -- filter=31 channel=7
    0, -7, 20, 19, -1, -7, 16, -18, 16,
    -- filter=31 channel=8
    -19, 0, -10, 18, 15, 5, -11, 0, -9,
    -- filter=31 channel=9
    6, 19, -15, 1, 3, -14, -7, -11, 6,
    -- filter=31 channel=10
    12, -12, 16, 0, 15, 11, -3, -1, 10,
    -- filter=31 channel=11
    18, 20, -11, -12, 12, -6, -16, -8, 11,
    -- filter=31 channel=12
    7, 10, 18, -9, -12, -20, 3, 15, 0,
    -- filter=31 channel=13
    -18, -7, -19, -15, 14, -4, 24, -6, 3,
    -- filter=31 channel=14
    6, 2, 7, 17, 3, -9, 4, 18, 16,
    -- filter=31 channel=15
    12, -11, 0, 13, 15, -6, -19, -1, -5,

    -- ifmap
    -- channel=0
    146, 126, 125, 126, 125, 123, 125, 127, 129, 125, 123, 122, 128, 124, 126, 213, 
    119, 117, 112, 113, 116, 120, 112, 122, 120, 104, 104, 92, 97, 117, 123, 218, 
    108, 111, 123, 121, 114, 91, 144, 104, 131, 82, 74, 86, 94, 87, 120, 222, 
    138, 91, 118, 119, 118, 103, 129, 125, 90, 31, 98, 65, 109, 111, 103, 225, 
    128, 57, 106, 110, 137, 94, 72, 105, 87, 77, 107, 105, 104, 122, 103, 231, 
    74, 38, 120, 135, 27, 92, 105, 98, 128, 56, 40, 96, 78, 108, 130, 202, 
    97, 58, 112, 157, 26, 78, 97, 95, 143, 0, 82, 103, 74, 85, 98, 197, 
    93, 101, 125, 159, 68, 25, 56, 70, 109, 0, 82, 92, 70, 48, 107, 218, 
    45, 43, 133, 107, 132, 40, 102, 84, 94, 75, 91, 105, 87, 99, 104, 231, 
    24, 0, 108, 25, 99, 132, 82, 96, 90, 124, 111, 130, 89, 85, 105, 237, 
    33, 13, 97, 13, 106, 110, 43, 57, 118, 99, 128, 114, 41, 66, 95, 216, 
    0, 19, 102, 0, 46, 69, 26, 32, 66, 94, 57, 22, 29, 17, 33, 166, 
    11, 0, 34, 0, 81, 95, 41, 37, 37, 36, 25, 23, 12, 15, 16, 172, 
    27, 22, 0, 102, 102, 25, 40, 35, 36, 27, 15, 7, 23, 11, 0, 191, 
    18, 16, 18, 107, 82, 27, 36, 35, 28, 20, 17, 22, 24, 0, 55, 174, 
    36, 14, 31, 35, 59, 37, 36, 32, 15, 19, 29, 29, 0, 27, 51, 149, 
    
    -- channel=1
    156, 159, 161, 165, 163, 161, 166, 168, 166, 155, 130, 120, 130, 133, 127, 116, 
    159, 164, 164, 171, 168, 214, 238, 171, 167, 138, 127, 113, 107, 126, 132, 125, 
    155, 156, 168, 168, 168, 199, 193, 122, 79, 122, 161, 136, 114, 86, 126, 132, 
    130, 106, 176, 172, 180, 163, 171, 144, 84, 136, 170, 144, 107, 64, 93, 122, 
    215, 203, 221, 197, 293, 276, 197, 165, 98, 98, 211, 180, 102, 94, 53, 84, 
    233, 241, 256, 167, 243, 279, 241, 219, 134, 138, 240, 181, 102, 102, 73, 48, 
    250, 237, 246, 163, 143, 231, 273, 261, 168, 152, 241, 167, 105, 121, 118, 97, 
    278, 249, 222, 171, 151, 260, 298, 228, 155, 158, 215, 171, 107, 125, 125, 127, 
    297, 273, 244, 174, 189, 177, 194, 160, 147, 149, 153, 154, 60, 106, 149, 147, 
    295, 284, 260, 182, 206, 148, 160, 223, 195, 163, 141, 77, 68, 140, 163, 158, 
    254, 296, 255, 246, 341, 270, 239, 264, 242, 120, 65, 71, 91, 148, 153, 140, 
    192, 270, 262, 327, 374, 281, 133, 142, 127, 101, 78, 81, 97, 110, 108, 99, 
    111, 186, 258, 350, 335, 147, 86, 76, 75, 78, 88, 107, 113, 114, 134, 152, 
    107, 92, 214, 310, 259, 97, 97, 86, 77, 85, 93, 100, 102, 118, 147, 136, 
    115, 92, 103, 164, 152, 78, 99, 94, 95, 111, 112, 87, 135, 160, 139, 94, 
    113, 95, 84, 84, 75, 49, 58, 63, 84, 120, 116, 95, 147, 168, 126, 65, 
    
    -- channel=2
    66, 32, 30, 26, 26, 31, 23, 29, 33, 31, 26, 32, 29, 20, 23, 21, 
    69, 34, 33, 27, 34, 71, 16, 35, 36, 46, 23, 25, 32, 30, 27, 20, 
    79, 49, 34, 28, 36, 80, 0, 21, 31, 62, 2, 0, 0, 35, 45, 14, 
    79, 65, 32, 37, 39, 47, 42, 7, 10, 49, 0, 0, 0, 12, 55, 22, 
    70, 27, 0, 91, 97, 16, 22, 0, 0, 85, 43, 0, 2, 0, 56, 54, 
    66, 36, 0, 88, 123, 0, 21, 0, 0, 122, 16, 0, 5, 0, 11, 45, 
    36, 50, 0, 12, 108, 36, 38, 0, 0, 108, 0, 0, 10, 8, 0, 0, 
    63, 33, 0, 25, 54, 97, 0, 0, 0, 61, 0, 0, 15, 13, 0, 7, 
    96, 0, 0, 19, 36, 67, 0, 4, 10, 18, 26, 0, 24, 16, 10, 13, 
    128, 0, 0, 28, 0, 31, 36, 42, 14, 0, 3, 10, 44, 30, 14, 22, 
    180, 0, 0, 83, 0, 2, 30, 16, 0, 0, 1, 19, 27, 25, 20, 25, 
    175, 0, 0, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    100, 7, 42, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    82, 0, 72, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    82, 0, 23, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    83, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=3
    163, 154, 140, 144, 146, 144, 151, 160, 158, 149, 143, 142, 137, 132, 139, 132, 
    165, 154, 145, 146, 147, 126, 154, 155, 152, 143, 134, 149, 150, 158, 138, 132, 
    156, 179, 158, 156, 159, 201, 188, 159, 150, 112, 53, 62, 77, 153, 153, 130, 
    125, 197, 178, 155, 147, 156, 133, 58, 63, 120, 92, 96, 95, 93, 150, 137, 
    74, 33, 138, 152, 77, 63, 50, 67, 86, 119, 123, 70, 91, 59, 150, 167, 
    84, 74, 126, 138, 166, 113, 58, 60, 72, 77, 47, 83, 85, 76, 67, 135, 
    78, 67, 166, 153, 129, 125, 88, 57, 63, 72, 81, 83, 89, 96, 56, 80, 
    68, 49, 120, 147, 104, 95, 106, 111, 107, 97, 106, 83, 89, 85, 106, 109, 
    72, 49, 34, 96, 99, 155, 178, 110, 99, 130, 157, 128, 115, 114, 111, 121, 
    123, 58, 50, 89, 79, 109, 104, 44, 93, 135, 104, 130, 77, 100, 137, 138, 
    133, 61, 58, 53, 0, 62, 30, 64, 46, 149, 148, 74, 66, 121, 127, 129, 
    132, 137, 46, 21, 118, 130, 140, 164, 135, 88, 38, 32, 30, 47, 45, 31, 
    80, 137, 125, 67, 119, 90, 27, 34, 36, 39, 35, 27, 19, 28, 13, 0, 
    24, 61, 105, 148, 77, 31, 29, 35, 30, 19, 21, 42, 38, 48, 40, 73, 
    14, 16, 72, 171, 102, 67, 63, 41, 21, 20, 22, 36, 32, 0, 47, 63, 
    108, 90, 100, 101, 98, 93, 96, 117, 129, 125, 113, 98, 128, 139, 105, 90, 
    
    -- channel=4
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 22, 68, 0, 0, 10, 52, 48, 15, 0, 0, 0, 
    0, 0, 0, 0, 0, 18, 80, 16, 9, 34, 104, 94, 62, 22, 0, 0, 
    92, 47, 0, 0, 0, 7, 64, 82, 34, 35, 116, 87, 61, 37, 0, 2, 
    180, 98, 111, 0, 159, 198, 143, 124, 48, 29, 121, 121, 44, 46, 13, 0, 
    187, 156, 169, 0, 160, 243, 169, 154, 74, 33, 176, 138, 47, 51, 50, 0, 
    197, 177, 180, 4, 35, 149, 173, 197, 102, 53, 192, 133, 55, 49, 66, 25, 
    214, 205, 210, 54, 27, 107, 204, 173, 104, 49, 165, 123, 56, 54, 69, 6, 
    244, 204, 231, 90, 116, 92, 155, 84, 80, 52, 74, 108, 30, 42, 36, 8, 
    233, 209, 223, 134, 148, 107, 71, 145, 168, 80, 53, 54, 5, 4, 7, 15, 
    164, 225, 204, 141, 284, 215, 120, 190, 212, 98, 45, 54, 77, 81, 93, 103, 
    129, 215, 213, 156, 300, 277, 128, 152, 158, 113, 97, 106, 123, 128, 132, 156, 
    145, 139, 182, 243, 301, 195, 111, 106, 95, 95, 110, 125, 136, 137, 153, 201, 
    163, 140, 115, 273, 289, 114, 123, 110, 102, 114, 124, 133, 141, 134, 167, 197, 
    169, 142, 136, 187, 194, 98, 121, 120, 112, 132, 137, 123, 131, 190, 196, 137, 
    172, 141, 131, 110, 99, 72, 83, 91, 98, 133, 144, 119, 131, 204, 194, 119, 
    
    -- channel=5
    165, 165, 167, 165, 165, 160, 170, 173, 167, 154, 143, 141, 143, 139, 136, 123, 
    165, 167, 167, 173, 172, 189, 159, 166, 157, 142, 122, 108, 123, 143, 141, 130, 
    149, 170, 176, 170, 177, 229, 195, 139, 126, 140, 137, 116, 95, 117, 139, 133, 
    123, 129, 170, 173, 167, 174, 143, 98, 99, 152, 165, 116, 105, 80, 125, 136, 
    147, 165, 168, 184, 223, 185, 175, 115, 93, 157, 158, 120, 98, 72, 92, 128, 
    163, 201, 176, 198, 268, 199, 204, 140, 101, 183, 191, 131, 103, 102, 56, 87, 
    159, 198, 182, 166, 180, 202, 232, 183, 138, 208, 201, 123, 105, 105, 99, 86, 
    187, 206, 131, 159, 149, 231, 239, 168, 145, 199, 190, 138, 100, 132, 124, 126, 
    208, 209, 144, 156, 160, 236, 183, 144, 121, 158, 180, 122, 104, 127, 145, 153, 
    232, 219, 185, 156, 156, 142, 158, 176, 131, 141, 131, 78, 77, 161, 164, 157, 
    229, 219, 193, 223, 197, 158, 208, 225, 154, 115, 76, 61, 88, 139, 141, 124, 
    203, 229, 196, 307, 303, 198, 181, 181, 133, 77, 82, 88, 90, 99, 98, 87, 
    128, 181, 231, 298, 250, 107, 78, 77, 77, 78, 83, 90, 103, 103, 109, 109, 
    83, 115, 213, 303, 144, 95, 87, 75, 78, 85, 96, 107, 106, 106, 122, 132, 
    92, 80, 160, 199, 137, 98, 95, 92, 92, 98, 86, 90, 113, 131, 115, 80, 
    93, 94, 85, 89, 70, 73, 79, 83, 106, 115, 107, 103, 151, 154, 99, 64, 
    
    -- channel=6
    58, 60, 56, 58, 60, 56, 57, 60, 62, 55, 53, 51, 56, 55, 59, 110, 
    57, 60, 56, 60, 58, 82, 68, 60, 63, 47, 43, 40, 36, 53, 60, 115, 
    57, 54, 62, 62, 60, 60, 73, 52, 49, 29, 34, 40, 41, 35, 59, 115, 
    67, 24, 61, 60, 71, 53, 61, 59, 39, 6, 50, 29, 42, 39, 34, 118, 
    65, 32, 60, 59, 86, 80, 42, 50, 38, 17, 43, 55, 35, 47, 44, 122, 
    53, 19, 63, 72, 30, 55, 65, 45, 64, 0, 40, 53, 28, 38, 49, 83, 
    57, 45, 46, 87, 5, 24, 57, 58, 67, 0, 40, 44, 24, 30, 38, 100, 
    49, 47, 70, 82, 52, 24, 50, 30, 45, 1, 42, 39, 23, 21, 41, 112, 
    28, 17, 75, 53, 69, 12, 39, 47, 27, 48, 30, 54, 23, 34, 47, 128, 
    21, 3, 58, 0, 51, 60, 35, 64, 58, 50, 51, 39, 33, 32, 45, 122, 
    23, 14, 49, 0, 74, 54, 4, 33, 59, 40, 25, 32, 11, 16, 34, 110, 
    0, 10, 40, 0, 41, 43, 0, 0, 8, 22, 18, 3, 1, 0, 9, 70, 
    1, 0, 17, 31, 41, 23, 6, 4, 3, 0, 0, 0, 0, 0, 0, 82, 
    0, 0, 0, 63, 36, 3, 5, 1, 1, 0, 0, 0, 0, 0, 0, 70, 
    0, 0, 0, 29, 23, 0, 3, 8, 0, 0, 1, 0, 0, 0, 3, 58, 
    5, 2, 1, 8, 13, 8, 9, 6, 0, 1, 6, 5, 0, 6, 12, 43, 
    
    -- channel=7
    142, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    138, 0, 0, 0, 0, 1, 0, 0, 0, 23, 13, 6, 12, 10, 0, 0, 
    141, 15, 0, 0, 0, 16, 0, 0, 20, 81, 30, 17, 18, 22, 45, 0, 
    177, 75, 28, 0, 0, 0, 23, 0, 37, 93, 62, 23, 22, 19, 65, 18, 
    233, 86, 0, 0, 77, 0, 28, 0, 28, 89, 103, 0, 35, 14, 51, 66, 
    247, 102, 0, 0, 110, 0, 51, 0, 7, 159, 98, 0, 46, 28, 16, 50, 
    252, 117, 0, 0, 115, 41, 62, 0, 4, 165, 53, 0, 37, 47, 25, 18, 
    268, 104, 0, 53, 64, 93, 0, 12, 6, 129, 37, 0, 52, 49, 18, 5, 
    297, 54, 0, 72, 0, 83, 38, 25, 44, 39, 42, 0, 58, 61, 7, 0, 
    297, 37, 8, 99, 28, 0, 84, 72, 32, 63, 2, 39, 76, 37, 0, 0, 
    261, 16, 10, 146, 81, 12, 66, 67, 0, 6, 56, 66, 74, 78, 41, 46, 
    227, 95, 27, 144, 46, 9, 75, 73, 72, 75, 84, 89, 95, 87, 81, 84, 
    214, 121, 103, 131, 0, 76, 75, 78, 78, 86, 95, 95, 97, 88, 104, 98, 
    221, 100, 135, 178, 34, 82, 85, 81, 85, 89, 91, 98, 89, 115, 117, 84, 
    228, 102, 106, 139, 64, 97, 93, 84, 87, 89, 87, 95, 120, 110, 84, 71, 
    228, 98, 90, 79, 77, 97, 91, 87, 98, 94, 68, 88, 118, 99, 68, 89, 
    
    -- channel=8
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    
    -- channel=9
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 68, 62, 33, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 12, 29, 40, 42, 34, 31, 25, 0, 0, 
    96, 83, 0, 0, 0, 0, 16, 18, 30, 14, 30, 19, 23, 30, 0, 0, 
    125, 133, 0, 0, 28, 36, 15, 16, 25, 34, 57, 40, 32, 42, 37, 0, 
    125, 131, 0, 0, 0, 2, 49, 37, 40, 64, 76, 46, 40, 48, 47, 0, 
    115, 132, 77, 0, 0, 52, 77, 50, 27, 55, 68, 47, 44, 40, 16, 0, 
    152, 161, 141, 82, 0, 37, 48, 20, 38, 0, 7, 23, 30, 23, 0, 0, 
    145, 164, 152, 111, 92, 25, 21, 76, 64, 7, 18, 34, 43, 0, 0, 0, 
    145, 134, 122, 133, 168, 129, 144, 157, 144, 86, 140, 175, 195, 168, 140, 149, 
    291, 239, 157, 133, 191, 218, 228, 232, 245, 257, 285, 302, 321, 326, 324, 332, 
    363, 311, 214, 160, 228, 275, 277, 269, 274, 295, 325, 339, 340, 346, 371, 372, 
    394, 371, 287, 237, 245, 288, 288, 279, 289, 315, 344, 358, 361, 394, 403, 374, 
    395, 384, 348, 273, 265, 286, 293, 288, 295, 319, 341, 349, 365, 406, 410, 343, 
    368, 356, 345, 288, 272, 279, 284, 279, 286, 313, 316, 313, 340, 377, 377, 329, 
    
    -- channel=10
    148, 102, 96, 98, 92, 96, 97, 91, 86, 81, 70, 77, 82, 78, 68, 53, 
    147, 99, 100, 101, 106, 184, 111, 96, 90, 102, 109, 91, 73, 81, 81, 62, 
    145, 100, 105, 98, 103, 171, 93, 57, 67, 184, 168, 126, 100, 77, 96, 71, 
    171, 139, 133, 104, 115, 123, 157, 82, 93, 206, 184, 120, 103, 40, 103, 93, 
    235, 228, 144, 185, 282, 204, 207, 110, 90, 183, 220, 119, 100, 74, 77, 100, 
    248, 276, 158, 149, 295, 211, 261, 139, 113, 282, 257, 128, 115, 99, 53, 64, 
    231, 302, 138, 121, 225, 253, 300, 172, 144, 306, 249, 121, 107, 136, 111, 70, 
    280, 305, 135, 163, 170, 329, 276, 170, 136, 269, 223, 131, 118, 147, 110, 95, 
    346, 297, 180, 200, 148, 235, 166, 150, 152, 163, 161, 98, 95, 117, 113, 103, 
    358, 296, 237, 245, 185, 119, 193, 254, 158, 160, 112, 42, 100, 141, 122, 94, 
    333, 283, 239, 375, 359, 186, 260, 304, 152, 110, 85, 113, 141, 158, 134, 124, 
    308, 293, 253, 436, 411, 167, 197, 188, 144, 123, 136, 151, 165, 172, 162, 162, 
    198, 273, 322, 426, 256, 142, 138, 130, 129, 138, 160, 175, 178, 178, 212, 218, 
    177, 180, 341, 425, 130, 158, 152, 135, 139, 153, 164, 181, 174, 203, 216, 207, 
    186, 159, 220, 277, 120, 152, 158, 144, 165, 177, 161, 159, 233, 249, 194, 139, 
    189, 155, 153, 142, 106, 121, 126, 125, 166, 183, 162, 164, 252, 249, 146, 121, 
    
    -- channel=11
    42, 44, 42, 41, 42, 45, 40, 43, 44, 44, 46, 46, 45, 45, 48, 87, 
    20, 25, 23, 25, 23, 9, 18, 36, 59, 39, 32, 39, 42, 39, 32, 89, 
    53, 47, 27, 25, 22, 55, 57, 61, 54, 17, 29, 36, 45, 39, 33, 89, 
    62, 23, 22, 22, 27, 28, 32, 43, 38, 14, 38, 34, 53, 56, 30, 89, 
    45, 0, 27, 24, 16, 28, 30, 44, 49, 35, 36, 36, 41, 54, 49, 100, 
    39, 14, 38, 30, 31, 43, 26, 40, 58, 11, 22, 52, 33, 43, 53, 87, 
    46, 37, 46, 49, 23, 19, 38, 45, 64, 0, 34, 48, 35, 33, 38, 76, 
    35, 41, 51, 43, 23, 12, 63, 35, 49, 0, 33, 53, 37, 32, 45, 86, 
    6, 8, 62, 22, 34, 26, 54, 31, 30, 35, 45, 70, 46, 34, 24, 92, 
    8, 0, 48, 18, 38, 72, 34, 27, 35, 55, 75, 60, 40, 15, 31, 100, 
    9, 1, 58, 4, 14, 7, 11, 43, 70, 54, 52, 35, 24, 26, 39, 109, 
    15, 24, 26, 0, 57, 80, 40, 47, 60, 45, 38, 29, 31, 23, 29, 105, 
    43, 7, 32, 10, 71, 60, 34, 33, 35, 32, 27, 24, 29, 32, 24, 120, 
    43, 30, 9, 77, 61, 31, 32, 33, 34, 30, 29, 30, 34, 27, 47, 129, 
    44, 30, 28, 89, 60, 42, 41, 43, 27, 24, 31, 31, 23, 18, 50, 110, 
    93, 82, 82, 82, 83, 76, 76, 70, 72, 89, 95, 86, 79, 110, 102, 110, 
    
    -- channel=12
    26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 
    28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 8, 0, 
    1, 20, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 24, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    
    -- channel=13
    204, 214, 215, 213, 208, 217, 219, 205, 193, 188, 176, 167, 178, 175, 154, 132, 
    190, 206, 215, 218, 221, 324, 333, 208, 199, 193, 228, 209, 159, 163, 159, 149, 
    191, 201, 211, 214, 215, 348, 342, 178, 136, 303, 365, 322, 243, 137, 166, 171, 
    220, 178, 223, 215, 237, 230, 304, 267, 198, 332, 389, 314, 256, 137, 149, 172, 
    436, 415, 379, 314, 545, 510, 435, 341, 218, 262, 423, 347, 227, 193, 92, 132, 
    510, 534, 464, 292, 611, 608, 508, 431, 274, 335, 516, 384, 232, 230, 160, 91, 
    526, 527, 464, 232, 382, 478, 576, 518, 357, 415, 529, 358, 230, 263, 260, 173, 
    589, 572, 439, 274, 289, 559, 629, 486, 357, 414, 504, 367, 231, 289, 277, 189, 
    665, 643, 539, 380, 354, 497, 480, 336, 298, 301, 359, 319, 182, 241, 232, 223, 
    671, 655, 593, 423, 433, 289, 359, 464, 401, 298, 263, 186, 153, 234, 251, 224, 
    593, 651, 583, 571, 714, 540, 502, 579, 483, 270, 171, 199, 266, 309, 299, 270, 
    539, 630, 595, 775, 852, 624, 444, 458, 400, 269, 285, 310, 343, 364, 358, 348, 
    396, 513, 604, 805, 771, 394, 303, 287, 275, 283, 321, 357, 377, 377, 424, 444, 
    376, 343, 552, 743, 586, 329, 326, 298, 293, 322, 348, 373, 379, 394, 449, 460, 
    388, 354, 392, 495, 408, 308, 331, 318, 334, 369, 362, 339, 424, 495, 449, 331, 
    386, 352, 335, 305, 258, 237, 261, 269, 328, 385, 379, 332, 464, 518, 426, 275, 
    
    -- channel=14
    174, 174, 173, 175, 182, 174, 176, 192, 190, 168, 137, 133, 140, 149, 152, 144, 
    179, 181, 176, 181, 180, 190, 179, 188, 175, 144, 134, 113, 120, 146, 152, 147, 
    156, 167, 183, 187, 189, 202, 164, 138, 125, 94, 69, 60, 67, 114, 141, 148, 
    103, 154, 175, 190, 182, 170, 152, 81, 56, 78, 81, 78, 67, 69, 113, 131, 
    70, 82, 169, 192, 197, 163, 93, 73, 61, 113, 101, 84, 72, 44, 92, 108, 
    90, 99, 165, 161, 186, 108, 111, 94, 68, 92, 96, 76, 65, 60, 53, 89, 
    98, 94, 145, 152, 147, 148, 131, 97, 80, 92, 103, 85, 74, 76, 55, 69, 
    94, 88, 128, 142, 143, 136, 134, 109, 88, 113, 106, 98, 67, 65, 109, 117, 
    90, 88, 77, 107, 140, 128, 127, 113, 90, 153, 168, 70, 67, 95, 127, 146, 
    106, 100, 84, 94, 89, 104, 112, 100, 91, 81, 81, 83, 59, 118, 154, 157, 
    104, 106, 89, 114, 135, 112, 116, 87, 73, 94, 88, 47, 61, 96, 117, 108, 
    58, 95, 90, 120, 124, 105, 62, 70, 54, 29, 0, 0, 0, 9, 10, 2, 
    43, 65, 125, 128, 97, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 21, 71, 98, 91, 4, 0, 0, 0, 0, 0, 0, 0, 7, 0, 7, 
    0, 0, 34, 76, 48, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 11, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    109, 91, 88, 89, 89, 88, 92, 99, 97, 80, 63, 68, 72, 82, 85, 77, 
    111, 97, 95, 91, 90, 84, 87, 95, 89, 62, 38, 47, 60, 74, 81, 76, 
    107, 86, 95, 97, 94, 89, 52, 65, 52, 21, 0, 0, 14, 55, 66, 72, 
    80, 62, 84, 98, 91, 73, 40, 10, 11, 14, 0, 0, 4, 28, 69, 63, 
    38, 8, 67, 84, 60, 18, 6, 0, 2, 29, 10, 2, 2, 8, 66, 70, 
    29, 0, 35, 73, 75, 0, 0, 0, 0, 18, 0, 0, 2, 0, 21, 63, 
    31, 0, 25, 72, 54, 0, 0, 0, 0, 8, 0, 0, 2, 0, 0, 32, 
    34, 0, 12, 46, 46, 13, 0, 0, 0, 27, 0, 0, 0, 0, 30, 50, 
    31, 0, 0, 7, 34, 20, 0, 0, 0, 26, 17, 0, 17, 32, 63, 75, 
    47, 0, 0, 0, 0, 8, 17, 0, 0, 12, 18, 10, 15, 54, 71, 72, 
    53, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 2, 2, 0, 
    19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end inmem_package;
