library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 0, 0, 13, 36, 23, 20, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 18, 22, 16, 43, 28, 27, 11, 0, 
    35, 7, 0, 0, 0, 26, 37, 29, 27, 6, 19, 26, 11, 10, 0, 
    71, 48, 8, 34, 51, 60, 46, 17, 18, 0, 64, 40, 13, 17, 7, 
    63, 71, 3, 0, 9, 30, 45, 44, 22, 21, 58, 29, 20, 15, 20, 
    75, 51, 19, 0, 0, 30, 80, 50, 26, 28, 57, 32, 17, 31, 11, 
    84, 66, 75, 24, 28, 45, 25, 19, 2, 23, 15, 40, 18, 3, 0, 
    78, 75, 66, 33, 27, 34, 17, 26, 35, 32, 36, 3, 0, 0, 0, 
    52, 67, 67, 17, 68, 20, 58, 77, 56, 23, 4, 19, 33, 20, 20, 
    66, 79, 52, 60, 131, 90, 66, 63, 56, 48, 55, 61, 65, 70, 69, 
    80, 69, 60, 101, 89, 59, 61, 58, 55, 55, 59, 62, 74, 74, 67, 
    82, 68, 66, 107, 65, 59, 63, 57, 60, 64, 75, 77, 78, 70, 106, 
    90, 76, 84, 52, 61, 63, 67, 63, 61, 66, 71, 66, 60, 86, 80, 
    
    -- channel=1
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 31, 0, 0, 0, 10, 1, 
    0, 61, 0, 1, 0, 4, 0, 0, 0, 48, 0, 0, 0, 0, 38, 
    0, 46, 0, 61, 0, 12, 0, 0, 0, 65, 0, 0, 0, 0, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 125, 0, 0, 7, 0, 0, 
    0, 0, 0, 0, 29, 26, 0, 0, 0, 87, 0, 0, 0, 10, 0, 
    0, 0, 7, 0, 44, 42, 0, 0, 0, 52, 0, 0, 14, 0, 0, 
    0, 0, 0, 12, 0, 0, 0, 0, 26, 0, 0, 0, 0, 15, 16, 
    0, 0, 0, 38, 0, 0, 21, 0, 1, 0, 0, 0, 32, 28, 0, 
    13, 0, 0, 117, 0, 17, 25, 0, 0, 0, 14, 19, 20, 0, 0, 
    28, 0, 0, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 29, 45, 0, 0, 0, 0, 0, 0, 0, 3, 7, 0, 0, 9, 
    0, 0, 82, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 33, 0, 0, 
    
    -- channel=2
    92, 96, 96, 97, 97, 90, 100, 113, 104, 77, 61, 67, 74, 80, 84, 
    94, 105, 99, 100, 97, 80, 77, 85, 57, 24, 0, 2, 29, 59, 77, 
    60, 74, 106, 107, 105, 84, 55, 27, 1, 0, 0, 0, 0, 6, 58, 
    0, 10, 88, 104, 87, 53, 5, 0, 0, 0, 0, 0, 0, 0, 26, 
    0, 0, 59, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 54, 78, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 31, 86, 13, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 28, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 
    0, 0, 0, 0, 6, 0, 0, 0, 0, 15, 5, 0, 0, 12, 50, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 67, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=3
    186, 193, 189, 194, 191, 188, 198, 194, 187, 181, 165, 159, 167, 170, 158, 
    181, 189, 194, 201, 191, 227, 227, 193, 172, 134, 161, 143, 126, 139, 163, 
    182, 136, 192, 195, 194, 234, 191, 126, 97, 162, 222, 174, 167, 105, 142, 
    200, 104, 200, 191, 208, 158, 213, 163, 146, 160, 239, 173, 142, 98, 94, 
    259, 237, 242, 176, 324, 303, 277, 181, 138, 98, 247, 206, 140, 125, 86, 
    286, 280, 259, 219, 240, 277, 299, 210, 168, 122, 326, 199, 144, 151, 112, 
    275, 325, 192, 198, 172, 237, 336, 259, 204, 190, 295, 186, 140, 150, 167, 
    313, 313, 222, 208, 172, 292, 326, 222, 176, 205, 262, 192, 133, 184, 160, 
    354, 326, 276, 196, 226, 204, 198, 189, 153, 236, 168, 158, 97, 132, 183, 
    329, 329, 298, 202, 245, 168, 179, 279, 213, 182, 155, 67, 97, 178, 200, 
    265, 326, 302, 212, 397, 265, 271, 311, 233, 145, 88, 111, 145, 173, 170, 
    204, 270, 296, 377, 456, 199, 163, 156, 137, 131, 138, 147, 154, 171, 166, 
    178, 181, 229, 448, 255, 149, 151, 140, 135, 133, 143, 161, 180, 170, 176, 
    174, 149, 187, 362, 172, 154, 159, 143, 139, 150, 162, 163, 158, 158, 219, 
    193, 149, 163, 174, 139, 124, 143, 146, 157, 173, 170, 144, 167, 243, 175, 
    
    -- channel=4
    118, 126, 120, 123, 119, 116, 130, 133, 123, 112, 98, 98, 98, 106, 103, 
    117, 125, 126, 128, 119, 111, 121, 121, 95, 52, 38, 46, 63, 91, 101, 
    110, 99, 125, 129, 125, 132, 98, 55, 31, 22, 50, 33, 37, 47, 89, 
    64, 28, 124, 124, 119, 66, 69, 33, 24, 38, 65, 48, 35, 29, 58, 
    50, 52, 116, 80, 98, 49, 79, 46, 33, 0, 64, 49, 29, 27, 21, 
    39, 78, 119, 78, 111, 86, 93, 57, 39, 3, 81, 54, 34, 25, 13, 
    31, 84, 105, 117, 61, 64, 114, 57, 64, 19, 79, 41, 19, 26, 41, 
    45, 73, 44, 87, 46, 96, 80, 67, 60, 49, 73, 51, 27, 47, 66, 
    60, 64, 45, 61, 48, 57, 69, 50, 40, 54, 85, 49, 17, 60, 95, 
    75, 63, 70, 12, 84, 21, 28, 66, 36, 80, 41, 10, 23, 78, 108, 
    57, 64, 70, 14, 62, 36, 33, 76, 51, 1, 0, 0, 0, 15, 20, 
    11, 40, 60, 59, 115, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 110, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 101, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=5
    0, 2, 0, 5, 5, 0, 0, 4, 8, 5, 3, 0, 0, 6, 12, 
    1, 0, 0, 6, 0, 0, 26, 9, 10, 0, 11, 8, 0, 0, 6, 
    26, 0, 0, 6, 0, 0, 43, 18, 0, 0, 23, 17, 31, 0, 0, 
    90, 0, 0, 0, 24, 0, 14, 22, 7, 0, 53, 2, 34, 22, 0, 
    72, 0, 30, 0, 5, 6, 52, 48, 27, 0, 13, 51, 4, 39, 0, 
    50, 0, 44, 5, 0, 6, 50, 36, 66, 0, 60, 64, 0, 24, 20, 
    49, 30, 0, 58, 0, 0, 12, 39, 66, 0, 69, 45, 0, 0, 25, 
    35, 34, 18, 21, 0, 0, 84, 11, 39, 0, 41, 54, 0, 0, 18, 
    45, 0, 93, 0, 22, 0, 24, 16, 0, 18, 0, 64, 0, 0, 0, 
    14, 0, 101, 0, 40, 6, 0, 21, 15, 13, 51, 0, 0, 0, 11, 
    0, 0, 90, 0, 86, 19, 0, 14, 62, 34, 0, 0, 0, 0, 0, 
    0, 0, 19, 0, 97, 57, 0, 0, 12, 0, 0, 0, 0, 0, 5, 
    11, 0, 0, 12, 127, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 0, 0, 81, 33, 0, 11, 0, 0, 0, 0, 0, 1, 0, 8, 
    32, 0, 0, 1, 11, 0, 0, 0, 0, 0, 10, 0, 0, 18, 44, 
    
    -- channel=6
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 7, 0, 0, 
    0, 0, 0, 0, 0, 4, 4, 30, 8, 0, 0, 0, 0, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 14, 20, 0, 0, 0, 52, 3, 7, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 5, 0, 16, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 6, 
    25, 0, 0, 0, 0, 63, 42, 49, 28, 2, 0, 0, 0, 0, 0, 
    0, 14, 0, 0, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 0, 3, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 
    0, 0, 0, 63, 9, 17, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=7
    0, 2, 4, 0, 0, 7, 0, 0, 2, 0, 3, 11, 7, 0, 0, 
    2, 3, 4, 0, 7, 31, 0, 1, 0, 31, 0, 0, 11, 15, 0, 
    0, 38, 1, 0, 2, 7, 0, 0, 11, 42, 0, 0, 0, 4, 21, 
    0, 57, 0, 10, 0, 28, 0, 0, 0, 44, 0, 0, 0, 0, 46, 
    0, 15, 0, 58, 0, 0, 0, 0, 0, 75, 0, 0, 1, 0, 9, 
    0, 12, 0, 0, 73, 0, 0, 0, 0, 129, 0, 0, 8, 0, 0, 
    0, 0, 0, 0, 58, 47, 0, 0, 0, 96, 0, 0, 3, 12, 0, 
    0, 0, 0, 0, 27, 43, 0, 0, 0, 50, 0, 0, 17, 0, 0, 
    0, 0, 0, 35, 0, 1, 0, 0, 24, 0, 11, 0, 17, 17, 0, 
    0, 0, 0, 44, 0, 0, 36, 0, 0, 0, 0, 4, 34, 20, 0, 
    58, 0, 0, 114, 0, 0, 26, 0, 0, 0, 7, 13, 16, 13, 0, 
    31, 33, 0, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 26, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 22, 0, 0, 
    
    -- channel=8
    63, 69, 68, 70, 67, 65, 71, 75, 67, 52, 42, 45, 53, 61, 59, 
    67, 72, 73, 72, 68, 69, 65, 56, 34, 17, 14, 14, 21, 39, 56, 
    43, 37, 68, 73, 71, 49, 32, 14, 13, 13, 21, 17, 15, 16, 41, 
    28, 25, 60, 67, 58, 30, 35, 21, 11, 12, 25, 17, 10, 12, 25, 
    22, 34, 58, 46, 59, 44, 32, 21, 10, 4, 29, 26, 15, 15, 14, 
    9, 22, 60, 42, 17, 30, 38, 29, 20, 11, 27, 15, 13, 12, 16, 
    14, 17, 35, 54, 27, 27, 31, 23, 24, 7, 20, 16, 8, 11, 25, 
    17, 17, 22, 35, 28, 31, 22, 13, 24, 23, 23, 15, 8, 20, 39, 
    15, 10, 12, 15, 23, 9, 21, 18, 17, 20, 18, 8, 8, 32, 58, 
    15, 14, 17, 0, 23, 15, 12, 27, 21, 18, 4, 0, 20, 45, 53, 
    0, 12, 14, 12, 35, 25, 5, 0, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 18, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=9
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 16, 21, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 6, 3, 2, 0, 0, 
    7, 0, 0, 0, 0, 2, 4, 4, 6, 10, 9, 5, 0, 0, 0, 
    6, 9, 0, 0, 0, 0, 3, 6, 7, 6, 3, 0, 3, 3, 0, 
    5, 10, 0, 0, 0, 0, 0, 2, 3, 0, 2, 4, 0, 0, 12, 
    
    -- channel=10
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=11
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 37, 0, 0, 0, 0, 28, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 10, 3, 11, 10, 0, 0, 
    37, 26, 0, 0, 0, 0, 30, 10, 0, 0, 0, 0, 0, 0, 0, 
    45, 56, 0, 0, 95, 54, 1, 7, 0, 0, 30, 22, 10, 19, 0, 
    0, 0, 0, 0, 0, 0, 25, 24, 29, 13, 0, 0, 0, 9, 34, 
    14, 0, 0, 0, 0, 2, 0, 6, 9, 0, 0, 9, 0, 12, 16, 
    9, 19, 24, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 2, 0, 0, 0, 0, 7, 6, 0, 0, 0, 0, 0, 3, 
    0, 0, 10, 2, 2, 0, 2, 53, 0, 0, 0, 0, 14, 0, 0, 
    0, 0, 0, 46, 128, 92, 0, 0, 0, 13, 41, 52, 19, 0, 0, 
    0, 0, 17, 11, 0, 0, 0, 0, 0, 0, 1, 0, 10, 5, 4, 
    10, 0, 0, 0, 0, 5, 2, 1, 5, 12, 19, 25, 0, 0, 35, 
    7, 3, 0, 0, 0, 6, 17, 6, 1, 7, 0, 0, 0, 21, 0, 
    9, 3, 0, 0, 0, 0, 0, 0, 20, 27, 10, 6, 44, 35, 14, 
    
    -- channel=12
    51, 50, 52, 52, 55, 48, 53, 57, 54, 44, 37, 40, 41, 45, 47, 
    55, 52, 56, 52, 55, 52, 41, 42, 32, 31, 19, 23, 33, 43, 45, 
    30, 53, 54, 55, 57, 56, 22, 26, 19, 33, 1, 10, 15, 33, 45, 
    0, 61, 50, 58, 43, 40, 19, 6, 15, 35, 0, 12, 4, 14, 55, 
    0, 37, 33, 62, 15, 10, 0, 0, 9, 43, 11, 0, 17, 9, 37, 
    0, 14, 18, 29, 24, 0, 0, 7, 3, 59, 0, 0, 20, 9, 12, 
    0, 4, 25, 24, 52, 23, 4, 0, 0, 57, 0, 0, 19, 17, 7, 
    0, 0, 13, 21, 45, 23, 0, 10, 0, 49, 0, 0, 20, 12, 25, 
    0, 0, 0, 25, 3, 19, 10, 15, 27, 32, 14, 0, 20, 38, 48, 
    0, 0, 0, 33, 0, 8, 25, 5, 5, 4, 2, 14, 32, 51, 41, 
    17, 0, 0, 40, 0, 0, 7, 0, 0, 4, 7, 4, 11, 21, 9, 
    10, 0, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 8, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=13
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 3, 15, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 8, 0, 7, 8, 7, 6, 0, 
    13, 0, 0, 0, 0, 0, 5, 0, 18, 0, 0, 2, 0, 5, 0, 
    32, 19, 0, 0, 14, 0, 0, 0, 12, 0, 24, 12, 2, 5, 0, 
    9, 55, 0, 0, 0, 0, 21, 0, 15, 0, 23, 5, 2, 0, 0, 
    17, 24, 3, 0, 0, 4, 37, 21, 0, 0, 14, 12, 4, 8, 0, 
    35, 35, 34, 0, 0, 17, 0, 0, 0, 0, 0, 23, 1, 0, 0, 
    25, 33, 41, 16, 17, 0, 0, 2, 13, 7, 32, 7, 0, 0, 0, 
    28, 22, 44, 0, 15, 11, 41, 60, 47, 24, 17, 31, 52, 49, 42, 
    103, 50, 17, 16, 113, 80, 77, 72, 70, 69, 79, 83, 81, 87, 84, 
    111, 89, 10, 69, 77, 72, 79, 73, 73, 74, 82, 83, 97, 96, 84, 
    111, 98, 68, 102, 65, 74, 75, 75, 77, 82, 97, 103, 101, 93, 138, 
    111, 103, 99, 90, 81, 83, 86, 75, 72, 78, 91, 84, 69, 109, 113, 
    
    -- channel=14
    56, 57, 57, 54, 52, 54, 62, 63, 52, 45, 44, 48, 47, 48, 44, 
    54, 59, 59, 57, 54, 28, 41, 51, 43, 11, 0, 3, 29, 48, 45, 
    39, 67, 60, 59, 60, 40, 22, 9, 8, 0, 0, 0, 0, 28, 46, 
    0, 28, 54, 55, 38, 24, 0, 0, 0, 15, 0, 0, 0, 0, 46, 
    0, 0, 33, 41, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 23, 
    0, 0, 31, 41, 29, 10, 0, 0, 0, 20, 0, 0, 0, 0, 0, 
    0, 0, 42, 25, 23, 7, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 15, 12, 0, 0, 0, 8, 0, 0, 0, 3, 13, 
    0, 0, 0, 0, 2, 7, 0, 0, 1, 0, 17, 0, 8, 18, 39, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 9, 28, 31, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    74, 68, 75, 75, 72, 66, 78, 81, 71, 55, 46, 51, 57, 64, 63, 
    73, 72, 77, 75, 78, 30, 76, 52, 38, 21, 7, 12, 24, 53, 61, 
    26, 53, 78, 76, 78, 25, 36, 24, 35, 0, 16, 16, 2, 34, 42, 
    6, 20, 76, 72, 45, 46, 18, 31, 8, 25, 9, 18, 10, 15, 32, 
    31, 0, 79, 89, 17, 44, 16, 18, 0, 31, 21, 26, 6, 7, 25, 
    51, 0, 86, 51, 0, 57, 4, 26, 0, 14, 20, 26, 12, 11, 18, 
    71, 0, 65, 49, 0, 27, 3, 23, 8, 0, 23, 18, 7, 14, 27, 
    49, 0, 47, 32, 45, 12, 14, 9, 28, 2, 15, 14, 13, 17, 53, 
    17, 0, 28, 1, 44, 17, 27, 0, 30, 0, 25, 10, 10, 34, 60, 
    4, 7, 2, 0, 37, 34, 26, 0, 27, 28, 0, 9, 8, 35, 57, 
    0, 13, 0, 14, 3, 31, 0, 0, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 28, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end gold_package;
