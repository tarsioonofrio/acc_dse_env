library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    146, 126, 125, 126, 125, 123, 125, 127, 129, 125, 123, 122, 128, 124, 126, 213, 
    119, 117, 112, 113, 116, 120, 112, 122, 120, 104, 104, 92, 97, 117, 123, 218, 
    108, 111, 123, 121, 114, 91, 144, 104, 131, 82, 74, 86, 94, 87, 120, 222, 
    138, 91, 118, 119, 118, 103, 129, 125, 90, 31, 98, 65, 109, 111, 103, 225, 
    128, 57, 106, 110, 137, 94, 72, 105, 87, 77, 107, 105, 104, 122, 103, 231, 
    74, 38, 120, 135, 27, 92, 105, 98, 128, 56, 40, 96, 78, 108, 130, 202, 
    97, 58, 112, 157, 26, 78, 97, 95, 143, 0, 82, 103, 74, 85, 98, 197, 
    93, 101, 125, 159, 68, 25, 56, 70, 109, 0, 82, 92, 70, 48, 107, 218, 
    45, 43, 133, 107, 132, 40, 102, 84, 94, 75, 91, 105, 87, 99, 104, 231, 
    24, 0, 108, 25, 99, 132, 82, 96, 90, 124, 111, 130, 89, 85, 105, 237, 
    33, 13, 97, 13, 106, 110, 43, 57, 118, 99, 128, 114, 41, 66, 95, 216, 
    0, 19, 102, 0, 46, 69, 26, 32, 66, 94, 57, 22, 29, 17, 33, 166, 
    11, 0, 34, 0, 81, 95, 41, 37, 37, 36, 25, 23, 12, 15, 16, 172, 
    27, 22, 0, 102, 102, 25, 40, 35, 36, 27, 15, 7, 23, 11, 0, 191, 
    18, 16, 18, 107, 82, 27, 36, 35, 28, 20, 17, 22, 24, 0, 55, 174, 
    36, 14, 31, 35, 59, 37, 36, 32, 15, 19, 29, 29, 0, 27, 51, 149, 
    
    -- channel=1
    156, 159, 161, 165, 163, 161, 166, 168, 166, 155, 130, 120, 130, 133, 127, 116, 
    159, 164, 164, 171, 168, 214, 238, 171, 167, 138, 127, 113, 107, 126, 132, 125, 
    155, 156, 168, 168, 168, 199, 193, 122, 79, 122, 161, 136, 114, 86, 126, 132, 
    130, 106, 176, 172, 180, 163, 171, 144, 84, 136, 170, 144, 107, 64, 93, 122, 
    215, 203, 221, 197, 293, 276, 197, 165, 98, 98, 211, 180, 102, 94, 53, 84, 
    233, 241, 256, 167, 243, 279, 241, 219, 134, 138, 240, 181, 102, 102, 73, 48, 
    250, 237, 246, 163, 143, 231, 273, 261, 168, 152, 241, 167, 105, 121, 118, 97, 
    278, 249, 222, 171, 151, 260, 298, 228, 155, 158, 215, 171, 107, 125, 125, 127, 
    297, 273, 244, 174, 189, 177, 194, 160, 147, 149, 153, 154, 60, 106, 149, 147, 
    295, 284, 260, 182, 206, 148, 160, 223, 195, 163, 141, 77, 68, 140, 163, 158, 
    254, 296, 255, 246, 341, 270, 239, 264, 242, 120, 65, 71, 91, 148, 153, 140, 
    192, 270, 262, 327, 374, 281, 133, 142, 127, 101, 78, 81, 97, 110, 108, 99, 
    111, 186, 258, 350, 335, 147, 86, 76, 75, 78, 88, 107, 113, 114, 134, 152, 
    107, 92, 214, 310, 259, 97, 97, 86, 77, 85, 93, 100, 102, 118, 147, 136, 
    115, 92, 103, 164, 152, 78, 99, 94, 95, 111, 112, 87, 135, 160, 139, 94, 
    113, 95, 84, 84, 75, 49, 58, 63, 84, 120, 116, 95, 147, 168, 126, 65, 
    
    -- channel=2
    66, 32, 30, 26, 26, 31, 23, 29, 33, 31, 26, 32, 29, 20, 23, 21, 
    69, 34, 33, 27, 34, 71, 16, 35, 36, 46, 23, 25, 32, 30, 27, 20, 
    79, 49, 34, 28, 36, 80, 0, 21, 31, 62, 2, 0, 0, 35, 45, 14, 
    79, 65, 32, 37, 39, 47, 42, 7, 10, 49, 0, 0, 0, 12, 55, 22, 
    70, 27, 0, 91, 97, 16, 22, 0, 0, 85, 43, 0, 2, 0, 56, 54, 
    66, 36, 0, 88, 123, 0, 21, 0, 0, 122, 16, 0, 5, 0, 11, 45, 
    36, 50, 0, 12, 108, 36, 38, 0, 0, 108, 0, 0, 10, 8, 0, 0, 
    63, 33, 0, 25, 54, 97, 0, 0, 0, 61, 0, 0, 15, 13, 0, 7, 
    96, 0, 0, 19, 36, 67, 0, 4, 10, 18, 26, 0, 24, 16, 10, 13, 
    128, 0, 0, 28, 0, 31, 36, 42, 14, 0, 3, 10, 44, 30, 14, 22, 
    180, 0, 0, 83, 0, 2, 30, 16, 0, 0, 1, 19, 27, 25, 20, 25, 
    175, 0, 0, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    100, 7, 42, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    82, 0, 72, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    82, 0, 23, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    83, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=3
    163, 154, 140, 144, 146, 144, 151, 160, 158, 149, 143, 142, 137, 132, 139, 132, 
    165, 154, 145, 146, 147, 126, 154, 155, 152, 143, 134, 149, 150, 158, 138, 132, 
    156, 179, 158, 156, 159, 201, 188, 159, 150, 112, 53, 62, 77, 153, 153, 130, 
    125, 197, 178, 155, 147, 156, 133, 58, 63, 120, 92, 96, 95, 93, 150, 137, 
    74, 33, 138, 152, 77, 63, 50, 67, 86, 119, 123, 70, 91, 59, 150, 167, 
    84, 74, 126, 138, 166, 113, 58, 60, 72, 77, 47, 83, 85, 76, 67, 135, 
    78, 67, 166, 153, 129, 125, 88, 57, 63, 72, 81, 83, 89, 96, 56, 80, 
    68, 49, 120, 147, 104, 95, 106, 111, 107, 97, 106, 83, 89, 85, 106, 109, 
    72, 49, 34, 96, 99, 155, 178, 110, 99, 130, 157, 128, 115, 114, 111, 121, 
    123, 58, 50, 89, 79, 109, 104, 44, 93, 135, 104, 130, 77, 100, 137, 138, 
    133, 61, 58, 53, 0, 62, 30, 64, 46, 149, 148, 74, 66, 121, 127, 129, 
    132, 137, 46, 21, 118, 130, 140, 164, 135, 88, 38, 32, 30, 47, 45, 31, 
    80, 137, 125, 67, 119, 90, 27, 34, 36, 39, 35, 27, 19, 28, 13, 0, 
    24, 61, 105, 148, 77, 31, 29, 35, 30, 19, 21, 42, 38, 48, 40, 73, 
    14, 16, 72, 171, 102, 67, 63, 41, 21, 20, 22, 36, 32, 0, 47, 63, 
    108, 90, 100, 101, 98, 93, 96, 117, 129, 125, 113, 98, 128, 139, 105, 90, 
    
    -- channel=4
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 22, 68, 0, 0, 10, 52, 48, 15, 0, 0, 0, 
    0, 0, 0, 0, 0, 18, 80, 16, 9, 34, 104, 94, 62, 22, 0, 0, 
    92, 47, 0, 0, 0, 7, 64, 82, 34, 35, 116, 87, 61, 37, 0, 2, 
    180, 98, 111, 0, 159, 198, 143, 124, 48, 29, 121, 121, 44, 46, 13, 0, 
    187, 156, 169, 0, 160, 243, 169, 154, 74, 33, 176, 138, 47, 51, 50, 0, 
    197, 177, 180, 4, 35, 149, 173, 197, 102, 53, 192, 133, 55, 49, 66, 25, 
    214, 205, 210, 54, 27, 107, 204, 173, 104, 49, 165, 123, 56, 54, 69, 6, 
    244, 204, 231, 90, 116, 92, 155, 84, 80, 52, 74, 108, 30, 42, 36, 8, 
    233, 209, 223, 134, 148, 107, 71, 145, 168, 80, 53, 54, 5, 4, 7, 15, 
    164, 225, 204, 141, 284, 215, 120, 190, 212, 98, 45, 54, 77, 81, 93, 103, 
    129, 215, 213, 156, 300, 277, 128, 152, 158, 113, 97, 106, 123, 128, 132, 156, 
    145, 139, 182, 243, 301, 195, 111, 106, 95, 95, 110, 125, 136, 137, 153, 201, 
    163, 140, 115, 273, 289, 114, 123, 110, 102, 114, 124, 133, 141, 134, 167, 197, 
    169, 142, 136, 187, 194, 98, 121, 120, 112, 132, 137, 123, 131, 190, 196, 137, 
    172, 141, 131, 110, 99, 72, 83, 91, 98, 133, 144, 119, 131, 204, 194, 119, 
    
    -- channel=5
    165, 165, 167, 165, 165, 160, 170, 173, 167, 154, 143, 141, 143, 139, 136, 123, 
    165, 167, 167, 173, 172, 189, 159, 166, 157, 142, 122, 108, 123, 143, 141, 130, 
    149, 170, 176, 170, 177, 229, 195, 139, 126, 140, 137, 116, 95, 117, 139, 133, 
    123, 129, 170, 173, 167, 174, 143, 98, 99, 152, 165, 116, 105, 80, 125, 136, 
    147, 165, 168, 184, 223, 185, 175, 115, 93, 157, 158, 120, 98, 72, 92, 128, 
    163, 201, 176, 198, 268, 199, 204, 140, 101, 183, 191, 131, 103, 102, 56, 87, 
    159, 198, 182, 166, 180, 202, 232, 183, 138, 208, 201, 123, 105, 105, 99, 86, 
    187, 206, 131, 159, 149, 231, 239, 168, 145, 199, 190, 138, 100, 132, 124, 126, 
    208, 209, 144, 156, 160, 236, 183, 144, 121, 158, 180, 122, 104, 127, 145, 153, 
    232, 219, 185, 156, 156, 142, 158, 176, 131, 141, 131, 78, 77, 161, 164, 157, 
    229, 219, 193, 223, 197, 158, 208, 225, 154, 115, 76, 61, 88, 139, 141, 124, 
    203, 229, 196, 307, 303, 198, 181, 181, 133, 77, 82, 88, 90, 99, 98, 87, 
    128, 181, 231, 298, 250, 107, 78, 77, 77, 78, 83, 90, 103, 103, 109, 109, 
    83, 115, 213, 303, 144, 95, 87, 75, 78, 85, 96, 107, 106, 106, 122, 132, 
    92, 80, 160, 199, 137, 98, 95, 92, 92, 98, 86, 90, 113, 131, 115, 80, 
    93, 94, 85, 89, 70, 73, 79, 83, 106, 115, 107, 103, 151, 154, 99, 64, 
    
    -- channel=6
    58, 60, 56, 58, 60, 56, 57, 60, 62, 55, 53, 51, 56, 55, 59, 110, 
    57, 60, 56, 60, 58, 82, 68, 60, 63, 47, 43, 40, 36, 53, 60, 115, 
    57, 54, 62, 62, 60, 60, 73, 52, 49, 29, 34, 40, 41, 35, 59, 115, 
    67, 24, 61, 60, 71, 53, 61, 59, 39, 6, 50, 29, 42, 39, 34, 118, 
    65, 32, 60, 59, 86, 80, 42, 50, 38, 17, 43, 55, 35, 47, 44, 122, 
    53, 19, 63, 72, 30, 55, 65, 45, 64, 0, 40, 53, 28, 38, 49, 83, 
    57, 45, 46, 87, 5, 24, 57, 58, 67, 0, 40, 44, 24, 30, 38, 100, 
    49, 47, 70, 82, 52, 24, 50, 30, 45, 1, 42, 39, 23, 21, 41, 112, 
    28, 17, 75, 53, 69, 12, 39, 47, 27, 48, 30, 54, 23, 34, 47, 128, 
    21, 3, 58, 0, 51, 60, 35, 64, 58, 50, 51, 39, 33, 32, 45, 122, 
    23, 14, 49, 0, 74, 54, 4, 33, 59, 40, 25, 32, 11, 16, 34, 110, 
    0, 10, 40, 0, 41, 43, 0, 0, 8, 22, 18, 3, 1, 0, 9, 70, 
    1, 0, 17, 31, 41, 23, 6, 4, 3, 0, 0, 0, 0, 0, 0, 82, 
    0, 0, 0, 63, 36, 3, 5, 1, 1, 0, 0, 0, 0, 0, 0, 70, 
    0, 0, 0, 29, 23, 0, 3, 8, 0, 0, 1, 0, 0, 0, 3, 58, 
    5, 2, 1, 8, 13, 8, 9, 6, 0, 1, 6, 5, 0, 6, 12, 43, 
    
    -- channel=7
    142, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    138, 0, 0, 0, 0, 1, 0, 0, 0, 23, 13, 6, 12, 10, 0, 0, 
    141, 15, 0, 0, 0, 16, 0, 0, 20, 81, 30, 17, 18, 22, 45, 0, 
    177, 75, 28, 0, 0, 0, 23, 0, 37, 93, 62, 23, 22, 19, 65, 18, 
    233, 86, 0, 0, 77, 0, 28, 0, 28, 89, 103, 0, 35, 14, 51, 66, 
    247, 102, 0, 0, 110, 0, 51, 0, 7, 159, 98, 0, 46, 28, 16, 50, 
    252, 117, 0, 0, 115, 41, 62, 0, 4, 165, 53, 0, 37, 47, 25, 18, 
    268, 104, 0, 53, 64, 93, 0, 12, 6, 129, 37, 0, 52, 49, 18, 5, 
    297, 54, 0, 72, 0, 83, 38, 25, 44, 39, 42, 0, 58, 61, 7, 0, 
    297, 37, 8, 99, 28, 0, 84, 72, 32, 63, 2, 39, 76, 37, 0, 0, 
    261, 16, 10, 146, 81, 12, 66, 67, 0, 6, 56, 66, 74, 78, 41, 46, 
    227, 95, 27, 144, 46, 9, 75, 73, 72, 75, 84, 89, 95, 87, 81, 84, 
    214, 121, 103, 131, 0, 76, 75, 78, 78, 86, 95, 95, 97, 88, 104, 98, 
    221, 100, 135, 178, 34, 82, 85, 81, 85, 89, 91, 98, 89, 115, 117, 84, 
    228, 102, 106, 139, 64, 97, 93, 84, 87, 89, 87, 95, 120, 110, 84, 71, 
    228, 98, 90, 79, 77, 97, 91, 87, 98, 94, 68, 88, 118, 99, 68, 89, 
    
    -- channel=8
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    
    -- channel=9
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 68, 62, 33, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 12, 29, 40, 42, 34, 31, 25, 0, 0, 
    96, 83, 0, 0, 0, 0, 16, 18, 30, 14, 30, 19, 23, 30, 0, 0, 
    125, 133, 0, 0, 28, 36, 15, 16, 25, 34, 57, 40, 32, 42, 37, 0, 
    125, 131, 0, 0, 0, 2, 49, 37, 40, 64, 76, 46, 40, 48, 47, 0, 
    115, 132, 77, 0, 0, 52, 77, 50, 27, 55, 68, 47, 44, 40, 16, 0, 
    152, 161, 141, 82, 0, 37, 48, 20, 38, 0, 7, 23, 30, 23, 0, 0, 
    145, 164, 152, 111, 92, 25, 21, 76, 64, 7, 18, 34, 43, 0, 0, 0, 
    145, 134, 122, 133, 168, 129, 144, 157, 144, 86, 140, 175, 195, 168, 140, 149, 
    291, 239, 157, 133, 191, 218, 228, 232, 245, 257, 285, 302, 321, 326, 324, 332, 
    363, 311, 214, 160, 228, 275, 277, 269, 274, 295, 325, 339, 340, 346, 371, 372, 
    394, 371, 287, 237, 245, 288, 288, 279, 289, 315, 344, 358, 361, 394, 403, 374, 
    395, 384, 348, 273, 265, 286, 293, 288, 295, 319, 341, 349, 365, 406, 410, 343, 
    368, 356, 345, 288, 272, 279, 284, 279, 286, 313, 316, 313, 340, 377, 377, 329, 
    
    -- channel=10
    148, 102, 96, 98, 92, 96, 97, 91, 86, 81, 70, 77, 82, 78, 68, 53, 
    147, 99, 100, 101, 106, 184, 111, 96, 90, 102, 109, 91, 73, 81, 81, 62, 
    145, 100, 105, 98, 103, 171, 93, 57, 67, 184, 168, 126, 100, 77, 96, 71, 
    171, 139, 133, 104, 115, 123, 157, 82, 93, 206, 184, 120, 103, 40, 103, 93, 
    235, 228, 144, 185, 282, 204, 207, 110, 90, 183, 220, 119, 100, 74, 77, 100, 
    248, 276, 158, 149, 295, 211, 261, 139, 113, 282, 257, 128, 115, 99, 53, 64, 
    231, 302, 138, 121, 225, 253, 300, 172, 144, 306, 249, 121, 107, 136, 111, 70, 
    280, 305, 135, 163, 170, 329, 276, 170, 136, 269, 223, 131, 118, 147, 110, 95, 
    346, 297, 180, 200, 148, 235, 166, 150, 152, 163, 161, 98, 95, 117, 113, 103, 
    358, 296, 237, 245, 185, 119, 193, 254, 158, 160, 112, 42, 100, 141, 122, 94, 
    333, 283, 239, 375, 359, 186, 260, 304, 152, 110, 85, 113, 141, 158, 134, 124, 
    308, 293, 253, 436, 411, 167, 197, 188, 144, 123, 136, 151, 165, 172, 162, 162, 
    198, 273, 322, 426, 256, 142, 138, 130, 129, 138, 160, 175, 178, 178, 212, 218, 
    177, 180, 341, 425, 130, 158, 152, 135, 139, 153, 164, 181, 174, 203, 216, 207, 
    186, 159, 220, 277, 120, 152, 158, 144, 165, 177, 161, 159, 233, 249, 194, 139, 
    189, 155, 153, 142, 106, 121, 126, 125, 166, 183, 162, 164, 252, 249, 146, 121, 
    
    -- channel=11
    42, 44, 42, 41, 42, 45, 40, 43, 44, 44, 46, 46, 45, 45, 48, 87, 
    20, 25, 23, 25, 23, 9, 18, 36, 59, 39, 32, 39, 42, 39, 32, 89, 
    53, 47, 27, 25, 22, 55, 57, 61, 54, 17, 29, 36, 45, 39, 33, 89, 
    62, 23, 22, 22, 27, 28, 32, 43, 38, 14, 38, 34, 53, 56, 30, 89, 
    45, 0, 27, 24, 16, 28, 30, 44, 49, 35, 36, 36, 41, 54, 49, 100, 
    39, 14, 38, 30, 31, 43, 26, 40, 58, 11, 22, 52, 33, 43, 53, 87, 
    46, 37, 46, 49, 23, 19, 38, 45, 64, 0, 34, 48, 35, 33, 38, 76, 
    35, 41, 51, 43, 23, 12, 63, 35, 49, 0, 33, 53, 37, 32, 45, 86, 
    6, 8, 62, 22, 34, 26, 54, 31, 30, 35, 45, 70, 46, 34, 24, 92, 
    8, 0, 48, 18, 38, 72, 34, 27, 35, 55, 75, 60, 40, 15, 31, 100, 
    9, 1, 58, 4, 14, 7, 11, 43, 70, 54, 52, 35, 24, 26, 39, 109, 
    15, 24, 26, 0, 57, 80, 40, 47, 60, 45, 38, 29, 31, 23, 29, 105, 
    43, 7, 32, 10, 71, 60, 34, 33, 35, 32, 27, 24, 29, 32, 24, 120, 
    43, 30, 9, 77, 61, 31, 32, 33, 34, 30, 29, 30, 34, 27, 47, 129, 
    44, 30, 28, 89, 60, 42, 41, 43, 27, 24, 31, 31, 23, 18, 50, 110, 
    93, 82, 82, 82, 83, 76, 76, 70, 72, 89, 95, 86, 79, 110, 102, 110, 
    
    -- channel=12
    26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 
    28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 8, 0, 
    1, 20, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 24, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    
    -- channel=13
    204, 214, 215, 213, 208, 217, 219, 205, 193, 188, 176, 167, 178, 175, 154, 132, 
    190, 206, 215, 218, 221, 324, 333, 208, 199, 193, 228, 209, 159, 163, 159, 149, 
    191, 201, 211, 214, 215, 348, 342, 178, 136, 303, 365, 322, 243, 137, 166, 171, 
    220, 178, 223, 215, 237, 230, 304, 267, 198, 332, 389, 314, 256, 137, 149, 172, 
    436, 415, 379, 314, 545, 510, 435, 341, 218, 262, 423, 347, 227, 193, 92, 132, 
    510, 534, 464, 292, 611, 608, 508, 431, 274, 335, 516, 384, 232, 230, 160, 91, 
    526, 527, 464, 232, 382, 478, 576, 518, 357, 415, 529, 358, 230, 263, 260, 173, 
    589, 572, 439, 274, 289, 559, 629, 486, 357, 414, 504, 367, 231, 289, 277, 189, 
    665, 643, 539, 380, 354, 497, 480, 336, 298, 301, 359, 319, 182, 241, 232, 223, 
    671, 655, 593, 423, 433, 289, 359, 464, 401, 298, 263, 186, 153, 234, 251, 224, 
    593, 651, 583, 571, 714, 540, 502, 579, 483, 270, 171, 199, 266, 309, 299, 270, 
    539, 630, 595, 775, 852, 624, 444, 458, 400, 269, 285, 310, 343, 364, 358, 348, 
    396, 513, 604, 805, 771, 394, 303, 287, 275, 283, 321, 357, 377, 377, 424, 444, 
    376, 343, 552, 743, 586, 329, 326, 298, 293, 322, 348, 373, 379, 394, 449, 460, 
    388, 354, 392, 495, 408, 308, 331, 318, 334, 369, 362, 339, 424, 495, 449, 331, 
    386, 352, 335, 305, 258, 237, 261, 269, 328, 385, 379, 332, 464, 518, 426, 275, 
    
    -- channel=14
    174, 174, 173, 175, 182, 174, 176, 192, 190, 168, 137, 133, 140, 149, 152, 144, 
    179, 181, 176, 181, 180, 190, 179, 188, 175, 144, 134, 113, 120, 146, 152, 147, 
    156, 167, 183, 187, 189, 202, 164, 138, 125, 94, 69, 60, 67, 114, 141, 148, 
    103, 154, 175, 190, 182, 170, 152, 81, 56, 78, 81, 78, 67, 69, 113, 131, 
    70, 82, 169, 192, 197, 163, 93, 73, 61, 113, 101, 84, 72, 44, 92, 108, 
    90, 99, 165, 161, 186, 108, 111, 94, 68, 92, 96, 76, 65, 60, 53, 89, 
    98, 94, 145, 152, 147, 148, 131, 97, 80, 92, 103, 85, 74, 76, 55, 69, 
    94, 88, 128, 142, 143, 136, 134, 109, 88, 113, 106, 98, 67, 65, 109, 117, 
    90, 88, 77, 107, 140, 128, 127, 113, 90, 153, 168, 70, 67, 95, 127, 146, 
    106, 100, 84, 94, 89, 104, 112, 100, 91, 81, 81, 83, 59, 118, 154, 157, 
    104, 106, 89, 114, 135, 112, 116, 87, 73, 94, 88, 47, 61, 96, 117, 108, 
    58, 95, 90, 120, 124, 105, 62, 70, 54, 29, 0, 0, 0, 9, 10, 2, 
    43, 65, 125, 128, 97, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 21, 71, 98, 91, 4, 0, 0, 0, 0, 0, 0, 0, 7, 0, 7, 
    0, 0, 34, 76, 48, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 11, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    109, 91, 88, 89, 89, 88, 92, 99, 97, 80, 63, 68, 72, 82, 85, 77, 
    111, 97, 95, 91, 90, 84, 87, 95, 89, 62, 38, 47, 60, 74, 81, 76, 
    107, 86, 95, 97, 94, 89, 52, 65, 52, 21, 0, 0, 14, 55, 66, 72, 
    80, 62, 84, 98, 91, 73, 40, 10, 11, 14, 0, 0, 4, 28, 69, 63, 
    38, 8, 67, 84, 60, 18, 6, 0, 2, 29, 10, 2, 2, 8, 66, 70, 
    29, 0, 35, 73, 75, 0, 0, 0, 0, 18, 0, 0, 2, 0, 21, 63, 
    31, 0, 25, 72, 54, 0, 0, 0, 0, 8, 0, 0, 2, 0, 0, 32, 
    34, 0, 12, 46, 46, 13, 0, 0, 0, 27, 0, 0, 0, 0, 30, 50, 
    31, 0, 0, 7, 34, 20, 0, 0, 0, 26, 17, 0, 17, 32, 63, 75, 
    47, 0, 0, 0, 0, 8, 17, 0, 0, 12, 18, 10, 15, 54, 71, 72, 
    53, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 2, 2, 0, 
    19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end ifmap_package;
