-- https://docs.xilinx.com/r/en-US/ug953-vivado-7series-libraries/BRAM_SINGLE_MACRO

library UNISIM;
use UNISIM.vcomponents.all;
library UNIMACRO;
use unimacro.Vcomponents.all;


-- BRAM_SINGLE_MACRO: Single Port RAM
--                    7 Series
-- Xilinx HDL Language Template, version 2021.2

-- Note -  This Unimacro model assumes the port directions to be "downto".
--         Simulation of this model with "to" in the port directions could lead to erroneous results.

---------------------------------------------------------------------
--  READ_WIDTH | BRAM_SIZE | READ Depth  | ADDR Width |            --
-- WRITE_WIDTH |           | WRITE Depth |            |  WE Width  --
-- ============|===========|=============|============|============--
--    37-72    |  "36Kb"   |      512    |    9-bit   |    8-bit   --
--    19-36    |  "36Kb"   |     1024    |   10-bit   |    4-bit   --
--    19-36    |  "18Kb"   |      512    |    9-bit   |    4-bit   --
--    10-18    |  "36Kb"   |     2048    |   11-bit   |    2-bit   --
--    10-18    |  "18Kb"   |     1024    |   10-bit   |    2-bit   --
--     5-9     |  "36Kb"   |     4096    |   12-bit   |    1-bit   --
--     5-9     |  "18Kb"   |     2048    |   11-bit   |    1-bit   --
--     3-4     |  "36Kb"   |     8192    |   13-bit   |    1-bit   --
--     3-4     |  "18Kb"   |     4096    |   12-bit   |    1-bit   --
--       2     |  "36Kb"   |    16384    |   14-bit   |    1-bit   --
--       2     |  "18Kb"   |     8192    |   13-bit   |    1-bit   --
--       1     |  "36Kb"   |    32768    |   15-bit   |    1-bit   --
--       1     |  "18Kb"   |    16384    |   14-bit   |    1-bit   --
---------------------------------------------------------------------

entity gold_18k_layer2_entity2 is
    generic (
        DEVICE: string := "7SERIES"
        );
  
    port (
        RST  : in std_logic;
        CLK  : in std_logic;
        EN   : in std_logic;
        WE   : in std_logic_vector(2-1 downto 0);;
        DI   : in std_logic_vector(16-1 downto 0);
        ADDR : in std_logic_vector(10-1 downto 0);
        DO   : out std_logic_vector(16-1 downto 0)
    );
  end gold_18k_layer2_entity2;

  architecture a1 of bram is

    begin

    BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
    generic map (
       BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
       DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
       DO_REG => 0,                     -- Optional output register (0 or 1)
       INIT => X"000000000000000000",   -- Initial values on output port
       INIT_FILE => "NONE",
       WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       SRVAL => X"000000000000000000",  -- Set/Reset value for port output
       WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
       -- The following INIT_xx declarations specify the initial contents of the RAM
       INIT_00 => X"009c0000000000000000000000000000000000000000000000000000000f0071",
       INIT_01 => X"00000000000000000000002d00000000000a002b000000000072004f003200c7",
       INIT_02 => X"003a000000530000000001db01760128008300cc009e002c003f0104008c0000",
       INIT_03 => X"0000012900640000007b0000008a007e005c000a000000000000004300000051",
       INIT_04 => X"0000000000000021002b00000000017800f100010024008d0079004200580060",
       INIT_05 => X"0000000000000000000000000000000000000000000000000000000000030044",
       INIT_06 => X"000e00000096002b000000100008000000000000001f00000000000000000000",
       INIT_07 => X"000000000000000000000000000000000000000000000000000000000000003b",
       INIT_08 => X"00000000000000000050005a00f800620000000000e200000000000000000000",
       INIT_09 => X"00000000000000000000000000000000000000000000000000000051008700ae",
       INIT_0A => X"0000009000cf011a00e3010d00000000000000000091000000000052013800ae",
       INIT_0B => X"0047005000000197007c006a007f00f9002b00bc010100ef0000000000000098",
       INIT_0C => X"00e30000003d00210000017b010a003301c30162013b00890059013b00e70030",
       INIT_0D => X"01150113017f0000000000000000000000000063009b01320000000000000000",
       INIT_0E => X"00a50000000f0027000801aa00ca000001620000000000000000000001380164",
       INIT_0F => X"01580000009501920032002d015400420114007c0049015e00da012e0212026d",
       INIT_10 => X"003f000000000014000000000000007600000000000000000000000000000000",
       INIT_11 => X"0000000b00000009005500000036004900000000009c00000000000000000000",
       INIT_12 => X"00000000000000000000000000000000002b001c00000000000000aa010d0000",
       INIT_13 => X"00e000cf0074010e00b1004e0000000000000000000000000000000000710000",
       INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_15 => X"00000034006100590000006e017c00320000010000c500a001d300ee009c00e8",
       INIT_16 => X"0190014e007500ed006900ff00fc00e6002e005500de000000d4006501260084",
       INIT_17 => X"0094007b00520000000000000000000000000000000000000000000000540000",
       INIT_18 => X"000000000000003e0000000000080083004f000300000000004c007300000000",
       INIT_19 => X"0000001600000000008300800032000000000069000000f5007700bf00ad0078",
       INIT_1A => X"005a0079000000fb0011000000a900760037000000000000001a000000000000",
       INIT_1B => X"00000008000000000000000000000000000000000000005a002a000800070000",
       INIT_1C => X"001a00000000001b000000000044008d0000003e000000000000006000000000",
       INIT_1D => X"001000000000001f001b00660010004800000000000000000000000000000000",
       INIT_1E => X"000000970037003d0059014a00be0086007300e100000000000000000000001c",
       INIT_1F => X"00000000002e0000000000000000000000000000000000000000000000000000",
       INIT_20 => X"00000000000000000000002c002a00890048003700810039000100f800000000",
       INIT_21 => X"00000000000000000000000000000000003700000000003e0000003000000000",
       INIT_22 => X"00000000000000000000000000000000000000ee00d100b2015200d900ec001b",
       INIT_23 => X"008e009b00a600de006f0068000000420000000000000000000000000000000d",
       INIT_24 => X"00be0000003b00d300000000000000000000000000000000000000dd0151015c",
       INIT_25 => X"015600e600a90115009c0000000000000000000000000042000000000012010e",
       INIT_26 => X"00520078010f0000000000af0008002b00070000000000000000001700000055",
       INIT_27 => X"00b800000037000000000047000000390054000000000000000e003f00000000",
       INIT_28 => X"0000000000190000000000000000000000000000000000390047000000ad0075",
       INIT_29 => X"0000000c003f00f0000000000000000000000000000000000000000000f4010e",
       INIT_2A => X"019101530000000001a20166000000d100000017003b00000000000400150039",
       INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_2C => X"0000000000000000000000000000000000290000000000000000000000000000",
       INIT_2D => X"00000000000000000066000000000085003f0000000500a30000000000450000",
       INIT_2E => X"000000000060003c0000000000280005000000000000009200000000006d0000",
       INIT_2F => X"000000220095003e0000004a00a2000000000000000000000000000000000000",
       INIT_30 => X"0000000001110000003c00ab001600ce0000000000c7007f002b009600a50043",
       INIT_31 => X"00ba00dd001e0026015b00ab00d7003f000000f400da00000161015a013900f2",
       INIT_32 => X"00b2011b0190007b011400000000000000980000000000000044000000000000",
       INIT_33 => X"0000000000370000002300a60000000000000000000000000000000000000000",
       INIT_34 => X"007000a5010e00c6000000e000de0089008300190086007800a0005100540000",
       INIT_35 => X"0000000000000000000000000000003100000000000000000000000000000000",
       INIT_36 => X"000000000000000000e4011800cd002d00c40000003b00910096007d00000000",
       INIT_37 => X"0076002600000000000000000000000000560000000000d4003d0000002c0000",
       INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_39 => X"000000000048008a00be005d009700000056004e004d0003005c0000000100dd",
       INIT_3A => X"001a0000002a0020000000000055000000000000000000000000000000410000",
       INIT_3B => X"0000000000be002f002b000000000000001c0000000000000000000000000000",
       INIT_3C => X"00000026000000550000004900b00000000000000000001e0022003e00930025",
       INIT_3D => X"00340054003d004c00be0000000000290000006d000000000000000000000000",
       INIT_3E => X"000000000000000000000000000000000000000000000000002b0000000000df",
       INIT_3F => X"00000000005a000000cf00860000006d001e0000000000320000000000000000",

       -- The next set of INITP_xx are for the parity bits
       INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

    port map (
       DO => DO,      -- Output data, width defined by READ_WIDTH parameter
       ADDR => ADDR,  -- Input address, width defined by read/write port depth
       CLK => CLK,    -- 1-bit input clock
       DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
       EN => EN,      -- 1-bit input RAM enable
       REGCE => REGCE, -- 1-bit input output register enable
       RST => RST,    -- 1-bit input reset
       WE => WE       -- Input write enable, width defined by write port depth
    );


-- End of BRAM_SINGLE_MACRO_inst instantiation
