library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package inmem_package is
  type mem is array(0 to 4000000) of integer;

  constant input_mem : mem := (
    -- bias
    2441, -1091, -2467, -412, 1901, -841, -1714, -667, -2181, -484, -2046, 1445, 91, -4220, -2420, -152, -1273, -1126, -1144, -2006, -4584, -1398, 2058, -6835, -764, 853, 3991, 2784, -548, 481, 54, -104, -1167, 2470, -633, -1106, -269, 2793, 2087, -817, -4994, -1170, -3141, -4656, -3850, 1422, 644, 1301, -1510, 992, -3068, -1605, 782, -2150, -1237, -403, -1374, -676, -1302, 3453, 94, -2445, 155, -3076, -1728, -2924, -425, 2497, 160, 1145, -814, -492, 99, 1339, 5045, 3540, 973, -196, 194, -54, -2736, 3663, -820, -2413, -87, -2793, 313, -112, 1317, -531, 450, 722, -1988, -4829, 1940, -1390, 1499, 1366, -737, -1283, 1671, 1503, -1265, 11, 1307, 934, 3812, -3462, 635, -3735, -2560, -2834, 3573, 3935, 3667, -5375, -1141, 537, 1612, -890, 1165, 1584, 1690, 2232, 1209, 1250, -1031, 1291, -1327, 1098, 196, 3340, 1579, -2069, 2305, -1543, 5650, -549, 708, -945, -1542, -2385, -1649, -1619, -429, 4556, 3134, -1918, -1750, 912, -134, 710, 1112, 622, -1035, 960, 5342, -167, 658, -822, -2449, -2586, -2175, 685, -228, 1337, -1899, -1142, -1861, 887, 4081, 1116, -1413, -2622, 2474, -1431, -323, 3630, -1875, 998, 3325, 2450, 3251, 1868, 3086, 1841, 791, 3495, 886, -1721, 3242, 465, 1867, -1127, 652, -2009, 3091, -1693, -1080, 2650, 1456, 782, -1015, -60, -1424, 280, 2343, -1513, 44, -1421, -398, 90, 1596, 2916, 4044, -95, -2766, 942, 1436, -1522, -144, -2813, -80, -992, 2328, -588, -1044, -2847, -4653, -31, 1988, -59, -295, -3775, -236, 1658, -1773, -139, -1796, -3957, -317, -1976, 109, 1558, 2293, -1953, -92, -896, 966, 2827, 384, 1481, 2243, 3076, -1018, 586,

    -- weights
    -- filter=0 channel=0
    10, 11, 2, -1, 7, 11, -9, 0, -7,
    -- filter=0 channel=1
    2, 12, 8, -8, -4, 9, -19, -12, 4,
    -- filter=0 channel=2
    5, 3, 7, -6, -6, -8, -5, 0, -11,
    -- filter=0 channel=3
    10, -6, -1, 0, -5, -7, -1, 0, -3,
    -- filter=0 channel=4
    3, 3, 3, -3, -15, -11, -3, -19, -12,
    -- filter=0 channel=5
    3, 2, 3, 5, 2, 4, 6, -12, -1,
    -- filter=0 channel=6
    -7, 7, 4, 0, -4, 1, 0, 1, -2,
    -- filter=0 channel=7
    0, -4, 0, -4, -2, -4, -2, 4, -3,
    -- filter=0 channel=8
    0, -1, -3, 5, 2, -4, -5, -2, -3,
    -- filter=0 channel=9
    -3, -1, 0, 5, 6, 0, 4, -2, 3,
    -- filter=0 channel=10
    0, -3, 0, 0, 11, 2, -7, 8, 3,
    -- filter=0 channel=11
    -3, -2, 2, -3, 3, 0, -4, 3, 8,
    -- filter=0 channel=12
    -4, -2, 0, -4, 11, 8, -10, 6, -5,
    -- filter=0 channel=13
    -7, 7, -4, -14, 18, 2, -5, 14, -1,
    -- filter=0 channel=14
    2, -3, 0, -4, 4, 0, -5, 2, 0,
    -- filter=0 channel=15
    -9, 10, 0, -4, 1, 8, -17, 7, -4,
    -- filter=0 channel=16
    -1, -4, -4, 4, -5, -8, 0, 3, 5,
    -- filter=0 channel=17
    2, -3, 0, 3, 4, -5, 7, 0, 2,
    -- filter=0 channel=18
    -13, 19, 8, -21, 8, 1, -16, 1, -2,
    -- filter=0 channel=19
    -3, 3, 1, 2, 0, -3, 5, 4, -4,
    -- filter=0 channel=20
    -14, -8, -9, -14, -2, 0, -1, 0, -2,
    -- filter=0 channel=21
    3, -12, 0, 10, 4, -5, 19, 4, -7,
    -- filter=0 channel=22
    -4, -1, 5, 2, 1, 2, -10, -2, -2,
    -- filter=0 channel=23
    -5, 5, 7, -1, 4, 9, -6, 10, 0,
    -- filter=0 channel=24
    2, 7, -5, -7, 3, -2, -1, 5, 4,
    -- filter=0 channel=25
    1, 14, 9, -13, 14, 0, -10, 1, 1,
    -- filter=0 channel=26
    4, 3, 0, 13, -5, -7, 6, -5, -7,
    -- filter=0 channel=27
    3, 10, 9, -1, 5, 5, -9, 0, 0,
    -- filter=0 channel=28
    0, -6, 7, -5, -6, 1, 2, 4, 1,
    -- filter=0 channel=29
    -12, -6, -3, -1, 0, -5, -7, -2, -2,
    -- filter=0 channel=30
    7, 2, -5, 1, 1, 2, -3, -11, -2,
    -- filter=0 channel=31
    -4, -10, 0, 17, 5, -13, 18, 11, -3,
    -- filter=0 channel=32
    -8, 15, 3, -22, 6, 6, -20, 5, 2,
    -- filter=0 channel=33
    -7, 11, -1, -9, 16, 10, -17, 4, 0,
    -- filter=0 channel=34
    1, 5, 5, 0, -7, 9, -1, 2, 5,
    -- filter=0 channel=35
    -3, 7, 5, -5, 5, -6, 1, -4, 5,
    -- filter=0 channel=36
    -8, 0, -5, 4, 6, -12, 5, -5, -1,
    -- filter=0 channel=37
    12, 6, 5, 1, -6, 8, -7, -12, -7,
    -- filter=0 channel=38
    -6, 0, 0, 1, 8, -3, 5, -1, 3,
    -- filter=0 channel=39
    -5, -5, -4, -2, -3, -1, -4, 6, 4,
    -- filter=0 channel=40
    -6, 0, -4, 6, 5, 6, 8, 6, 6,
    -- filter=0 channel=41
    -15, 21, 8, -26, 7, -2, -30, 1, 0,
    -- filter=0 channel=42
    4, 0, -2, -1, 1, -1, 3, -3, -9,
    -- filter=0 channel=43
    3, 1, 5, -12, -8, -6, -2, 0, 0,
    -- filter=0 channel=44
    4, 7, 1, 0, -5, 9, 2, -5, 1,
    -- filter=0 channel=45
    5, 2, 2, 1, 5, 2, 1, 2, -3,
    -- filter=0 channel=46
    -5, -2, 0, -8, -4, 0, 0, 0, 6,
    -- filter=0 channel=47
    4, 1, 0, 12, -3, -2, 6, 1, -9,
    -- filter=0 channel=48
    -2, 2, -4, 0, -5, 6, 5, -14, -9,
    -- filter=0 channel=49
    6, 14, 12, -15, 1, 5, -10, -2, -4,
    -- filter=0 channel=50
    9, -4, 1, 3, 7, 0, 0, 0, 3,
    -- filter=0 channel=51
    1, -5, -3, -2, -3, 0, 7, 6, -5,
    -- filter=0 channel=52
    -3, 0, -7, -5, -4, 3, -2, 0, -2,
    -- filter=0 channel=53
    -10, -2, -3, 1, 7, -1, -3, -5, -1,
    -- filter=0 channel=54
    -6, 5, 2, 1, 2, 1, -1, -3, 6,
    -- filter=0 channel=55
    -13, 0, -2, -7, 7, -2, -12, 6, -2,
    -- filter=0 channel=56
    5, -5, 2, -1, -1, 8, -4, 2, -3,
    -- filter=0 channel=57
    4, 6, 8, 2, 4, 2, -8, -5, -4,
    -- filter=0 channel=58
    11, 1, -6, 3, -6, 2, -6, -3, -2,
    -- filter=0 channel=59
    -8, 11, 0, -11, 7, 9, -4, -7, 3,
    -- filter=0 channel=60
    2, 2, 0, 2, -4, -5, 4, -4, 1,
    -- filter=0 channel=61
    -6, -1, -1, 0, -4, 5, 5, 6, 0,
    -- filter=0 channel=62
    2, 0, 3, -4, -3, -6, -3, -1, -3,
    -- filter=0 channel=63
    6, 2, -3, 2, 0, -11, 4, -2, -6,
    -- filter=0 channel=64
    -6, -9, -5, -1, -4, -6, 3, -3, 6,
    -- filter=0 channel=65
    3, -5, -1, -3, -5, -3, 1, 5, -1,
    -- filter=0 channel=66
    -8, 3, -6, -5, 14, 0, -6, 3, 2,
    -- filter=0 channel=67
    -6, 3, 7, -6, 4, 3, 3, -4, 0,
    -- filter=0 channel=68
    -7, -1, 4, -8, -5, -10, 0, -3, -3,
    -- filter=0 channel=69
    -5, -8, -5, 2, -2, 6, -5, 1, 2,
    -- filter=0 channel=70
    2, 4, 2, -1, 1, 12, -3, 5, 2,
    -- filter=0 channel=71
    9, -2, 3, 0, 0, -3, 5, 4, 5,
    -- filter=0 channel=72
    0, -5, -7, 4, 0, -2, 9, 5, 4,
    -- filter=0 channel=73
    -5, 0, 8, -11, 3, -3, -10, 0, -6,
    -- filter=0 channel=74
    8, 3, 1, 0, 0, 2, 7, -3, 0,
    -- filter=0 channel=75
    8, 7, 1, -9, 9, 9, -17, -2, -8,
    -- filter=0 channel=76
    -7, 1, 1, -9, 10, -6, -4, 15, 4,
    -- filter=0 channel=77
    -6, 6, 0, 5, -1, 2, -6, 0, 0,
    -- filter=0 channel=78
    0, -2, -4, 1, -4, -3, 0, -6, -4,
    -- filter=0 channel=79
    -12, 19, 9, -23, 16, 8, -31, -1, -1,
    -- filter=0 channel=80
    -3, -3, 1, -5, 2, 3, 9, -3, -7,
    -- filter=0 channel=81
    1, 2, 1, 6, 3, 2, 0, -6, 7,
    -- filter=0 channel=82
    0, -4, -2, 0, -2, -5, 4, -2, -3,
    -- filter=0 channel=83
    0, -4, 6, 8, -3, -7, -4, -1, -5,
    -- filter=0 channel=84
    -5, 12, 10, -7, -1, 3, -14, -7, -5,
    -- filter=0 channel=85
    6, -5, 4, 1, 7, 6, 5, -6, -5,
    -- filter=0 channel=86
    3, 0, 6, 0, -4, -3, -7, -3, 2,
    -- filter=0 channel=87
    -9, -6, 0, 2, 3, 8, -1, -1, 5,
    -- filter=0 channel=88
    -2, -8, 1, 3, -6, -1, 16, -2, 6,
    -- filter=0 channel=89
    -6, 7, 0, -20, 7, 2, -3, 6, -6,
    -- filter=0 channel=90
    4, 1, -5, 6, -8, 0, 17, 4, 4,
    -- filter=0 channel=91
    1, 4, 4, -8, 1, 4, -11, 1, 5,
    -- filter=0 channel=92
    6, 0, 2, 9, -5, -2, -7, -4, 2,
    -- filter=0 channel=93
    9, -3, -2, -1, -7, 0, 0, -8, -9,
    -- filter=0 channel=94
    -2, -6, -5, 1, 7, 5, 7, -6, 6,
    -- filter=0 channel=95
    -3, 1, 6, -2, -2, -6, 5, 3, -5,
    -- filter=0 channel=96
    -2, -4, -3, -6, -6, -6, 0, -2, 5,
    -- filter=0 channel=97
    10, -1, -2, 4, -4, 6, -6, 0, 0,
    -- filter=0 channel=98
    -6, 8, 4, -7, 4, 0, -13, -2, -2,
    -- filter=0 channel=99
    -14, 0, -12, 6, 3, 0, 9, 5, -5,
    -- filter=0 channel=100
    2, -6, 0, -1, 0, -4, -3, 3, -7,
    -- filter=0 channel=101
    -2, 0, 0, -9, -11, -5, -3, -1, -9,
    -- filter=0 channel=102
    -5, 0, -6, 7, -5, -1, -1, 5, 0,
    -- filter=0 channel=103
    -1, -9, 4, 2, -7, 3, -1, -10, -4,
    -- filter=0 channel=104
    -5, -8, -9, 3, 3, -3, 12, 0, -2,
    -- filter=0 channel=105
    -10, -7, -2, 0, -3, 3, -5, 0, -3,
    -- filter=0 channel=106
    -6, 4, -3, -3, 3, -2, -3, 6, -5,
    -- filter=0 channel=107
    -6, 5, 2, 0, 0, 1, -14, -2, -5,
    -- filter=0 channel=108
    -6, 2, 1, -9, -4, 5, -8, 0, -8,
    -- filter=0 channel=109
    -6, 14, 5, -19, 9, 12, -6, 1, 3,
    -- filter=0 channel=110
    -7, -5, -2, 1, 3, -4, 1, 10, -3,
    -- filter=0 channel=111
    -3, 0, 1, -2, -7, -6, -1, -1, 7,
    -- filter=0 channel=112
    8, -2, -3, 0, -2, 9, -6, -5, 0,
    -- filter=0 channel=113
    -2, 2, 4, -3, 6, 0, -5, 7, 4,
    -- filter=0 channel=114
    -10, 15, 12, -20, 2, 0, -26, -15, 0,
    -- filter=0 channel=115
    5, 6, 6, 2, 6, 0, -1, -6, -2,
    -- filter=0 channel=116
    -3, 0, 3, -11, -2, -10, -12, -10, 0,
    -- filter=0 channel=117
    0, -1, 4, -4, -2, 3, -3, 0, 4,
    -- filter=0 channel=118
    6, 1, 2, 1, 7, -5, -3, -2, 1,
    -- filter=0 channel=119
    9, 0, -1, 5, -5, -2, 0, 0, 8,
    -- filter=0 channel=120
    1, 7, 3, 0, -5, 3, 0, -2, -8,
    -- filter=0 channel=121
    -4, -1, 0, -7, -1, 5, -9, 6, 3,
    -- filter=0 channel=122
    0, -8, -5, 16, 0, -6, 25, -7, 4,
    -- filter=0 channel=123
    -1, -3, 3, 8, 3, -1, 5, -4, 8,
    -- filter=0 channel=124
    -3, 0, 3, -10, 2, -6, -6, 4, 0,
    -- filter=0 channel=125
    -3, -3, 3, 2, 8, -3, 7, -5, 0,
    -- filter=0 channel=126
    -13, 6, -1, -14, -1, 0, -9, -4, -5,
    -- filter=0 channel=127
    0, -3, -3, 0, 2, 3, 1, 3, -7,
    -- filter=1 channel=0
    -7, -7, -15, 1, -4, -13, 2, 4, 0,
    -- filter=1 channel=1
    -14, -15, -20, -7, -5, -9, -1, 1, 2,
    -- filter=1 channel=2
    0, 1, 10, -5, 6, 2, 7, 3, 4,
    -- filter=1 channel=3
    -3, -4, 4, -7, -6, -7, -9, -3, -4,
    -- filter=1 channel=4
    -3, 9, 7, 0, -5, -3, 0, 8, 9,
    -- filter=1 channel=5
    -4, -9, -9, 6, 5, 5, -5, 0, 13,
    -- filter=1 channel=6
    1, 5, 4, 0, 0, 6, -6, -8, -2,
    -- filter=1 channel=7
    1, -2, 1, 2, 0, -6, 0, 4, 0,
    -- filter=1 channel=8
    -5, -3, 6, -7, -5, 6, -4, 7, 1,
    -- filter=1 channel=9
    -7, -2, 2, -6, 3, 3, 3, 7, 9,
    -- filter=1 channel=10
    -2, -5, -2, -4, -6, -3, 2, -4, 1,
    -- filter=1 channel=11
    -1, 10, 12, 5, 6, 7, -14, -4, -13,
    -- filter=1 channel=12
    2, -5, 0, 8, 6, 2, -2, 8, 5,
    -- filter=1 channel=13
    8, -5, 6, 0, -5, 1, 0, -8, -9,
    -- filter=1 channel=14
    0, 5, 4, 0, 5, 2, -4, 2, -2,
    -- filter=1 channel=15
    -2, 11, 9, -10, -1, -2, 0, -12, -6,
    -- filter=1 channel=16
    -5, -16, 0, 4, -4, -6, -6, 5, 8,
    -- filter=1 channel=17
    0, 3, 0, 7, 2, 4, 3, 1, -3,
    -- filter=1 channel=18
    0, 0, -4, -2, 0, 0, -6, 7, -2,
    -- filter=1 channel=19
    7, -6, 6, 0, -1, 0, -3, 0, 1,
    -- filter=1 channel=20
    -1, 18, 17, 7, 15, 15, -17, -15, -7,
    -- filter=1 channel=21
    -9, -15, -2, -10, -11, 4, 0, -2, 7,
    -- filter=1 channel=22
    -3, 3, -1, 2, -5, -7, 0, 3, -4,
    -- filter=1 channel=23
    2, 6, 13, -2, -8, 0, -6, -8, -4,
    -- filter=1 channel=24
    1, 0, 3, 0, -6, -4, 1, -2, 3,
    -- filter=1 channel=25
    -4, 0, 0, -5, -4, 0, 10, 4, -1,
    -- filter=1 channel=26
    2, 0, 0, -3, 3, -3, -8, 0, -2,
    -- filter=1 channel=27
    -4, -4, -4, -5, -9, 0, 3, 6, 8,
    -- filter=1 channel=28
    0, 0, 2, -2, -6, 4, 3, 0, 0,
    -- filter=1 channel=29
    10, 22, 16, 0, 8, 14, -17, -15, -5,
    -- filter=1 channel=30
    -5, -3, 2, -12, 0, -4, 1, 6, 11,
    -- filter=1 channel=31
    -6, -13, 2, -11, -8, 0, 5, 0, 12,
    -- filter=1 channel=32
    -3, 1, -5, 0, 2, -5, -4, 0, -8,
    -- filter=1 channel=33
    0, 0, -1, -6, -4, 0, -2, -3, -5,
    -- filter=1 channel=34
    7, 1, -3, 4, 6, -4, 0, 12, 0,
    -- filter=1 channel=35
    7, 6, -6, -2, 3, -6, -2, -5, 4,
    -- filter=1 channel=36
    -2, -5, 9, 0, -5, 2, 5, 1, -1,
    -- filter=1 channel=37
    -13, -17, -19, -8, -5, 0, 2, -3, 1,
    -- filter=1 channel=38
    1, -7, 5, -9, -6, 4, 1, -6, 3,
    -- filter=1 channel=39
    2, 8, 9, 0, 0, 11, 0, -8, 2,
    -- filter=1 channel=40
    2, 1, 6, -3, -3, 4, 0, -3, -2,
    -- filter=1 channel=41
    1, 10, 5, 5, 14, -12, -1, 6, 1,
    -- filter=1 channel=42
    -5, -10, 3, -3, 3, -8, -1, -5, -3,
    -- filter=1 channel=43
    0, 0, 5, -5, -8, -5, -3, 1, -1,
    -- filter=1 channel=44
    -10, -14, -14, -1, -6, -8, 2, 2, 12,
    -- filter=1 channel=45
    -4, 0, 5, -5, -2, 3, 0, -5, 4,
    -- filter=1 channel=46
    5, 3, 5, -2, 0, -8, -6, 1, 1,
    -- filter=1 channel=47
    -19, -24, -16, -9, -11, -3, -9, -9, 10,
    -- filter=1 channel=48
    -14, -13, 0, -10, -11, 0, 1, 7, 9,
    -- filter=1 channel=49
    6, 7, 9, 0, -2, 5, 1, 3, 2,
    -- filter=1 channel=50
    3, -8, -3, 4, -5, -3, 8, 9, 7,
    -- filter=1 channel=51
    -1, -2, -7, -6, 0, 2, -7, -4, 6,
    -- filter=1 channel=52
    2, 6, 0, -4, -5, 0, -5, -7, -4,
    -- filter=1 channel=53
    -4, 8, 5, -3, 1, 6, -2, -10, -8,
    -- filter=1 channel=54
    -3, -6, -3, 5, 0, 5, -5, -2, 4,
    -- filter=1 channel=55
    6, 7, 14, 4, -1, 4, -2, -8, -6,
    -- filter=1 channel=56
    7, -3, 2, 1, -5, -2, 7, -1, -3,
    -- filter=1 channel=57
    4, 2, 2, 2, 0, -3, -6, -5, -5,
    -- filter=1 channel=58
    0, 0, -7, 2, -3, 6, -9, 2, 7,
    -- filter=1 channel=59
    -4, 0, 1, 0, -8, 2, 9, 10, 3,
    -- filter=1 channel=60
    -2, 0, 0, -2, 5, -4, 1, 7, -6,
    -- filter=1 channel=61
    7, 0, 8, 0, 1, 7, -3, 6, 4,
    -- filter=1 channel=62
    1, 5, 4, -6, 1, -4, 3, -4, 3,
    -- filter=1 channel=63
    -3, -2, -3, 3, 2, 7, 6, -1, 9,
    -- filter=1 channel=64
    2, 2, 0, -3, -2, -1, 4, -2, -2,
    -- filter=1 channel=65
    1, 3, 6, -6, -3, 5, -1, -6, 3,
    -- filter=1 channel=66
    3, 0, -6, -1, 0, -3, 9, 10, 1,
    -- filter=1 channel=67
    6, 8, 4, 0, 8, 3, 0, -1, -2,
    -- filter=1 channel=68
    8, -3, 4, 7, 4, -4, 7, 7, 1,
    -- filter=1 channel=69
    -7, 3, 7, 4, 1, 2, -4, 0, 6,
    -- filter=1 channel=70
    -3, 1, 5, 5, -4, 4, 1, 2, -3,
    -- filter=1 channel=71
    -5, 4, 0, 1, -3, -5, -6, -9, -4,
    -- filter=1 channel=72
    0, 1, 2, 5, 1, 4, 9, -7, 0,
    -- filter=1 channel=73
    -1, 7, -1, 0, 1, 6, 5, -3, -4,
    -- filter=1 channel=74
    4, -3, -6, -5, -1, 6, -6, 10, 5,
    -- filter=1 channel=75
    -1, -8, -9, -5, -12, -3, -1, 2, 12,
    -- filter=1 channel=76
    5, 20, 15, -4, 14, 3, -9, -10, -12,
    -- filter=1 channel=77
    -2, -1, 3, 0, 1, 6, 0, -2, -1,
    -- filter=1 channel=78
    0, -8, -6, -6, -5, 6, -6, -1, 0,
    -- filter=1 channel=79
    0, 9, -3, 2, 0, 1, 2, -4, -5,
    -- filter=1 channel=80
    -8, -11, -7, -3, -17, 7, 2, -4, 13,
    -- filter=1 channel=81
    -6, 4, -4, 0, 3, -3, 5, -2, 5,
    -- filter=1 channel=82
    -6, 8, 1, 4, 2, -4, 3, 4, 3,
    -- filter=1 channel=83
    -10, 1, 0, -7, -6, 2, 5, 5, 1,
    -- filter=1 channel=84
    8, 0, 4, 7, 2, 8, 0, 8, 0,
    -- filter=1 channel=85
    6, -2, -3, -4, -1, -4, 6, -3, 0,
    -- filter=1 channel=86
    5, -5, -1, 0, 2, 8, -2, 4, 1,
    -- filter=1 channel=87
    3, 8, 9, 7, 9, 1, -2, -6, 0,
    -- filter=1 channel=88
    8, 6, 5, 1, -2, 4, -5, -4, 1,
    -- filter=1 channel=89
    2, 6, -3, -6, -2, -3, 4, -9, -4,
    -- filter=1 channel=90
    -2, -2, -7, 3, 0, -4, -5, 3, -2,
    -- filter=1 channel=91
    4, 6, 3, 4, -1, -3, -5, 9, 6,
    -- filter=1 channel=92
    7, 3, 0, -2, 0, 5, -6, 1, -5,
    -- filter=1 channel=93
    -11, -19, -2, -14, -14, 0, -3, 0, 5,
    -- filter=1 channel=94
    -1, 2, 5, 0, -2, -4, -7, -1, -1,
    -- filter=1 channel=95
    0, -6, -5, -6, -4, 0, -6, 4, 2,
    -- filter=1 channel=96
    -2, 5, 2, 6, -3, -7, 3, 0, 2,
    -- filter=1 channel=97
    -1, 0, 5, -11, -13, -7, -1, -3, 5,
    -- filter=1 channel=98
    -4, -10, 0, -2, -4, -2, 0, 2, 2,
    -- filter=1 channel=99
    5, 4, 0, 3, -1, 16, 1, 0, 2,
    -- filter=1 channel=100
    9, 4, 0, 7, 2, -2, -3, 2, -2,
    -- filter=1 channel=101
    0, 7, 11, -8, -10, 5, 6, 0, -3,
    -- filter=1 channel=102
    -6, 0, 4, -2, 6, -2, 5, 4, 7,
    -- filter=1 channel=103
    -18, -7, -9, -17, -19, -3, 1, 1, 1,
    -- filter=1 channel=104
    -14, -18, 2, -10, -12, 3, 7, -2, 6,
    -- filter=1 channel=105
    -2, 12, 11, -1, 10, 10, -17, -13, -3,
    -- filter=1 channel=106
    3, 9, -4, 5, -3, 7, -1, -11, -10,
    -- filter=1 channel=107
    8, 12, 2, -5, 7, 9, -1, -7, -5,
    -- filter=1 channel=108
    2, -6, -3, 5, 4, 4, -3, 3, 2,
    -- filter=1 channel=109
    5, 3, -6, -1, -7, -2, 11, 8, 4,
    -- filter=1 channel=110
    -5, -6, -5, 0, -9, 8, -4, -3, 0,
    -- filter=1 channel=111
    7, 1, 2, -4, -2, -3, -6, -5, 4,
    -- filter=1 channel=112
    -5, -11, -4, -2, -2, 0, 2, 5, 8,
    -- filter=1 channel=113
    -5, 2, 1, 4, -3, -3, 9, -7, -6,
    -- filter=1 channel=114
    6, 3, 0, 0, -1, -4, -3, 6, -6,
    -- filter=1 channel=115
    3, -1, 2, -2, 0, 0, 6, 0, -5,
    -- filter=1 channel=116
    5, 5, 6, -4, 3, 0, 2, 3, 9,
    -- filter=1 channel=117
    5, -2, 5, 5, 2, 3, 1, 4, -1,
    -- filter=1 channel=118
    6, 7, 2, 3, 4, 3, 3, -6, 5,
    -- filter=1 channel=119
    2, -3, -6, 3, 6, 6, 2, 1, -2,
    -- filter=1 channel=120
    5, 2, 9, -4, 1, 9, -14, 0, -4,
    -- filter=1 channel=121
    -3, 6, -3, 0, -1, -4, 8, 5, 6,
    -- filter=1 channel=122
    -31, -24, -27, -21, -17, 0, -2, -4, 12,
    -- filter=1 channel=123
    6, 6, -2, 4, -6, 0, 3, 0, 4,
    -- filter=1 channel=124
    -6, 4, 5, 4, -1, 11, -9, -3, -1,
    -- filter=1 channel=125
    -6, 4, 0, -4, 0, -2, 0, 3, 11,
    -- filter=1 channel=126
    -3, 5, -6, -4, -4, -2, -3, -8, -4,
    -- filter=1 channel=127
    -3, 0, 3, 2, 7, 3, -5, 0, -6,
    -- filter=2 channel=0
    7, 10, 5, -2, -3, -3, 8, -5, -8,
    -- filter=2 channel=1
    4, -5, -4, 12, -4, -3, 13, -10, -14,
    -- filter=2 channel=2
    -7, -6, 0, 3, 3, 5, 8, -1, 0,
    -- filter=2 channel=3
    7, 9, 0, 0, -5, 1, 0, 10, 3,
    -- filter=2 channel=4
    -3, 1, 5, 12, 21, 6, 5, -4, 1,
    -- filter=2 channel=5
    0, 4, 3, 2, 4, 2, 7, 0, 4,
    -- filter=2 channel=6
    8, 6, 0, 9, 6, 0, 0, -3, -7,
    -- filter=2 channel=7
    0, -6, -1, 1, -4, 1, -4, -7, 3,
    -- filter=2 channel=8
    0, -4, -4, 9, 1, -7, -1, 0, -8,
    -- filter=2 channel=9
    -6, -4, 3, 0, 1, 11, 0, -3, 5,
    -- filter=2 channel=10
    -1, -10, -16, -13, -1, 8, 10, 1, 10,
    -- filter=2 channel=11
    3, -8, 0, 0, 10, 14, 2, -2, 7,
    -- filter=2 channel=12
    5, -9, -4, 0, 3, -2, 2, -7, -10,
    -- filter=2 channel=13
    -2, -17, -11, -8, 3, 7, 1, -5, -9,
    -- filter=2 channel=14
    6, -7, 4, -5, -3, 2, -1, -1, 5,
    -- filter=2 channel=15
    -14, -14, -3, -15, 2, 4, 0, 2, -5,
    -- filter=2 channel=16
    7, 1, -1, -1, 0, -4, 0, 6, -3,
    -- filter=2 channel=17
    -6, -5, 1, -3, -6, -7, 6, -3, 7,
    -- filter=2 channel=18
    -12, -24, -8, -10, 11, 21, 15, 10, -3,
    -- filter=2 channel=19
    0, 1, 2, -3, -5, 6, -4, -4, -2,
    -- filter=2 channel=20
    -2, -7, 2, -2, 5, 7, 2, -3, -1,
    -- filter=2 channel=21
    1, -4, 0, -10, -9, -1, -3, 0, 2,
    -- filter=2 channel=22
    -1, -5, -6, -1, -7, 0, 5, -3, 0,
    -- filter=2 channel=23
    -4, -13, -15, -18, 7, 7, -3, 9, -6,
    -- filter=2 channel=24
    0, 2, 2, -6, -3, -2, -1, 0, 1,
    -- filter=2 channel=25
    -2, -17, -5, 1, 5, 6, 6, 1, -2,
    -- filter=2 channel=26
    6, 1, 0, -1, 6, 7, 5, 3, 0,
    -- filter=2 channel=27
    -24, -20, -19, -11, 15, 11, 6, 0, -7,
    -- filter=2 channel=28
    0, 3, 3, 5, 2, 4, 0, 4, -2,
    -- filter=2 channel=29
    -2, 2, 15, -4, 12, 23, 2, 4, 3,
    -- filter=2 channel=30
    -8, -1, -8, 0, 9, 3, -2, 5, -8,
    -- filter=2 channel=31
    -5, -4, -23, -3, -1, 2, 8, 4, 8,
    -- filter=2 channel=32
    -12, -23, -14, -3, 2, 8, 0, 10, -6,
    -- filter=2 channel=33
    -9, -10, -16, -6, -7, -1, 8, 11, -6,
    -- filter=2 channel=34
    1, 3, -3, 0, 11, -9, 6, -10, 1,
    -- filter=2 channel=35
    -4, -5, -7, 6, -1, -5, 0, -6, 5,
    -- filter=2 channel=36
    1, -8, -3, 8, 1, 6, 0, -5, 0,
    -- filter=2 channel=37
    3, -4, 1, 9, 2, -1, 12, 0, -7,
    -- filter=2 channel=38
    2, -7, -6, -7, -4, 5, -1, -1, 6,
    -- filter=2 channel=39
    -6, -1, 7, 0, 8, 5, 1, -7, -7,
    -- filter=2 channel=40
    -3, 0, 1, -4, -8, 5, -10, 0, -4,
    -- filter=2 channel=41
    0, -7, -10, 6, -7, -9, 7, 1, 0,
    -- filter=2 channel=42
    2, -2, 0, -2, 0, 5, -2, 1, 0,
    -- filter=2 channel=43
    6, -8, 0, 1, -2, -2, -2, 1, -1,
    -- filter=2 channel=44
    0, -6, 0, 1, -3, -6, 7, -2, -2,
    -- filter=2 channel=45
    -4, 2, -5, 1, 2, 6, -4, -2, 4,
    -- filter=2 channel=46
    -6, -4, -1, -4, -5, -3, -5, 5, -7,
    -- filter=2 channel=47
    -4, -7, -9, -1, -4, 0, 0, 1, 7,
    -- filter=2 channel=48
    -7, -14, -5, 6, 0, 7, 15, -4, -3,
    -- filter=2 channel=49
    -15, -10, 0, 10, 17, 11, 7, -4, 2,
    -- filter=2 channel=50
    -6, -4, -4, -13, 8, 2, -2, -5, 3,
    -- filter=2 channel=51
    4, -4, 6, 2, 7, 5, 5, 2, 0,
    -- filter=2 channel=52
    -10, -7, -7, -3, 2, -3, -3, -3, 3,
    -- filter=2 channel=53
    -6, 2, -2, -5, 1, 2, 5, 7, 3,
    -- filter=2 channel=54
    3, -4, 5, -7, 6, 5, 4, -6, -3,
    -- filter=2 channel=55
    -8, -7, -14, -3, 3, 15, 12, 11, 5,
    -- filter=2 channel=56
    0, 4, -1, -2, 4, 2, -6, 1, 0,
    -- filter=2 channel=57
    -6, -3, 1, -5, -1, 4, 8, 5, 0,
    -- filter=2 channel=58
    3, 0, 6, 9, -6, 7, 8, -5, 7,
    -- filter=2 channel=59
    -3, -11, -2, -1, -1, 2, 7, 12, 7,
    -- filter=2 channel=60
    6, -5, -4, 0, 5, 0, 0, 0, 3,
    -- filter=2 channel=61
    4, 4, 4, 1, 3, 3, -2, 4, -1,
    -- filter=2 channel=62
    -3, 1, -7, 4, 2, -3, -5, 0, -4,
    -- filter=2 channel=63
    7, 12, 3, 2, -3, 5, 2, -1, 4,
    -- filter=2 channel=64
    4, 6, -2, 6, 1, -6, -2, 1, -5,
    -- filter=2 channel=65
    2, -4, 6, 4, 5, 6, 7, 7, -6,
    -- filter=2 channel=66
    1, -4, -2, 4, 1, 1, -3, -4, -13,
    -- filter=2 channel=67
    5, -6, -5, -5, -6, -4, -4, 2, 0,
    -- filter=2 channel=68
    -2, 4, 2, 7, 0, 6, 7, 0, -7,
    -- filter=2 channel=69
    7, 3, 0, -6, 3, -6, -5, -2, 0,
    -- filter=2 channel=70
    -13, -23, -19, -7, 1, 0, -2, 2, -2,
    -- filter=2 channel=71
    8, 4, -5, 0, -7, -3, -1, -5, 4,
    -- filter=2 channel=72
    -6, -16, -16, -2, 0, 2, 0, 4, 2,
    -- filter=2 channel=73
    -8, -11, -7, -6, 5, 6, 11, 8, -6,
    -- filter=2 channel=74
    -9, -1, -6, -4, 15, -1, -5, -9, -4,
    -- filter=2 channel=75
    7, 5, -9, -9, -9, -7, 9, 11, 2,
    -- filter=2 channel=76
    8, -5, -4, -11, 9, 3, -4, 4, -6,
    -- filter=2 channel=77
    0, 0, -3, -5, 6, -4, 0, -5, 5,
    -- filter=2 channel=78
    0, 3, -2, 0, 4, 3, 4, 1, 7,
    -- filter=2 channel=79
    -7, -28, -6, -3, 0, 8, 15, 0, -13,
    -- filter=2 channel=80
    -8, -18, -12, -12, -3, 5, 8, 12, 0,
    -- filter=2 channel=81
    -4, 3, 1, -7, 2, 0, -5, 0, 3,
    -- filter=2 channel=82
    5, -1, -4, -2, -4, 5, -7, -3, 1,
    -- filter=2 channel=83
    -8, 5, 2, 4, 0, 7, 7, -2, -4,
    -- filter=2 channel=84
    -14, -5, -2, 2, 8, 12, 6, 4, 0,
    -- filter=2 channel=85
    6, -5, 6, -5, -5, 3, 7, -3, 0,
    -- filter=2 channel=86
    1, 4, 2, -1, 7, -5, 3, 2, -11,
    -- filter=2 channel=87
    -6, 4, 7, 2, 9, 3, 2, -4, -7,
    -- filter=2 channel=88
    5, 5, -5, 5, 2, -7, 2, -8, -2,
    -- filter=2 channel=89
    1, -23, -7, -8, -2, 16, 8, 10, 5,
    -- filter=2 channel=90
    7, 1, -11, -5, 0, -3, -4, -4, -1,
    -- filter=2 channel=91
    -21, -4, -4, 5, 12, 14, 8, -1, -3,
    -- filter=2 channel=92
    4, 2, -3, 0, -1, -5, -5, -4, -3,
    -- filter=2 channel=93
    -4, -5, 4, -1, 0, 4, 7, 0, -5,
    -- filter=2 channel=94
    -5, -4, -3, 4, -3, 5, -1, 2, 3,
    -- filter=2 channel=95
    -5, -1, 0, 0, 4, 0, 0, -3, 0,
    -- filter=2 channel=96
    -4, 6, -5, -1, 4, 2, 1, 5, -3,
    -- filter=2 channel=97
    7, 6, -5, -5, -8, 0, 0, 5, 0,
    -- filter=2 channel=98
    -11, -12, -9, -10, 1, 16, 15, 8, 6,
    -- filter=2 channel=99
    0, -7, -8, -5, 9, 14, 1, 10, 8,
    -- filter=2 channel=100
    0, 6, 0, -2, -5, 0, 6, -4, -8,
    -- filter=2 channel=101
    -9, 0, 14, 10, 17, 0, 0, 5, -4,
    -- filter=2 channel=102
    -1, 2, -6, 0, 6, -2, 5, 7, 2,
    -- filter=2 channel=103
    -3, 4, -2, -8, -6, -7, 9, 6, 14,
    -- filter=2 channel=104
    1, -13, -5, -4, 3, -1, 7, 1, 1,
    -- filter=2 channel=105
    3, 4, 0, 2, 7, 9, -1, 7, 5,
    -- filter=2 channel=106
    4, 6, 3, 6, 3, 0, 7, -5, -3,
    -- filter=2 channel=107
    0, -10, 5, -1, 8, 3, -8, -1, -3,
    -- filter=2 channel=108
    1, 9, 1, 9, 2, 0, 7, 7, -2,
    -- filter=2 channel=109
    -8, -13, -14, -10, 19, 11, 9, 9, -2,
    -- filter=2 channel=110
    7, -6, -9, -8, 1, 2, 2, 9, 8,
    -- filter=2 channel=111
    5, 0, 0, -4, -2, -5, 2, -1, -1,
    -- filter=2 channel=112
    2, 0, -7, -8, 8, -6, -3, -6, -4,
    -- filter=2 channel=113
    -5, -16, -20, -11, -11, -7, 0, 1, -1,
    -- filter=2 channel=114
    -14, -18, 8, 10, 24, 21, 16, 3, -8,
    -- filter=2 channel=115
    5, 4, 0, 3, -5, -6, -2, 7, 2,
    -- filter=2 channel=116
    -13, -16, -6, 2, 11, 14, 9, -6, 5,
    -- filter=2 channel=117
    -5, -1, -4, -5, -3, -2, 0, 1, 0,
    -- filter=2 channel=118
    5, -5, 5, 6, -6, 7, -3, -4, -7,
    -- filter=2 channel=119
    -5, 0, -4, -1, 6, -1, 5, -10, -1,
    -- filter=2 channel=120
    -23, -19, 4, 5, 30, 17, 0, 6, 0,
    -- filter=2 channel=121
    -1, -12, -6, -11, -4, 6, 4, 2, 3,
    -- filter=2 channel=122
    -6, -1, -16, -1, -13, -10, 1, 4, 3,
    -- filter=2 channel=123
    -4, -8, -6, -9, 0, -7, -3, 0, 2,
    -- filter=2 channel=124
    -4, 5, 7, -5, 0, 3, 3, 5, 4,
    -- filter=2 channel=125
    0, -7, -7, -3, 2, 1, 2, 4, -3,
    -- filter=2 channel=126
    5, -14, -2, -12, -12, 9, -2, 14, 4,
    -- filter=2 channel=127
    7, -6, 3, 1, 4, 0, 4, -3, -2,
    -- filter=3 channel=0
    0, -4, 2, 4, -2, -13, 8, 13, 8,
    -- filter=3 channel=1
    1, 2, -1, 7, -7, -3, 1, 11, 0,
    -- filter=3 channel=2
    -4, 1, 0, 7, 10, 0, -5, 6, 0,
    -- filter=3 channel=3
    10, 14, 3, 4, -3, 1, 8, 8, 0,
    -- filter=3 channel=4
    11, 10, 8, 11, 20, -3, -8, -7, -6,
    -- filter=3 channel=5
    4, 4, 3, -5, -15, -7, 8, -2, -3,
    -- filter=3 channel=6
    2, -4, 2, 0, -2, 0, 7, -3, -5,
    -- filter=3 channel=7
    2, -3, 7, -1, 1, -5, 0, 2, -6,
    -- filter=3 channel=8
    7, -7, 0, -2, 5, -1, -5, 6, 0,
    -- filter=3 channel=9
    -7, -2, -6, -1, 2, 0, 0, -6, 5,
    -- filter=3 channel=10
    3, 11, 9, -1, -4, 1, -2, -2, -1,
    -- filter=3 channel=11
    -6, -3, 7, -4, -1, 2, -3, -1, -2,
    -- filter=3 channel=12
    6, 2, 0, -2, -8, -9, 4, 1, 5,
    -- filter=3 channel=13
    2, 7, 7, 2, -3, -4, 0, 1, -5,
    -- filter=3 channel=14
    -4, 5, 0, -3, 0, -2, 6, 2, -7,
    -- filter=3 channel=15
    -6, 9, -3, -2, -1, 1, 7, 5, -7,
    -- filter=3 channel=16
    -2, 3, 2, -2, -12, -2, 8, 3, -3,
    -- filter=3 channel=17
    0, 1, 3, 1, 1, 5, -4, -1, 3,
    -- filter=3 channel=18
    -9, 0, -3, 6, -8, -4, 5, 2, -7,
    -- filter=3 channel=19
    -5, 0, -2, 0, 6, 1, 6, -6, -6,
    -- filter=3 channel=20
    2, 1, 7, 1, -2, -4, -2, -6, 5,
    -- filter=3 channel=21
    1, -4, 1, -3, 0, 3, 0, 1, -2,
    -- filter=3 channel=22
    3, 1, 1, 6, -9, 2, -1, 10, 3,
    -- filter=3 channel=23
    3, 19, 11, -12, -6, 1, 7, 11, 5,
    -- filter=3 channel=24
    7, 0, -3, -6, 3, -2, 1, 7, -6,
    -- filter=3 channel=25
    -7, 4, 3, -7, -15, -11, 7, 8, -4,
    -- filter=3 channel=26
    4, -10, 2, -1, 5, -6, -2, 1, -7,
    -- filter=3 channel=27
    -3, 3, -3, -6, -19, -13, 0, -2, 6,
    -- filter=3 channel=28
    2, 5, 5, -1, -4, -5, 2, -1, 2,
    -- filter=3 channel=29
    -1, -4, -4, -4, 0, -1, -8, 4, -2,
    -- filter=3 channel=30
    0, 4, 7, 4, -8, -2, -2, 9, 3,
    -- filter=3 channel=31
    6, 12, 10, -14, -13, 4, 2, -4, 4,
    -- filter=3 channel=32
    -7, 9, 0, 0, -11, -1, 8, -1, 4,
    -- filter=3 channel=33
    6, 2, 11, 0, -17, -9, 0, 13, -3,
    -- filter=3 channel=34
    3, 6, -6, -1, 0, 4, 2, -6, -4,
    -- filter=3 channel=35
    1, 5, 0, -3, 5, -6, -1, -6, -2,
    -- filter=3 channel=36
    3, 3, 4, 6, -4, 0, 5, 0, 4,
    -- filter=3 channel=37
    5, 0, -1, 1, 3, -5, -3, 4, 6,
    -- filter=3 channel=38
    -5, 8, 0, 0, -4, 1, -2, 4, -2,
    -- filter=3 channel=39
    -2, -1, -3, -2, -6, -2, -7, 5, -3,
    -- filter=3 channel=40
    4, 10, -1, 1, -4, 1, 0, -1, 4,
    -- filter=3 channel=41
    1, -10, -2, 10, -2, 1, 3, 5, 3,
    -- filter=3 channel=42
    0, 5, -5, -3, -2, 0, 5, 0, 3,
    -- filter=3 channel=43
    -3, 0, 9, 1, -6, 3, 1, 12, 5,
    -- filter=3 channel=44
    -3, 1, 1, -3, 0, -5, 10, 2, 7,
    -- filter=3 channel=45
    2, -5, -5, -5, 3, 3, -5, 4, 5,
    -- filter=3 channel=46
    -5, 1, 0, 3, -1, 4, 1, -4, 2,
    -- filter=3 channel=47
    -1, 3, -4, -7, -7, -10, 10, 4, -3,
    -- filter=3 channel=48
    5, -5, 5, -7, -6, -6, 6, 0, 4,
    -- filter=3 channel=49
    -6, 3, -2, -1, 5, 0, -1, -3, -5,
    -- filter=3 channel=50
    -4, 9, 6, -6, -6, 1, -3, 1, -5,
    -- filter=3 channel=51
    0, 0, 3, 3, -5, 1, -6, 1, 0,
    -- filter=3 channel=52
    -4, -3, -5, 0, 7, 5, 11, 7, 0,
    -- filter=3 channel=53
    0, 0, -1, -4, -2, 0, 2, 0, -6,
    -- filter=3 channel=54
    0, 2, 6, 5, 0, -3, -5, -2, -1,
    -- filter=3 channel=55
    -8, 1, 2, -6, -8, -4, 5, -4, -3,
    -- filter=3 channel=56
    -7, -4, -2, -1, 5, 5, 5, 4, 0,
    -- filter=3 channel=57
    0, 3, -5, 6, 9, -1, -2, -6, -6,
    -- filter=3 channel=58
    2, -6, 4, 6, 2, -3, -5, 0, 6,
    -- filter=3 channel=59
    0, -2, 2, 2, -1, -6, 0, 4, 0,
    -- filter=3 channel=60
    5, 0, 0, 3, -4, -1, 4, 2, -7,
    -- filter=3 channel=61
    0, 2, -4, 0, -1, 0, 0, 0, 3,
    -- filter=3 channel=62
    1, -1, -1, -6, 7, 0, -3, 2, 3,
    -- filter=3 channel=63
    -2, 0, 2, 5, -5, -4, -6, 2, -7,
    -- filter=3 channel=64
    -6, -2, -3, 2, -2, 3, 5, 2, -4,
    -- filter=3 channel=65
    4, -2, -5, -4, -6, -4, 0, -4, 7,
    -- filter=3 channel=66
    0, -9, -7, 9, -2, 2, 7, 9, 3,
    -- filter=3 channel=67
    4, 1, -4, 6, 3, 5, -1, 5, 6,
    -- filter=3 channel=68
    -6, -4, 5, -1, -2, 6, -5, 2, -4,
    -- filter=3 channel=69
    0, -5, -8, 1, 5, -2, 1, 8, 4,
    -- filter=3 channel=70
    4, 5, 5, 4, 0, -3, 9, -3, -4,
    -- filter=3 channel=71
    0, 8, 4, 2, 4, -1, 2, 5, -3,
    -- filter=3 channel=72
    -2, 9, 2, -8, -5, -8, 0, -3, 0,
    -- filter=3 channel=73
    3, 3, -4, 0, 4, -2, -6, -2, 2,
    -- filter=3 channel=74
    8, 2, -4, 2, 5, 5, 9, 1, 4,
    -- filter=3 channel=75
    4, -2, -5, -3, -12, -15, 3, 13, -2,
    -- filter=3 channel=76
    -8, 1, -2, 7, 5, 4, 4, -5, -7,
    -- filter=3 channel=77
    2, 3, -5, 2, 1, 5, -4, 1, -2,
    -- filter=3 channel=78
    -3, -5, -1, -6, 4, -2, 0, -2, -1,
    -- filter=3 channel=79
    -5, 11, 0, -6, -8, -9, -1, 15, -6,
    -- filter=3 channel=80
    0, 10, -2, -8, -20, -7, 2, -3, -1,
    -- filter=3 channel=81
    5, 1, 0, -2, -3, 2, -7, 2, -2,
    -- filter=3 channel=82
    1, 8, -4, 6, -2, 1, -2, -1, 0,
    -- filter=3 channel=83
    -6, -7, 4, -4, 6, -1, 5, -4, 1,
    -- filter=3 channel=84
    -3, -6, 3, 4, -3, 3, -3, -2, 0,
    -- filter=3 channel=85
    5, -7, -5, 6, -2, 4, 1, -5, 1,
    -- filter=3 channel=86
    7, 3, -9, 1, 5, 0, -4, 8, 2,
    -- filter=3 channel=87
    1, 0, 0, 7, -5, -2, 7, 4, 1,
    -- filter=3 channel=88
    -5, -4, -1, -4, 2, 7, 5, -7, 4,
    -- filter=3 channel=89
    1, 0, 8, -6, -7, -9, 1, 3, -1,
    -- filter=3 channel=90
    1, 2, 2, 6, -2, 0, -1, 1, -4,
    -- filter=3 channel=91
    -7, 3, -1, -3, -2, -5, 3, 0, 3,
    -- filter=3 channel=92
    7, -3, -2, -3, -5, 1, 9, 0, 3,
    -- filter=3 channel=93
    4, 0, -9, 2, -10, 2, 4, 2, -4,
    -- filter=3 channel=94
    4, 7, -7, -4, 4, -6, -6, 3, -4,
    -- filter=3 channel=95
    -6, -1, -3, -4, 0, 0, -5, 8, -5,
    -- filter=3 channel=96
    6, 1, -5, 0, 2, -7, 6, -1, 0,
    -- filter=3 channel=97
    3, 2, 5, 6, -6, 2, 7, 10, -5,
    -- filter=3 channel=98
    5, 8, 3, -12, -19, 0, -5, 8, -2,
    -- filter=3 channel=99
    0, -2, -3, -12, -10, -4, -1, -2, -1,
    -- filter=3 channel=100
    -1, -1, 4, -6, 5, -5, -2, -3, -2,
    -- filter=3 channel=101
    2, 5, 1, 6, 3, 4, -4, -5, 0,
    -- filter=3 channel=102
    -4, -6, -6, -6, 4, -5, 1, 3, -4,
    -- filter=3 channel=103
    7, 3, 9, -9, -10, -4, 4, 7, -3,
    -- filter=3 channel=104
    -8, 0, 7, -9, -11, -1, 4, -4, 0,
    -- filter=3 channel=105
    -7, 6, 5, -3, -2, -4, 4, 1, 0,
    -- filter=3 channel=106
    -1, 7, 5, 5, 7, 4, -3, 1, -2,
    -- filter=3 channel=107
    -3, 3, -1, -2, 8, -2, 5, 9, -6,
    -- filter=3 channel=108
    -4, -1, -6, -3, -7, 2, -1, 9, 3,
    -- filter=3 channel=109
    -4, -5, 1, -4, -1, -7, 1, 5, 0,
    -- filter=3 channel=110
    -5, -2, 1, -2, -2, 6, -5, -4, 5,
    -- filter=3 channel=111
    -2, 5, -2, 0, 4, -1, 3, -1, 3,
    -- filter=3 channel=112
    5, 4, 6, -3, -2, -6, 5, 8, 3,
    -- filter=3 channel=113
    0, 1, 2, 0, -7, 3, 10, 11, 0,
    -- filter=3 channel=114
    3, -9, -10, 6, -4, -5, 2, 0, -5,
    -- filter=3 channel=115
    2, -7, -7, 0, 4, -5, -6, -5, 2,
    -- filter=3 channel=116
    -3, 1, -4, -6, -10, 1, -8, -2, -7,
    -- filter=3 channel=117
    1, -5, 1, -1, 3, 0, -3, -6, -1,
    -- filter=3 channel=118
    2, -6, 0, 4, 0, -6, -3, -1, 7,
    -- filter=3 channel=119
    4, -6, 3, 2, -6, -1, 4, 4, 2,
    -- filter=3 channel=120
    6, -7, -6, -3, -11, 0, 6, 0, -7,
    -- filter=3 channel=121
    0, 2, 8, -4, -10, -3, -4, 9, 5,
    -- filter=3 channel=122
    0, -4, 0, -2, -6, -2, 8, 7, 1,
    -- filter=3 channel=123
    0, 3, 8, -6, 6, 2, 9, 0, 0,
    -- filter=3 channel=124
    -5, 2, 7, -4, -6, 7, 5, 0, -7,
    -- filter=3 channel=125
    4, 6, 4, 0, -2, -9, -3, 4, -5,
    -- filter=3 channel=126
    5, 6, 3, 1, -13, -7, 9, 10, 5,
    -- filter=3 channel=127
    -5, -4, -2, -6, 6, 0, 5, 1, 1,
    -- filter=4 channel=0
    -1, -6, -24, 11, -23, -30, 0, -13, -13,
    -- filter=4 channel=1
    0, -5, -20, -2, -10, -20, -4, -6, -4,
    -- filter=4 channel=2
    5, -3, 7, -2, -3, 6, 1, 3, -2,
    -- filter=4 channel=3
    6, -1, -2, 4, 0, -11, 12, 11, 6,
    -- filter=4 channel=4
    1, 4, -7, 9, 0, -5, 5, 0, -3,
    -- filter=4 channel=5
    0, -9, -10, 1, -15, -12, 0, -10, -8,
    -- filter=4 channel=6
    5, 0, -8, -7, 0, 0, 2, -3, -11,
    -- filter=4 channel=7
    0, -6, 2, 2, -2, -6, -5, 4, -2,
    -- filter=4 channel=8
    2, -1, 1, 7, -1, -3, 5, 5, 3,
    -- filter=4 channel=9
    0, 0, -8, 2, -5, 4, 2, 3, 0,
    -- filter=4 channel=10
    0, 0, 13, -2, 1, 17, -10, 3, -5,
    -- filter=4 channel=11
    5, 5, -4, 5, -1, -5, 0, 2, -2,
    -- filter=4 channel=12
    0, 4, 2, 6, 2, 13, -3, 3, 0,
    -- filter=4 channel=13
    2, 2, 3, 5, 2, 8, -4, 0, -5,
    -- filter=4 channel=14
    6, 0, 5, -6, -2, 1, 0, -3, -1,
    -- filter=4 channel=15
    0, 2, -14, 3, 2, -16, -1, 1, -14,
    -- filter=4 channel=16
    -4, -2, 16, -7, -3, 13, 0, 6, 10,
    -- filter=4 channel=17
    3, 7, -7, 5, 0, 2, 4, -7, 2,
    -- filter=4 channel=18
    -3, -6, -18, 9, -12, -20, 7, 0, -15,
    -- filter=4 channel=19
    2, -1, -1, 3, -7, -6, 2, -3, 2,
    -- filter=4 channel=20
    5, 6, 0, 0, -3, -2, -8, -3, -13,
    -- filter=4 channel=21
    -8, 3, 20, -12, 13, 15, -5, -1, 10,
    -- filter=4 channel=22
    8, -6, -5, 7, -10, -13, -1, -1, -9,
    -- filter=4 channel=23
    9, 0, -9, 8, 7, -6, 0, -10, -7,
    -- filter=4 channel=24
    -6, 2, -1, -6, -2, -4, 1, 2, -6,
    -- filter=4 channel=25
    -7, -7, -2, 8, -4, -6, 0, 4, 1,
    -- filter=4 channel=26
    5, -4, -2, 4, -5, 12, -5, 0, 2,
    -- filter=4 channel=27
    8, -6, -17, 4, -16, -26, 1, -17, -19,
    -- filter=4 channel=28
    -2, 0, 4, -3, 6, 6, -4, -5, 6,
    -- filter=4 channel=29
    -3, 12, 5, 3, 7, -6, -8, -4, -6,
    -- filter=4 channel=30
    4, -3, -8, 7, -5, -9, 5, -8, -2,
    -- filter=4 channel=31
    -6, -5, 16, 0, 8, 16, -7, -7, 13,
    -- filter=4 channel=32
    3, -7, -7, 6, -10, -15, 5, 0, -8,
    -- filter=4 channel=33
    -1, -8, -8, 5, -2, -9, 9, -6, -14,
    -- filter=4 channel=34
    4, -4, 10, 4, 5, -1, 11, 1, 8,
    -- filter=4 channel=35
    -4, 1, 4, -7, -1, 3, 4, -7, 4,
    -- filter=4 channel=36
    -1, 3, 21, -8, 12, 16, -1, 6, 9,
    -- filter=4 channel=37
    10, 2, -15, -3, -8, -22, 2, -7, -13,
    -- filter=4 channel=38
    3, -8, -3, 3, -8, 0, 5, -10, 5,
    -- filter=4 channel=39
    0, 2, 2, 2, 0, -7, -8, 0, 0,
    -- filter=4 channel=40
    -1, -1, 3, 3, -3, -5, 4, -8, -3,
    -- filter=4 channel=41
    7, 11, 4, 15, 11, 2, 1, 15, 11,
    -- filter=4 channel=42
    3, -2, 0, 1, -7, -9, 7, -7, -5,
    -- filter=4 channel=43
    7, -7, -15, 4, 0, -15, 9, 5, -9,
    -- filter=4 channel=44
    -5, -8, -6, -6, -9, -6, 0, -6, 6,
    -- filter=4 channel=45
    -8, 4, 0, -5, 0, 1, 0, 4, -10,
    -- filter=4 channel=46
    0, -4, 5, -4, -6, 4, -3, 0, -5,
    -- filter=4 channel=47
    -11, -10, 7, -4, -7, 13, -2, -3, 8,
    -- filter=4 channel=48
    0, -6, -4, -4, -8, -1, 1, 0, -4,
    -- filter=4 channel=49
    -2, -4, -8, 1, -1, -19, -2, -6, -16,
    -- filter=4 channel=50
    4, -5, -5, 4, 4, -8, 0, -3, -5,
    -- filter=4 channel=51
    5, -6, -1, -3, -4, 0, -1, -6, 2,
    -- filter=4 channel=52
    10, 3, 10, 8, 6, -4, 5, -8, 9,
    -- filter=4 channel=53
    6, -2, 7, 0, 0, 6, 3, 1, 0,
    -- filter=4 channel=54
    -4, 6, 6, 6, 4, 2, 5, 3, 0,
    -- filter=4 channel=55
    0, 2, 0, 0, 10, 4, -1, 3, -5,
    -- filter=4 channel=56
    5, -6, 6, 8, -7, 4, 0, -2, 7,
    -- filter=4 channel=57
    4, 9, -4, -2, -3, 0, -2, 3, -2,
    -- filter=4 channel=58
    4, 1, -9, 8, 0, -7, 2, -8, -7,
    -- filter=4 channel=59
    1, 2, 5, -3, 1, 12, -5, -2, 6,
    -- filter=4 channel=60
    0, -3, 1, 6, -1, -2, 3, 2, -2,
    -- filter=4 channel=61
    1, 4, 5, -4, 0, 9, -4, 5, 8,
    -- filter=4 channel=62
    1, -1, -5, -6, 0, 3, 8, -1, 0,
    -- filter=4 channel=63
    -6, -1, 0, -6, 3, -4, -3, -4, 6,
    -- filter=4 channel=64
    4, -2, 10, 1, 0, 4, -4, 0, 6,
    -- filter=4 channel=65
    -6, -1, 5, 3, 4, 0, -3, -5, 5,
    -- filter=4 channel=66
    5, 13, 4, -3, 0, 7, -8, 8, 16,
    -- filter=4 channel=67
    -2, -5, 6, 2, 3, 5, 3, -5, 7,
    -- filter=4 channel=68
    -1, 3, -1, -2, 0, -4, -2, 7, 6,
    -- filter=4 channel=69
    6, 6, 1, -5, -1, 8, -2, 0, -2,
    -- filter=4 channel=70
    2, -6, -15, 10, -10, -15, 12, -11, -14,
    -- filter=4 channel=71
    -2, 3, -1, 9, 6, 4, -1, 9, 6,
    -- filter=4 channel=72
    0, 5, 12, 0, 17, 10, 1, -3, 1,
    -- filter=4 channel=73
    9, 5, 1, 10, 4, -1, 8, -4, -8,
    -- filter=4 channel=74
    -7, 1, 6, -3, -6, -6, 0, 0, -1,
    -- filter=4 channel=75
    1, -2, -14, 4, -13, -21, 0, -1, -10,
    -- filter=4 channel=76
    1, 6, 8, 6, 6, 6, -6, -2, -4,
    -- filter=4 channel=77
    -5, -7, 5, -3, 0, -3, 6, 0, -1,
    -- filter=4 channel=78
    -4, -1, 4, -1, -7, 0, 2, -7, -4,
    -- filter=4 channel=79
    1, 0, -17, 12, -10, -32, 3, -7, -16,
    -- filter=4 channel=80
    -2, -7, 17, -1, 2, 20, -9, 4, 4,
    -- filter=4 channel=81
    -2, -3, -3, -5, 0, -1, -2, -1, -5,
    -- filter=4 channel=82
    1, 0, -6, -1, 0, 2, 2, 3, -6,
    -- filter=4 channel=83
    -3, 4, 0, -6, 0, 4, -2, -1, -6,
    -- filter=4 channel=84
    5, 0, -7, 8, 0, -15, 0, -1, -13,
    -- filter=4 channel=85
    -5, 1, 4, 0, 6, 2, 3, -4, 1,
    -- filter=4 channel=86
    -3, -4, -8, -1, -1, 3, 5, 2, 5,
    -- filter=4 channel=87
    -3, -2, 0, -3, -5, -3, 6, -7, -3,
    -- filter=4 channel=88
    0, -1, 7, 2, 7, 16, 3, 1, 11,
    -- filter=4 channel=89
    1, 2, 8, -1, 15, 0, -4, 10, -5,
    -- filter=4 channel=90
    1, -1, 8, 5, 12, 10, -1, -4, 5,
    -- filter=4 channel=91
    -2, -2, -12, 0, -8, -12, 6, 2, -3,
    -- filter=4 channel=92
    -1, 3, 2, 5, -6, 2, 4, 3, -3,
    -- filter=4 channel=93
    -5, -5, 3, -2, -6, -2, 0, -14, -4,
    -- filter=4 channel=94
    4, 2, 2, 2, -4, -2, 2, -6, -5,
    -- filter=4 channel=95
    2, -3, 3, 0, 4, -4, 0, 7, -1,
    -- filter=4 channel=96
    -5, 1, 4, 3, 0, 1, 6, -5, -8,
    -- filter=4 channel=97
    6, 1, 7, 9, 6, -5, 8, 1, 2,
    -- filter=4 channel=98
    6, -1, 1, -2, 5, -2, 4, 0, -6,
    -- filter=4 channel=99
    -4, 4, 15, -4, 12, 14, -12, 1, 10,
    -- filter=4 channel=100
    1, 0, 3, -2, 5, 4, -6, 5, 0,
    -- filter=4 channel=101
    0, 9, 7, -3, -3, -7, -2, 7, 1,
    -- filter=4 channel=102
    2, 5, 0, -1, -7, 5, 2, 1, 3,
    -- filter=4 channel=103
    -10, -9, 2, 0, -4, 16, 0, 0, 8,
    -- filter=4 channel=104
    -7, 2, 14, -1, 0, 23, -3, -8, 11,
    -- filter=4 channel=105
    -8, -4, -10, 0, 0, -6, 6, 4, -11,
    -- filter=4 channel=106
    0, 2, -2, 2, 1, -3, -3, -2, -7,
    -- filter=4 channel=107
    -7, -10, -8, 6, -3, -19, 1, -4, -18,
    -- filter=4 channel=108
    6, 0, 0, 0, -6, -6, -4, 6, -6,
    -- filter=4 channel=109
    8, -5, -2, 0, -7, -7, -1, -5, -11,
    -- filter=4 channel=110
    3, 10, 15, 0, 14, 11, -3, 3, 1,
    -- filter=4 channel=111
    -2, -2, 7, 5, 1, 8, -6, -2, 8,
    -- filter=4 channel=112
    5, -12, -5, 7, -5, -13, 3, -5, -4,
    -- filter=4 channel=113
    0, -7, -3, 6, 3, 0, -3, 0, 6,
    -- filter=4 channel=114
    -1, -19, -21, 13, -27, -41, 8, -11, -21,
    -- filter=4 channel=115
    2, -2, 5, -1, 7, 4, 6, 2, -2,
    -- filter=4 channel=116
    1, -3, 0, 5, -4, -3, 3, -7, -6,
    -- filter=4 channel=117
    -4, 1, -3, -6, -1, -3, -5, 7, 2,
    -- filter=4 channel=118
    -5, 0, 2, 0, -3, -6, -5, -4, 2,
    -- filter=4 channel=119
    2, -2, -1, 0, -6, 0, 2, -3, 12,
    -- filter=4 channel=120
    9, 0, -10, -1, -6, -17, 9, -15, -7,
    -- filter=4 channel=121
    5, -2, 13, 7, 7, 10, -2, 0, 1,
    -- filter=4 channel=122
    -10, 5, 25, 0, 0, 38, -15, 1, 17,
    -- filter=4 channel=123
    5, -4, 4, 0, 6, -2, 0, -3, 9,
    -- filter=4 channel=124
    -3, 2, -5, 6, 0, -6, -2, 2, -8,
    -- filter=4 channel=125
    -3, -5, 6, -1, 6, 10, -7, -9, -3,
    -- filter=4 channel=126
    2, 1, 1, 0, 5, -4, 7, 4, -3,
    -- filter=4 channel=127
    0, -2, 8, 7, -2, 8, 8, 8, 7,
    -- filter=5 channel=0
    0, -1, -8, -1, 2, 1, 4, -1, 0,
    -- filter=5 channel=1
    -6, -6, -7, -2, -6, -1, -5, -10, -1,
    -- filter=5 channel=2
    5, -5, -1, 4, 2, -1, -4, 3, 4,
    -- filter=5 channel=3
    -9, -7, 4, -2, 1, -1, -7, -1, 5,
    -- filter=5 channel=4
    -3, 0, 1, 0, -6, 9, -8, -6, -5,
    -- filter=5 channel=5
    -6, 4, -5, -5, 0, -4, 5, -2, 5,
    -- filter=5 channel=6
    -3, 0, -1, 6, -1, 4, 0, 1, -3,
    -- filter=5 channel=7
    -3, 5, 2, -1, 0, 4, -1, 0, 4,
    -- filter=5 channel=8
    0, -2, -4, -4, -4, -10, -3, 4, -9,
    -- filter=5 channel=9
    5, 6, -7, 2, -2, 0, 7, 0, 2,
    -- filter=5 channel=10
    0, 1, 1, -6, 8, 3, -4, -2, 5,
    -- filter=5 channel=11
    -1, 0, 4, 4, 6, -7, 5, -5, 4,
    -- filter=5 channel=12
    -6, 1, 0, -8, -9, -3, -6, -7, -9,
    -- filter=5 channel=13
    -3, -10, -6, -7, 1, 8, -7, -10, 0,
    -- filter=5 channel=14
    -5, 7, 1, 1, 1, 7, 1, -2, -5,
    -- filter=5 channel=15
    6, 0, -8, 0, 8, -12, 4, 6, -4,
    -- filter=5 channel=16
    0, -4, -5, -3, 3, -7, 0, 3, 1,
    -- filter=5 channel=17
    5, -4, -5, -3, -5, 2, -2, 5, 6,
    -- filter=5 channel=18
    12, -5, -8, 6, 9, -3, 0, 2, 9,
    -- filter=5 channel=19
    6, 3, 0, 3, -5, -4, 0, 5, -1,
    -- filter=5 channel=20
    4, -5, -9, -7, -5, 2, 2, 0, -6,
    -- filter=5 channel=21
    -10, 2, -4, -6, 4, -6, 2, 0, 2,
    -- filter=5 channel=22
    1, -2, -4, 0, 7, -11, 4, 3, -5,
    -- filter=5 channel=23
    5, -10, -20, 4, 14, -10, 4, 11, -8,
    -- filter=5 channel=24
    1, 6, -2, -6, 7, -6, -4, -6, 4,
    -- filter=5 channel=25
    10, 3, -3, -4, 3, 0, -8, -8, 10,
    -- filter=5 channel=26
    1, 1, 0, -1, -4, -1, -4, 3, 7,
    -- filter=5 channel=27
    0, -3, -16, -2, 16, -7, -7, 13, 4,
    -- filter=5 channel=28
    4, 4, 5, -4, -6, -6, 5, -4, -1,
    -- filter=5 channel=29
    -3, 0, 2, 6, 8, -2, -7, -5, -6,
    -- filter=5 channel=30
    -1, -4, -4, -2, 0, -6, -3, 6, 3,
    -- filter=5 channel=31
    -7, -2, -1, -6, 6, -7, -1, 7, 7,
    -- filter=5 channel=32
    11, -9, -3, 8, 4, 0, -4, -4, 7,
    -- filter=5 channel=33
    0, -4, -14, 10, 10, -2, 7, 6, 1,
    -- filter=5 channel=34
    -3, -8, -9, 0, -7, 0, 3, 7, -3,
    -- filter=5 channel=35
    4, 5, 0, 6, 7, -5, 6, -1, 0,
    -- filter=5 channel=36
    -5, -7, -1, -1, -9, 0, -1, -4, -3,
    -- filter=5 channel=37
    -3, -5, -8, -11, -9, 0, -3, -9, -5,
    -- filter=5 channel=38
    8, -1, 2, -3, 11, -2, -4, 2, 8,
    -- filter=5 channel=39
    3, 4, -5, 2, 1, 5, -4, -6, 0,
    -- filter=5 channel=40
    -1, -8, -8, -6, -5, -10, 0, 0, -4,
    -- filter=5 channel=41
    -1, -1, 11, 5, -3, 5, -8, -3, 6,
    -- filter=5 channel=42
    2, 0, 7, 0, -4, 0, 4, 0, 9,
    -- filter=5 channel=43
    3, -9, 0, -5, -1, -1, 3, 3, -2,
    -- filter=5 channel=44
    -1, -2, 2, -7, -8, -5, -1, 6, 3,
    -- filter=5 channel=45
    -2, 5, -6, 0, 2, -2, 3, -3, -2,
    -- filter=5 channel=46
    4, -3, -7, 5, -7, 6, 2, 3, 2,
    -- filter=5 channel=47
    -8, -9, -7, -7, 1, 5, -3, 0, 2,
    -- filter=5 channel=48
    -3, -1, -7, -4, 0, 0, -6, -4, 4,
    -- filter=5 channel=49
    -2, 1, -1, 0, 1, 7, -6, 6, 0,
    -- filter=5 channel=50
    8, -2, 0, 6, 8, -3, -8, 10, -6,
    -- filter=5 channel=51
    -4, -5, -1, 0, -4, 6, -2, 6, 3,
    -- filter=5 channel=52
    4, -4, -1, -2, 2, -7, 4, -7, 0,
    -- filter=5 channel=53
    5, -3, 1, -4, 6, 0, 2, -4, 0,
    -- filter=5 channel=54
    -1, -5, 0, 0, -1, -2, -7, 0, 6,
    -- filter=5 channel=55
    12, 1, -2, 8, 2, -10, 4, 0, -7,
    -- filter=5 channel=56
    -2, -5, -9, -1, -3, -7, 3, 5, -3,
    -- filter=5 channel=57
    -5, 1, 7, -5, 6, 5, 0, 3, 3,
    -- filter=5 channel=58
    5, 7, -2, 0, 0, 7, 1, 0, 0,
    -- filter=5 channel=59
    1, 5, -7, 5, 1, 11, 5, -7, 6,
    -- filter=5 channel=60
    -1, 1, 1, -6, -7, 4, 7, 6, 0,
    -- filter=5 channel=61
    2, -2, -6, -8, -3, 0, -8, 5, 1,
    -- filter=5 channel=62
    -4, -7, -2, 4, -2, -7, 2, -1, -3,
    -- filter=5 channel=63
    1, 8, 5, 1, 6, 4, 1, 0, 6,
    -- filter=5 channel=64
    -9, -7, -5, -4, 2, -3, 1, 2, -1,
    -- filter=5 channel=65
    7, 2, 1, 7, -2, -5, -1, 6, -6,
    -- filter=5 channel=66
    -4, -2, -4, 3, -12, 6, 5, -2, 7,
    -- filter=5 channel=67
    -6, -2, -5, 1, -2, -5, 7, 4, -6,
    -- filter=5 channel=68
    5, -5, 0, -6, 5, -3, -1, -8, 2,
    -- filter=5 channel=69
    -2, -2, 3, 0, 3, 2, -5, 2, 4,
    -- filter=5 channel=70
    4, -4, -11, 0, 6, -4, 2, 8, -2,
    -- filter=5 channel=71
    -8, -3, 4, -6, 3, -3, 2, -4, -1,
    -- filter=5 channel=72
    5, 1, 0, 2, 2, -5, 5, 3, 0,
    -- filter=5 channel=73
    -2, -1, -5, 9, 3, 0, 1, 4, -5,
    -- filter=5 channel=74
    0, -3, -4, -4, 4, -5, -7, 5, -11,
    -- filter=5 channel=75
    -5, 0, 4, -6, 2, 1, 1, 3, 8,
    -- filter=5 channel=76
    -3, -6, -7, -3, -8, -10, -1, 0, -1,
    -- filter=5 channel=77
    6, -6, -6, 0, -7, -3, -5, -2, 4,
    -- filter=5 channel=78
    -1, -5, -6, 3, -4, -6, 8, 8, -6,
    -- filter=5 channel=79
    14, -9, -20, 7, 2, 1, 2, -3, 8,
    -- filter=5 channel=80
    0, -8, 0, -6, 12, 7, 0, -1, 14,
    -- filter=5 channel=81
    -6, 4, 0, 0, 6, 1, 6, 0, 3,
    -- filter=5 channel=82
    -3, -1, -7, 2, 4, 2, -5, 0, -1,
    -- filter=5 channel=83
    0, -2, -6, 0, 4, -2, 1, -3, 0,
    -- filter=5 channel=84
    5, 0, -12, 0, 8, 0, 4, 0, 2,
    -- filter=5 channel=85
    -6, 1, 6, 3, 0, 7, 0, 3, 0,
    -- filter=5 channel=86
    -6, -10, 2, 0, -7, 1, -1, 1, -1,
    -- filter=5 channel=87
    -4, -5, -6, -5, -7, -12, -7, 4, -11,
    -- filter=5 channel=88
    -2, -8, -8, -4, -7, -10, -4, 6, -7,
    -- filter=5 channel=89
    5, -3, -11, 8, 0, 2, 0, -7, 9,
    -- filter=5 channel=90
    0, 0, -7, -7, -8, -10, -2, 0, -8,
    -- filter=5 channel=91
    0, 2, -6, -3, 5, -8, -3, -1, -3,
    -- filter=5 channel=92
    -2, -1, -6, 5, -1, 3, 5, 1, 0,
    -- filter=5 channel=93
    -10, 3, 5, -11, 0, -6, -3, 2, 6,
    -- filter=5 channel=94
    4, 5, 4, 4, -2, 0, -3, 3, 5,
    -- filter=5 channel=95
    5, 5, -3, -1, -5, -1, -6, 0, -3,
    -- filter=5 channel=96
    2, -5, 2, -2, 1, -5, -5, 1, 0,
    -- filter=5 channel=97
    -8, -2, -7, -5, -7, 2, -6, 5, 5,
    -- filter=5 channel=98
    11, -4, -2, 5, 7, 3, 5, -4, 14,
    -- filter=5 channel=99
    -4, -1, -10, 7, 14, -17, -7, 13, -1,
    -- filter=5 channel=100
    -5, 0, -7, -1, 5, 5, -1, 0, -6,
    -- filter=5 channel=101
    2, 4, 2, -8, 2, -1, -12, 2, 0,
    -- filter=5 channel=102
    -4, 7, 4, 4, 4, 4, 5, 0, 3,
    -- filter=5 channel=103
    1, -8, -1, -11, -2, 7, 1, 7, 10,
    -- filter=5 channel=104
    -8, 7, 2, 0, -1, 0, -8, -3, 2,
    -- filter=5 channel=105
    -1, -7, 3, 4, -3, -6, 3, 0, 3,
    -- filter=5 channel=106
    0, 0, 0, 1, -6, 1, 1, -1, 2,
    -- filter=5 channel=107
    5, -4, 1, 2, 0, -13, -7, 8, 2,
    -- filter=5 channel=108
    -2, -5, 6, 0, 2, 6, -1, -2, 0,
    -- filter=5 channel=109
    5, -6, -3, 8, 9, -6, -3, 4, -1,
    -- filter=5 channel=110
    2, -6, -3, 2, 3, -5, -1, 0, 3,
    -- filter=5 channel=111
    3, 7, 0, -6, -7, -5, -5, 1, -2,
    -- filter=5 channel=112
    -4, -8, -7, 1, 4, -1, -3, 11, 0,
    -- filter=5 channel=113
    0, 0, -2, 2, 2, -1, 8, -2, 0,
    -- filter=5 channel=114
    11, 3, -16, 7, 3, -2, 3, 0, -2,
    -- filter=5 channel=115
    3, 6, 4, -6, 7, -3, -4, -4, 6,
    -- filter=5 channel=116
    9, 5, 2, 3, 3, 3, -6, 5, 12,
    -- filter=5 channel=117
    -2, 5, -1, 1, 0, 0, -6, -8, 2,
    -- filter=5 channel=118
    -2, -4, -2, 5, -3, 3, -1, -2, -5,
    -- filter=5 channel=119
    -8, 3, -9, -2, -7, -11, 4, 9, -1,
    -- filter=5 channel=120
    1, -4, -11, 1, 8, -13, -1, 16, -4,
    -- filter=5 channel=121
    0, -8, 0, -5, -8, -2, 8, -9, -3,
    -- filter=5 channel=122
    -19, -5, -7, -14, -3, -10, -14, 4, -2,
    -- filter=5 channel=123
    -5, -1, -5, -3, -1, 3, -1, 3, -9,
    -- filter=5 channel=124
    3, -4, -5, -2, 1, -4, 6, -4, 0,
    -- filter=5 channel=125
    -5, 2, -9, 5, 10, 4, 1, 3, 0,
    -- filter=5 channel=126
    3, 0, 4, 5, 7, 4, 4, 0, 2,
    -- filter=5 channel=127
    -5, -7, 7, -1, 1, 5, -5, 1, -3,
    -- filter=6 channel=0
    6, -5, 0, -2, 5, 8, 9, 7, 3,
    -- filter=6 channel=1
    -6, -1, 3, 3, -12, 2, -3, -4, -3,
    -- filter=6 channel=2
    3, -4, 0, 6, -7, -3, -6, -1, 0,
    -- filter=6 channel=3
    5, 11, 1, 6, 1, 10, -2, 0, 7,
    -- filter=6 channel=4
    -1, 3, 0, -3, -8, -5, 1, -3, -10,
    -- filter=6 channel=5
    2, -1, 5, 9, 0, 12, 4, 11, 2,
    -- filter=6 channel=6
    2, 7, -5, -3, 6, 5, 2, 6, -3,
    -- filter=6 channel=7
    -3, -5, 2, 5, 5, 4, 6, -2, -2,
    -- filter=6 channel=8
    -3, 2, 7, 0, -6, -1, -7, -8, -7,
    -- filter=6 channel=9
    -8, -1, 9, -1, 1, -2, 2, 5, -2,
    -- filter=6 channel=10
    2, 7, 14, -8, -5, 8, -8, -10, 0,
    -- filter=6 channel=11
    -2, 4, 5, 5, 7, 7, 1, -6, -1,
    -- filter=6 channel=12
    -6, 0, -6, -3, -7, -7, -3, -5, -6,
    -- filter=6 channel=13
    -11, -4, 11, -7, -6, -2, -10, -11, 0,
    -- filter=6 channel=14
    2, -1, 6, -6, 3, 0, 0, 0, -1,
    -- filter=6 channel=15
    0, 14, 17, -14, 5, 13, -21, -1, 7,
    -- filter=6 channel=16
    -8, -8, -5, -6, -8, 0, 3, -8, -7,
    -- filter=6 channel=17
    6, -5, -5, 2, -2, 5, 1, 4, 7,
    -- filter=6 channel=18
    -17, 9, 10, -18, -2, 9, -25, -2, 1,
    -- filter=6 channel=19
    -3, -3, 3, 0, -7, 1, 3, 6, -2,
    -- filter=6 channel=20
    0, 14, 7, 0, 11, 14, -10, -1, 4,
    -- filter=6 channel=21
    -13, -9, 5, -4, -1, -1, -4, -4, -3,
    -- filter=6 channel=22
    2, 9, -2, 3, 10, 7, 0, 8, 11,
    -- filter=6 channel=23
    -7, 22, 19, -5, 7, 10, -17, -5, 6,
    -- filter=6 channel=24
    -5, 5, 7, -6, 6, 4, 1, 7, -4,
    -- filter=6 channel=25
    -14, 6, 14, -18, -6, 4, -10, -4, -2,
    -- filter=6 channel=26
    -6, -4, -3, 6, 0, 5, 1, 1, 0,
    -- filter=6 channel=27
    -20, 16, 22, -14, 1, 14, -19, -13, -8,
    -- filter=6 channel=28
    -7, -2, 3, 1, 1, 7, -4, 4, 4,
    -- filter=6 channel=29
    0, 10, 8, -5, 14, 13, -6, -4, 10,
    -- filter=6 channel=30
    -7, 0, 15, -12, -2, 2, -7, -8, 7,
    -- filter=6 channel=31
    -20, 0, 17, -10, 2, 11, -2, -15, -10,
    -- filter=6 channel=32
    -13, 6, 7, -19, 0, 3, -10, -5, 5,
    -- filter=6 channel=33
    -12, 15, 7, -14, 0, 14, -1, -12, 1,
    -- filter=6 channel=34
    -2, 10, 3, -2, 12, 8, 3, 1, 10,
    -- filter=6 channel=35
    2, -6, 3, 0, -3, 2, 1, -7, 4,
    -- filter=6 channel=36
    0, -4, 3, -5, -1, -3, 0, -9, -10,
    -- filter=6 channel=37
    -1, -4, -4, 6, 3, 0, 12, 0, -1,
    -- filter=6 channel=38
    0, 1, 12, -5, -2, 0, 0, 1, 2,
    -- filter=6 channel=39
    4, 1, 0, 0, 6, -1, 2, -4, 4,
    -- filter=6 channel=40
    -2, 0, -2, 2, 2, 1, -1, -3, 1,
    -- filter=6 channel=41
    3, -4, 11, -2, -1, 8, -17, -10, 4,
    -- filter=6 channel=42
    -5, 0, 0, 5, -5, 0, 9, 0, 0,
    -- filter=6 channel=43
    0, 8, -3, -8, 4, 4, -3, 9, 5,
    -- filter=6 channel=44
    -12, 5, 5, -8, -8, -4, 6, -12, -6,
    -- filter=6 channel=45
    -3, 2, 2, -4, 0, 7, 6, 0, 2,
    -- filter=6 channel=46
    0, 0, -1, -3, -1, -6, -1, 1, -2,
    -- filter=6 channel=47
    -14, -12, 3, -4, -15, 4, -2, -1, -14,
    -- filter=6 channel=48
    -10, -4, 5, -8, -9, 1, 2, -9, -10,
    -- filter=6 channel=49
    0, 12, 11, -6, 4, 8, -2, 1, -5,
    -- filter=6 channel=50
    -5, 0, 5, -9, 2, 13, -3, -5, 0,
    -- filter=6 channel=51
    -3, -3, 2, -5, -3, 2, -3, -4, 0,
    -- filter=6 channel=52
    -5, 9, 7, -5, 0, 4, -12, -2, 6,
    -- filter=6 channel=53
    2, 0, 2, -2, 8, -3, -9, 0, -3,
    -- filter=6 channel=54
    3, -3, -3, 3, -3, -4, -4, -2, 5,
    -- filter=6 channel=55
    -18, 8, 13, -10, 10, 11, -21, -15, 0,
    -- filter=6 channel=56
    8, 1, -4, 3, 5, -4, -3, 0, -4,
    -- filter=6 channel=57
    1, -6, 9, 6, 4, 6, -5, 0, -4,
    -- filter=6 channel=58
    0, -5, 8, 10, 7, 0, 6, 2, 10,
    -- filter=6 channel=59
    -18, 2, 15, -9, -9, 7, -10, -16, -2,
    -- filter=6 channel=60
    6, 0, 7, 1, -1, 0, -6, 6, 0,
    -- filter=6 channel=61
    1, 6, -7, -1, -1, 0, -5, 3, -5,
    -- filter=6 channel=62
    -2, -4, 1, 5, 5, 4, 5, -4, 2,
    -- filter=6 channel=63
    -1, -4, -3, 11, 9, 8, 11, 7, 1,
    -- filter=6 channel=64
    -7, -8, 0, 1, 4, 4, 4, -7, 0,
    -- filter=6 channel=65
    -1, -6, 2, 0, 0, 6, -6, -6, -2,
    -- filter=6 channel=66
    0, -5, 6, 0, -3, 6, 0, 5, 2,
    -- filter=6 channel=67
    7, 0, 0, -5, -1, 5, -3, -6, -3,
    -- filter=6 channel=68
    3, -7, -5, 5, -5, -6, -2, 5, 0,
    -- filter=6 channel=69
    4, -6, 3, 8, 6, -2, 5, 4, 5,
    -- filter=6 channel=70
    0, 14, 6, -5, 3, 12, -14, -10, -5,
    -- filter=6 channel=71
    -3, 7, 3, -2, -2, -2, -5, -5, -4,
    -- filter=6 channel=72
    -16, -3, 11, -14, -3, 9, 1, -10, -8,
    -- filter=6 channel=73
    -12, 7, 12, -9, 6, 10, -10, -1, -1,
    -- filter=6 channel=74
    3, 20, 12, -4, 10, 2, -10, -10, 2,
    -- filter=6 channel=75
    0, 0, 5, 3, -7, 10, 0, -3, -2,
    -- filter=6 channel=76
    4, 0, 2, -7, -2, 7, -7, -5, 0,
    -- filter=6 channel=77
    5, -3, -7, 4, -6, 0, 0, 7, -4,
    -- filter=6 channel=78
    -5, 4, -2, 6, 8, 7, 2, 9, 0,
    -- filter=6 channel=79
    -8, 10, 11, -21, 0, 18, -17, -18, 0,
    -- filter=6 channel=80
    -22, -8, 17, -8, -6, 7, -5, -9, -5,
    -- filter=6 channel=81
    5, 4, 6, 0, 1, 5, -3, 7, -1,
    -- filter=6 channel=82
    6, 4, 5, -4, 7, 3, 8, 1, 0,
    -- filter=6 channel=83
    -10, -8, 10, -4, -2, -1, -3, 3, 1,
    -- filter=6 channel=84
    -7, 5, 4, -8, 6, 0, -3, -3, -2,
    -- filter=6 channel=85
    -5, 5, 0, 6, 5, -5, 5, -6, 0,
    -- filter=6 channel=86
    1, 7, 0, -6, 7, 4, -5, 0, 3,
    -- filter=6 channel=87
    5, -1, 4, 5, 7, 0, -4, 0, -4,
    -- filter=6 channel=88
    -5, -5, -4, 3, 0, 0, 0, 5, -1,
    -- filter=6 channel=89
    -8, 0, 13, -16, -5, 3, -13, -15, -3,
    -- filter=6 channel=90
    5, 8, -5, 8, 0, 0, 4, -5, -1,
    -- filter=6 channel=91
    -3, 13, 18, -11, 3, 3, -14, -19, -10,
    -- filter=6 channel=92
    1, 5, 6, 3, -3, 10, -2, -3, 0,
    -- filter=6 channel=93
    0, -4, -2, -6, -11, -9, 4, 0, 0,
    -- filter=6 channel=94
    -6, -5, 0, -3, -3, 3, -3, 0, -2,
    -- filter=6 channel=95
    -4, -6, -1, 5, -4, -1, 3, -5, 0,
    -- filter=6 channel=96
    -6, -4, 4, 3, -8, -1, 0, -4, 5,
    -- filter=6 channel=97
    8, 0, -4, 7, -6, -4, -4, 3, 7,
    -- filter=6 channel=98
    -15, 2, 18, -17, 3, 7, -9, -7, 1,
    -- filter=6 channel=99
    -19, 18, 16, -11, 13, 13, -12, -8, 0,
    -- filter=6 channel=100
    2, -4, -5, 1, 3, -3, 3, -4, -4,
    -- filter=6 channel=101
    -4, -1, 2, -4, -6, 0, -3, -7, -6,
    -- filter=6 channel=102
    2, 1, 5, 0, 0, -1, 7, -3, 3,
    -- filter=6 channel=103
    0, -2, 8, -6, -14, 0, -4, 1, -12,
    -- filter=6 channel=104
    -6, -7, 8, -4, -7, -7, -2, -5, -10,
    -- filter=6 channel=105
    6, 0, 7, 4, 11, 6, -7, 8, 4,
    -- filter=6 channel=106
    3, 4, 5, -4, 4, -3, -4, -2, 4,
    -- filter=6 channel=107
    1, 18, 6, -3, 10, 13, 0, 8, 12,
    -- filter=6 channel=108
    0, 3, 0, 6, -7, -4, 5, 0, 1,
    -- filter=6 channel=109
    -20, 17, 22, -20, 5, 8, -11, -19, -11,
    -- filter=6 channel=110
    -8, 7, 3, 2, 5, -5, 6, -4, 7,
    -- filter=6 channel=111
    2, 4, 6, -2, -6, 7, 4, 7, 3,
    -- filter=6 channel=112
    1, 12, 4, -9, 2, 0, -1, -7, -2,
    -- filter=6 channel=113
    0, 0, 14, -2, 4, 8, -9, -12, -5,
    -- filter=6 channel=114
    -10, 12, 14, -18, 5, 11, -6, -4, 7,
    -- filter=6 channel=115
    -5, 7, -4, -6, -2, -6, 7, -2, 4,
    -- filter=6 channel=116
    -11, 4, 18, -15, -6, 5, -1, -16, -4,
    -- filter=6 channel=117
    -3, 0, -2, 0, 4, -6, 4, -1, 2,
    -- filter=6 channel=118
    1, 2, -5, -1, -2, 0, -1, -1, 1,
    -- filter=6 channel=119
    9, 6, 6, -9, 9, 5, 0, -2, 1,
    -- filter=6 channel=120
    -12, 21, 26, -12, 8, 4, -6, -8, -2,
    -- filter=6 channel=121
    -1, -7, 2, -4, -9, 1, 0, -12, -9,
    -- filter=6 channel=122
    -14, -7, -10, 2, -10, -7, 3, -10, -11,
    -- filter=6 channel=123
    6, 8, -2, -7, 0, 7, -8, 0, 7,
    -- filter=6 channel=124
    -1, 11, 3, -4, 7, 0, 0, 2, 8,
    -- filter=6 channel=125
    -13, 6, 15, -8, -6, 3, -1, -9, -2,
    -- filter=6 channel=126
    -4, 5, 1, -10, 1, 11, -7, -11, 0,
    -- filter=6 channel=127
    -4, -3, 8, 5, -6, 3, 0, -3, -1,
    -- filter=7 channel=0
    16, 3, 2, 2, 2, -1, -7, -10, -2,
    -- filter=7 channel=1
    0, -5, 4, 3, 14, 6, -3, -12, -12,
    -- filter=7 channel=2
    -6, 0, -8, -2, 19, 5, 7, 0, -2,
    -- filter=7 channel=3
    20, 39, 24, 16, 15, 21, -3, -2, 0,
    -- filter=7 channel=4
    4, -4, 11, 23, 37, 26, 17, 31, 7,
    -- filter=7 channel=5
    11, 1, 5, -1, 4, -8, -9, 0, 7,
    -- filter=7 channel=6
    -6, -6, -7, 3, 0, 4, 6, 0, 2,
    -- filter=7 channel=7
    2, 7, 2, 3, 0, -6, 0, 0, -7,
    -- filter=7 channel=8
    2, 1, -4, 0, 12, -1, 9, 0, 6,
    -- filter=7 channel=9
    -2, 0, -9, 7, 19, 12, -13, -16, -6,
    -- filter=7 channel=10
    -1, 3, 2, 6, 14, 10, -2, -11, -9,
    -- filter=7 channel=11
    -12, -5, 1, 8, 10, 2, 3, 1, 6,
    -- filter=7 channel=12
    5, -9, -2, -8, 1, -3, 1, 1, -2,
    -- filter=7 channel=13
    -11, -10, -8, 23, 29, 17, -9, -21, -4,
    -- filter=7 channel=14
    -7, -3, 7, -3, 0, 6, 2, 0, 0,
    -- filter=7 channel=15
    -4, 1, -6, 18, 11, 12, -4, -1, -6,
    -- filter=7 channel=16
    -9, -1, -4, -4, 7, 0, -5, -5, -4,
    -- filter=7 channel=17
    4, -1, -4, 0, -6, -1, 5, 7, 0,
    -- filter=7 channel=18
    -10, -14, -6, 15, 19, 17, -3, -22, -9,
    -- filter=7 channel=19
    -4, 0, -4, 0, -6, 0, 5, -4, 3,
    -- filter=7 channel=20
    -14, -9, 0, -1, 15, 9, 1, -2, -3,
    -- filter=7 channel=21
    -8, 1, -5, -4, 10, 5, -9, -1, -2,
    -- filter=7 channel=22
    3, 5, 0, -3, -3, -4, -1, 2, 6,
    -- filter=7 channel=23
    -8, 6, -13, 24, 32, 16, -15, -20, -1,
    -- filter=7 channel=24
    4, 1, 5, 4, 2, -3, -2, 0, 1,
    -- filter=7 channel=25
    -19, -23, -13, 24, 31, 26, -14, -19, -10,
    -- filter=7 channel=26
    -5, -5, 3, -8, -2, 3, -4, -7, -4,
    -- filter=7 channel=27
    -22, -34, -27, 49, 58, 34, -33, -40, -23,
    -- filter=7 channel=28
    0, -1, 0, -5, 6, -6, 4, 0, 2,
    -- filter=7 channel=29
    -12, -12, -12, 5, 9, 11, -5, -6, -5,
    -- filter=7 channel=30
    -9, -21, -5, 21, 33, 24, -20, -20, -6,
    -- filter=7 channel=31
    -21, -15, -7, 26, 33, 18, -26, -21, -3,
    -- filter=7 channel=32
    -6, -24, -8, 33, 36, 13, -16, -23, -7,
    -- filter=7 channel=33
    -2, 6, -10, 13, 14, 6, -8, -11, 0,
    -- filter=7 channel=34
    -3, -10, -10, 0, -9, -8, -10, 0, 4,
    -- filter=7 channel=35
    -2, -3, -6, 6, 6, -1, 3, -3, 7,
    -- filter=7 channel=36
    -1, -6, 1, 6, 8, 2, 6, -1, 0,
    -- filter=7 channel=37
    -2, -15, -4, -4, 9, 4, 4, 1, -8,
    -- filter=7 channel=38
    -3, 0, 0, 14, 18, 3, -16, -20, 0,
    -- filter=7 channel=39
    -13, 0, -10, -2, 11, 12, -8, -7, 1,
    -- filter=7 channel=40
    -6, 5, -7, -8, 0, 4, 2, 0, 4,
    -- filter=7 channel=41
    -4, -12, -17, -18, -3, -3, 4, 3, -9,
    -- filter=7 channel=42
    -6, 0, -5, 4, 14, 10, -4, -11, -6,
    -- filter=7 channel=43
    17, 22, 5, 4, 6, 0, -4, -5, 9,
    -- filter=7 channel=44
    -9, -9, 3, 13, 12, 5, -3, -12, -2,
    -- filter=7 channel=45
    3, 9, -2, 4, -6, 4, -9, 5, 6,
    -- filter=7 channel=46
    8, 5, -6, -8, 3, -2, 7, 0, 0,
    -- filter=7 channel=47
    4, 2, 0, 3, 13, 2, -12, -10, 0,
    -- filter=7 channel=48
    -17, -28, -2, 34, 45, 25, -7, -19, -8,
    -- filter=7 channel=49
    -16, -16, -5, 23, 29, 16, -5, 0, -6,
    -- filter=7 channel=50
    -11, -14, -5, 23, 25, 13, -11, -23, -11,
    -- filter=7 channel=51
    4, -6, -6, 0, 3, 6, 7, 1, 6,
    -- filter=7 channel=52
    -4, -1, -8, 8, -6, 0, 5, 8, 8,
    -- filter=7 channel=53
    0, -2, -8, -2, 8, 7, 0, 0, -3,
    -- filter=7 channel=54
    -5, 0, 1, 0, 5, 5, -1, 3, 2,
    -- filter=7 channel=55
    -8, -13, -12, 14, 29, 18, 0, -2, -6,
    -- filter=7 channel=56
    -9, -8, 0, -1, -2, 5, 3, 1, 3,
    -- filter=7 channel=57
    3, -10, -3, 5, 9, 1, 3, 0, 8,
    -- filter=7 channel=58
    4, 0, 4, -4, 1, -9, 2, -1, -4,
    -- filter=7 channel=59
    -7, -18, -9, 13, 17, 15, -3, -14, -5,
    -- filter=7 channel=60
    -3, 3, 2, -4, -3, -2, 0, 5, -4,
    -- filter=7 channel=61
    0, -10, -1, 0, 2, -1, -4, 6, -4,
    -- filter=7 channel=62
    -2, 9, 3, 4, 1, 3, 0, 8, 4,
    -- filter=7 channel=63
    6, -2, -5, 3, 0, -3, -5, 0, 4,
    -- filter=7 channel=64
    -1, -5, -6, 6, 0, 6, 5, 0, -2,
    -- filter=7 channel=65
    -7, 2, -6, -4, -5, -3, 4, -1, 1,
    -- filter=7 channel=66
    -2, -5, -10, -12, 2, -12, 6, 2, 6,
    -- filter=7 channel=67
    -4, 5, 8, 0, -8, 5, -3, 3, -1,
    -- filter=7 channel=68
    0, -8, 1, -3, 10, 3, 2, 1, 8,
    -- filter=7 channel=69
    0, -7, -1, 0, 3, 4, -7, -8, -4,
    -- filter=7 channel=70
    -6, -2, 0, 23, 13, 13, -7, -6, 0,
    -- filter=7 channel=71
    5, 22, 6, -5, -4, -1, 0, 9, 10,
    -- filter=7 channel=72
    -4, -5, -11, 16, 18, 10, -4, -10, -1,
    -- filter=7 channel=73
    -7, -22, -8, 14, 22, 9, -2, -8, -12,
    -- filter=7 channel=74
    -13, -16, -6, 7, 9, 3, -4, -2, -2,
    -- filter=7 channel=75
    5, 9, 6, 10, -2, 0, -11, -17, 4,
    -- filter=7 channel=76
    0, 2, 0, -8, 5, 5, 3, -5, 4,
    -- filter=7 channel=77
    1, -4, -3, -7, 0, 0, 1, 0, -5,
    -- filter=7 channel=78
    4, -3, 4, -8, 2, -1, -6, -6, -7,
    -- filter=7 channel=79
    -14, -19, -17, 21, 40, 13, -20, -22, -12,
    -- filter=7 channel=80
    -16, -20, -7, 25, 34, 21, -20, -22, -16,
    -- filter=7 channel=81
    3, 2, -5, -3, -1, 5, 3, -3, -2,
    -- filter=7 channel=82
    -4, 12, 6, 0, -7, -5, 6, 5, 10,
    -- filter=7 channel=83
    -5, -6, -2, 11, 7, 6, -3, 1, 3,
    -- filter=7 channel=84
    -12, -24, -14, 8, 21, 17, -6, -11, -8,
    -- filter=7 channel=85
    2, -2, 0, -5, -2, 5, 1, -3, 7,
    -- filter=7 channel=86
    -3, -6, 1, -4, -4, -2, -9, 5, -7,
    -- filter=7 channel=87
    -1, 0, 1, 3, 1, 2, 3, -2, 1,
    -- filter=7 channel=88
    0, -10, -3, 10, 11, 5, -8, -3, 4,
    -- filter=7 channel=89
    6, -12, -11, 15, 23, 19, -4, -28, -2,
    -- filter=7 channel=90
    0, 13, 1, 3, -12, -7, 2, 9, 6,
    -- filter=7 channel=91
    -27, -28, -6, 29, 36, 24, 0, -12, -11,
    -- filter=7 channel=92
    7, 7, 1, -1, -7, 0, 10, 6, 1,
    -- filter=7 channel=93
    -5, -20, -3, 23, 21, 12, -3, -7, -11,
    -- filter=7 channel=94
    -1, -5, -6, -6, -3, -6, 0, -4, 0,
    -- filter=7 channel=95
    2, 8, -1, 3, -5, 5, -4, -1, -2,
    -- filter=7 channel=96
    4, 6, -1, 0, 7, 5, 3, -1, 0,
    -- filter=7 channel=97
    15, 32, 8, 4, -1, 4, -1, 12, 1,
    -- filter=7 channel=98
    -5, -15, -13, 32, 37, 17, -18, -24, -14,
    -- filter=7 channel=99
    -20, -13, -14, 19, 26, 12, -14, -13, -5,
    -- filter=7 channel=100
    -3, -10, 4, 0, -1, -6, -1, 3, 4,
    -- filter=7 channel=101
    7, -5, 2, 11, 30, 16, 10, 12, 12,
    -- filter=7 channel=102
    -6, -5, 5, 1, 7, -2, -4, -4, -2,
    -- filter=7 channel=103
    10, 16, 2, 0, -7, 6, -6, -5, 11,
    -- filter=7 channel=104
    -12, -1, 2, 8, 15, 5, -8, -15, 0,
    -- filter=7 channel=105
    -2, -5, -2, -3, 7, 7, 7, -8, -2,
    -- filter=7 channel=106
    0, 2, -3, 1, -2, -1, -3, 0, 5,
    -- filter=7 channel=107
    -7, -10, 0, 0, 3, 9, -7, 2, 2,
    -- filter=7 channel=108
    4, -3, 1, -4, -7, 5, 8, -6, -6,
    -- filter=7 channel=109
    -19, -36, -13, 24, 43, 29, -8, -26, -6,
    -- filter=7 channel=110
    5, 9, 5, 4, 7, 2, -3, 5, 3,
    -- filter=7 channel=111
    0, 5, 4, 3, -7, -1, 6, 4, 0,
    -- filter=7 channel=112
    -1, -2, -2, 16, 2, 0, -12, -3, 5,
    -- filter=7 channel=113
    -1, 15, -6, 1, 3, -2, -10, -12, 0,
    -- filter=7 channel=114
    -8, -32, -18, 30, 31, 30, -11, -33, -7,
    -- filter=7 channel=115
    5, 0, -2, 0, -4, -5, 5, -7, -4,
    -- filter=7 channel=116
    -23, -43, -21, 29, 50, 33, -15, -25, -8,
    -- filter=7 channel=117
    -5, -16, 0, 7, 9, 9, 0, -9, 0,
    -- filter=7 channel=118
    2, -1, 2, 2, -4, -7, 1, 1, 0,
    -- filter=7 channel=119
    -8, -15, -7, -6, -8, -7, -2, 0, 10,
    -- filter=7 channel=120
    -19, -40, -23, 29, 35, 21, -21, -27, -17,
    -- filter=7 channel=121
    0, -2, -8, 0, 7, 8, -3, -4, 5,
    -- filter=7 channel=122
    -8, -5, -7, 8, 1, 8, -10, -17, 2,
    -- filter=7 channel=123
    3, 1, 0, 5, -13, 0, 10, 0, 1,
    -- filter=7 channel=124
    0, -4, -4, 0, -3, -2, 5, -7, 1,
    -- filter=7 channel=125
    -17, -27, -11, 13, 30, 18, -13, -18, -12,
    -- filter=7 channel=126
    9, 8, -6, 6, 0, -1, -8, -8, -3,
    -- filter=7 channel=127
    -3, -9, -10, -10, -3, -6, 4, -2, 3,
    -- filter=8 channel=0
    -10, -10, -5, -9, 1, -4, 0, -4, 0,
    -- filter=8 channel=1
    -12, 0, -7, -13, -10, 1, -6, -1, 5,
    -- filter=8 channel=2
    -2, 1, 6, -7, -7, 4, 2, 1, 8,
    -- filter=8 channel=3
    -2, 1, 7, 2, 7, 3, 0, -4, -1,
    -- filter=8 channel=4
    -10, 3, -4, -9, 0, 3, -2, -6, 12,
    -- filter=8 channel=5
    -7, -6, 8, 0, -9, -3, 0, 0, 8,
    -- filter=8 channel=6
    7, -3, -8, 9, 0, -4, 4, -5, 2,
    -- filter=8 channel=7
    6, 1, 0, 0, 3, -7, -2, 6, 0,
    -- filter=8 channel=8
    2, 1, 7, 6, -7, -4, -5, -3, 6,
    -- filter=8 channel=9
    3, -5, -3, 3, 0, 1, -4, 1, -1,
    -- filter=8 channel=10
    10, 12, 15, -4, -6, -6, 0, -7, -11,
    -- filter=8 channel=11
    10, -2, 0, 9, 7, 0, 5, 3, -1,
    -- filter=8 channel=12
    -2, 0, -4, -4, 1, 0, 0, -1, -6,
    -- filter=8 channel=13
    0, 13, 1, -6, -4, -11, -4, -7, -8,
    -- filter=8 channel=14
    0, 2, -1, 1, 5, -5, -5, 0, 1,
    -- filter=8 channel=15
    4, 0, -2, -1, 0, 3, -6, -4, -9,
    -- filter=8 channel=16
    -10, 4, 7, -7, -1, 4, -10, -5, -2,
    -- filter=8 channel=17
    5, 5, -5, -3, 6, 0, 4, 2, 7,
    -- filter=8 channel=18
    8, 13, 4, -3, 7, -5, -2, 0, -1,
    -- filter=8 channel=19
    -6, 2, 2, -3, -3, 0, -3, -1, -4,
    -- filter=8 channel=20
    2, 0, -7, 12, -5, -10, 6, -9, -2,
    -- filter=8 channel=21
    -9, 1, -1, -4, -5, -6, -13, -5, 0,
    -- filter=8 channel=22
    7, 2, 9, 1, 5, -5, 3, 5, 0,
    -- filter=8 channel=23
    18, 19, 19, 10, 3, 3, 0, -14, 1,
    -- filter=8 channel=24
    3, 2, 7, 0, 2, -1, -4, 2, -3,
    -- filter=8 channel=25
    -7, 12, 2, -13, -3, 1, 1, 0, -3,
    -- filter=8 channel=26
    -4, 0, -6, 0, -5, -7, -8, 2, 4,
    -- filter=8 channel=27
    5, 9, 16, -5, 4, -7, 2, -1, 9,
    -- filter=8 channel=28
    7, 6, 0, -1, -5, 3, -6, -7, -2,
    -- filter=8 channel=29
    -1, -2, -12, 8, 3, -10, 0, 2, -8,
    -- filter=8 channel=30
    -2, -5, 2, -2, 2, -3, -7, -6, 6,
    -- filter=8 channel=31
    3, 15, 14, -12, 2, -2, -17, -3, 8,
    -- filter=8 channel=32
    5, 11, 2, -1, 5, -9, -8, -3, -8,
    -- filter=8 channel=33
    6, 9, 16, -2, -4, 5, -2, -9, 0,
    -- filter=8 channel=34
    -4, 1, 0, -3, -5, 7, -4, 0, 0,
    -- filter=8 channel=35
    -4, 7, 0, 2, 1, 4, -7, -3, -5,
    -- filter=8 channel=36
    -1, 4, -1, 0, 1, -1, -3, -3, -7,
    -- filter=8 channel=37
    -16, 0, -2, -14, 0, -11, 0, -7, 0,
    -- filter=8 channel=38
    0, 11, 11, -6, 0, -4, -8, -5, -7,
    -- filter=8 channel=39
    5, -2, -4, 8, 0, -2, 3, -4, -9,
    -- filter=8 channel=40
    8, 8, -8, -4, 6, -5, 0, 2, -11,
    -- filter=8 channel=41
    -6, -2, -5, -7, -8, -12, -11, -5, -1,
    -- filter=8 channel=42
    2, -7, 5, 1, -1, -1, 1, -3, 6,
    -- filter=8 channel=43
    11, -2, 2, 11, -1, 2, 5, -8, 2,
    -- filter=8 channel=44
    -13, -1, 0, -4, -9, -1, -4, -8, 7,
    -- filter=8 channel=45
    3, 5, 4, -3, -2, -4, 3, 1, 0,
    -- filter=8 channel=46
    -5, -4, 4, 6, 2, 6, -7, 0, 5,
    -- filter=8 channel=47
    0, -7, 1, -14, 0, 0, -6, 0, 4,
    -- filter=8 channel=48
    -3, -5, 9, -7, -1, 0, -3, 2, 11,
    -- filter=8 channel=49
    -1, 5, -1, -3, -2, -3, 7, 7, 3,
    -- filter=8 channel=50
    6, 12, 13, 1, 0, 4, 1, -8, 7,
    -- filter=8 channel=51
    2, 5, -5, -4, 0, 1, 6, -2, -3,
    -- filter=8 channel=52
    7, 1, -1, -5, -3, 0, 3, -4, 3,
    -- filter=8 channel=53
    8, 0, -2, 4, 6, -3, -3, -6, 4,
    -- filter=8 channel=54
    -4, 1, 3, 1, 2, 4, -5, -7, 0,
    -- filter=8 channel=55
    17, 14, -2, 10, 6, 2, 3, -10, -7,
    -- filter=8 channel=56
    -2, 3, 5, 4, -4, 2, -4, -3, 2,
    -- filter=8 channel=57
    -8, -6, -8, -4, -4, 4, 2, -1, -6,
    -- filter=8 channel=58
    -8, 5, -3, -6, -7, -3, -6, 4, 3,
    -- filter=8 channel=59
    6, 13, 3, -9, -10, 0, 0, 2, -1,
    -- filter=8 channel=60
    6, -2, 4, -3, -1, 7, 0, -1, -3,
    -- filter=8 channel=61
    1, 0, -4, -7, -5, -4, 0, 0, 2,
    -- filter=8 channel=62
    -2, 6, 7, 7, 5, 1, -2, -2, -3,
    -- filter=8 channel=63
    5, -5, -5, -8, -6, -4, 5, -6, 3,
    -- filter=8 channel=64
    0, -8, -2, 3, 6, 4, -8, 4, 2,
    -- filter=8 channel=65
    -5, -2, -6, 1, 1, -2, -5, 5, 2,
    -- filter=8 channel=66
    -3, -4, -2, -8, 0, -5, -8, 2, -11,
    -- filter=8 channel=67
    -7, 3, 5, -5, 0, 5, 0, -3, -4,
    -- filter=8 channel=68
    -6, -1, -4, 0, -3, -2, 2, 1, -6,
    -- filter=8 channel=69
    2, -5, 3, -5, -5, 0, -7, 2, -3,
    -- filter=8 channel=70
    12, 12, 4, -2, -1, 4, 1, -5, 0,
    -- filter=8 channel=71
    7, 0, 3, -1, 0, 4, -9, -5, -8,
    -- filter=8 channel=72
    0, 15, 1, -8, 1, 3, -12, -9, -4,
    -- filter=8 channel=73
    9, 1, 0, 3, -5, -4, 2, 0, 1,
    -- filter=8 channel=74
    0, 6, 0, 3, -9, -5, 0, -6, 1,
    -- filter=8 channel=75
    0, -6, 5, -5, -7, 2, -4, -11, -4,
    -- filter=8 channel=76
    2, -5, -6, 14, 0, -10, 1, -2, -5,
    -- filter=8 channel=77
    2, 2, -1, -7, -2, -7, 0, -6, -1,
    -- filter=8 channel=78
    -1, -3, -3, -8, -1, 1, -5, -6, 8,
    -- filter=8 channel=79
    13, 7, 7, -7, 0, -13, 3, -12, -16,
    -- filter=8 channel=80
    -4, 11, 9, -18, -4, -4, -14, -10, -1,
    -- filter=8 channel=81
    0, -5, 4, 0, -3, 3, -2, 1, 6,
    -- filter=8 channel=82
    4, 0, 1, 3, 0, -6, 3, 0, 4,
    -- filter=8 channel=83
    -4, 5, 3, 0, 0, -4, -6, 1, 5,
    -- filter=8 channel=84
    0, -7, 4, -5, 0, -2, -1, -8, 2,
    -- filter=8 channel=85
    -7, -3, 0, 7, -4, -7, -4, 3, 6,
    -- filter=8 channel=86
    -6, -9, 2, -9, 3, -8, -1, -4, 2,
    -- filter=8 channel=87
    -5, -9, 1, 5, 0, 6, 0, -4, -3,
    -- filter=8 channel=88
    -4, -2, 5, -8, -3, -3, 6, -4, -4,
    -- filter=8 channel=89
    11, 21, 14, 0, -2, -7, -9, -6, -14,
    -- filter=8 channel=90
    6, -7, 0, 4, -6, 10, 3, -8, 0,
    -- filter=8 channel=91
    9, -2, 5, -7, -7, -4, 2, -7, -5,
    -- filter=8 channel=92
    -3, -2, 4, -4, -8, 7, 0, 0, -3,
    -- filter=8 channel=93
    -9, 1, -4, -17, -8, -4, -1, -1, 9,
    -- filter=8 channel=94
    0, 3, 0, -1, 1, 4, 0, 1, -3,
    -- filter=8 channel=95
    -6, 5, 5, -1, 6, -1, -8, -2, 4,
    -- filter=8 channel=96
    -6, 4, 7, 1, 0, -7, 2, 2, -2,
    -- filter=8 channel=97
    6, 1, 6, 0, 5, 1, 0, -1, -3,
    -- filter=8 channel=98
    8, 17, 9, -10, -7, -6, -2, -9, -9,
    -- filter=8 channel=99
    12, 9, 7, -7, -4, 5, -9, -3, 1,
    -- filter=8 channel=100
    0, -2, -3, 0, 4, 1, -3, 5, 1,
    -- filter=8 channel=101
    1, 3, -4, -6, 1, 5, 2, 0, 5,
    -- filter=8 channel=102
    -6, 0, 6, 1, 5, 0, -5, 2, 6,
    -- filter=8 channel=103
    -10, -1, 8, -14, -8, 5, -11, -6, -8,
    -- filter=8 channel=104
    -3, 6, 5, -9, -1, -8, -1, -8, 7,
    -- filter=8 channel=105
    7, 1, -6, 10, 7, -2, 0, 2, -5,
    -- filter=8 channel=106
    -5, 1, -2, 5, 4, -1, -2, 2, 1,
    -- filter=8 channel=107
    5, 0, -2, 5, -2, 3, -2, -2, 1,
    -- filter=8 channel=108
    3, 0, 0, 0, -2, 0, -2, 5, -1,
    -- filter=8 channel=109
    0, 3, 10, -6, -1, 2, -3, -9, 3,
    -- filter=8 channel=110
    5, 7, 5, 1, -1, 6, -9, -3, -2,
    -- filter=8 channel=111
    2, 3, -3, -3, -8, 2, 4, -5, -1,
    -- filter=8 channel=112
    1, 7, 3, -7, 1, 3, -9, -4, 5,
    -- filter=8 channel=113
    7, 16, 15, -5, -4, 1, -1, -2, 2,
    -- filter=8 channel=114
    4, 1, 2, 3, -6, -4, -2, -1, 4,
    -- filter=8 channel=115
    -1, 0, -3, 2, 6, -1, 4, -2, -5,
    -- filter=8 channel=116
    4, 5, -2, -13, -7, -2, -6, -10, -7,
    -- filter=8 channel=117
    5, 0, 3, -3, 5, 1, 4, 2, -6,
    -- filter=8 channel=118
    -6, -3, 0, -3, -7, 5, -1, 1, 3,
    -- filter=8 channel=119
    1, -9, 10, 0, -12, 2, 1, -2, -3,
    -- filter=8 channel=120
    13, 10, 3, 3, -4, -10, -2, -6, 2,
    -- filter=8 channel=121
    -5, 7, 2, 1, 1, 3, -6, 1, 0,
    -- filter=8 channel=122
    -15, 0, 6, -22, -11, -10, -8, -14, 0,
    -- filter=8 channel=123
    1, -4, 5, 3, 5, 9, 0, 4, 5,
    -- filter=8 channel=124
    8, 4, -8, 6, 6, 0, 0, -7, -10,
    -- filter=8 channel=125
    5, 3, 5, -14, -3, -2, -1, 1, -6,
    -- filter=8 channel=126
    12, 8, 6, 6, 5, -8, -2, -7, -7,
    -- filter=8 channel=127
    -2, 2, -7, 5, 0, -6, -3, -1, -4,
    -- filter=9 channel=0
    -5, -3, 3, -5, 7, -1, 3, 0, 3,
    -- filter=9 channel=1
    2, 0, 0, 8, -5, -2, 2, 9, 6,
    -- filter=9 channel=2
    7, -1, -6, 1, 0, 5, 6, -6, -2,
    -- filter=9 channel=3
    2, 2, -5, 0, -5, -2, 1, 7, 5,
    -- filter=9 channel=4
    -5, -6, 0, 0, 0, -1, 5, -2, -5,
    -- filter=9 channel=5
    3, -5, 0, 0, 0, -1, -3, 1, 0,
    -- filter=9 channel=6
    0, -4, -2, -5, -6, 1, -3, -2, -6,
    -- filter=9 channel=7
    4, 4, -5, -1, 2, 0, 3, 3, 2,
    -- filter=9 channel=8
    2, 0, -7, 0, 5, 6, -7, -7, -6,
    -- filter=9 channel=9
    3, -7, -5, -7, -6, -7, -3, -4, 4,
    -- filter=9 channel=10
    -8, 3, -3, -2, -7, -2, 4, 1, 4,
    -- filter=9 channel=11
    -3, 4, 3, -7, -2, -1, 4, -1, 2,
    -- filter=9 channel=12
    4, -2, 2, -4, -4, -4, 0, 1, 2,
    -- filter=9 channel=13
    -3, 1, 6, -5, 4, -2, -3, -4, -4,
    -- filter=9 channel=14
    2, 2, 2, 4, 4, -2, 0, 0, 6,
    -- filter=9 channel=15
    6, 4, -4, 4, 5, 4, 4, 1, 6,
    -- filter=9 channel=16
    1, 3, -6, -3, 0, -7, -5, -3, -7,
    -- filter=9 channel=17
    0, -7, 5, 0, -3, 2, 4, 4, 3,
    -- filter=9 channel=18
    -5, -7, -2, -4, -5, -4, -3, -3, 3,
    -- filter=9 channel=19
    0, 1, -1, 0, -6, -6, 7, 3, 2,
    -- filter=9 channel=20
    1, 4, -4, 5, -7, 3, -6, 7, 7,
    -- filter=9 channel=21
    -1, 3, -5, 4, 0, -3, 1, 4, 1,
    -- filter=9 channel=22
    4, 6, 0, 0, -5, 1, 7, -5, 5,
    -- filter=9 channel=23
    5, 1, 6, 6, -2, 5, 2, -3, 2,
    -- filter=9 channel=24
    -2, -7, 0, 1, -3, 7, -1, 2, 0,
    -- filter=9 channel=25
    -5, 4, 0, -4, -1, 3, 7, -7, -9,
    -- filter=9 channel=26
    0, -1, -2, 7, 3, 2, 7, -4, 6,
    -- filter=9 channel=27
    0, 0, -6, -8, -3, -9, 2, 5, 2,
    -- filter=9 channel=28
    0, -2, 0, -1, -2, -6, -7, -1, -2,
    -- filter=9 channel=29
    1, 1, 1, -5, 4, 1, -4, -6, 7,
    -- filter=9 channel=30
    0, 1, -4, 1, 0, -1, 0, -3, -4,
    -- filter=9 channel=31
    1, 5, 2, 0, -8, -7, 0, -5, -8,
    -- filter=9 channel=32
    1, -6, 0, -3, -6, 3, -3, -7, 5,
    -- filter=9 channel=33
    -4, 4, 0, -1, -3, -1, 5, -3, -1,
    -- filter=9 channel=34
    -1, 2, 7, 1, -3, 5, -4, 5, -7,
    -- filter=9 channel=35
    3, 3, 4, 2, 6, -7, 1, 5, -1,
    -- filter=9 channel=36
    -5, 0, -2, -5, 5, -2, 4, 1, -2,
    -- filter=9 channel=37
    2, -4, 6, 3, -3, 5, 9, 8, -2,
    -- filter=9 channel=38
    4, 4, -4, -1, -5, 4, 3, 2, -5,
    -- filter=9 channel=39
    -7, 3, 7, -1, 6, -2, -5, 6, 4,
    -- filter=9 channel=40
    3, 0, -3, -2, 2, 4, 1, 2, 0,
    -- filter=9 channel=41
    4, -1, -4, 10, -3, -5, 5, 0, -3,
    -- filter=9 channel=42
    5, 6, -7, -1, -1, -7, 6, 0, -2,
    -- filter=9 channel=43
    0, -2, 0, 2, 7, 1, -3, -2, -1,
    -- filter=9 channel=44
    2, -7, 0, -4, -5, -2, 2, 3, 5,
    -- filter=9 channel=45
    -1, -4, 0, -2, -4, -4, -2, 2, 1,
    -- filter=9 channel=46
    -4, -6, 5, 2, -5, 0, -1, 8, -3,
    -- filter=9 channel=47
    0, -4, -1, 5, 5, 6, 3, 5, 4,
    -- filter=9 channel=48
    0, -1, 1, -7, 3, -2, 0, -4, 5,
    -- filter=9 channel=49
    -1, 2, 1, 2, 4, -1, -3, -4, 4,
    -- filter=9 channel=50
    -3, 3, 1, 2, 2, -4, -3, 4, 2,
    -- filter=9 channel=51
    -6, -1, 4, 1, -1, 2, 0, 0, -6,
    -- filter=9 channel=52
    0, -6, 3, 2, 2, 7, -1, -6, -1,
    -- filter=9 channel=53
    -5, 5, 1, -5, -3, 0, -2, 7, -6,
    -- filter=9 channel=54
    4, -6, 3, -5, 6, 4, -4, -7, 5,
    -- filter=9 channel=55
    0, 1, 4, 4, -7, -4, -1, 5, 4,
    -- filter=9 channel=56
    3, 7, 0, -5, -6, 0, -2, 6, -7,
    -- filter=9 channel=57
    -7, -6, 6, 0, 2, -6, 3, 4, 2,
    -- filter=9 channel=58
    -5, 3, 0, 0, -2, 2, 5, -1, 3,
    -- filter=9 channel=59
    -2, -2, -7, -1, -5, 2, 0, 2, 4,
    -- filter=9 channel=60
    6, 1, 2, 1, -4, 0, 6, -2, -4,
    -- filter=9 channel=61
    -1, 2, -2, -7, -3, -1, -4, -7, 2,
    -- filter=9 channel=62
    -6, -2, 6, 5, -1, 2, -7, -5, 5,
    -- filter=9 channel=63
    0, -6, 4, 3, 0, -5, -6, 3, 0,
    -- filter=9 channel=64
    3, 6, 6, 0, -2, -3, 0, -6, 3,
    -- filter=9 channel=65
    1, -1, -5, 3, -3, -1, 6, -7, 0,
    -- filter=9 channel=66
    -5, -3, 1, 3, 1, -2, 1, -3, -5,
    -- filter=9 channel=67
    -5, 6, 3, 4, -1, 7, -2, 1, -4,
    -- filter=9 channel=68
    0, -1, 1, 4, -3, 0, -2, -3, 2,
    -- filter=9 channel=69
    3, 1, 2, -5, -6, 0, 0, 7, 1,
    -- filter=9 channel=70
    -1, -2, 3, 2, -5, -8, -3, -2, -7,
    -- filter=9 channel=71
    -6, 4, 1, 3, 7, -5, -2, 0, 2,
    -- filter=9 channel=72
    6, 5, 0, -2, -6, 6, -6, 2, -7,
    -- filter=9 channel=73
    -2, 2, -5, 4, -4, 0, -5, -5, -2,
    -- filter=9 channel=74
    -3, -3, 6, -6, 2, -5, -5, -2, -6,
    -- filter=9 channel=75
    -5, 0, 5, 8, -4, 0, 5, -1, 1,
    -- filter=9 channel=76
    3, -2, -2, 4, 1, 0, 4, -6, -6,
    -- filter=9 channel=77
    0, 0, -1, -1, 2, 1, 7, 6, 5,
    -- filter=9 channel=78
    4, -5, 1, 7, 4, 5, -2, -4, 7,
    -- filter=9 channel=79
    6, -1, 3, -6, -6, -7, 2, -5, -6,
    -- filter=9 channel=80
    5, -6, 1, 0, 1, -8, 1, 4, 0,
    -- filter=9 channel=81
    3, 5, -1, -4, 0, -5, -5, 0, 2,
    -- filter=9 channel=82
    -7, -6, 3, -1, 2, 1, 2, 6, 1,
    -- filter=9 channel=83
    -7, -5, -4, -5, 5, 5, 7, 5, 3,
    -- filter=9 channel=84
    6, 0, 6, 5, 0, -4, 4, 1, 4,
    -- filter=9 channel=85
    -4, 3, -6, 0, -5, -2, 0, 6, 0,
    -- filter=9 channel=86
    4, 4, 0, -5, 3, 0, 4, -1, -1,
    -- filter=9 channel=87
    5, 6, -2, -3, 0, 5, 1, 5, -4,
    -- filter=9 channel=88
    4, -2, 7, -6, -5, 0, -4, 1, 2,
    -- filter=9 channel=89
    0, 4, 0, -3, -7, -6, 0, 0, 0,
    -- filter=9 channel=90
    4, -5, -1, -2, 3, 0, 2, 2, -5,
    -- filter=9 channel=91
    -5, -5, -3, 0, -6, -1, 1, 1, -7,
    -- filter=9 channel=92
    1, 3, -1, -3, -7, -7, 6, -6, 3,
    -- filter=9 channel=93
    4, 0, -4, 3, 2, -1, 4, -1, -8,
    -- filter=9 channel=94
    -4, -5, -5, -2, -1, 1, 4, -2, 5,
    -- filter=9 channel=95
    -4, 6, -4, 2, -3, -2, -5, 3, -2,
    -- filter=9 channel=96
    1, 0, 0, 1, -1, 3, -5, -5, -5,
    -- filter=9 channel=97
    -6, 6, -3, 8, 6, 2, 3, 5, -5,
    -- filter=9 channel=98
    4, -3, -5, -5, 0, -8, -1, 5, 0,
    -- filter=9 channel=99
    -5, -6, -1, -2, -8, -3, 6, -6, -4,
    -- filter=9 channel=100
    -5, 6, 0, -4, -6, -6, 1, 0, -4,
    -- filter=9 channel=101
    -4, 6, 3, -4, -1, -5, -4, 6, 0,
    -- filter=9 channel=102
    5, 7, -2, -5, -1, -2, -2, 5, 0,
    -- filter=9 channel=103
    3, 0, -7, 2, -3, 3, -5, -3, -1,
    -- filter=9 channel=104
    -3, 5, -8, -7, 4, -2, 0, 3, -8,
    -- filter=9 channel=105
    -5, 5, 0, -7, -7, 2, 7, -2, 7,
    -- filter=9 channel=106
    1, 1, 6, 7, 7, 2, -5, -2, -5,
    -- filter=9 channel=107
    6, -5, -4, -5, 8, 1, 7, -6, 8,
    -- filter=9 channel=108
    -3, -2, 1, 4, 1, -3, 0, 8, 5,
    -- filter=9 channel=109
    -6, 0, -3, -2, 2, -7, 5, 3, -7,
    -- filter=9 channel=110
    4, -1, 0, -1, 1, 3, 4, -3, 0,
    -- filter=9 channel=111
    5, 0, 7, 6, 0, -5, 7, 7, 5,
    -- filter=9 channel=112
    5, 2, 2, 6, -7, 0, 1, -5, -2,
    -- filter=9 channel=113
    0, 4, 2, -3, 0, 0, 0, 3, -3,
    -- filter=9 channel=114
    -1, 4, -3, -1, -4, 0, 1, 0, -4,
    -- filter=9 channel=115
    7, 0, -6, 2, 2, 0, 2, -1, 0,
    -- filter=9 channel=116
    -1, 2, -6, -5, 3, 4, 1, 6, -2,
    -- filter=9 channel=117
    5, 0, 0, -3, 3, -7, 7, 1, -5,
    -- filter=9 channel=118
    5, 5, -6, -4, 6, -5, -2, -1, -2,
    -- filter=9 channel=119
    5, -4, 4, -6, -4, -5, 5, -1, 3,
    -- filter=9 channel=120
    -2, -5, -7, -3, -3, -8, 3, -5, 0,
    -- filter=9 channel=121
    -4, -6, 3, 7, 1, 3, 0, -3, 5,
    -- filter=9 channel=122
    -3, 1, 6, 3, 0, -3, -1, 2, 2,
    -- filter=9 channel=123
    -2, 0, -2, 4, -6, -5, -3, -3, -4,
    -- filter=9 channel=124
    -6, 6, -1, 1, 7, 4, 0, 0, 7,
    -- filter=9 channel=125
    4, -2, 0, 2, 2, -2, -5, 0, 2,
    -- filter=9 channel=126
    0, 0, -5, 4, -5, 2, 2, -3, -4,
    -- filter=9 channel=127
    -6, -5, 5, 6, 3, 2, 6, 5, 3,
    -- filter=10 channel=0
    -17, -3, 6, -18, -3, 15, -4, 0, 16,
    -- filter=10 channel=1
    -12, -8, 9, -16, -4, 17, -10, 4, 14,
    -- filter=10 channel=2
    5, 4, 2, -3, -3, 1, 4, 4, -8,
    -- filter=10 channel=3
    -3, 0, 11, 1, 5, 10, -3, 4, 3,
    -- filter=10 channel=4
    0, -4, -7, 0, -9, -7, -12, -1, 7,
    -- filter=10 channel=5
    -9, 0, 9, -14, 1, 0, -5, -3, 0,
    -- filter=10 channel=6
    -2, 3, -6, -2, 4, -2, -4, 0, -2,
    -- filter=10 channel=7
    -4, 2, 1, -4, 0, -7, 5, 6, -1,
    -- filter=10 channel=8
    0, -2, -2, 6, 0, -6, 2, 4, 3,
    -- filter=10 channel=9
    5, 2, -4, 2, 4, 0, 7, -7, -4,
    -- filter=10 channel=10
    0, 0, -4, 15, 14, -1, 10, 5, -7,
    -- filter=10 channel=11
    4, 4, -10, 8, 13, -10, 2, -2, -13,
    -- filter=10 channel=12
    -7, 6, -2, 0, 4, 0, -2, -6, -2,
    -- filter=10 channel=13
    -1, -1, -4, -1, 3, 3, 8, -4, -12,
    -- filter=10 channel=14
    6, -5, -1, 2, 2, 3, -5, 0, 0,
    -- filter=10 channel=15
    -13, 2, -1, 5, 0, 0, -7, -6, 0,
    -- filter=10 channel=16
    -5, 0, 3, -3, 5, -9, 2, -2, -4,
    -- filter=10 channel=17
    -4, -3, 0, 7, 5, 2, 5, 6, 4,
    -- filter=10 channel=18
    -23, -5, 6, -5, 10, 3, -1, 2, 1,
    -- filter=10 channel=19
    2, 1, 3, 0, 3, 3, 2, 7, 5,
    -- filter=10 channel=20
    6, 2, -5, 13, 11, 0, 7, 5, -11,
    -- filter=10 channel=21
    12, 5, 0, 12, 13, -7, 6, 4, -17,
    -- filter=10 channel=22
    -7, -9, -3, -7, 2, 11, -6, 3, 0,
    -- filter=10 channel=23
    -2, 1, -7, 15, 5, -5, 4, -6, 0,
    -- filter=10 channel=24
    -2, -5, 6, -3, -6, -3, 1, 6, 2,
    -- filter=10 channel=25
    -10, 3, 4, 3, 11, -4, -7, -4, -3,
    -- filter=10 channel=26
    -3, -1, 1, -2, -5, 4, -3, 1, 4,
    -- filter=10 channel=27
    -11, -7, 11, 3, -6, 0, -11, -16, -6,
    -- filter=10 channel=28
    -6, 1, 3, 3, 2, 4, 6, 5, 3,
    -- filter=10 channel=29
    3, 4, -8, 6, 10, -10, 12, 6, -11,
    -- filter=10 channel=30
    -5, 4, -3, 1, -3, 3, -4, -5, 3,
    -- filter=10 channel=31
    15, 9, -5, 28, 0, -11, 5, -10, -27,
    -- filter=10 channel=32
    -6, -8, 9, -4, 5, -2, -3, -4, 4,
    -- filter=10 channel=33
    -9, -2, 1, -1, -2, 5, -5, -3, -3,
    -- filter=10 channel=34
    1, -5, 1, 2, -10, -1, -3, -3, 0,
    -- filter=10 channel=35
    3, -1, 0, -6, -4, 3, 1, -5, 4,
    -- filter=10 channel=36
    20, 1, -11, 19, 0, -13, -4, 0, -12,
    -- filter=10 channel=37
    -14, -2, 8, -13, -9, 13, -9, 0, 7,
    -- filter=10 channel=38
    2, 0, -2, 0, -1, 5, 0, 1, 3,
    -- filter=10 channel=39
    6, 5, -11, 12, 5, -5, 3, 4, -2,
    -- filter=10 channel=40
    6, 4, 0, 5, 5, -7, 0, -2, 4,
    -- filter=10 channel=41
    -5, -8, -1, 0, 8, 1, -10, 6, -5,
    -- filter=10 channel=42
    1, 3, 6, -6, 3, -3, -5, -3, -5,
    -- filter=10 channel=43
    -13, -10, 5, -8, -4, 1, 6, -5, 5,
    -- filter=10 channel=44
    -8, 3, 11, 3, 4, -2, -3, -5, -6,
    -- filter=10 channel=45
    -3, -8, -6, 2, 0, 2, -4, 3, 8,
    -- filter=10 channel=46
    -4, -6, -4, 3, -6, 3, -2, 4, 4,
    -- filter=10 channel=47
    -8, -2, 7, 10, 4, -6, 7, 4, -9,
    -- filter=10 channel=48
    8, 0, 2, 9, 3, -4, 2, -11, -6,
    -- filter=10 channel=49
    -6, -1, -9, -2, -1, 1, -7, 1, -3,
    -- filter=10 channel=50
    -4, -5, -4, 0, -4, -6, 7, -5, -4,
    -- filter=10 channel=51
    0, -4, 0, 4, -4, 4, -2, -2, -3,
    -- filter=10 channel=52
    -3, 4, 1, 2, 0, -8, -5, -7, -6,
    -- filter=10 channel=53
    0, 0, -9, 9, 10, -8, -2, 1, -3,
    -- filter=10 channel=54
    -2, 0, 7, 7, 2, 4, 1, 1, -5,
    -- filter=10 channel=55
    -6, 3, 3, 12, 11, -7, 10, -1, -3,
    -- filter=10 channel=56
    7, 1, -1, 6, -6, -3, 1, -4, -5,
    -- filter=10 channel=57
    0, -6, 2, 2, 3, 4, 3, 3, -7,
    -- filter=10 channel=58
    -4, -8, 3, -7, -2, 2, -1, -1, 0,
    -- filter=10 channel=59
    -4, 6, 4, 6, 0, 0, 3, 2, -15,
    -- filter=10 channel=60
    1, -2, -2, 3, 5, 3, -1, -4, -1,
    -- filter=10 channel=61
    0, -1, -7, 7, 3, -1, 7, -4, 2,
    -- filter=10 channel=62
    0, -1, -3, 0, 4, 6, 8, -5, -5,
    -- filter=10 channel=63
    3, 4, -7, -1, 6, 4, 4, 0, 0,
    -- filter=10 channel=64
    5, 7, -11, 12, -4, 0, 5, 4, -8,
    -- filter=10 channel=65
    -6, 0, -5, 6, -3, 1, 2, 7, 5,
    -- filter=10 channel=66
    2, -10, -7, 5, -2, 5, -2, -5, 0,
    -- filter=10 channel=67
    -1, -3, 0, 5, 4, 2, -3, 3, -4,
    -- filter=10 channel=68
    9, -3, -5, 3, 2, -1, -6, -4, 3,
    -- filter=10 channel=69
    -2, 1, -8, 2, 2, -7, 0, 7, 6,
    -- filter=10 channel=70
    -8, 2, -5, -3, 1, 3, -1, -10, 0,
    -- filter=10 channel=71
    3, 1, 2, 5, 2, 7, 5, 0, 2,
    -- filter=10 channel=72
    6, 11, 0, 15, 13, -14, 13, -5, -24,
    -- filter=10 channel=73
    2, 5, 5, 9, 1, -2, -4, -2, -7,
    -- filter=10 channel=74
    11, 0, -6, 10, -6, -3, 0, -5, -8,
    -- filter=10 channel=75
    -15, -14, 16, -15, 8, 13, -3, 13, 8,
    -- filter=10 channel=76
    9, 12, 0, 14, 18, -9, 12, 4, -7,
    -- filter=10 channel=77
    5, -1, 0, 7, 7, -2, 0, -2, -3,
    -- filter=10 channel=78
    -1, 0, -2, 6, 0, -1, 0, -2, 3,
    -- filter=10 channel=79
    -24, -5, 7, -2, 9, 6, -9, -8, -5,
    -- filter=10 channel=80
    2, 4, 0, 19, 16, -13, 6, -7, -27,
    -- filter=10 channel=81
    3, 0, -6, 1, -4, 4, 0, -1, -2,
    -- filter=10 channel=82
    -4, 2, 3, -6, -3, 5, -3, 5, 6,
    -- filter=10 channel=83
    7, 9, 5, 4, -1, -3, 3, 2, -11,
    -- filter=10 channel=84
    -4, -3, -3, 0, 5, 4, -2, -2, 1,
    -- filter=10 channel=85
    0, -4, -5, 0, 5, 5, -5, 7, -3,
    -- filter=10 channel=86
    -6, 1, 6, -2, 5, 6, 2, -5, 7,
    -- filter=10 channel=87
    1, 2, -1, 7, 0, 5, 2, 9, -5,
    -- filter=10 channel=88
    12, 0, -2, 8, 4, -4, 9, -5, -16,
    -- filter=10 channel=89
    -5, -4, 5, 7, 16, -4, 2, 1, -14,
    -- filter=10 channel=90
    9, 0, -2, 8, -2, -3, 10, -4, -16,
    -- filter=10 channel=91
    3, 3, -7, 6, 3, -5, -9, -7, -4,
    -- filter=10 channel=92
    -8, -5, -2, -7, 0, 1, 5, 0, -6,
    -- filter=10 channel=93
    -9, 0, 2, 5, -6, -8, -4, 2, 1,
    -- filter=10 channel=94
    6, -6, -1, 5, -1, -2, -1, -4, -7,
    -- filter=10 channel=95
    6, -1, 8, 6, -4, 7, 1, -3, -4,
    -- filter=10 channel=96
    5, 4, -5, 1, -6, -5, -6, -4, -6,
    -- filter=10 channel=97
    -5, -4, 0, -2, -5, 8, 7, 3, -5,
    -- filter=10 channel=98
    -17, -8, 7, 10, 0, 3, 2, -3, -8,
    -- filter=10 channel=99
    14, 12, -9, 35, 8, -22, 15, -12, -24,
    -- filter=10 channel=100
    4, -6, -7, 0, 1, -8, -2, -2, 1,
    -- filter=10 channel=101
    2, 8, -6, 4, 0, 1, -2, -6, 0,
    -- filter=10 channel=102
    3, 2, 7, 0, -5, 5, 5, 0, -1,
    -- filter=10 channel=103
    -11, -7, 5, 7, 10, -4, 9, -3, -12,
    -- filter=10 channel=104
    15, 3, 2, 18, 1, -14, 0, -2, -24,
    -- filter=10 channel=105
    2, 9, -8, 2, 7, 0, 10, 6, 0,
    -- filter=10 channel=106
    6, 3, 0, 4, 5, 4, 0, 7, 0,
    -- filter=10 channel=107
    -2, -2, 1, -4, -4, -6, -4, -7, 4,
    -- filter=10 channel=108
    -9, 2, -6, -7, 0, 0, 1, 7, 6,
    -- filter=10 channel=109
    -11, 2, 0, 5, 7, 0, 3, -15, -6,
    -- filter=10 channel=110
    6, 1, 0, 14, 6, -12, 2, -6, -16,
    -- filter=10 channel=111
    -4, -1, 2, -5, -1, -1, 5, 0, 1,
    -- filter=10 channel=112
    -10, -1, 2, -6, 0, 6, 3, -8, 0,
    -- filter=10 channel=113
    -9, -8, -2, -3, 4, -5, 4, -2, 0,
    -- filter=10 channel=114
    -25, -5, -1, -20, -4, 7, -19, -5, 0,
    -- filter=10 channel=115
    4, -2, 0, 4, 7, 7, 2, 6, 4,
    -- filter=10 channel=116
    0, 11, -8, 13, 7, -11, -3, -12, -16,
    -- filter=10 channel=117
    -4, 1, -1, 7, 8, 4, 4, 4, -9,
    -- filter=10 channel=118
    -5, -1, -4, -1, 1, 1, 5, 6, 2,
    -- filter=10 channel=119
    -2, -2, -3, -2, 5, -5, 1, 5, 4,
    -- filter=10 channel=120
    4, 11, 0, 17, -1, -10, 4, -7, 1,
    -- filter=10 channel=121
    -3, -4, -4, -4, -2, -2, 1, 5, 0,
    -- filter=10 channel=122
    10, 11, 2, 12, 2, -8, 10, -5, -21,
    -- filter=10 channel=123
    -6, -6, -8, -5, 0, -8, 5, -3, -2,
    -- filter=10 channel=124
    -7, -3, -7, 3, 9, 0, 8, -4, 4,
    -- filter=10 channel=125
    10, 2, 5, 25, 6, -13, 1, -14, -21,
    -- filter=10 channel=126
    -15, -12, 1, 0, 5, 5, -2, 1, 3,
    -- filter=10 channel=127
    -2, 4, -3, 2, -2, -6, 0, -2, 0,
    -- filter=11 channel=0
    5, 3, 11, -7, 15, 3, -4, 0, -12,
    -- filter=11 channel=1
    3, 6, 3, 3, 9, 4, 0, -7, -17,
    -- filter=11 channel=2
    -5, -3, 2, -5, 8, -9, 2, 0, -1,
    -- filter=11 channel=3
    -4, -11, -4, -9, 4, 15, -8, 5, -4,
    -- filter=11 channel=4
    -14, -4, -15, 3, -4, -9, -2, -11, 21,
    -- filter=11 channel=5
    1, 1, -3, 4, 0, -9, 0, 2, -16,
    -- filter=11 channel=6
    -4, 0, 6, 2, 0, -9, 5, 4, 2,
    -- filter=11 channel=7
    -4, -7, -6, 6, 0, -4, 0, 0, 4,
    -- filter=11 channel=8
    -6, 3, 0, 8, 8, -5, 3, -8, 7,
    -- filter=11 channel=9
    -8, -5, -5, -7, -1, -9, -3, 4, 5,
    -- filter=11 channel=10
    -3, -5, 1, 0, 2, 13, 0, 13, -13,
    -- filter=11 channel=11
    -6, -4, -7, 1, 8, -8, 4, -3, -6,
    -- filter=11 channel=12
    7, 0, 1, 5, 11, -1, 0, 3, -13,
    -- filter=11 channel=13
    6, -1, -1, -9, 8, 0, -9, 10, -16,
    -- filter=11 channel=14
    2, 1, -3, 4, -7, -2, -5, 0, -7,
    -- filter=11 channel=15
    0, 1, 2, 2, 6, 2, 1, -5, -5,
    -- filter=11 channel=16
    -1, -3, 2, 3, -3, 3, 6, -2, -3,
    -- filter=11 channel=17
    1, 4, 0, -6, -2, 2, 2, 0, 0,
    -- filter=11 channel=18
    5, -3, 10, -8, 19, 1, 1, 12, -23,
    -- filter=11 channel=19
    -4, 0, 6, -3, -4, 6, -3, -5, 6,
    -- filter=11 channel=20
    0, 3, -9, -4, 3, -1, -5, 5, 0,
    -- filter=11 channel=21
    -5, -11, 3, 5, -7, 4, -1, 8, -2,
    -- filter=11 channel=22
    0, 0, -3, 6, -2, -1, -7, 5, -3,
    -- filter=11 channel=23
    -12, 4, 0, -13, 14, -21, -2, 0, -5,
    -- filter=11 channel=24
    1, -5, -5, 0, 2, 3, 3, -2, -6,
    -- filter=11 channel=25
    1, -11, 12, -3, 9, -12, 0, 6, -10,
    -- filter=11 channel=26
    -6, 5, -5, 1, 0, -3, -1, -6, 5,
    -- filter=11 channel=27
    -6, 8, 6, -3, 17, -27, 4, -9, -7,
    -- filter=11 channel=28
    -2, 6, -1, 0, 5, -4, -1, 0, 6,
    -- filter=11 channel=29
    -8, -4, -6, -5, 11, -5, 10, -2, -8,
    -- filter=11 channel=30
    -7, -5, 0, 1, 9, -10, -1, -7, -7,
    -- filter=11 channel=31
    -7, -4, 6, -1, 5, -6, 5, -9, 1,
    -- filter=11 channel=32
    -4, -3, 10, -2, 14, -8, 3, 6, -23,
    -- filter=11 channel=33
    1, -10, 5, -1, 2, -6, -3, 11, -25,
    -- filter=11 channel=34
    -10, 10, -5, 5, 9, -5, -7, -8, 16,
    -- filter=11 channel=35
    -6, 2, -3, 0, -3, -7, -4, 6, 3,
    -- filter=11 channel=36
    -3, 2, -5, 0, 5, -3, 7, 5, 3,
    -- filter=11 channel=37
    -2, 5, -2, -4, 15, -1, 11, -5, 0,
    -- filter=11 channel=38
    3, -1, -3, -1, 13, -10, 0, -2, -14,
    -- filter=11 channel=39
    -5, 4, -3, -1, -4, -3, 3, 1, 2,
    -- filter=11 channel=40
    2, -5, -6, -5, 3, 6, -6, 5, 2,
    -- filter=11 channel=41
    4, -18, -1, -5, -17, 21, -3, 20, -9,
    -- filter=11 channel=42
    -4, 6, 0, -8, -4, -7, 5, 1, -3,
    -- filter=11 channel=43
    -1, -1, -5, 0, 4, -1, -13, -1, -16,
    -- filter=11 channel=44
    -2, 5, 1, -2, 6, -8, 13, -10, -3,
    -- filter=11 channel=45
    6, 0, 6, -2, -6, -7, 7, -7, -6,
    -- filter=11 channel=46
    -2, 3, 5, -6, -3, 6, 1, 2, 0,
    -- filter=11 channel=47
    4, -9, 0, -6, -3, -4, 12, 3, 1,
    -- filter=11 channel=48
    -5, -5, 6, -8, 17, -13, 9, -8, -6,
    -- filter=11 channel=49
    -2, 6, -1, -1, 0, -5, 9, -4, 0,
    -- filter=11 channel=50
    2, 7, -2, -9, 0, -9, 3, -4, -6,
    -- filter=11 channel=51
    -4, -5, -5, -3, 0, 7, -1, -2, 3,
    -- filter=11 channel=52
    -3, 14, -6, 6, 9, -6, -1, -1, 1,
    -- filter=11 channel=53
    0, -2, 2, 0, 6, -10, 2, -5, -2,
    -- filter=11 channel=54
    -5, 5, 7, 0, 2, -4, 6, 1, -2,
    -- filter=11 channel=55
    -5, -2, 9, -7, 18, 3, -4, 4, -5,
    -- filter=11 channel=56
    1, 7, -3, 4, 8, -2, 2, 7, 15,
    -- filter=11 channel=57
    -5, -8, 2, 0, -1, 3, 0, -3, 4,
    -- filter=11 channel=58
    2, 4, 2, -2, -7, 5, -5, 6, 0,
    -- filter=11 channel=59
    4, -6, 7, -5, 7, -1, 4, 3, -10,
    -- filter=11 channel=60
    3, 5, 5, -4, 6, 1, 4, 3, 3,
    -- filter=11 channel=61
    -2, 0, 0, -1, 3, 2, -6, -7, -3,
    -- filter=11 channel=62
    -4, 0, 0, -5, 7, 8, -1, 0, 5,
    -- filter=11 channel=63
    -3, -4, 3, -5, -8, -1, -1, -6, -2,
    -- filter=11 channel=64
    6, -3, 0, 0, 1, -2, 5, 3, 5,
    -- filter=11 channel=65
    -4, 0, -5, 6, -1, -7, 5, -6, -2,
    -- filter=11 channel=66
    3, -7, 1, 1, 1, 1, -6, 9, -7,
    -- filter=11 channel=67
    4, 5, 5, 4, 4, 5, 7, 1, 2,
    -- filter=11 channel=68
    2, -2, -6, -4, -1, -8, -1, 1, -1,
    -- filter=11 channel=69
    -4, 2, -1, -1, 2, 3, -6, 6, -9,
    -- filter=11 channel=70
    -5, 6, 1, 4, 16, -12, 5, -11, 11,
    -- filter=11 channel=71
    -1, -9, -3, 0, -7, -1, -3, -2, 5,
    -- filter=11 channel=72
    2, -2, 7, -5, 10, 3, -1, -4, -1,
    -- filter=11 channel=73
    -5, 8, 3, -9, 20, -6, 13, -7, 0,
    -- filter=11 channel=74
    -10, 4, -7, 3, 13, -21, 6, -15, 15,
    -- filter=11 channel=75
    2, -3, 1, 1, 5, 16, -3, 15, -24,
    -- filter=11 channel=76
    -3, -8, 6, -8, 9, 8, -7, 7, -7,
    -- filter=11 channel=77
    -4, 1, -6, -5, 0, -5, 1, 7, 2,
    -- filter=11 channel=78
    -4, 1, -2, -6, -2, -3, 0, 1, 3,
    -- filter=11 channel=79
    6, -3, 13, -5, 22, 0, -1, 8, -28,
    -- filter=11 channel=80
    -5, -16, 7, -18, 11, -3, 7, 9, -14,
    -- filter=11 channel=81
    2, 4, -5, -4, 5, -4, -2, 0, 0,
    -- filter=11 channel=82
    -1, 0, 3, 3, -4, 0, 4, -6, -4,
    -- filter=11 channel=83
    -10, 0, -1, 7, 6, -5, 0, -3, 4,
    -- filter=11 channel=84
    -2, 10, -5, -2, 15, -6, 1, -4, 4,
    -- filter=11 channel=85
    -5, 2, 0, -4, 0, 0, 2, 6, 0,
    -- filter=11 channel=86
    7, 6, 0, -1, 12, -13, 2, -8, -1,
    -- filter=11 channel=87
    1, 0, 0, 0, 4, -9, 0, 0, 6,
    -- filter=11 channel=88
    -6, 0, 0, 5, 10, 0, 6, 2, 5,
    -- filter=11 channel=89
    -7, -19, 3, -4, 10, 8, -5, 16, -29,
    -- filter=11 channel=90
    -8, 6, -2, 3, -6, 0, -5, -6, 21,
    -- filter=11 channel=91
    -1, 6, -1, 3, 12, -21, 0, -12, -3,
    -- filter=11 channel=92
    -1, -6, -9, -1, -9, 5, 0, -4, 6,
    -- filter=11 channel=93
    0, 1, 5, 3, 1, -7, 16, -12, -12,
    -- filter=11 channel=94
    1, 2, -7, -2, -5, 0, 7, 4, 5,
    -- filter=11 channel=95
    0, 3, 0, -5, 0, 0, 4, -1, 2,
    -- filter=11 channel=96
    0, -2, -8, -6, -5, 6, 1, 0, 0,
    -- filter=11 channel=97
    5, -2, -6, 5, 2, 5, -2, 10, -1,
    -- filter=11 channel=98
    -11, -15, 3, -13, 16, -1, 7, 0, -25,
    -- filter=11 channel=99
    -8, 0, 6, -11, 18, -14, -1, -5, 4,
    -- filter=11 channel=100
    0, 3, -7, 1, 0, 0, 5, -4, 9,
    -- filter=11 channel=101
    -5, -1, -3, 2, 1, -6, 0, -6, 15,
    -- filter=11 channel=102
    -1, -1, -6, 3, 6, 3, 0, -4, -2,
    -- filter=11 channel=103
    -1, -16, 5, -11, 0, -7, 4, 1, -16,
    -- filter=11 channel=104
    0, -6, 6, 0, 4, -9, 10, 0, -1,
    -- filter=11 channel=105
    0, -6, 7, -8, 10, 5, 4, 1, -9,
    -- filter=11 channel=106
    2, -3, 4, -5, -4, 11, -2, -2, 7,
    -- filter=11 channel=107
    -8, 2, -2, -6, 7, -7, 2, -1, -9,
    -- filter=11 channel=108
    -2, -5, -3, 5, -9, 13, 1, 1, 0,
    -- filter=11 channel=109
    -14, -3, 4, 0, 20, -25, 19, -14, -2,
    -- filter=11 channel=110
    -7, 3, -3, -10, 6, 7, -1, 6, 4,
    -- filter=11 channel=111
    -4, 3, 0, 3, -4, 5, -4, 6, 2,
    -- filter=11 channel=112
    -9, 9, -3, -2, 1, -4, -5, -6, 0,
    -- filter=11 channel=113
    -5, 0, 10, -6, 6, -1, -9, 6, -2,
    -- filter=11 channel=114
    -9, 5, 9, -7, 23, -16, 17, -9, -21,
    -- filter=11 channel=115
    -3, -2, -2, 0, -5, 6, -7, 5, 1,
    -- filter=11 channel=116
    -6, -1, 0, -10, 14, -16, 3, -6, -15,
    -- filter=11 channel=117
    1, -2, -5, -2, 6, -4, 5, -7, 1,
    -- filter=11 channel=118
    -5, 4, 2, -3, -2, 0, 0, 3, -1,
    -- filter=11 channel=119
    -6, 17, 0, -1, 11, -1, -6, 1, 13,
    -- filter=11 channel=120
    -9, 17, -8, -2, 27, -33, 11, -17, 2,
    -- filter=11 channel=121
    -2, -2, 3, -6, -1, 11, -6, 3, 0,
    -- filter=11 channel=122
    -4, -8, 10, 5, 0, 3, 7, 8, 7,
    -- filter=11 channel=123
    -2, -3, -5, 2, -3, -7, -9, 5, 11,
    -- filter=11 channel=124
    6, 3, 4, -7, -3, -8, 3, -5, -3,
    -- filter=11 channel=125
    0, 6, 3, -6, 4, -13, 7, -10, -3,
    -- filter=11 channel=126
    -2, -9, 10, -9, 7, 8, 0, 4, -14,
    -- filter=11 channel=127
    -1, -9, 5, -5, -6, 3, -1, -1, -1,
    -- filter=12 channel=0
    -4, 2, 13, -7, -3, 0, -8, -9, 10,
    -- filter=12 channel=1
    4, 5, 5, 2, -4, 2, -9, 3, 10,
    -- filter=12 channel=2
    1, -4, -5, -3, -5, 5, 8, -2, 2,
    -- filter=12 channel=3
    -2, -7, 1, -12, -6, 2, 0, -6, 0,
    -- filter=12 channel=4
    -4, 4, -12, 7, -12, 1, 1, -1, -4,
    -- filter=12 channel=5
    0, 1, 16, -5, -1, 12, -14, -7, 1,
    -- filter=12 channel=6
    3, -2, -6, 3, 4, -13, 2, -2, -2,
    -- filter=12 channel=7
    5, 0, 0, 7, 2, 4, 6, 1, 6,
    -- filter=12 channel=8
    0, -5, 2, -5, -6, -8, -1, -9, 2,
    -- filter=12 channel=9
    -3, 0, 0, -2, -4, 3, 2, 1, -3,
    -- filter=12 channel=10
    1, -2, 2, 0, -5, 5, -1, -7, -4,
    -- filter=12 channel=11
    -4, 0, 2, 9, 2, -11, 15, 10, -14,
    -- filter=12 channel=12
    5, -5, -2, -4, -7, 3, -3, 7, 5,
    -- filter=12 channel=13
    4, -13, 0, 11, -12, -6, 15, 0, 2,
    -- filter=12 channel=14
    -1, -1, 5, 3, -5, 0, -2, -7, 4,
    -- filter=12 channel=15
    0, -14, 1, 12, -6, -21, 23, 5, -15,
    -- filter=12 channel=16
    -5, 2, 14, -13, 5, 7, -12, 4, 2,
    -- filter=12 channel=17
    2, 6, 0, -2, 6, -5, 2, 6, 5,
    -- filter=12 channel=18
    3, -17, -5, 10, -13, -22, 31, 4, -19,
    -- filter=12 channel=19
    1, 0, 1, 4, -3, 1, -3, 0, -5,
    -- filter=12 channel=20
    1, -12, -5, 16, -6, -12, 21, 7, -13,
    -- filter=12 channel=21
    -2, 10, 5, -13, -2, 6, -12, -3, 8,
    -- filter=12 channel=22
    4, 0, 4, -2, -8, 0, -1, -1, 4,
    -- filter=12 channel=23
    -5, -7, 0, 8, -14, -13, 21, -9, -6,
    -- filter=12 channel=24
    -3, 3, -5, -2, -1, -3, -4, 4, 6,
    -- filter=12 channel=25
    -10, 0, 0, -3, 3, 0, 9, 0, 8,
    -- filter=12 channel=26
    -9, 1, 7, -8, -4, 7, -9, 5, 5,
    -- filter=12 channel=27
    -9, -3, 1, 4, -8, -6, 14, 0, 1,
    -- filter=12 channel=28
    -6, -1, 5, -3, -7, 0, -4, -5, -6,
    -- filter=12 channel=29
    -5, -2, -6, 15, 7, -12, 15, 5, -5,
    -- filter=12 channel=30
    -5, 7, 0, -8, -7, -1, 2, -4, 1,
    -- filter=12 channel=31
    -5, 8, 11, -5, 0, 5, -13, -13, -7,
    -- filter=12 channel=32
    0, -8, -2, 13, -14, -13, 28, 10, -8,
    -- filter=12 channel=33
    -11, -2, 12, 1, -1, -3, 2, -5, 2,
    -- filter=12 channel=34
    6, -2, 1, -2, 2, -5, 1, -5, 8,
    -- filter=12 channel=35
    0, -3, 3, -3, 1, -7, -1, -5, 6,
    -- filter=12 channel=36
    -5, -7, -3, 4, 3, -4, -3, -6, -7,
    -- filter=12 channel=37
    0, -1, 1, -9, -2, 17, -18, 0, 13,
    -- filter=12 channel=38
    -1, 0, 9, 4, -2, 2, -3, 0, 0,
    -- filter=12 channel=39
    4, 0, -3, 11, -4, -4, 10, -3, -12,
    -- filter=12 channel=40
    -2, -8, -2, 0, 1, -5, 0, -5, -8,
    -- filter=12 channel=41
    3, -8, -5, 15, -10, -8, 9, 9, -2,
    -- filter=12 channel=42
    -6, -3, 0, 5, -5, -4, 1, -6, 7,
    -- filter=12 channel=43
    -3, -6, -4, 5, -12, -6, 5, -8, -11,
    -- filter=12 channel=44
    -2, 1, 6, -6, -8, 12, -10, -1, 13,
    -- filter=12 channel=45
    5, -5, 4, 4, -1, 2, -1, -7, -6,
    -- filter=12 channel=46
    3, 1, -8, 9, 5, -4, -3, 0, -4,
    -- filter=12 channel=47
    -1, 15, 11, -9, 6, 16, -13, -3, 4,
    -- filter=12 channel=48
    -5, 4, 10, -1, 4, 2, 0, -5, 9,
    -- filter=12 channel=49
    -4, 1, 0, 14, -13, -11, 9, -5, -16,
    -- filter=12 channel=50
    -9, 2, 9, 0, -4, -5, 12, -2, -1,
    -- filter=12 channel=51
    -1, 0, 6, 1, -3, 0, 0, 6, -3,
    -- filter=12 channel=52
    -1, 2, 0, 2, -8, -1, 8, -7, 5,
    -- filter=12 channel=53
    -5, -6, 5, 0, 2, -1, 12, 0, -4,
    -- filter=12 channel=54
    -4, -5, 3, -2, 4, 0, -5, 0, 4,
    -- filter=12 channel=55
    0, -16, -1, 10, 0, -19, 31, 5, -10,
    -- filter=12 channel=56
    8, 0, 2, 0, 4, -1, -3, -2, -5,
    -- filter=12 channel=57
    -5, -6, -3, -3, -7, -7, 0, 2, 2,
    -- filter=12 channel=58
    -4, 8, -3, -1, -1, 4, -12, 2, -3,
    -- filter=12 channel=59
    3, -6, 6, 9, 9, -4, 7, -2, -2,
    -- filter=12 channel=60
    0, 0, -7, 2, -1, -4, -2, 1, 3,
    -- filter=12 channel=61
    2, 0, 2, -3, 1, 0, -1, -4, -2,
    -- filter=12 channel=62
    3, 3, -3, -4, -5, 3, -4, -3, -5,
    -- filter=12 channel=63
    0, 1, -2, -8, -1, 3, -6, 5, -2,
    -- filter=12 channel=64
    4, 0, -8, 6, 3, -1, 2, 5, -4,
    -- filter=12 channel=65
    -1, -3, 3, -7, -6, 0, 5, 5, -6,
    -- filter=12 channel=66
    -6, -3, 10, 5, 0, 2, 4, -3, 4,
    -- filter=12 channel=67
    -5, -4, -4, -2, 0, 4, 6, -2, -3,
    -- filter=12 channel=68
    7, -6, 3, 0, -5, 2, 11, -3, -6,
    -- filter=12 channel=69
    -2, 6, -2, 2, 2, 7, -4, -3, 1,
    -- filter=12 channel=70
    -8, -3, 1, 8, -15, -10, 8, -5, -10,
    -- filter=12 channel=71
    2, 2, -3, -1, -2, 0, 5, -2, -2,
    -- filter=12 channel=72
    -3, -5, 10, 4, 6, 8, 10, -7, 3,
    -- filter=12 channel=73
    -3, 0, -10, 15, -7, -10, 22, 6, -5,
    -- filter=12 channel=74
    -8, 0, -6, 6, -6, 0, 1, -11, 4,
    -- filter=12 channel=75
    1, -9, 7, -17, -5, 11, -3, -10, 7,
    -- filter=12 channel=76
    -5, -1, -10, 18, -3, -10, 23, 14, -9,
    -- filter=12 channel=77
    6, 6, -3, 7, 4, 0, 3, -4, 3,
    -- filter=12 channel=78
    2, 5, 5, 0, -6, -5, -3, -6, 2,
    -- filter=12 channel=79
    -4, -14, -2, 20, -7, -23, 37, 4, -10,
    -- filter=12 channel=80
    -9, -4, 5, -9, 2, 14, 4, -5, 0,
    -- filter=12 channel=81
    2, 1, 4, -5, 0, 0, -4, -6, 0,
    -- filter=12 channel=82
    -2, 6, 0, 0, -5, 3, -6, -8, -3,
    -- filter=12 channel=83
    1, 0, 2, 3, -3, 7, 4, -5, -1,
    -- filter=12 channel=84
    -2, -1, -3, 4, -1, -13, 6, 9, -7,
    -- filter=12 channel=85
    -1, -1, -4, 5, -3, -2, 4, -5, -3,
    -- filter=12 channel=86
    -3, 5, 8, 3, 0, 0, -8, -9, 0,
    -- filter=12 channel=87
    -5, -5, -2, 4, -4, -7, 3, 7, -3,
    -- filter=12 channel=88
    0, -5, -9, -3, -4, -5, -4, -5, -8,
    -- filter=12 channel=89
    -8, -2, 0, 8, 4, -10, 12, 7, -1,
    -- filter=12 channel=90
    -4, 3, 7, -13, 4, 6, -8, -7, -2,
    -- filter=12 channel=91
    1, -2, 2, 16, -12, -9, 19, -7, -4,
    -- filter=12 channel=92
    5, 0, 7, 2, -5, -8, 0, 3, 4,
    -- filter=12 channel=93
    -2, 7, 2, -12, 5, 2, -8, 3, 9,
    -- filter=12 channel=94
    5, 5, -4, -4, 0, 3, 0, -6, 2,
    -- filter=12 channel=95
    4, -8, 6, -5, 0, 3, 0, 0, -3,
    -- filter=12 channel=96
    6, -4, 1, -5, 0, 0, 0, 7, -6,
    -- filter=12 channel=97
    -1, 6, 6, -11, -3, -1, 0, -12, 0,
    -- filter=12 channel=98
    -4, 0, 2, 0, 1, -6, 7, -7, 1,
    -- filter=12 channel=99
    -13, -1, 0, 2, 4, -1, 12, 0, -9,
    -- filter=12 channel=100
    -1, 5, -5, 2, -7, 5, 2, -3, 1,
    -- filter=12 channel=101
    2, 4, -6, -2, -8, 3, 4, 0, 2,
    -- filter=12 channel=102
    3, 1, -6, 2, 2, 2, -5, -2, -1,
    -- filter=12 channel=103
    -6, 13, 8, -12, 6, 12, -17, -6, 5,
    -- filter=12 channel=104
    2, 0, 2, 3, 2, 3, 2, -8, -5,
    -- filter=12 channel=105
    -2, 2, 0, 11, -2, -7, 9, 10, -7,
    -- filter=12 channel=106
    7, -8, -2, 3, -1, 1, 11, 3, -10,
    -- filter=12 channel=107
    0, -5, -10, 2, -12, -9, 18, 1, -12,
    -- filter=12 channel=108
    -3, 4, -6, 6, -5, -5, 4, -4, 7,
    -- filter=12 channel=109
    -10, -1, 0, 10, -4, -2, 23, 2, 2,
    -- filter=12 channel=110
    -7, -7, -3, -9, 5, 0, -2, 1, -7,
    -- filter=12 channel=111
    10, -4, -7, 0, 4, -7, -1, -3, 6,
    -- filter=12 channel=112
    -1, 3, 9, 3, -7, 2, 3, -11, 2,
    -- filter=12 channel=113
    -11, -10, 0, -7, 0, -5, 6, -1, 5,
    -- filter=12 channel=114
    -4, -12, -10, 14, -15, -8, 29, 9, -1,
    -- filter=12 channel=115
    -3, -6, -2, 3, -3, 0, 1, -6, 7,
    -- filter=12 channel=116
    -4, -9, -1, 14, 7, -2, 22, 0, -7,
    -- filter=12 channel=117
    -7, 4, 2, -2, 2, -2, 5, -5, -1,
    -- filter=12 channel=118
    2, -2, -1, -3, 7, -6, -3, 3, 0,
    -- filter=12 channel=119
    1, -2, -5, -7, -7, -6, -9, 0, 4,
    -- filter=12 channel=120
    -9, -8, -5, 8, -6, -6, 16, -2, 1,
    -- filter=12 channel=121
    2, 2, 5, 4, -1, -4, -3, -6, -1,
    -- filter=12 channel=122
    -5, 11, 15, -26, 8, 15, -26, -13, 5,
    -- filter=12 channel=123
    0, -1, -4, 0, 0, 4, 0, 5, 0,
    -- filter=12 channel=124
    0, 4, 0, 0, -1, -8, 14, -1, 3,
    -- filter=12 channel=125
    -2, 1, 8, -4, 1, -5, 3, 1, 0,
    -- filter=12 channel=126
    0, -7, -5, -1, -1, -9, 13, -4, 0,
    -- filter=12 channel=127
    6, -4, -3, -1, 3, 3, -2, -1, 7,
    -- filter=13 channel=0
    13, 10, 13, -11, -5, 2, -17, -6, -2,
    -- filter=13 channel=1
    14, 13, 2, -5, -5, 9, -22, -11, -13,
    -- filter=13 channel=2
    -3, 0, -1, 0, 4, -5, 0, -2, -3,
    -- filter=13 channel=3
    -14, -11, -8, -11, 0, -8, 2, 6, 14,
    -- filter=13 channel=4
    0, 1, 5, -11, 0, -3, 0, 3, 4,
    -- filter=13 channel=5
    1, 5, 11, -1, -1, -1, -16, -7, -1,
    -- filter=13 channel=6
    2, -6, -4, -5, 2, 3, -1, 9, 8,
    -- filter=13 channel=7
    0, 0, 5, -3, 4, 6, -7, -6, -3,
    -- filter=13 channel=8
    4, 0, -8, -12, -12, -11, 0, 0, -6,
    -- filter=13 channel=9
    7, 8, 2, 7, 11, -3, 7, 2, -4,
    -- filter=13 channel=10
    4, -6, -10, 7, 7, -9, 0, 10, -1,
    -- filter=13 channel=11
    -8, -11, -8, 8, 5, 1, 15, 8, 13,
    -- filter=13 channel=12
    3, -11, -8, -6, -4, 0, -7, 3, -10,
    -- filter=13 channel=13
    -4, -16, -18, 9, -2, -5, 12, 11, -8,
    -- filter=13 channel=14
    0, 2, -1, 4, 7, -5, 7, -2, 6,
    -- filter=13 channel=15
    -4, -12, -17, 8, -6, -5, 13, 13, 5,
    -- filter=13 channel=16
    -3, -2, 2, -9, -2, 1, -12, 1, -6,
    -- filter=13 channel=17
    0, -2, 7, -2, -6, 0, -7, 3, -1,
    -- filter=13 channel=18
    1, -2, -17, 6, 8, -4, 18, 3, 4,
    -- filter=13 channel=19
    2, -3, -3, 6, 7, -1, 4, -2, 5,
    -- filter=13 channel=20
    -3, -6, -1, 2, -6, -2, 23, 7, 13,
    -- filter=13 channel=21
    0, 9, 10, 3, 8, 1, -15, 2, -9,
    -- filter=13 channel=22
    -1, -2, 0, -2, -5, -13, 0, 1, -5,
    -- filter=13 channel=23
    -13, -31, -27, 7, -12, -22, 22, 6, -14,
    -- filter=13 channel=24
    5, -1, 0, 2, 2, 1, 4, -7, -1,
    -- filter=13 channel=25
    14, -1, -7, 11, 16, 1, -5, 7, -10,
    -- filter=13 channel=26
    2, 7, 10, -1, -2, -2, 0, -1, 0,
    -- filter=13 channel=27
    8, -11, -29, 22, 9, -7, 15, 13, -10,
    -- filter=13 channel=28
    0, -5, 0, 3, 5, 1, -4, -7, -6,
    -- filter=13 channel=29
    6, -12, 1, 12, -6, 6, 24, 18, 11,
    -- filter=13 channel=30
    6, 4, 4, -4, 12, 4, -4, 8, 3,
    -- filter=13 channel=31
    -12, -21, -14, 15, 9, -6, 5, 8, -3,
    -- filter=13 channel=32
    -2, -10, -19, 12, 4, -8, 14, 13, 2,
    -- filter=13 channel=33
    -4, -18, -10, 4, 3, -3, 9, 2, -2,
    -- filter=13 channel=34
    -14, -23, -15, -6, -26, -7, 4, -5, -6,
    -- filter=13 channel=35
    2, 6, 5, 1, 0, -6, 7, 5, -7,
    -- filter=13 channel=36
    -5, -13, -6, -3, 1, -2, 0, -8, -11,
    -- filter=13 channel=37
    11, 18, 17, -4, -3, 1, -26, -14, -2,
    -- filter=13 channel=38
    -1, -9, -5, 13, -1, -1, 5, 12, -3,
    -- filter=13 channel=39
    -5, -2, 5, -5, 5, 4, 5, 6, 12,
    -- filter=13 channel=40
    -11, -13, 0, 5, -5, -9, 6, 2, 2,
    -- filter=13 channel=41
    5, 0, -1, -3, -10, -16, 0, -6, -11,
    -- filter=13 channel=42
    0, 12, -2, 2, -1, 6, -7, -3, 3,
    -- filter=13 channel=43
    -1, -11, 0, -2, -12, -10, -3, 4, 1,
    -- filter=13 channel=44
    -1, 9, 4, 0, 7, -4, -15, -13, -6,
    -- filter=13 channel=45
    0, 5, 3, -4, -1, 5, -8, 3, -1,
    -- filter=13 channel=46
    0, 4, -4, -6, -7, -1, -3, 2, 6,
    -- filter=13 channel=47
    -3, 7, 7, 6, 17, 4, -20, -7, 0,
    -- filter=13 channel=48
    18, 10, -3, 11, 21, 0, -7, 2, -9,
    -- filter=13 channel=49
    0, 1, -8, 4, -2, -3, 10, 0, 4,
    -- filter=13 channel=50
    5, -1, -16, 16, 9, -7, 6, -1, -1,
    -- filter=13 channel=51
    6, 1, -4, -4, 6, 6, 2, -3, 4,
    -- filter=13 channel=52
    -2, -8, -5, -7, -10, -14, -7, 3, -7,
    -- filter=13 channel=53
    1, -12, 1, 2, 2, -5, 10, 4, -2,
    -- filter=13 channel=54
    -6, -1, -3, 4, 2, 6, 0, 5, -4,
    -- filter=13 channel=55
    3, -23, -22, 11, 0, -18, 18, 7, 1,
    -- filter=13 channel=56
    -8, -6, -4, 0, -1, -5, 6, 1, -7,
    -- filter=13 channel=57
    -4, 0, 0, -4, 2, 4, -3, 4, -5,
    -- filter=13 channel=58
    -4, 10, 16, -13, 1, 0, -15, -9, 6,
    -- filter=13 channel=59
    10, 7, -18, 7, 20, -4, -3, 6, -10,
    -- filter=13 channel=60
    1, 0, 7, 0, -6, -7, -5, -3, -3,
    -- filter=13 channel=61
    -3, -6, 0, -8, 0, -4, -3, 4, -6,
    -- filter=13 channel=62
    -1, -7, -5, 4, 5, 1, 3, 0, 6,
    -- filter=13 channel=63
    -1, 4, 17, 0, 8, 12, -8, -3, 5,
    -- filter=13 channel=64
    1, -13, 0, -8, 3, -10, -4, -4, -2,
    -- filter=13 channel=65
    -4, 1, -4, -1, 2, 1, -3, 3, -6,
    -- filter=13 channel=66
    -6, -2, -5, -5, 0, -10, 2, -8, -6,
    -- filter=13 channel=67
    4, 0, 3, -2, 0, -9, -5, -5, 2,
    -- filter=13 channel=68
    0, 0, 3, 1, -7, -2, 8, 0, 4,
    -- filter=13 channel=69
    8, 8, 3, -6, 6, 0, 0, 5, -5,
    -- filter=13 channel=70
    -6, -23, -12, 1, -8, -17, 0, 1, -10,
    -- filter=13 channel=71
    -2, -6, -2, -6, -8, -3, 4, -7, 0,
    -- filter=13 channel=72
    -1, -16, -20, 14, 10, -8, 3, 14, 3,
    -- filter=13 channel=73
    0, 0, -12, 11, 1, -9, 10, 1, 1,
    -- filter=13 channel=74
    -10, -10, -8, 2, -4, -4, 4, -4, -12,
    -- filter=13 channel=75
    -7, -2, 10, -3, -5, 0, -25, -1, 4,
    -- filter=13 channel=76
    -6, -9, -12, -6, -13, 0, 15, 7, 8,
    -- filter=13 channel=77
    6, -6, -4, 0, 1, 3, 1, 0, 2,
    -- filter=13 channel=78
    -4, 9, 5, 1, 4, -2, 1, 5, -4,
    -- filter=13 channel=79
    0, -9, -24, 13, 2, -14, 18, 15, 0,
    -- filter=13 channel=80
    6, 2, -7, 10, 27, 6, -4, 11, -10,
    -- filter=13 channel=81
    -3, 1, 3, -4, -3, 5, -1, -3, -3,
    -- filter=13 channel=82
    -2, 4, -6, 1, 0, 1, -1, -6, 3,
    -- filter=13 channel=83
    7, 9, -8, 13, 10, -3, 6, 3, -3,
    -- filter=13 channel=84
    2, -3, -2, 8, 0, -6, 5, -2, -5,
    -- filter=13 channel=85
    1, -5, 0, 0, 1, 3, -3, -4, 6,
    -- filter=13 channel=86
    0, 1, 2, -6, -7, -1, -11, -2, -5,
    -- filter=13 channel=87
    -9, -13, 0, -1, -7, -10, 1, -4, 1,
    -- filter=13 channel=88
    -12, -7, -1, -9, -5, -2, 7, -5, -3,
    -- filter=13 channel=89
    0, -21, -25, 12, 0, -9, 16, 12, 2,
    -- filter=13 channel=90
    -16, -17, -5, -7, -13, -2, -7, 0, -8,
    -- filter=13 channel=91
    8, -8, -17, 10, -2, -12, 5, 5, -8,
    -- filter=13 channel=92
    -9, 1, -6, -8, -1, -6, 0, -2, -3,
    -- filter=13 channel=93
    3, 10, 16, -5, 13, 14, -10, -13, -5,
    -- filter=13 channel=94
    -5, -4, 5, -2, 5, 2, 3, 2, -3,
    -- filter=13 channel=95
    2, -5, 5, -7, 4, -2, -2, -3, -4,
    -- filter=13 channel=96
    2, 6, 0, -1, 8, 2, -1, 2, -3,
    -- filter=13 channel=97
    -15, -3, -2, -4, -3, -4, 2, -1, 0,
    -- filter=13 channel=98
    -1, -6, -17, 19, 22, 3, 10, 10, -8,
    -- filter=13 channel=99
    -4, -29, -25, 14, -2, -16, 16, 1, -8,
    -- filter=13 channel=100
    -2, -6, -5, 5, 0, 0, -3, 1, -10,
    -- filter=13 channel=101
    5, -6, 6, -10, 1, 2, 5, 1, 7,
    -- filter=13 channel=102
    -1, 3, 1, -2, -2, 3, 2, 2, 0,
    -- filter=13 channel=103
    -8, 2, 10, -5, 16, 11, -7, 4, 0,
    -- filter=13 channel=104
    9, 0, -5, 5, 12, 8, -2, 10, -5,
    -- filter=13 channel=105
    6, 3, 0, -2, 3, -3, 12, 7, 8,
    -- filter=13 channel=106
    -8, 0, -1, 0, -3, -6, 11, 1, 0,
    -- filter=13 channel=107
    -1, -3, 4, -5, -8, -1, 8, 6, 9,
    -- filter=13 channel=108
    0, -3, 9, 3, 0, -6, -8, 1, 1,
    -- filter=13 channel=109
    10, -6, -26, 23, 15, -4, 17, 1, -5,
    -- filter=13 channel=110
    -12, -4, 2, 4, -6, 4, 7, 1, 0,
    -- filter=13 channel=111
    6, 4, 1, -3, -7, -2, 8, 4, 4,
    -- filter=13 channel=112
    5, -10, -2, 0, -6, 1, 2, -2, -9,
    -- filter=13 channel=113
    -6, -17, -22, 1, 0, -8, 8, 8, -1,
    -- filter=13 channel=114
    20, 1, 0, 1, -1, -1, 1, 1, -1,
    -- filter=13 channel=115
    0, 3, 4, -4, 6, -3, -5, -2, 2,
    -- filter=13 channel=116
    13, 0, -6, 8, 6, 1, 14, 6, 2,
    -- filter=13 channel=117
    -7, -3, -6, 0, 8, 2, -4, 0, 2,
    -- filter=13 channel=118
    5, -6, 1, 1, 3, -6, 3, -4, -6,
    -- filter=13 channel=119
    -2, -15, -16, -8, -9, -12, -5, -7, -18,
    -- filter=13 channel=120
    -4, -27, -25, 17, -4, -10, 19, 9, -16,
    -- filter=13 channel=121
    2, -12, -10, 9, 0, -9, 7, -4, 2,
    -- filter=13 channel=122
    2, 4, 12, 0, 18, -1, -18, -15, -19,
    -- filter=13 channel=123
    -5, -14, -13, -2, -15, -4, -4, -5, -9,
    -- filter=13 channel=124
    7, -5, -7, -4, 5, -6, 0, 12, 2,
    -- filter=13 channel=125
    1, -15, -15, 15, 15, -2, 11, 12, -8,
    -- filter=13 channel=126
    -7, -4, -14, 8, -3, -4, 9, 5, 8,
    -- filter=13 channel=127
    -5, 0, -5, 4, -3, -8, 0, 3, 0,
    -- filter=14 channel=0
    3, 0, 3, -7, -18, 12, -11, -13, 7,
    -- filter=14 channel=1
    -3, -2, 11, -9, -15, 7, 0, -13, 4,
    -- filter=14 channel=2
    6, -2, -4, 2, -1, -7, 1, -2, -1,
    -- filter=14 channel=3
    -6, 8, -7, -3, -2, -4, 0, 3, 0,
    -- filter=14 channel=4
    -2, -6, -3, 4, -4, 0, 8, 0, 7,
    -- filter=14 channel=5
    -1, -6, 4, 1, -5, 6, 7, -12, 8,
    -- filter=14 channel=6
    -1, 0, -1, -4, -2, 1, -7, -6, 0,
    -- filter=14 channel=7
    7, -2, -7, -3, -1, -6, 0, -5, 0,
    -- filter=14 channel=8
    4, 9, -3, -5, -4, -4, 2, 0, 4,
    -- filter=14 channel=9
    4, -3, 0, 3, -4, -1, -1, 0, 6,
    -- filter=14 channel=10
    1, -4, -5, -4, 6, 3, 0, 0, 0,
    -- filter=14 channel=11
    -6, 0, 2, 1, 8, 0, -7, 0, 2,
    -- filter=14 channel=12
    -6, 7, 5, -2, 0, -2, 0, 10, 6,
    -- filter=14 channel=13
    0, 0, 1, -2, -2, -5, -5, 4, 2,
    -- filter=14 channel=14
    4, 4, -6, 4, 1, 6, 1, 3, 3,
    -- filter=14 channel=15
    -9, -5, 13, -11, 4, 0, -7, 0, -3,
    -- filter=14 channel=16
    7, -3, -2, 0, 1, 5, 5, -4, -5,
    -- filter=14 channel=17
    6, 1, 0, -2, 3, 3, -7, 3, -2,
    -- filter=14 channel=18
    -10, 0, 12, -4, -10, 0, -8, -6, 4,
    -- filter=14 channel=19
    0, 2, -1, -4, -5, 4, 2, -4, 0,
    -- filter=14 channel=20
    -1, 8, 11, -2, 5, 4, -6, 2, -7,
    -- filter=14 channel=21
    8, -7, 3, 5, 0, -2, 8, 4, -5,
    -- filter=14 channel=22
    -5, 8, 8, -3, 4, 3, -3, 1, 4,
    -- filter=14 channel=23
    -2, 12, 14, -12, -3, 4, -4, 4, -4,
    -- filter=14 channel=24
    0, 3, 0, -5, 3, 5, 6, -3, 0,
    -- filter=14 channel=25
    -6, -8, 11, 0, -11, 5, 5, 1, 7,
    -- filter=14 channel=26
    9, 5, -1, 2, -4, 2, 1, -5, 1,
    -- filter=14 channel=27
    -14, -13, 27, -14, -20, 4, 3, -8, 9,
    -- filter=14 channel=28
    1, -1, 6, -1, -6, 5, -3, 4, 4,
    -- filter=14 channel=29
    -1, 9, 0, 4, 14, -9, -1, 5, 2,
    -- filter=14 channel=30
    2, -8, 2, -1, -11, 7, 6, 0, 8,
    -- filter=14 channel=31
    -4, 0, 1, -5, -9, -5, 4, -6, 3,
    -- filter=14 channel=32
    -10, -7, 7, -5, -12, 10, 3, -7, 3,
    -- filter=14 channel=33
    -4, -3, 3, -8, -12, 0, 0, -5, 6,
    -- filter=14 channel=34
    2, 11, 12, 4, 0, 20, -8, -2, 13,
    -- filter=14 channel=35
    0, 0, -2, -4, 2, 4, 3, -6, 4,
    -- filter=14 channel=36
    8, 5, -10, -2, 7, -6, 9, 8, 2,
    -- filter=14 channel=37
    -2, -8, -3, -1, -19, -1, -3, -14, 7,
    -- filter=14 channel=38
    -6, 3, 9, -8, 3, 1, 3, -7, 0,
    -- filter=14 channel=39
    3, 2, -7, 5, 7, -5, 4, 7, -7,
    -- filter=14 channel=40
    -5, -3, 0, -6, 9, 8, -1, 6, -4,
    -- filter=14 channel=41
    8, 2, 1, -2, -1, 6, 9, 14, 13,
    -- filter=14 channel=42
    3, -8, 6, 1, -10, 1, 5, 0, -8,
    -- filter=14 channel=43
    -7, 7, -3, -8, -6, 8, -3, -4, 1,
    -- filter=14 channel=44
    -6, -11, 9, -3, -8, 3, -7, -10, 3,
    -- filter=14 channel=45
    7, 7, -1, -2, 0, -4, -7, 3, -1,
    -- filter=14 channel=46
    -1, 0, -1, 6, 0, -3, 0, 2, 2,
    -- filter=14 channel=47
    0, -11, -3, 4, -14, -1, 7, -5, -6,
    -- filter=14 channel=48
    -6, -12, 0, 3, 0, -1, -1, -3, 7,
    -- filter=14 channel=49
    -3, 5, 5, -1, -8, -1, 2, 8, 9,
    -- filter=14 channel=50
    -6, -8, 11, -7, -11, 1, 3, -7, 8,
    -- filter=14 channel=51
    0, -5, -6, -6, -6, 3, 3, 0, -3,
    -- filter=14 channel=52
    -5, 1, -2, -1, 3, 10, -11, 0, -2,
    -- filter=14 channel=53
    -4, 9, -1, -1, 7, 2, -6, 0, -2,
    -- filter=14 channel=54
    6, -6, 4, 1, 6, -3, -3, -7, 0,
    -- filter=14 channel=55
    -9, -4, 4, -5, 3, -1, -5, 5, -6,
    -- filter=14 channel=56
    -3, 0, 3, 4, -3, 8, 6, 4, 4,
    -- filter=14 channel=57
    4, 3, -4, 4, 8, 2, -2, 8, 1,
    -- filter=14 channel=58
    7, 1, -1, 2, -9, -2, -1, -8, 7,
    -- filter=14 channel=59
    0, -13, 11, 7, -2, 2, 10, -3, 5,
    -- filter=14 channel=60
    6, -1, 2, 4, 0, 0, 2, -4, -3,
    -- filter=14 channel=61
    -1, -1, -7, 0, -2, -2, -2, 7, 2,
    -- filter=14 channel=62
    2, -5, 5, 5, 6, 0, -3, -6, 2,
    -- filter=14 channel=63
    5, 2, 9, 9, -2, 2, 9, 2, 7,
    -- filter=14 channel=64
    -5, 0, 0, 4, 5, -1, 0, -2, -4,
    -- filter=14 channel=65
    0, 2, 0, -5, 6, -2, -1, 2, -5,
    -- filter=14 channel=66
    -4, 2, 0, 0, 2, 9, 2, 6, 8,
    -- filter=14 channel=67
    2, 4, 2, 3, -1, -5, 3, -1, -3,
    -- filter=14 channel=68
    5, -4, -2, 6, 0, -3, 8, -4, 4,
    -- filter=14 channel=69
    4, -2, 2, -6, 4, 7, 0, -2, -1,
    -- filter=14 channel=70
    -10, 4, 7, -11, -2, 9, -10, -5, 5,
    -- filter=14 channel=71
    8, -4, -8, 2, 3, -7, -3, -4, 3,
    -- filter=14 channel=72
    -1, -1, 4, 9, 3, 0, 3, -1, 0,
    -- filter=14 channel=73
    1, 0, 1, -2, -4, -5, 2, -3, 3,
    -- filter=14 channel=74
    -3, 7, 16, -9, -10, 5, -3, 0, 14,
    -- filter=14 channel=75
    -10, -3, 6, 1, -12, 0, 6, -7, -2,
    -- filter=14 channel=76
    1, 7, -6, 1, 15, -5, -8, -1, 0,
    -- filter=14 channel=77
    7, -3, 5, 5, 8, -3, -3, 1, 0,
    -- filter=14 channel=78
    8, -3, 3, 3, 3, -4, -3, 0, 6,
    -- filter=14 channel=79
    -11, 0, 20, -2, -9, 10, -7, -6, 5,
    -- filter=14 channel=80
    -6, -9, -5, 5, -1, -2, 10, -9, -3,
    -- filter=14 channel=81
    -5, -6, -4, -4, -1, 3, -4, 7, -4,
    -- filter=14 channel=82
    3, 3, -3, 1, -3, 6, -7, -1, 2,
    -- filter=14 channel=83
    5, -3, -1, 7, -2, -3, 0, -5, 4,
    -- filter=14 channel=84
    -6, 5, 8, -1, 5, -2, -1, 0, 3,
    -- filter=14 channel=85
    -5, 1, 3, 4, -6, -5, 1, -2, -3,
    -- filter=14 channel=86
    -6, 0, 6, 1, -2, 4, -7, 7, 2,
    -- filter=14 channel=87
    4, 9, 2, -1, -3, 6, -6, 5, 5,
    -- filter=14 channel=88
    2, 7, -2, -2, 11, 1, 8, -1, 8,
    -- filter=14 channel=89
    1, -11, 7, 5, -2, 0, 9, 6, -11,
    -- filter=14 channel=90
    0, 6, 0, 4, 12, -1, 3, 1, -4,
    -- filter=14 channel=91
    -8, -8, 15, -7, 1, -1, 0, -7, -1,
    -- filter=14 channel=92
    -3, 8, 4, -7, 6, 1, -7, -1, 0,
    -- filter=14 channel=93
    3, -14, 0, -3, -12, -8, 5, -2, 3,
    -- filter=14 channel=94
    2, 6, -6, -5, 1, 1, 4, -6, -6,
    -- filter=14 channel=95
    5, 1, 1, 5, 1, -4, -1, -1, -3,
    -- filter=14 channel=96
    2, -6, 6, 6, -3, 4, 1, 0, -4,
    -- filter=14 channel=97
    5, 3, -8, -6, -5, 0, 0, -6, -8,
    -- filter=14 channel=98
    -5, -4, 14, -2, -15, -2, 2, -12, 4,
    -- filter=14 channel=99
    -5, 2, -2, 3, 1, -2, 0, 4, 7,
    -- filter=14 channel=100
    -5, 10, 8, 0, -4, -2, 3, 0, 7,
    -- filter=14 channel=101
    7, 0, -5, 2, 0, 2, 8, 2, 0,
    -- filter=14 channel=102
    -5, 2, 2, 4, 6, 5, -3, -2, -3,
    -- filter=14 channel=103
    -4, -11, 6, 7, -11, 4, 0, -4, -5,
    -- filter=14 channel=104
    5, -13, -5, 2, 3, -1, 11, 1, 5,
    -- filter=14 channel=105
    3, 8, 8, -3, 1, 4, -4, 5, -10,
    -- filter=14 channel=106
    -1, -4, 1, -5, -3, 3, -3, 4, 0,
    -- filter=14 channel=107
    -9, 5, 8, -8, 2, 11, -3, 2, 1,
    -- filter=14 channel=108
    5, 7, -2, -3, 3, -2, -5, -5, -3,
    -- filter=14 channel=109
    -4, 1, 10, -3, -8, 10, -6, 3, 6,
    -- filter=14 channel=110
    -6, 5, -6, 5, -4, -1, 2, 2, -10,
    -- filter=14 channel=111
    6, 6, -3, -1, -1, 9, 6, -3, 0,
    -- filter=14 channel=112
    -3, -5, 16, -3, -8, 5, -1, 3, 0,
    -- filter=14 channel=113
    -10, 0, 6, 3, 1, 10, -1, -6, -5,
    -- filter=14 channel=114
    -7, -9, 19, -12, -15, 2, -6, -11, 11,
    -- filter=14 channel=115
    0, 0, -1, 0, -3, -6, 3, -5, 1,
    -- filter=14 channel=116
    2, -7, 0, 2, 0, 0, 7, 4, 0,
    -- filter=14 channel=117
    -1, -7, 5, 5, -6, -9, 7, 0, -1,
    -- filter=14 channel=118
    -6, -4, 5, -5, -3, 3, -6, -1, 0,
    -- filter=14 channel=119
    -5, 14, 14, -6, 0, 17, -7, 8, 13,
    -- filter=14 channel=120
    -11, 8, 11, -11, -6, 0, 0, 0, 11,
    -- filter=14 channel=121
    -6, 0, 3, 5, -6, -6, 0, 8, 4,
    -- filter=14 channel=122
    4, -15, 0, 1, -7, -2, 3, -7, 0,
    -- filter=14 channel=123
    1, -1, 5, 1, 5, 13, 1, 7, -2,
    -- filter=14 channel=124
    0, -1, 6, 4, 7, 2, -1, -3, -2,
    -- filter=14 channel=125
    -6, -4, 8, 8, 1, -9, 0, -2, -4,
    -- filter=14 channel=126
    7, -5, 5, 7, -5, 0, 3, -1, 1,
    -- filter=14 channel=127
    -4, 0, -5, -4, 6, 8, 0, 8, -1,
    -- filter=15 channel=0
    14, 11, -5, 3, 4, -12, 0, -5, -17,
    -- filter=15 channel=1
    7, 9, 2, 2, 3, -8, -2, -5, -16,
    -- filter=15 channel=2
    0, -9, -6, 3, -3, -5, 8, 11, -1,
    -- filter=15 channel=3
    3, 0, 4, 0, -1, 1, -2, 3, -3,
    -- filter=15 channel=4
    -12, 0, 2, -4, 0, -2, 14, 9, 17,
    -- filter=15 channel=5
    1, 5, -4, 1, 12, -7, -8, -6, -6,
    -- filter=15 channel=6
    -6, -10, -4, -2, 2, 4, 1, 1, 4,
    -- filter=15 channel=7
    -5, -4, -5, 0, 5, 1, 5, -6, -2,
    -- filter=15 channel=8
    -6, -8, 4, 1, -1, -3, -1, 6, -3,
    -- filter=15 channel=9
    4, -4, -7, -4, 11, 0, -5, 5, -1,
    -- filter=15 channel=10
    3, 1, -5, -7, 0, 6, -3, -1, 6,
    -- filter=15 channel=11
    -4, -8, 0, -2, 0, 2, 7, 1, 2,
    -- filter=15 channel=12
    6, 1, 9, -1, -1, 2, -6, -4, 4,
    -- filter=15 channel=13
    0, -17, 1, -8, -11, -7, -3, 3, 5,
    -- filter=15 channel=14
    6, -5, 3, -4, -1, -3, -7, 0, -3,
    -- filter=15 channel=15
    5, -15, -3, 4, -5, -6, 14, 7, 3,
    -- filter=15 channel=16
    0, -1, 5, -5, -4, 4, -11, -1, -1,
    -- filter=15 channel=17
    0, 5, -3, 1, -7, 2, 4, -7, 0,
    -- filter=15 channel=18
    -2, -3, -9, -2, -9, 0, 9, 6, 17,
    -- filter=15 channel=19
    -7, 0, -5, -6, 3, 0, -7, 0, 4,
    -- filter=15 channel=20
    -8, -7, -8, 2, -1, 3, 4, 4, 4,
    -- filter=15 channel=21
    7, 11, 7, -4, 3, 0, -10, -2, -9,
    -- filter=15 channel=22
    6, 3, -4, -1, -9, -9, 0, -2, -4,
    -- filter=15 channel=23
    -3, -18, -18, -11, -4, -12, 5, 13, 4,
    -- filter=15 channel=24
    7, -2, 4, 0, 0, -6, 1, 7, -7,
    -- filter=15 channel=25
    2, -12, -2, 4, 4, 2, 9, 3, 2,
    -- filter=15 channel=26
    3, 11, 0, 2, 8, -4, -2, -2, -1,
    -- filter=15 channel=27
    -4, -7, -7, 7, -3, -6, 14, 18, 12,
    -- filter=15 channel=28
    -2, -5, -4, 2, -5, 6, -5, 3, 2,
    -- filter=15 channel=29
    -6, -10, -3, -10, -3, -1, 0, 15, 17,
    -- filter=15 channel=30
    0, 0, 1, 9, 5, -1, 2, 11, 3,
    -- filter=15 channel=31
    -11, 1, -8, -4, 9, 3, -3, 7, 0,
    -- filter=15 channel=32
    -2, -17, -11, 4, -1, -6, 6, 11, 4,
    -- filter=15 channel=33
    -3, -6, -2, 0, -2, -8, 4, 5, 3,
    -- filter=15 channel=34
    1, 0, -2, 0, -6, -13, -2, -10, -16,
    -- filter=15 channel=35
    6, -5, 4, -4, -4, -3, -3, -4, 3,
    -- filter=15 channel=36
    -2, -8, 3, 0, -2, 8, 0, 0, -3,
    -- filter=15 channel=37
    4, 2, -3, 0, 4, 3, 2, -3, -18,
    -- filter=15 channel=38
    4, -10, -3, -1, -4, -5, 4, 8, 6,
    -- filter=15 channel=39
    1, -1, 1, 2, -3, 3, 4, 0, 3,
    -- filter=15 channel=40
    -7, 3, 4, -2, 1, -5, -6, 0, -1,
    -- filter=15 channel=41
    5, -4, -7, 0, -11, 0, 0, -10, 1,
    -- filter=15 channel=42
    -1, -3, -1, 0, 7, -1, 1, 1, -3,
    -- filter=15 channel=43
    2, -5, -6, 5, -2, -4, 3, 8, 0,
    -- filter=15 channel=44
    -5, 10, 8, -1, 3, 0, -10, 2, -12,
    -- filter=15 channel=45
    3, 7, -6, 3, 2, 6, -7, 4, 5,
    -- filter=15 channel=46
    7, 0, -6, 0, 3, 1, -2, 3, -2,
    -- filter=15 channel=47
    -4, 11, 1, 2, 3, 5, -10, -2, -6,
    -- filter=15 channel=48
    -9, 4, -3, 0, 17, 1, -5, 3, 6,
    -- filter=15 channel=49
    1, 0, -2, 3, 4, 3, 8, 15, 12,
    -- filter=15 channel=50
    -9, -8, -7, 4, -2, 1, -1, 13, -3,
    -- filter=15 channel=51
    5, 4, 2, 0, -1, 5, 6, -3, 5,
    -- filter=15 channel=52
    -5, -7, -8, -1, -6, -2, 8, 0, 2,
    -- filter=15 channel=53
    4, -6, 0, 0, 3, -2, 8, 4, 12,
    -- filter=15 channel=54
    -6, 1, 1, 0, 5, -7, -4, 5, -5,
    -- filter=15 channel=55
    -7, -10, -2, 1, -15, -10, 14, 16, 18,
    -- filter=15 channel=56
    5, 0, -10, -5, 0, -10, 4, -8, -6,
    -- filter=15 channel=57
    -2, 1, 4, -5, 6, 6, 1, 0, 8,
    -- filter=15 channel=58
    -4, 2, 1, 2, -2, 2, -4, 2, -10,
    -- filter=15 channel=59
    -1, 3, -1, -2, 9, 2, 1, 8, 1,
    -- filter=15 channel=60
    -3, 0, 6, 6, 0, 6, 5, -1, 1,
    -- filter=15 channel=61
    -6, 0, 5, 0, 1, -7, 0, -3, 0,
    -- filter=15 channel=62
    -3, 1, -3, 0, -4, -7, -6, 2, 3,
    -- filter=15 channel=63
    4, 0, -2, -3, 10, -2, -2, 0, 0,
    -- filter=15 channel=64
    0, 3, 4, -6, -7, 4, 6, -1, 4,
    -- filter=15 channel=65
    3, 5, -1, -5, 0, -3, 0, 6, -3,
    -- filter=15 channel=66
    2, -4, 3, 9, -5, -3, 6, 1, 4,
    -- filter=15 channel=67
    3, -5, 0, 3, 0, -3, -6, -3, -8,
    -- filter=15 channel=68
    0, -4, -3, 3, 2, 3, -1, 0, 0,
    -- filter=15 channel=69
    7, -5, 3, 1, -1, -4, 3, 4, 2,
    -- filter=15 channel=70
    -3, -3, -3, -1, -4, -15, 2, 10, -5,
    -- filter=15 channel=71
    -2, -2, 0, 4, 2, 0, -2, -4, 1,
    -- filter=15 channel=72
    -4, 5, -4, 0, 6, 5, 6, 11, 12,
    -- filter=15 channel=73
    3, -6, -10, -4, -6, -5, 2, 12, 3,
    -- filter=15 channel=74
    -11, 0, -6, 0, -3, -7, 3, 0, 0,
    -- filter=15 channel=75
    1, 8, -8, 11, 6, 3, -7, -11, -14,
    -- filter=15 channel=76
    2, -4, -3, -5, -7, -8, -4, 1, 8,
    -- filter=15 channel=77
    3, 2, -3, 3, 0, 3, -7, 0, -7,
    -- filter=15 channel=78
    5, 8, -1, 7, 3, 3, -7, 4, -6,
    -- filter=15 channel=79
    -5, -18, -12, -5, -5, -6, 11, 3, 7,
    -- filter=15 channel=80
    -3, 6, 8, -6, 13, 2, 3, 4, 11,
    -- filter=15 channel=81
    -2, 6, 0, 3, 5, 6, 2, -2, 1,
    -- filter=15 channel=82
    -3, 3, -7, -6, 0, -1, 2, 5, 0,
    -- filter=15 channel=83
    0, 3, 3, -5, 12, 1, 9, 8, 11,
    -- filter=15 channel=84
    -3, 0, -2, 6, -8, -8, 8, 14, 13,
    -- filter=15 channel=85
    5, 4, 3, 0, 5, -6, 2, -6, -3,
    -- filter=15 channel=86
    4, -7, -2, 6, 2, -1, -8, -3, -13,
    -- filter=15 channel=87
    4, -1, -6, 0, 1, -12, 7, 6, 3,
    -- filter=15 channel=88
    -4, 0, 4, 0, 8, -6, -5, 4, -1,
    -- filter=15 channel=89
    0, -13, -2, 2, -12, 6, 12, 2, 12,
    -- filter=15 channel=90
    0, -2, -9, -10, 3, -8, -7, 0, -7,
    -- filter=15 channel=91
    0, -5, -5, 3, -4, -5, 15, 18, 3,
    -- filter=15 channel=92
    0, -3, 2, -1, 3, -5, 3, -3, -8,
    -- filter=15 channel=93
    4, 14, 5, 3, 17, 7, -9, -7, -7,
    -- filter=15 channel=94
    6, 4, 0, 2, -2, -5, 4, -4, 0,
    -- filter=15 channel=95
    3, -1, 3, -6, 3, 1, 3, -2, -2,
    -- filter=15 channel=96
    6, 0, -3, 8, 2, -3, 7, 0, 5,
    -- filter=15 channel=97
    1, -4, -6, -4, 2, 0, -6, 4, -8,
    -- filter=15 channel=98
    0, -10, -9, 4, 7, 4, 6, 14, 15,
    -- filter=15 channel=99
    -14, -11, -11, -2, 8, -10, 2, 7, 9,
    -- filter=15 channel=100
    0, 0, 1, -3, 4, 2, 4, 6, 3,
    -- filter=15 channel=101
    -9, -9, -6, -4, -4, 0, 2, 15, 14,
    -- filter=15 channel=102
    -6, 5, -5, 0, 6, 0, -6, 5, -6,
    -- filter=15 channel=103
    0, 0, -2, -1, 8, 9, -14, -9, -10,
    -- filter=15 channel=104
    -1, 3, -3, -7, 15, 11, 3, 7, 6,
    -- filter=15 channel=105
    0, 4, 3, -5, -6, -7, -4, -3, 10,
    -- filter=15 channel=106
    0, 0, 3, -2, 1, 0, 1, -4, 2,
    -- filter=15 channel=107
    1, -13, -3, -3, -1, -14, 3, 1, 6,
    -- filter=15 channel=108
    7, 7, -1, -1, 4, 4, 5, -1, -6,
    -- filter=15 channel=109
    0, -11, -5, 6, 6, 1, 19, 8, 4,
    -- filter=15 channel=110
    -1, 0, 3, -1, 0, -6, 5, 0, 2,
    -- filter=15 channel=111
    -4, -1, -4, 6, -1, -5, 3, -4, -4,
    -- filter=15 channel=112
    5, 1, -3, -2, -3, -5, 9, 2, -9,
    -- filter=15 channel=113
    -3, -11, -7, 1, 2, -2, -1, 4, -4,
    -- filter=15 channel=114
    4, -10, -12, 8, -12, -10, 14, 11, -1,
    -- filter=15 channel=115
    6, -4, -2, 4, 4, -1, -3, 0, -6,
    -- filter=15 channel=116
    0, -1, 1, -2, 2, 10, 12, 11, 17,
    -- filter=15 channel=117
    4, -5, 7, 0, -2, 5, -4, 1, 3,
    -- filter=15 channel=118
    -1, 6, -5, -3, 6, 0, 3, -5, -1,
    -- filter=15 channel=119
    4, -9, -12, -1, -6, -9, 7, -11, -7,
    -- filter=15 channel=120
    -7, -17, -17, -1, 1, -4, 11, 29, 6,
    -- filter=15 channel=121
    -3, 0, 0, -3, -5, 4, -6, 3, 2,
    -- filter=15 channel=122
    7, 11, 3, -5, 8, 3, -23, 0, -14,
    -- filter=15 channel=123
    -7, -4, 1, -2, -4, -10, -3, -4, 0,
    -- filter=15 channel=124
    5, -5, -1, -5, 0, -1, 8, 1, 6,
    -- filter=15 channel=125
    -1, -10, -2, -1, 4, 1, 5, 16, 16,
    -- filter=15 channel=126
    9, 1, -3, -3, -2, 0, 6, 3, 0,
    -- filter=15 channel=127
    -2, -7, 2, 5, -8, 2, 6, -3, 0,
    -- filter=16 channel=0
    3, 6, 0, -10, 3, 1, 0, 0, 7,
    -- filter=16 channel=1
    3, -4, 9, -6, -10, 7, 0, -2, 7,
    -- filter=16 channel=2
    -5, 3, -3, -7, -1, 2, -5, 7, 3,
    -- filter=16 channel=3
    1, -7, -5, 6, 0, 4, -2, 0, 0,
    -- filter=16 channel=4
    -6, -8, 3, 7, 3, 2, 12, 8, 0,
    -- filter=16 channel=5
    8, 2, 3, -11, 0, 0, -4, 0, 0,
    -- filter=16 channel=6
    6, 0, 2, 1, -3, -5, -4, 7, -5,
    -- filter=16 channel=7
    0, 3, 7, 4, -2, -5, -4, -2, 2,
    -- filter=16 channel=8
    -2, 1, 1, 4, 8, 0, 3, 1, 3,
    -- filter=16 channel=9
    -6, -2, 2, -4, 2, -5, 1, 5, 3,
    -- filter=16 channel=10
    -9, -10, 3, -3, 7, 5, -5, 3, 4,
    -- filter=16 channel=11
    2, -9, 6, -3, -9, -3, 7, -7, 0,
    -- filter=16 channel=12
    2, 0, -3, 3, 2, -4, -4, -1, -4,
    -- filter=16 channel=13
    0, -3, 3, -13, 2, 6, 0, 1, 1,
    -- filter=16 channel=14
    4, 7, -4, 4, 0, 0, 2, 0, 4,
    -- filter=16 channel=15
    2, -4, -2, -5, -6, 1, 2, 1, 9,
    -- filter=16 channel=16
    -2, 4, 6, -13, 6, -2, -8, 8, 7,
    -- filter=16 channel=17
    4, -2, -6, 4, -5, 4, 2, -2, 3,
    -- filter=16 channel=18
    -1, -10, 2, -13, -13, 7, -4, -9, 3,
    -- filter=16 channel=19
    0, 3, 0, 6, -3, -1, -4, -2, -1,
    -- filter=16 channel=20
    0, -8, 3, 0, -8, 1, 6, 0, 0,
    -- filter=16 channel=21
    0, -8, 3, -11, 10, 7, 2, -5, -2,
    -- filter=16 channel=22
    -2, 6, 7, -4, 0, 1, -1, 1, 4,
    -- filter=16 channel=23
    -10, 2, 5, -4, 4, -1, -9, 0, 0,
    -- filter=16 channel=24
    -2, 1, -5, -3, 5, 5, 2, -2, -2,
    -- filter=16 channel=25
    -11, -8, 10, -13, 5, 4, -6, -1, -1,
    -- filter=16 channel=26
    -1, 6, -4, -8, 7, -4, 1, 5, -1,
    -- filter=16 channel=27
    -10, 0, 11, -15, 5, 1, -11, 4, -8,
    -- filter=16 channel=28
    1, 2, 0, 3, -5, 5, 0, -1, -7,
    -- filter=16 channel=29
    0, 2, 5, 9, -6, 0, -1, -3, 3,
    -- filter=16 channel=30
    0, 6, 9, -9, 7, -3, 0, 0, -1,
    -- filter=16 channel=31
    -7, 1, 12, -13, 8, 10, 3, 6, 2,
    -- filter=16 channel=32
    0, -2, 7, -10, -11, 2, -6, -3, 6,
    -- filter=16 channel=33
    -1, 0, 6, -16, 2, 10, -1, 2, 6,
    -- filter=16 channel=34
    2, 15, 0, -7, 8, 8, -5, 11, -6,
    -- filter=16 channel=35
    1, -1, -1, -4, -6, 2, 3, 3, -3,
    -- filter=16 channel=36
    -8, -2, 1, 6, 8, 0, 1, 6, -2,
    -- filter=16 channel=37
    0, 5, 12, -7, -2, 11, 7, -9, 4,
    -- filter=16 channel=38
    -1, 3, 0, -1, 2, 1, 2, 7, 4,
    -- filter=16 channel=39
    3, -8, 0, 4, 4, 1, 5, 4, 5,
    -- filter=16 channel=40
    3, -4, -9, -3, 4, 0, -1, 1, -2,
    -- filter=16 channel=41
    -8, -7, -5, -5, -1, 6, -17, -4, 7,
    -- filter=16 channel=42
    -2, 2, -3, 3, -5, 2, 0, -8, 2,
    -- filter=16 channel=43
    0, 6, 0, -6, -7, 3, 4, 6, -1,
    -- filter=16 channel=44
    -6, 0, 12, -6, 5, 5, 2, 0, -2,
    -- filter=16 channel=45
    0, -1, 3, 6, 2, -1, 2, -2, -7,
    -- filter=16 channel=46
    3, 2, 6, -5, 0, 2, 5, -7, 0,
    -- filter=16 channel=47
    -9, 0, 3, -18, 0, 17, 1, 7, 8,
    -- filter=16 channel=48
    -6, -4, 0, -5, 11, 0, 1, 4, 4,
    -- filter=16 channel=49
    -5, -9, -5, -9, 0, -1, 1, -4, 8,
    -- filter=16 channel=50
    -8, -6, 9, -9, 0, 7, 1, -1, 0,
    -- filter=16 channel=51
    -6, -1, 5, -4, 5, -3, -2, -3, -6,
    -- filter=16 channel=52
    4, 2, 2, 8, 8, 6, 1, 6, 4,
    -- filter=16 channel=53
    6, 4, -2, 3, 4, -1, -3, 6, 1,
    -- filter=16 channel=54
    2, 1, -3, -3, 6, 0, -3, -2, 7,
    -- filter=16 channel=55
    0, -3, -4, -1, -2, -5, -2, -5, 0,
    -- filter=16 channel=56
    1, -2, 7, 7, 8, -4, 4, 3, 1,
    -- filter=16 channel=57
    -4, 0, 6, 0, 2, 3, -1, -2, -2,
    -- filter=16 channel=58
    0, 5, 8, -6, -8, -2, 2, 0, -6,
    -- filter=16 channel=59
    -3, -11, 9, -20, 0, 6, -11, 2, -4,
    -- filter=16 channel=60
    1, 2, 0, 4, 4, 4, 5, -6, -1,
    -- filter=16 channel=61
    5, 6, -7, -4, 0, -8, -1, 5, -8,
    -- filter=16 channel=62
    0, -7, 0, -2, 2, 0, 1, -2, -2,
    -- filter=16 channel=63
    -2, 3, 7, -2, -3, 6, 3, 5, -1,
    -- filter=16 channel=64
    2, -3, 0, 3, 0, -4, -6, 5, -1,
    -- filter=16 channel=65
    5, 0, 2, -1, -4, 5, 5, 5, 5,
    -- filter=16 channel=66
    5, -4, 4, 0, -2, -6, -2, 2, 1,
    -- filter=16 channel=67
    4, 4, -5, -3, 1, 6, 5, -6, -5,
    -- filter=16 channel=68
    2, -2, 0, -3, -8, 0, 2, 7, 4,
    -- filter=16 channel=69
    3, 1, 0, -1, -3, 7, -3, 2, -5,
    -- filter=16 channel=70
    -14, -5, -2, -12, 1, -3, -3, 0, -2,
    -- filter=16 channel=71
    9, 5, -2, 3, 0, 4, -4, -3, 0,
    -- filter=16 channel=72
    -15, -9, 10, -13, 4, 12, -12, 5, 6,
    -- filter=16 channel=73
    -2, -2, 0, -1, -1, 0, -3, 8, 1,
    -- filter=16 channel=74
    -7, 6, 7, -9, 17, 1, -2, 6, -3,
    -- filter=16 channel=75
    0, -4, 7, -10, -3, 10, 1, -6, 0,
    -- filter=16 channel=76
    -4, -1, -5, 1, -2, -4, -1, -1, 5,
    -- filter=16 channel=77
    3, -6, 2, 3, -6, -2, 4, -2, 6,
    -- filter=16 channel=78
    -7, -3, 0, 0, -2, -2, 7, 7, 6,
    -- filter=16 channel=79
    -3, -14, -5, -15, -3, 5, -16, -6, 0,
    -- filter=16 channel=80
    -17, -13, 6, -22, 5, 7, -14, -3, 5,
    -- filter=16 channel=81
    0, 7, 1, 5, 2, 0, 6, 5, 4,
    -- filter=16 channel=82
    4, 3, 3, 3, 2, 3, 0, 3, -6,
    -- filter=16 channel=83
    1, -6, -2, -6, 4, 2, -7, 6, 0,
    -- filter=16 channel=84
    -4, -6, 8, -7, 0, -2, -4, 4, -1,
    -- filter=16 channel=85
    2, 0, -2, 2, 1, 6, -6, -3, -7,
    -- filter=16 channel=86
    0, 8, 1, -1, 7, 4, 4, 8, 1,
    -- filter=16 channel=87
    -3, -3, -7, -1, 4, -2, 7, 7, -3,
    -- filter=16 channel=88
    -2, 4, 2, 1, 4, -2, 5, 1, -6,
    -- filter=16 channel=89
    -8, -18, 6, -15, -7, 10, -7, 6, 5,
    -- filter=16 channel=90
    -9, 1, 2, 3, 10, -6, -4, 7, -7,
    -- filter=16 channel=91
    -13, -9, 0, -5, -4, 4, -1, 1, 3,
    -- filter=16 channel=92
    -5, 5, -6, 3, 4, -5, 3, 4, 5,
    -- filter=16 channel=93
    -10, 5, 13, -7, -2, 3, -1, 5, 0,
    -- filter=16 channel=94
    0, 0, 2, 5, -2, -2, 0, 1, 2,
    -- filter=16 channel=95
    2, -3, 1, 0, -5, 6, -7, -3, 5,
    -- filter=16 channel=96
    3, -6, -6, 0, 4, 5, -3, -2, 4,
    -- filter=16 channel=97
    0, -5, -3, -5, -7, 5, -2, -5, 4,
    -- filter=16 channel=98
    -4, -3, 6, -13, 8, 0, -11, 7, 7,
    -- filter=16 channel=99
    -8, 8, 3, -7, 16, 7, -6, 8, -10,
    -- filter=16 channel=100
    1, 2, -1, -2, 2, -2, 5, 5, -5,
    -- filter=16 channel=101
    4, -3, 2, 2, 4, -4, 3, -4, 4,
    -- filter=16 channel=102
    -2, 3, 1, -7, 6, -2, -5, 5, 3,
    -- filter=16 channel=103
    -10, -6, 7, -9, -1, 5, 0, -1, 2,
    -- filter=16 channel=104
    -5, 1, 5, -8, 14, 12, -2, 5, 0,
    -- filter=16 channel=105
    0, 0, -7, 8, 2, -4, 2, -6, 0,
    -- filter=16 channel=106
    -2, -2, 4, 7, 4, -6, -1, 2, 7,
    -- filter=16 channel=107
    -4, 4, 0, -4, -3, 5, 4, 1, -3,
    -- filter=16 channel=108
    0, -2, 2, 0, -7, 4, -3, -8, 2,
    -- filter=16 channel=109
    -19, 0, 1, -15, 11, 12, -10, 0, -7,
    -- filter=16 channel=110
    2, 0, -5, 0, -1, 3, -1, -2, -5,
    -- filter=16 channel=111
    2, 1, 1, -1, -7, 6, 0, -5, 0,
    -- filter=16 channel=112
    -4, 1, 3, -8, 8, 9, -5, 5, -5,
    -- filter=16 channel=113
    -6, -2, 1, -9, 0, 7, -5, 0, 0,
    -- filter=16 channel=114
    -12, -3, 9, -17, -1, -1, -1, 1, 3,
    -- filter=16 channel=115
    -1, 0, 5, 3, -5, 0, 0, 2, 1,
    -- filter=16 channel=116
    -1, -1, 1, -10, -3, 4, -2, 3, -3,
    -- filter=16 channel=117
    2, 2, 5, -7, 1, 5, 0, 3, -5,
    -- filter=16 channel=118
    2, 4, -2, 1, 1, -5, -6, 2, -7,
    -- filter=16 channel=119
    -8, 11, 2, 8, 11, 6, -1, 0, 3,
    -- filter=16 channel=120
    -15, 6, 7, -11, 15, 6, -8, 1, -10,
    -- filter=16 channel=121
    -4, -4, -6, -6, -8, 1, -8, 4, -5,
    -- filter=16 channel=122
    -17, 2, 14, -19, 7, 10, -2, 11, -1,
    -- filter=16 channel=123
    -5, 8, 0, -1, 7, 8, 6, 0, 0,
    -- filter=16 channel=124
    -4, -5, 0, 3, -1, 2, -6, 1, -7,
    -- filter=16 channel=125
    -16, -8, 6, -9, 3, 12, -7, 4, -8,
    -- filter=16 channel=126
    -2, -7, 1, -9, -7, 4, -10, -2, 2,
    -- filter=16 channel=127
    -8, -4, 5, 1, 3, -1, 0, -7, -4,
    -- filter=17 channel=0
    -1, -15, 1, -12, -16, 12, -2, -17, 8,
    -- filter=17 channel=1
    2, -7, 14, -2, -13, 11, 0, -8, 12,
    -- filter=17 channel=2
    -1, 2, -2, 2, 2, -2, 1, -4, -4,
    -- filter=17 channel=3
    -7, -2, 0, -5, -1, 1, -3, -2, 6,
    -- filter=17 channel=4
    10, 3, 8, -3, -4, -5, -18, -6, -7,
    -- filter=17 channel=5
    -10, -2, 13, -1, -9, 7, -3, -9, 3,
    -- filter=17 channel=6
    6, -7, -2, 0, 4, -3, 0, 0, 0,
    -- filter=17 channel=7
    -7, -4, -2, -4, 3, -6, 3, -4, -6,
    -- filter=17 channel=8
    0, 0, -3, -7, -6, 2, -5, -8, -7,
    -- filter=17 channel=9
    -4, 3, 2, -4, 5, 0, -1, -1, 2,
    -- filter=17 channel=10
    0, -5, 1, 4, 9, 4, 2, 3, -3,
    -- filter=17 channel=11
    7, -2, -10, 7, 13, 0, 9, 6, -3,
    -- filter=17 channel=12
    -6, 0, 0, -4, -3, 5, -7, 0, 3,
    -- filter=17 channel=13
    5, -1, 4, 1, -5, -2, 4, -4, 1,
    -- filter=17 channel=14
    2, 0, 4, 0, 7, 4, -4, -6, 0,
    -- filter=17 channel=15
    0, -8, -7, 10, 3, -4, -5, 3, -6,
    -- filter=17 channel=16
    -9, -6, 6, -2, 0, 12, 5, -6, 0,
    -- filter=17 channel=17
    -3, -6, -7, 1, -2, 4, 4, 3, -4,
    -- filter=17 channel=18
    4, -11, -14, 11, 1, 3, -9, -8, 0,
    -- filter=17 channel=19
    -3, 0, 7, 1, -3, -4, 6, 2, 4,
    -- filter=17 channel=20
    8, 9, -19, 5, 18, -11, -1, 5, -2,
    -- filter=17 channel=21
    -5, 1, 11, 1, 4, 9, 7, 2, -10,
    -- filter=17 channel=22
    -3, -1, -2, -1, -8, 7, 2, 0, 2,
    -- filter=17 channel=23
    -1, 0, -7, -2, 3, 2, -2, 12, -10,
    -- filter=17 channel=24
    4, 1, 0, -5, 4, 0, -4, -4, -1,
    -- filter=17 channel=25
    7, 0, 7, 2, -3, 5, -5, -10, 0,
    -- filter=17 channel=26
    -4, 4, 7, -10, 2, 4, -9, 0, 0,
    -- filter=17 channel=27
    -4, -6, 11, -10, 4, 5, -3, 0, -1,
    -- filter=17 channel=28
    0, -7, 2, -6, 2, 6, 5, 5, 1,
    -- filter=17 channel=29
    2, 9, -14, 11, 3, -5, 0, 3, 3,
    -- filter=17 channel=30
    -7, 5, 3, 3, -6, 1, -9, -1, -8,
    -- filter=17 channel=31
    -11, -4, -1, 8, 19, 2, -2, 7, -14,
    -- filter=17 channel=32
    -7, -6, 4, 1, 4, 14, -7, -3, 1,
    -- filter=17 channel=33
    -6, -4, 1, 1, -6, 6, -3, 5, 0,
    -- filter=17 channel=34
    -17, -8, 12, -15, -16, 8, -17, -4, 9,
    -- filter=17 channel=35
    -5, 2, 3, -6, -1, -1, 1, 3, 5,
    -- filter=17 channel=36
    1, 2, 4, -1, 6, -10, -3, -2, -16,
    -- filter=17 channel=37
    -11, 2, 10, -6, -14, 12, 0, -16, 0,
    -- filter=17 channel=38
    0, 0, 3, -1, 2, 2, 4, 2, -3,
    -- filter=17 channel=39
    5, -2, 0, 5, 5, 1, 1, 2, -8,
    -- filter=17 channel=40
    7, -4, 0, 7, 5, -8, 8, -1, 3,
    -- filter=17 channel=41
    -1, -4, 15, 0, -26, 12, -17, -24, 11,
    -- filter=17 channel=42
    5, -2, 5, 1, 4, 3, -4, -7, 3,
    -- filter=17 channel=43
    2, 0, -7, -2, -11, 1, -9, -1, 2,
    -- filter=17 channel=44
    -4, -3, 9, -4, -8, 5, 1, -6, -6,
    -- filter=17 channel=45
    -3, -7, 6, 5, 0, -6, -2, -4, 2,
    -- filter=17 channel=46
    -4, 4, 8, 3, 3, 0, -6, -5, -1,
    -- filter=17 channel=47
    -1, 2, 12, 3, -2, 4, -1, 6, 8,
    -- filter=17 channel=48
    3, -2, 13, -5, 0, 13, -6, -5, -13,
    -- filter=17 channel=49
    0, -2, 3, 0, -6, -5, -1, -2, -5,
    -- filter=17 channel=50
    -1, 2, -6, 1, 1, 5, 7, 0, -9,
    -- filter=17 channel=51
    -4, -2, 1, -3, 7, 0, 0, 6, 6,
    -- filter=17 channel=52
    2, 1, 1, -5, -5, -3, -2, -8, -8,
    -- filter=17 channel=53
    -6, 4, 1, 8, 4, 2, 1, -1, -9,
    -- filter=17 channel=54
    -3, 1, 3, -2, -2, -3, 0, 5, 1,
    -- filter=17 channel=55
    10, 0, -16, 13, 2, -7, 1, -2, 2,
    -- filter=17 channel=56
    1, -6, 1, 0, 4, -4, 2, 0, 2,
    -- filter=17 channel=57
    6, 6, 6, 0, -7, -4, -4, 0, 0,
    -- filter=17 channel=58
    1, -4, -3, 2, -8, -6, 3, -1, -4,
    -- filter=17 channel=59
    6, -5, 1, 8, 7, 13, 0, 1, 1,
    -- filter=17 channel=60
    -3, 0, -1, -6, 4, -5, 0, 7, 4,
    -- filter=17 channel=61
    5, 0, 0, 3, 0, 2, 3, -7, -4,
    -- filter=17 channel=62
    -5, 6, 0, -2, -1, 2, 1, -1, 1,
    -- filter=17 channel=63
    -7, 1, 3, 2, 4, 7, 5, -5, -6,
    -- filter=17 channel=64
    -5, 0, -8, 8, 3, 0, 7, -4, 0,
    -- filter=17 channel=65
    -7, 0, 7, 4, 0, 5, -4, 6, 3,
    -- filter=17 channel=66
    -5, -6, 3, -5, -3, 9, -10, -16, 9,
    -- filter=17 channel=67
    6, -5, -3, 6, -2, -7, -1, 1, -1,
    -- filter=17 channel=68
    4, -1, 0, -1, -5, 3, 2, 2, -2,
    -- filter=17 channel=69
    -5, -7, 1, 6, 0, 2, 2, 2, 4,
    -- filter=17 channel=70
    2, 3, 1, 0, 7, 0, -6, -9, -3,
    -- filter=17 channel=71
    -5, 1, -6, 0, -7, 2, 8, 8, 3,
    -- filter=17 channel=72
    3, 2, -10, 1, 10, -2, 8, 8, -11,
    -- filter=17 channel=73
    -2, -1, -4, 5, 6, 1, -6, -1, -9,
    -- filter=17 channel=74
    -11, -4, 10, -12, -1, 12, -9, 0, -1,
    -- filter=17 channel=75
    -5, -10, 7, -3, -11, 8, -5, -6, 7,
    -- filter=17 channel=76
    7, 6, -18, 16, 11, -3, 6, 9, -4,
    -- filter=17 channel=77
    6, 2, 5, 0, -6, -2, 4, 2, 0,
    -- filter=17 channel=78
    -8, 0, -1, -8, -4, 7, -2, 1, 2,
    -- filter=17 channel=79
    -5, -5, -7, 4, -5, 6, -8, -2, 8,
    -- filter=17 channel=80
    -3, -4, -6, 12, 13, 12, 10, 6, -10,
    -- filter=17 channel=81
    0, 3, -3, 2, 5, 3, 0, -1, 3,
    -- filter=17 channel=82
    -2, 2, -5, -1, 4, -5, 5, -2, 4,
    -- filter=17 channel=83
    7, 0, 8, 5, 6, -7, 3, -1, -5,
    -- filter=17 channel=84
    4, 0, 1, -2, 4, 1, -4, -3, 0,
    -- filter=17 channel=85
    5, -5, 1, 3, 6, -6, 7, -2, -1,
    -- filter=17 channel=86
    -1, 0, 11, -3, -14, 11, -6, -10, 0,
    -- filter=17 channel=87
    -2, -8, -9, -2, -7, 0, -8, 4, 0,
    -- filter=17 channel=88
    7, 3, -9, 5, 12, -2, -3, -2, -15,
    -- filter=17 channel=89
    -1, 0, -10, 9, 9, 3, 1, 1, -9,
    -- filter=17 channel=90
    -12, 6, -2, -8, 6, 0, 4, 3, -3,
    -- filter=17 channel=91
    1, 3, 1, -6, 10, -4, 0, -4, -4,
    -- filter=17 channel=92
    -9, 5, 6, -2, 2, 5, 1, -6, 4,
    -- filter=17 channel=93
    0, 0, 19, 1, -10, 14, -3, -2, -9,
    -- filter=17 channel=94
    -6, 2, -7, 0, 0, -2, 4, 3, -4,
    -- filter=17 channel=95
    -1, 0, 0, 5, -3, -2, -1, -4, 7,
    -- filter=17 channel=96
    5, 0, -6, -5, 5, 2, 2, 3, 6,
    -- filter=17 channel=97
    -9, -2, 1, 4, -8, 0, 0, -4, 5,
    -- filter=17 channel=98
    -2, -1, 2, -3, 1, 12, -5, 3, -8,
    -- filter=17 channel=99
    0, 7, 0, 4, 12, 2, -4, 0, -16,
    -- filter=17 channel=100
    -6, 0, 0, -4, -5, -3, -5, -9, 3,
    -- filter=17 channel=101
    3, 0, -2, -11, -11, -9, -11, -7, -7,
    -- filter=17 channel=102
    -7, -3, 0, 4, 2, -1, 0, -4, -2,
    -- filter=17 channel=103
    -7, 0, 7, 1, -1, 14, 10, 3, 10,
    -- filter=17 channel=104
    -3, 6, 6, 3, 10, 5, 3, 4, -4,
    -- filter=17 channel=105
    -1, 3, -15, 12, 8, -7, -3, 1, 2,
    -- filter=17 channel=106
    5, 7, -9, 12, 7, -10, 7, -2, 1,
    -- filter=17 channel=107
    -3, -7, -14, 0, 5, -6, -12, 5, 4,
    -- filter=17 channel=108
    2, -1, 4, -8, -6, 5, 0, -1, 9,
    -- filter=17 channel=109
    0, -6, 10, -2, 9, 13, -6, -8, -1,
    -- filter=17 channel=110
    -8, -9, 0, 1, 4, -11, 8, -4, -2,
    -- filter=17 channel=111
    -4, 5, 3, 7, 1, 0, -1, 1, -4,
    -- filter=17 channel=112
    -5, -1, -1, -8, 4, 3, -12, 4, 2,
    -- filter=17 channel=113
    -4, -8, -1, 0, 0, 0, -3, 1, -2,
    -- filter=17 channel=114
    0, -8, 4, 0, -12, 4, -9, -22, -2,
    -- filter=17 channel=115
    -5, 2, 1, -3, 3, -2, 0, -3, 5,
    -- filter=17 channel=116
    13, -2, 3, -1, 4, -3, -5, -10, -11,
    -- filter=17 channel=117
    8, -7, 3, 1, -4, 4, 1, 0, -5,
    -- filter=17 channel=118
    5, -6, 0, -5, 0, -4, 2, 4, -5,
    -- filter=17 channel=119
    -12, -6, 10, -9, 0, 0, -13, -13, -4,
    -- filter=17 channel=120
    -4, 8, 4, -3, 5, 5, -14, 5, -2,
    -- filter=17 channel=121
    6, 0, 7, 5, 1, 2, 5, -6, 6,
    -- filter=17 channel=122
    -13, -6, 12, 2, 5, 6, 4, 7, -5,
    -- filter=17 channel=123
    0, 1, 0, 1, -7, 5, 2, 1, 9,
    -- filter=17 channel=124
    0, 6, -7, 9, 10, -2, 6, 5, -6,
    -- filter=17 channel=125
    -5, -6, 5, 4, 8, 0, -5, 0, -13,
    -- filter=17 channel=126
    -5, -4, 5, 1, 0, 1, -4, -3, 4,
    -- filter=17 channel=127
    -4, -6, -2, -4, 1, 3, -2, 1, 1,
    -- filter=18 channel=0
    0, -7, -6, 7, 1, 0, -1, 0, 4,
    -- filter=18 channel=1
    0, -7, -5, 1, -3, -4, -5, 7, 4,
    -- filter=18 channel=2
    1, -7, -1, -7, 0, -4, 0, 6, 2,
    -- filter=18 channel=3
    0, -2, -2, 7, -6, 4, 0, 0, -2,
    -- filter=18 channel=4
    -2, 1, 5, 7, 4, 6, -1, -5, -5,
    -- filter=18 channel=5
    0, -4, 1, 3, -5, 1, 2, -7, -2,
    -- filter=18 channel=6
    4, -7, 3, 5, -4, 2, -5, 5, -2,
    -- filter=18 channel=7
    3, 7, 0, -1, -5, 6, 2, 5, 0,
    -- filter=18 channel=8
    -3, 0, -3, -3, -3, 0, 0, 6, -5,
    -- filter=18 channel=9
    -1, -6, 3, -5, -2, 5, 2, 2, 3,
    -- filter=18 channel=10
    5, 5, 0, 6, -3, -4, -4, 4, -4,
    -- filter=18 channel=11
    -5, -6, 5, -5, -2, 7, -5, 0, 5,
    -- filter=18 channel=12
    -4, -5, -5, -2, -6, 7, 7, -4, 1,
    -- filter=18 channel=13
    -4, 1, 2, -4, 1, 0, -6, 2, -1,
    -- filter=18 channel=14
    0, 1, -1, -5, -3, -6, 0, -5, 0,
    -- filter=18 channel=15
    -6, 3, -1, -6, 3, 5, -2, 3, -1,
    -- filter=18 channel=16
    4, 0, 1, -7, -7, 0, 5, 3, -3,
    -- filter=18 channel=17
    1, 0, 0, 2, -4, -2, -1, -3, -1,
    -- filter=18 channel=18
    4, 2, 0, 2, -4, 0, 0, 0, -1,
    -- filter=18 channel=19
    -3, 4, -2, 4, 0, -1, -1, 1, 1,
    -- filter=18 channel=20
    4, -7, 4, -3, -6, -4, -2, 0, 6,
    -- filter=18 channel=21
    -7, -3, -1, 4, 3, 5, 0, -4, 3,
    -- filter=18 channel=22
    -3, -2, 3, 6, -1, 3, 0, 0, -6,
    -- filter=18 channel=23
    -5, 5, -3, -1, -7, -1, 6, 0, -2,
    -- filter=18 channel=24
    -2, 3, 5, 0, 2, -3, 4, 3, 1,
    -- filter=18 channel=25
    -1, 0, -7, 0, 7, -6, 6, -2, -6,
    -- filter=18 channel=26
    4, 6, 2, 2, -5, 5, 5, 4, 7,
    -- filter=18 channel=27
    1, 3, -5, -3, -4, 0, -3, -6, -1,
    -- filter=18 channel=28
    -1, 5, -3, -4, 5, 0, 0, -3, -3,
    -- filter=18 channel=29
    -2, 0, 6, -6, -1, -5, 4, 0, -4,
    -- filter=18 channel=30
    5, 4, 6, -1, 4, 0, 0, 4, -2,
    -- filter=18 channel=31
    -1, 5, -5, -5, 0, -4, 3, 0, -6,
    -- filter=18 channel=32
    -4, 4, -5, 0, -2, -2, 1, -3, -6,
    -- filter=18 channel=33
    -6, -2, 0, 2, 4, 0, -6, 0, -4,
    -- filter=18 channel=34
    -2, 6, 5, 2, 5, 6, 5, -5, -6,
    -- filter=18 channel=35
    3, 1, -6, 1, 5, 0, 6, 6, -2,
    -- filter=18 channel=36
    0, -3, 3, 4, -2, 0, -5, 6, -1,
    -- filter=18 channel=37
    4, 6, -1, 0, -4, -5, 3, 0, 2,
    -- filter=18 channel=38
    1, 6, -6, -7, -2, -4, 1, 4, -1,
    -- filter=18 channel=39
    0, 0, 7, 7, -3, 0, 6, -2, -3,
    -- filter=18 channel=40
    5, 1, 3, -6, -4, 0, 2, 0, 4,
    -- filter=18 channel=41
    -1, -1, -2, 5, -4, -2, -3, 4, -6,
    -- filter=18 channel=42
    5, 5, 1, -4, -6, -4, -6, 0, -3,
    -- filter=18 channel=43
    2, 4, 0, -7, -3, 4, -1, 1, -2,
    -- filter=18 channel=44
    -4, 3, -6, 7, 5, -5, -4, 2, 6,
    -- filter=18 channel=45
    3, 0, 4, 6, -4, 0, -5, 6, -5,
    -- filter=18 channel=46
    -3, 2, -3, -6, -3, -3, 2, -1, -5,
    -- filter=18 channel=47
    -4, 3, 5, -2, -4, -6, 2, -5, 0,
    -- filter=18 channel=48
    -3, -5, 0, -6, -1, -2, 5, -7, 3,
    -- filter=18 channel=49
    -4, 2, -1, -6, 1, -3, -3, 6, -5,
    -- filter=18 channel=50
    0, -2, 1, 0, -2, 4, 5, -2, 2,
    -- filter=18 channel=51
    -7, 3, 5, -2, 5, -7, -6, 7, 4,
    -- filter=18 channel=52
    -5, 5, 2, -7, -7, 6, 0, -3, 2,
    -- filter=18 channel=53
    -2, -3, 3, 1, 5, -3, 7, -7, 3,
    -- filter=18 channel=54
    0, 4, 2, -2, -1, 0, 3, 6, 0,
    -- filter=18 channel=55
    4, -1, -7, -5, -6, 6, -3, 2, -5,
    -- filter=18 channel=56
    -5, -5, 2, -4, 0, 6, 0, -7, -5,
    -- filter=18 channel=57
    1, 0, 5, -4, 0, -4, 7, -5, 1,
    -- filter=18 channel=58
    3, -2, 0, -1, 0, 0, 0, -1, 0,
    -- filter=18 channel=59
    -6, -6, -1, 6, 1, -4, 1, -3, 0,
    -- filter=18 channel=60
    -5, 0, 5, 4, -5, 0, -3, 2, 1,
    -- filter=18 channel=61
    1, -6, 7, -4, -5, 4, 3, 1, 2,
    -- filter=18 channel=62
    3, 1, -3, 3, -6, 6, -7, 0, 2,
    -- filter=18 channel=63
    6, -6, -2, 4, -3, 2, -4, 1, 2,
    -- filter=18 channel=64
    0, 0, 0, 4, 3, 1, 0, 1, 4,
    -- filter=18 channel=65
    7, 0, -6, 2, -5, 3, -3, 3, 1,
    -- filter=18 channel=66
    2, 4, 4, -3, -2, -5, -1, -2, -1,
    -- filter=18 channel=67
    1, -3, 5, 0, -3, -3, -4, 0, -5,
    -- filter=18 channel=68
    -2, -2, -3, 5, -6, -4, 0, -2, 7,
    -- filter=18 channel=69
    -4, 3, -4, 5, -2, 5, -3, 0, -7,
    -- filter=18 channel=70
    -7, -7, 3, -2, -1, -2, 0, -7, 2,
    -- filter=18 channel=71
    3, 6, -4, -6, 7, -5, -6, -5, -6,
    -- filter=18 channel=72
    0, -1, -2, -3, -6, 0, 0, 3, -3,
    -- filter=18 channel=73
    4, 5, -1, -1, 2, -6, -1, -6, -3,
    -- filter=18 channel=74
    0, 5, -3, 0, 5, 2, -4, 1, 2,
    -- filter=18 channel=75
    5, 3, -7, -5, -4, 3, -5, 4, 1,
    -- filter=18 channel=76
    1, -4, 2, 0, 6, 4, 0, 5, 5,
    -- filter=18 channel=77
    1, -6, 0, -1, 1, -3, -1, 3, 7,
    -- filter=18 channel=78
    -6, -6, 5, 0, 0, 0, 6, -1, 0,
    -- filter=18 channel=79
    -3, -2, -3, 0, -3, 1, 5, -1, -4,
    -- filter=18 channel=80
    3, 0, -2, 1, -3, -4, -3, -2, -1,
    -- filter=18 channel=81
    -2, 5, 5, 3, -3, 3, -2, 3, 0,
    -- filter=18 channel=82
    -4, 3, 7, 4, 5, 6, -7, 6, -1,
    -- filter=18 channel=83
    5, 6, 3, 0, -3, -2, 4, 7, -2,
    -- filter=18 channel=84
    -7, 4, 0, -3, -7, -5, 2, -1, -2,
    -- filter=18 channel=85
    1, 5, 0, 0, 3, 2, -2, 0, 0,
    -- filter=18 channel=86
    2, -6, 7, 6, -3, 0, 0, -6, 1,
    -- filter=18 channel=87
    -5, 0, -1, 0, -5, -7, -5, 5, -5,
    -- filter=18 channel=88
    -1, -7, -5, -4, -1, 0, 5, 3, 0,
    -- filter=18 channel=89
    0, 5, 5, 3, 0, 5, -3, -2, -5,
    -- filter=18 channel=90
    -2, -2, 7, -1, 4, -3, -2, 0, -7,
    -- filter=18 channel=91
    4, -6, 2, -6, 7, 6, 5, -3, -6,
    -- filter=18 channel=92
    7, 5, -5, 3, 6, 0, -4, 4, 1,
    -- filter=18 channel=93
    1, -5, 0, 6, 1, 7, -4, -3, -1,
    -- filter=18 channel=94
    -4, 0, 6, 0, 3, 0, -1, 3, -5,
    -- filter=18 channel=95
    -2, 1, 2, 6, 1, 2, -3, 0, -5,
    -- filter=18 channel=96
    2, -5, -4, 3, -5, 6, -5, 1, -6,
    -- filter=18 channel=97
    -4, 7, -2, 3, 0, 6, 6, -1, -3,
    -- filter=18 channel=98
    3, 3, -3, 2, 7, -1, -5, 7, 7,
    -- filter=18 channel=99
    -1, 6, 3, 0, 3, -6, 0, 0, 0,
    -- filter=18 channel=100
    3, 6, -4, -1, 5, -1, 0, -4, 1,
    -- filter=18 channel=101
    5, -3, -6, 1, 1, -2, 0, -6, -6,
    -- filter=18 channel=102
    -2, 4, -4, 4, 0, -5, 3, 4, 0,
    -- filter=18 channel=103
    -5, -6, 0, -3, 6, -5, 2, -4, -2,
    -- filter=18 channel=104
    -6, -5, 3, 2, 0, -5, 5, -5, 3,
    -- filter=18 channel=105
    7, 2, -4, 6, -4, -2, -5, -7, 6,
    -- filter=18 channel=106
    4, 6, 2, 0, 3, 5, -7, -3, -1,
    -- filter=18 channel=107
    7, -3, 0, -2, -5, 6, 0, 1, -2,
    -- filter=18 channel=108
    -1, 1, -6, -3, -6, 2, 5, 4, -5,
    -- filter=18 channel=109
    1, 3, 0, -5, 7, -2, 0, -6, 7,
    -- filter=18 channel=110
    -1, 1, 2, 6, -1, -2, 0, 0, 2,
    -- filter=18 channel=111
    1, 1, -4, 0, 6, -3, -2, 3, 1,
    -- filter=18 channel=112
    2, 0, -7, 0, 6, -2, 4, -2, 0,
    -- filter=18 channel=113
    6, 6, 2, -3, 0, -4, -3, -6, 4,
    -- filter=18 channel=114
    0, 0, -2, 4, -4, -1, 7, 0, -5,
    -- filter=18 channel=115
    -4, -4, 2, 0, -2, 0, -2, -7, 0,
    -- filter=18 channel=116
    -7, 4, 4, -2, -1, -1, -4, 6, -2,
    -- filter=18 channel=117
    6, -1, 0, 5, 0, 5, 0, 2, 0,
    -- filter=18 channel=118
    6, 2, 2, -5, 4, 3, -6, -2, 2,
    -- filter=18 channel=119
    -1, -4, -3, 3, -6, -6, 4, -4, -4,
    -- filter=18 channel=120
    3, 6, -4, 0, -2, -3, -2, 1, 1,
    -- filter=18 channel=121
    5, 6, -1, -3, -7, 2, -1, -6, 1,
    -- filter=18 channel=122
    0, 5, 1, 7, 0, 7, -2, -5, -4,
    -- filter=18 channel=123
    -1, 2, -6, -2, 5, 5, 1, -4, 5,
    -- filter=18 channel=124
    4, 3, 0, 3, 1, 4, 0, -2, 5,
    -- filter=18 channel=125
    -1, -1, 2, -4, -1, -2, 5, -6, -5,
    -- filter=18 channel=126
    -1, -5, 7, 7, 3, 1, -2, 3, 4,
    -- filter=18 channel=127
    2, -5, -2, 3, 0, -1, 6, -5, 5,
    -- filter=19 channel=0
    8, 6, 6, 1, -7, -3, 2, 5, -1,
    -- filter=19 channel=1
    -2, 10, 9, 1, -3, -4, -7, -7, -4,
    -- filter=19 channel=2
    0, -10, -6, -4, 11, 0, 7, 9, -5,
    -- filter=19 channel=3
    1, 7, -1, 0, 1, 3, -6, 10, 5,
    -- filter=19 channel=4
    3, -3, 5, 9, 30, 20, 9, 10, 9,
    -- filter=19 channel=5
    2, 14, 16, 5, -5, -3, 1, 6, -2,
    -- filter=19 channel=6
    0, -1, -3, -2, 9, 7, 8, 0, -1,
    -- filter=19 channel=7
    3, 1, -4, 5, -2, -7, 3, -1, 1,
    -- filter=19 channel=8
    -6, 1, -2, 6, 5, 2, 5, 7, -2,
    -- filter=19 channel=9
    1, 0, -10, 4, -1, 9, 0, 0, 9,
    -- filter=19 channel=10
    2, -8, -13, -11, -2, 0, 3, 7, 7,
    -- filter=19 channel=11
    0, -1, -2, 5, 1, 4, 0, -9, -7,
    -- filter=19 channel=12
    4, -11, 0, -5, -5, -8, 0, 2, -1,
    -- filter=19 channel=13
    6, -11, -18, -4, -15, 1, -10, 0, -6,
    -- filter=19 channel=14
    5, -2, -3, -3, -5, -4, 0, 3, 2,
    -- filter=19 channel=15
    4, -10, -11, 2, -13, 3, 3, 4, 3,
    -- filter=19 channel=16
    -3, 5, 6, -1, -2, -5, -7, 4, 3,
    -- filter=19 channel=17
    1, -6, -4, -3, -2, 2, 0, 0, -2,
    -- filter=19 channel=18
    6, -8, -14, 3, -1, 7, 4, 10, 6,
    -- filter=19 channel=19
    -1, 3, -2, 0, 2, 7, -5, -6, -4,
    -- filter=19 channel=20
    10, -5, 3, -5, 0, 2, 2, -1, -7,
    -- filter=19 channel=21
    -5, -5, -2, -6, -14, 4, 1, 5, 7,
    -- filter=19 channel=22
    2, 1, -5, -6, -6, 0, -5, -6, 4,
    -- filter=19 channel=23
    6, -14, -17, -9, -4, 5, 3, 16, 4,
    -- filter=19 channel=24
    2, -5, 8, 4, -6, -4, -6, 0, 1,
    -- filter=19 channel=25
    0, -16, -16, -10, -1, 13, -7, 0, 12,
    -- filter=19 channel=26
    -3, -3, -2, 4, 8, 9, -2, 0, -1,
    -- filter=19 channel=27
    4, -28, -23, -16, -1, 9, 0, 11, 15,
    -- filter=19 channel=28
    4, 4, -2, -6, -4, -6, -7, -2, 4,
    -- filter=19 channel=29
    12, 1, 1, -3, -1, 5, -1, -8, -10,
    -- filter=19 channel=30
    1, 0, 2, 1, 3, 13, 5, -1, 4,
    -- filter=19 channel=31
    -11, -22, -19, -20, -10, 8, 6, 19, 23,
    -- filter=19 channel=32
    8, -4, -11, 3, -7, 4, 2, 4, 5,
    -- filter=19 channel=33
    -2, -11, -16, -9, -18, 0, 2, 12, 13,
    -- filter=19 channel=34
    3, -7, -5, -5, 2, 0, 0, 6, 6,
    -- filter=19 channel=35
    3, -7, -3, 3, 5, -7, 0, -3, 4,
    -- filter=19 channel=36
    -3, -6, -14, 4, 3, 7, -3, -3, -2,
    -- filter=19 channel=37
    4, 3, 2, 2, 1, 1, -7, 1, -9,
    -- filter=19 channel=38
    -1, 2, -8, -7, -3, -2, -4, 3, 0,
    -- filter=19 channel=39
    -1, 1, 4, 6, 0, -3, 0, -7, -7,
    -- filter=19 channel=40
    6, -9, -4, -2, -14, 0, -8, 5, -4,
    -- filter=19 channel=41
    6, -3, 0, 2, 1, -7, -4, 12, 0,
    -- filter=19 channel=42
    -8, 2, 4, 0, -4, 10, -3, 2, 4,
    -- filter=19 channel=43
    6, 0, -1, 4, 2, -8, -8, 8, 5,
    -- filter=19 channel=44
    -10, -5, 3, -5, -3, 1, 1, 8, 1,
    -- filter=19 channel=45
    0, 6, 6, -1, 6, -2, 4, -2, 2,
    -- filter=19 channel=46
    -7, 8, -4, 1, -5, -8, -2, 1, -1,
    -- filter=19 channel=47
    -4, 7, -1, -12, -6, -5, -1, 10, 3,
    -- filter=19 channel=48
    -3, -7, -10, -4, 7, 11, 4, 0, 0,
    -- filter=19 channel=49
    -2, -13, -5, 1, 12, 7, 5, -7, -2,
    -- filter=19 channel=50
    -5, -15, -9, -3, -2, 4, 1, 6, 10,
    -- filter=19 channel=51
    0, 7, -6, -4, 1, 0, 0, 4, -6,
    -- filter=19 channel=52
    -2, -5, -8, -7, 2, 0, -3, 5, -2,
    -- filter=19 channel=53
    2, -5, -2, 0, -3, 8, 1, 0, 0,
    -- filter=19 channel=54
    -4, 3, 5, 3, -4, -1, 4, -6, 3,
    -- filter=19 channel=55
    2, -2, -16, 2, -14, -3, 5, 5, 3,
    -- filter=19 channel=56
    0, 4, 5, -3, 2, 4, -1, -4, 1,
    -- filter=19 channel=57
    -4, -3, 2, 5, -3, 1, -4, 7, 3,
    -- filter=19 channel=58
    3, 3, 6, -1, -4, -1, -2, -10, -5,
    -- filter=19 channel=59
    -6, -13, -6, -7, -11, 10, 8, 1, 11,
    -- filter=19 channel=60
    -5, 0, 7, 3, -2, -3, -1, 6, -6,
    -- filter=19 channel=61
    -6, -3, -8, 0, 7, -5, -4, -6, -7,
    -- filter=19 channel=62
    -2, -5, 2, -2, -5, -5, 1, 4, 5,
    -- filter=19 channel=63
    10, 11, 0, 0, 0, 4, 0, -1, 2,
    -- filter=19 channel=64
    -3, -6, -2, -4, -4, 6, 2, -7, -2,
    -- filter=19 channel=65
    1, 0, 5, 0, 2, 6, -2, 2, -4,
    -- filter=19 channel=66
    -3, 2, 1, 4, 1, -11, -9, 8, -9,
    -- filter=19 channel=67
    2, 0, -5, 1, 1, 2, -1, -2, -5,
    -- filter=19 channel=68
    0, -6, -4, 3, -3, 8, -7, 1, -5,
    -- filter=19 channel=69
    7, -4, 0, 6, -4, -7, -1, -5, 4,
    -- filter=19 channel=70
    0, -12, -15, 0, 5, 0, 2, 0, 11,
    -- filter=19 channel=71
    2, -2, 3, -4, -9, -5, 0, -1, 6,
    -- filter=19 channel=72
    2, -12, -8, -11, -13, 3, 2, 10, 16,
    -- filter=19 channel=73
    8, -11, 0, -2, 0, 15, 1, 9, -1,
    -- filter=19 channel=74
    -9, -8, 3, -5, 3, 0, 7, 0, -2,
    -- filter=19 channel=75
    8, 6, 0, -9, -16, -17, -7, 3, 4,
    -- filter=19 channel=76
    13, -1, -10, -7, -7, -12, -10, -3, -7,
    -- filter=19 channel=77
    2, -3, -5, 3, 6, 5, -5, -3, 3,
    -- filter=19 channel=78
    1, 7, 6, -7, 3, 3, 9, -1, 2,
    -- filter=19 channel=79
    5, -18, -14, 3, 0, 6, -2, 6, 8,
    -- filter=19 channel=80
    3, -9, -14, -13, -1, 1, -5, 7, 11,
    -- filter=19 channel=81
    7, 2, 4, 0, -6, -2, -1, 0, 6,
    -- filter=19 channel=82
    5, 5, 7, -6, -1, 1, -4, -5, 2,
    -- filter=19 channel=83
    -6, -3, 1, 4, 3, 4, 6, -3, 3,
    -- filter=19 channel=84
    0, -16, -5, 5, 15, 5, -4, 3, 1,
    -- filter=19 channel=85
    7, -2, 5, -6, -5, 3, -1, 6, 5,
    -- filter=19 channel=86
    6, -7, 2, 5, 1, 0, -1, 4, -6,
    -- filter=19 channel=87
    9, -8, 0, 0, 0, 1, 0, 5, -1,
    -- filter=19 channel=88
    0, -1, -5, -9, -2, 0, -8, 1, -4,
    -- filter=19 channel=89
    -3, -6, -17, -11, -16, 8, -4, 11, 8,
    -- filter=19 channel=90
    3, -11, -3, -3, 1, -2, 0, 1, 3,
    -- filter=19 channel=91
    -5, -11, -14, 1, 15, 10, 2, 8, 0,
    -- filter=19 channel=92
    0, 5, 6, 4, 2, 2, 5, 2, 3,
    -- filter=19 channel=93
    -7, 0, -2, -4, 14, 7, 3, -6, 1,
    -- filter=19 channel=94
    -1, -5, 1, -2, 7, 1, 3, -1, -1,
    -- filter=19 channel=95
    0, -5, 6, 0, -6, 0, 2, 5, 7,
    -- filter=19 channel=96
    -6, 4, -6, 2, -4, 4, 1, -3, -2,
    -- filter=19 channel=97
    5, -1, 3, -2, 0, -10, 4, 8, 7,
    -- filter=19 channel=98
    -1, -15, -8, -8, -4, 11, -6, 13, 7,
    -- filter=19 channel=99
    3, -21, -15, -4, -5, 3, 4, 18, 15,
    -- filter=19 channel=100
    -8, -6, -6, -3, -8, -10, 1, 4, -4,
    -- filter=19 channel=101
    -1, -5, 10, 0, 16, 11, 9, 4, 6,
    -- filter=19 channel=102
    5, -1, 0, -3, -2, 2, -5, -5, 6,
    -- filter=19 channel=103
    -3, 0, 1, -9, -14, -1, 0, 13, 4,
    -- filter=19 channel=104
    -8, -15, -4, 0, 6, 1, 0, 10, 17,
    -- filter=19 channel=105
    8, 2, 4, -4, 2, -4, -6, -5, -4,
    -- filter=19 channel=106
    6, -3, -2, -4, 0, 0, -8, -2, -11,
    -- filter=19 channel=107
    8, -4, -2, -1, 6, 9, -7, -6, 1,
    -- filter=19 channel=108
    8, 6, 1, 6, -3, 3, -6, 0, -3,
    -- filter=19 channel=109
    4, -13, -15, -4, 11, 18, 8, 14, 9,
    -- filter=19 channel=110
    6, -7, -9, 2, -1, -9, -6, 5, 1,
    -- filter=19 channel=111
    0, 2, 3, -1, 2, -2, -5, 3, -5,
    -- filter=19 channel=112
    -4, -11, -5, 4, -1, -4, 0, 7, 7,
    -- filter=19 channel=113
    -6, -3, -4, -11, -9, 0, -8, 8, 11,
    -- filter=19 channel=114
    7, 0, -5, 0, 13, 15, 4, 0, -7,
    -- filter=19 channel=115
    2, 3, 6, -4, 5, 4, 3, -6, -1,
    -- filter=19 channel=116
    2, -15, -19, -3, 13, 15, 3, 10, 1,
    -- filter=19 channel=117
    -2, 2, -12, -4, 2, -5, 0, 0, 3,
    -- filter=19 channel=118
    -7, 3, 6, 7, -1, -4, 5, -5, -6,
    -- filter=19 channel=119
    -2, -7, -4, -7, -1, -2, 4, 2, 1,
    -- filter=19 channel=120
    4, -20, -12, -9, 21, 20, 2, 8, 10,
    -- filter=19 channel=121
    -6, -3, -8, -5, -10, -10, -3, 5, -1,
    -- filter=19 channel=122
    -13, -1, -7, -18, -2, -4, -7, 5, 12,
    -- filter=19 channel=123
    0, -3, 5, 2, 4, -1, 6, 8, -2,
    -- filter=19 channel=124
    11, 3, 2, -5, 5, 5, 1, -5, 0,
    -- filter=19 channel=125
    4, -13, -17, -5, 0, 10, 5, 9, 18,
    -- filter=19 channel=126
    -2, 1, 0, -10, -17, -13, -3, 14, 10,
    -- filter=19 channel=127
    7, -2, 0, 6, 5, 0, -1, 4, -3,
    -- filter=20 channel=0
    6, -4, -20, 10, 0, -7, -9, 16, 8,
    -- filter=20 channel=1
    -5, -15, -26, 0, -2, -7, -8, 8, 5,
    -- filter=20 channel=2
    -1, 5, 3, -9, 1, 2, 3, 1, -8,
    -- filter=20 channel=3
    6, 1, 2, 0, -5, 6, -9, 1, 11,
    -- filter=20 channel=4
    -3, 1, -7, -6, -4, 1, -13, -6, 6,
    -- filter=20 channel=5
    0, -14, -13, 6, 2, 8, 13, 25, 17,
    -- filter=20 channel=6
    9, 12, 5, 8, 4, 4, -1, -13, -5,
    -- filter=20 channel=7
    0, -2, 7, -5, -4, -4, -2, 4, 6,
    -- filter=20 channel=8
    0, 0, -4, -9, 3, 2, -8, -6, -9,
    -- filter=20 channel=9
    0, -4, 0, 4, 1, 7, 10, 5, -2,
    -- filter=20 channel=10
    -5, 0, 9, -6, 9, 12, 0, 2, -3,
    -- filter=20 channel=11
    9, 20, 16, 6, -4, 6, -3, -13, -18,
    -- filter=20 channel=12
    0, -6, -5, 0, 3, 1, -12, -6, 0,
    -- filter=20 channel=13
    -2, 7, 1, 2, 3, 3, -5, -8, -15,
    -- filter=20 channel=14
    0, 0, -1, -1, 4, 4, -1, 1, -7,
    -- filter=20 channel=15
    4, 19, 15, -7, 1, 7, -14, -28, -20,
    -- filter=20 channel=16
    -6, -18, -17, -5, 4, -5, 7, 15, 16,
    -- filter=20 channel=17
    -7, 3, -1, 0, -6, 6, 7, 4, 4,
    -- filter=20 channel=18
    8, 15, 13, -4, 14, 1, -11, -21, -14,
    -- filter=20 channel=19
    -2, -3, 2, -2, 3, -1, -4, -5, -5,
    -- filter=20 channel=20
    8, 22, 26, 5, 2, 6, 0, -24, -25,
    -- filter=20 channel=21
    -8, -16, -17, -8, 0, 4, 12, 25, 19,
    -- filter=20 channel=22
    -3, 7, 7, 3, 4, 6, 2, -3, -12,
    -- filter=20 channel=23
    7, 19, 30, 0, 9, 17, -11, -22, -14,
    -- filter=20 channel=24
    0, -1, 1, 0, 0, -5, 5, 0, -2,
    -- filter=20 channel=25
    -1, -4, 5, -5, 6, 0, 3, -1, -11,
    -- filter=20 channel=26
    -5, -17, -20, -7, 2, 0, 0, 10, 9,
    -- filter=20 channel=27
    0, 15, 14, 2, -3, 4, -7, -13, -22,
    -- filter=20 channel=28
    -4, 6, 0, 3, 2, -5, 6, -6, 6,
    -- filter=20 channel=29
    7, 26, 27, 4, 6, 7, -6, -16, -7,
    -- filter=20 channel=30
    -10, -6, -2, -8, -4, 0, -4, 9, 0,
    -- filter=20 channel=31
    -10, 2, 2, -3, 0, 4, 12, 20, 8,
    -- filter=20 channel=32
    4, 5, 17, -5, 5, 4, -15, -9, -16,
    -- filter=20 channel=33
    2, 2, 2, -1, 0, 7, -7, 0, -2,
    -- filter=20 channel=34
    4, 3, -7, 1, 8, -2, -1, 11, -1,
    -- filter=20 channel=35
    2, 4, -7, 4, -3, 6, 5, -3, -4,
    -- filter=20 channel=36
    -6, -3, -1, -9, -12, -8, -8, -1, 4,
    -- filter=20 channel=37
    3, -17, -23, 6, 0, -1, 0, 22, 22,
    -- filter=20 channel=38
    1, 0, 8, 0, 11, 12, 0, 3, -9,
    -- filter=20 channel=39
    -2, 9, 8, -3, 0, 1, -3, -4, -4,
    -- filter=20 channel=40
    0, 5, 11, 2, 4, -1, -1, -4, -10,
    -- filter=20 channel=41
    0, 1, -6, -5, 8, -9, -16, 19, 0,
    -- filter=20 channel=42
    -4, 0, -2, 0, 3, -4, -2, 1, 7,
    -- filter=20 channel=43
    -2, 3, 6, -6, 2, 3, -8, -15, -7,
    -- filter=20 channel=44
    -6, -4, -14, -2, 7, 1, 5, 20, 6,
    -- filter=20 channel=45
    2, -1, 5, -2, -2, -3, 0, 4, 0,
    -- filter=20 channel=46
    -5, -1, -1, 0, 1, -1, 5, -3, 3,
    -- filter=20 channel=47
    -6, -20, -23, 4, 5, 0, 9, 36, 13,
    -- filter=20 channel=48
    -3, -11, -17, -3, 0, -4, 8, 8, -9,
    -- filter=20 channel=49
    5, 1, 1, -1, 0, 0, -4, -8, -7,
    -- filter=20 channel=50
    -6, 8, 8, 2, 8, 2, 2, -8, -14,
    -- filter=20 channel=51
    5, 0, -1, 0, -3, -3, -3, -5, 2,
    -- filter=20 channel=52
    0, 6, 12, -10, -8, 4, -2, -1, -9,
    -- filter=20 channel=53
    -2, 8, 18, 7, 2, 7, -5, -13, 0,
    -- filter=20 channel=54
    -5, -3, 3, 3, 1, 7, -6, -6, 1,
    -- filter=20 channel=55
    4, 13, 24, 0, 2, 13, -8, -24, -24,
    -- filter=20 channel=56
    -4, 4, -3, -10, 3, -6, 3, -3, -8,
    -- filter=20 channel=57
    -5, -2, -6, 2, 7, -6, 0, 0, 2,
    -- filter=20 channel=58
    -8, -2, -15, 1, -4, 0, 0, 5, 14,
    -- filter=20 channel=59
    -10, -5, 2, -7, -3, -2, 7, 11, -8,
    -- filter=20 channel=60
    4, -3, 0, -5, -3, -3, 1, -2, 8,
    -- filter=20 channel=61
    1, 0, 0, -4, -3, -3, 0, 1, -2,
    -- filter=20 channel=62
    -5, 0, 2, 5, 6, -2, -3, -1, 0,
    -- filter=20 channel=63
    0, -14, -15, 5, 5, 3, 6, 15, 16,
    -- filter=20 channel=64
    -2, -4, -2, -6, -6, 0, 2, -7, -5,
    -- filter=20 channel=65
    -6, -3, -2, 6, -6, -2, -5, -6, 1,
    -- filter=20 channel=66
    -2, 2, -4, -12, 7, 9, 0, 8, 6,
    -- filter=20 channel=67
    -5, -2, -4, -3, 4, -2, 7, 4, 0,
    -- filter=20 channel=68
    0, -7, -8, -5, 0, -9, 4, -7, 2,
    -- filter=20 channel=69
    3, -6, -2, 1, -5, -1, -4, 4, 9,
    -- filter=20 channel=70
    0, 9, 14, -1, 7, -4, -3, -20, -18,
    -- filter=20 channel=71
    0, -5, 2, -8, 5, 3, -4, 7, 3,
    -- filter=20 channel=72
    -7, 0, 6, 6, 2, 0, 12, -1, 2,
    -- filter=20 channel=73
    4, 7, 8, -9, 5, 6, -7, -15, -16,
    -- filter=20 channel=74
    2, 10, 8, -6, 2, -2, -4, -6, 0,
    -- filter=20 channel=75
    0, -14, -17, 7, 13, 9, -6, 19, 21,
    -- filter=20 channel=76
    4, 16, 22, -4, -2, -2, -5, -23, -10,
    -- filter=20 channel=77
    -1, 2, 0, 6, 7, 5, -5, 6, 7,
    -- filter=20 channel=78
    -3, 1, -8, 8, 0, 1, -4, 11, 12,
    -- filter=20 channel=79
    10, 7, 17, 7, 4, 4, -5, -26, -26,
    -- filter=20 channel=80
    -15, -11, -2, 4, 4, 7, 3, 26, 12,
    -- filter=20 channel=81
    0, 2, 0, -3, -4, 6, -6, 1, -3,
    -- filter=20 channel=82
    0, 3, -2, 2, -4, -2, -2, -2, 7,
    -- filter=20 channel=83
    1, -5, -2, -10, -7, 3, 4, 0, -2,
    -- filter=20 channel=84
    4, 9, 15, 1, -4, 1, -1, -12, -12,
    -- filter=20 channel=85
    4, -5, -2, -2, 2, 3, -5, -5, 4,
    -- filter=20 channel=86
    -1, -9, -4, -3, -5, 6, -2, 4, 7,
    -- filter=20 channel=87
    4, 0, 11, 0, -5, 6, -5, -12, -10,
    -- filter=20 channel=88
    -4, 4, -9, -4, 2, 0, 6, 7, -1,
    -- filter=20 channel=89
    -3, 0, 11, 3, 6, 8, -7, -13, -14,
    -- filter=20 channel=90
    -10, -4, -1, -12, -5, -3, -6, -2, -2,
    -- filter=20 channel=91
    -2, 7, 13, -8, -7, -7, -10, -21, -14,
    -- filter=20 channel=92
    8, -3, 0, -1, 0, 1, 1, 3, 0,
    -- filter=20 channel=93
    -1, -10, -27, -8, -8, -9, 0, 17, 6,
    -- filter=20 channel=94
    7, -6, 1, -2, 2, -6, -3, -3, -5,
    -- filter=20 channel=95
    -5, 2, 6, -1, 4, -2, 4, -2, 2,
    -- filter=20 channel=96
    -2, -2, -4, 2, -5, 3, -8, 4, 4,
    -- filter=20 channel=97
    3, 4, 2, 2, 4, -2, -4, 7, -2,
    -- filter=20 channel=98
    -2, -2, 8, 5, 11, 2, 12, 0, 0,
    -- filter=20 channel=99
    -7, 8, 18, -7, 7, 8, -6, -13, -7,
    -- filter=20 channel=100
    2, -4, 0, 2, 0, -5, -1, 1, 6,
    -- filter=20 channel=101
    -7, -4, 6, -5, -2, -5, -8, 4, -5,
    -- filter=20 channel=102
    0, 1, 0, 3, 6, 0, -6, 1, 4,
    -- filter=20 channel=103
    -4, -10, -20, 9, 9, -1, 12, 30, 13,
    -- filter=20 channel=104
    -6, -13, -4, 4, 8, 6, 2, 21, 5,
    -- filter=20 channel=105
    -1, 11, 17, -1, 1, 6, 2, -8, -11,
    -- filter=20 channel=106
    6, 1, -3, -3, 6, -7, -5, -1, -8,
    -- filter=20 channel=107
    5, 20, 20, -3, -1, 0, -4, -29, -14,
    -- filter=20 channel=108
    9, -4, -6, 6, -1, -3, -3, 14, 4,
    -- filter=20 channel=109
    0, 5, 14, -5, 7, 0, -6, -8, -13,
    -- filter=20 channel=110
    2, 4, 1, -8, 6, 6, -3, -2, 12,
    -- filter=20 channel=111
    -6, 6, -1, 0, -2, -7, 2, 2, 5,
    -- filter=20 channel=112
    -1, 5, -5, 2, -1, 0, 3, 9, 4,
    -- filter=20 channel=113
    0, 7, 4, -9, 0, 4, 4, -3, -3,
    -- filter=20 channel=114
    10, 16, 13, 6, 5, -1, -13, -15, -14,
    -- filter=20 channel=115
    -4, 5, -6, -5, 3, -2, 4, 0, -3,
    -- filter=20 channel=116
    -9, 2, 8, 4, -13, -10, 4, -9, -11,
    -- filter=20 channel=117
    5, 5, 0, 5, -6, -6, -6, 3, 2,
    -- filter=20 channel=118
    -4, 5, -2, -7, 4, 3, 2, -3, -2,
    -- filter=20 channel=119
    -5, 0, -4, -2, -8, 4, -5, 6, -7,
    -- filter=20 channel=120
    7, 19, 21, 3, 0, 3, -12, -25, -23,
    -- filter=20 channel=121
    -3, 4, -5, 0, 1, 8, -8, 6, 0,
    -- filter=20 channel=122
    -28, -37, -31, -6, -2, 0, 11, 43, 27,
    -- filter=20 channel=123
    6, 0, 1, -4, -4, -1, 4, 5, -10,
    -- filter=20 channel=124
    8, 0, 9, 6, 4, 0, 3, -14, -4,
    -- filter=20 channel=125
    -13, 0, 13, 0, 0, 3, 3, -8, -4,
    -- filter=20 channel=126
    4, 2, 8, 0, 3, 11, 5, -3, -9,
    -- filter=20 channel=127
    -2, 6, 3, 6, 2, 7, -4, 7, -6,
    -- filter=21 channel=0
    4, -10, 1, 10, -2, 3, 16, 4, 1,
    -- filter=21 channel=1
    0, -5, -7, 1, -5, -4, 6, -6, 9,
    -- filter=21 channel=2
    6, 6, 6, -3, 3, -7, 2, -3, 0,
    -- filter=21 channel=3
    -2, -9, 1, 19, 8, -4, 1, 9, -5,
    -- filter=21 channel=4
    3, 1, -5, -2, -12, -7, 10, 7, -2,
    -- filter=21 channel=5
    -5, -8, 7, -3, -7, 10, 7, 0, -2,
    -- filter=21 channel=6
    -8, 2, -7, -5, 8, -5, -5, 5, 3,
    -- filter=21 channel=7
    -1, -1, -1, -5, 4, 3, 6, 1, -3,
    -- filter=21 channel=8
    0, -2, -7, 0, -5, 0, -3, 5, -3,
    -- filter=21 channel=9
    7, -5, 2, 6, -6, 6, -1, 1, 0,
    -- filter=21 channel=10
    10, 7, 5, -1, 0, -3, -8, -5, -1,
    -- filter=21 channel=11
    2, 5, 6, -4, 1, 6, 4, 14, -1,
    -- filter=21 channel=12
    -3, -5, -3, -4, -6, -6, 0, -3, -1,
    -- filter=21 channel=13
    3, 5, 0, -2, 2, -5, -10, -1, 0,
    -- filter=21 channel=14
    6, -6, 2, 3, 0, -3, 2, 0, -4,
    -- filter=21 channel=15
    5, -1, -10, 9, 2, 2, -13, 4, 0,
    -- filter=21 channel=16
    3, 4, 6, -6, 3, -7, -9, -5, 0,
    -- filter=21 channel=17
    4, -3, -1, -4, 2, 0, -2, -4, -3,
    -- filter=21 channel=18
    9, 0, -8, 5, 9, -7, -11, 0, 0,
    -- filter=21 channel=19
    -7, -5, 5, 2, -4, -1, 3, 4, 6,
    -- filter=21 channel=20
    -11, 0, -9, -3, 5, 3, 1, 10, 9,
    -- filter=21 channel=21
    7, 9, 4, 1, -4, 5, -12, -17, -2,
    -- filter=21 channel=22
    0, 2, 2, 2, -3, -2, 7, 9, 0,
    -- filter=21 channel=23
    -2, -4, 0, 11, -3, -3, -5, 6, -9,
    -- filter=21 channel=24
    1, 2, 0, 5, 0, 0, 0, -2, 5,
    -- filter=21 channel=25
    10, 7, -4, -1, 0, -1, -6, -4, -7,
    -- filter=21 channel=26
    1, 5, 2, 0, -4, -1, 6, -5, -1,
    -- filter=21 channel=27
    15, 1, -5, 8, 5, 1, -18, -7, -10,
    -- filter=21 channel=28
    -4, 0, 0, -2, -7, -2, -6, 2, -2,
    -- filter=21 channel=29
    -3, -8, 2, -2, 0, 4, -3, 10, 4,
    -- filter=21 channel=30
    1, 3, 7, 1, 0, 5, -7, 4, 5,
    -- filter=21 channel=31
    14, 5, 0, 9, -2, -5, -10, -9, -10,
    -- filter=21 channel=32
    1, -7, -2, 0, 8, -1, -11, 3, 0,
    -- filter=21 channel=33
    13, 7, -1, 14, 5, -3, -11, 7, 3,
    -- filter=21 channel=34
    -4, -10, -1, 5, -3, 1, 2, -3, -6,
    -- filter=21 channel=35
    -5, -6, -2, -5, -2, 7, 6, -6, -2,
    -- filter=21 channel=36
    2, 0, 0, 0, 0, -7, -1, 0, -2,
    -- filter=21 channel=37
    0, -5, 8, 1, -2, 2, 3, 3, -3,
    -- filter=21 channel=38
    0, -1, 0, 5, 1, 1, -4, 0, -6,
    -- filter=21 channel=39
    -7, -3, 1, 4, -5, 0, -7, 10, 2,
    -- filter=21 channel=40
    5, 5, -2, -4, 0, -3, -6, 0, -5,
    -- filter=21 channel=41
    2, 1, -12, -2, -4, -7, 6, -7, -12,
    -- filter=21 channel=42
    5, -5, 3, 4, 4, 5, 6, -6, -6,
    -- filter=21 channel=43
    -4, -1, -4, 11, 3, -6, 4, 11, -3,
    -- filter=21 channel=44
    -1, 1, 10, 0, -3, 1, 2, -5, 4,
    -- filter=21 channel=45
    4, -3, 0, -6, -2, -1, 3, -3, 0,
    -- filter=21 channel=46
    6, -6, 1, -2, 5, 5, 5, 0, 1,
    -- filter=21 channel=47
    7, 5, 6, -2, -1, 5, 0, -10, -2,
    -- filter=21 channel=48
    2, 5, 0, -1, -1, 5, -10, -13, 0,
    -- filter=21 channel=49
    -4, -4, -2, -9, 6, -11, -12, 0, 4,
    -- filter=21 channel=50
    8, -5, 9, 4, -3, -7, -3, 2, 2,
    -- filter=21 channel=51
    -7, -4, 6, -6, 0, -4, -3, 3, -1,
    -- filter=21 channel=52
    2, -1, -4, 0, 0, -1, 6, -4, -5,
    -- filter=21 channel=53
    -1, -6, 1, 0, -3, -6, 0, 0, 3,
    -- filter=21 channel=54
    3, 0, 5, 7, 0, 7, -3, -2, 4,
    -- filter=21 channel=55
    4, -2, -2, -6, 13, -3, -12, 4, 3,
    -- filter=21 channel=56
    5, 3, -1, -1, -7, -3, -6, 3, 0,
    -- filter=21 channel=57
    -7, -3, -8, 5, -4, -2, 3, -2, 3,
    -- filter=21 channel=58
    -8, -1, 7, -4, 0, 0, 4, 0, -6,
    -- filter=21 channel=59
    12, 10, -1, 6, 5, 1, -14, -2, -10,
    -- filter=21 channel=60
    0, 3, 0, 1, 4, 0, 6, 2, 1,
    -- filter=21 channel=61
    7, 5, -6, -6, -1, -2, -7, -1, 4,
    -- filter=21 channel=62
    0, 0, -7, -4, 6, 4, -2, -6, 3,
    -- filter=21 channel=63
    1, -6, -2, 2, -6, -3, -2, 0, -2,
    -- filter=21 channel=64
    6, 3, -6, 4, 5, -5, -8, -2, -1,
    -- filter=21 channel=65
    5, 4, 0, 5, -6, 2, -1, -4, 0,
    -- filter=21 channel=66
    6, 6, 2, -2, -4, 0, 0, -3, -4,
    -- filter=21 channel=67
    -7, -1, 0, 2, -7, 7, 1, -4, -5,
    -- filter=21 channel=68
    4, 3, -4, -7, 5, -5, 0, -6, -3,
    -- filter=21 channel=69
    0, -4, 0, -1, -2, 1, 0, 4, -4,
    -- filter=21 channel=70
    5, -5, -7, 10, -8, -9, -6, 2, -11,
    -- filter=21 channel=71
    5, 0, -4, 3, -4, 3, -4, -3, -3,
    -- filter=21 channel=72
    13, 1, -4, 7, 8, 3, -3, -4, -4,
    -- filter=21 channel=73
    -2, -1, 3, -10, 3, 0, -5, -4, 0,
    -- filter=21 channel=74
    6, -8, 4, 1, -6, -9, -3, 0, -4,
    -- filter=21 channel=75
    0, -6, -5, 8, 4, -1, 6, -2, 1,
    -- filter=21 channel=76
    -7, 3, -3, 0, 6, 4, 0, 14, 5,
    -- filter=21 channel=77
    -7, 4, -3, 3, 0, -4, 0, 7, -5,
    -- filter=21 channel=78
    6, 0, -6, 1, -6, -5, 1, -7, -2,
    -- filter=21 channel=79
    7, -3, -11, 7, 7, -1, -12, 5, 3,
    -- filter=21 channel=80
    20, 4, 9, 11, 1, -3, -16, -13, -9,
    -- filter=21 channel=81
    0, 2, 0, 5, 0, 3, -6, -4, 2,
    -- filter=21 channel=82
    0, -1, 0, 6, 7, -3, 3, 5, 6,
    -- filter=21 channel=83
    -1, -2, 1, 1, -6, -2, -6, 0, 3,
    -- filter=21 channel=84
    6, -5, -7, -6, -7, -1, -1, -4, 0,
    -- filter=21 channel=85
    2, 6, -2, 1, 4, 7, -5, 0, 2,
    -- filter=21 channel=86
    0, -9, 4, 2, -6, -6, 1, -3, -1,
    -- filter=21 channel=87
    -3, 1, 1, -4, 0, -3, 0, 2, -8,
    -- filter=21 channel=88
    0, 4, -4, 2, 5, -8, 4, 2, -2,
    -- filter=21 channel=89
    6, 12, -4, 13, 11, -5, -6, -7, 0,
    -- filter=21 channel=90
    6, 2, 3, 7, -8, -2, 0, -5, -9,
    -- filter=21 channel=91
    -2, -4, 1, 0, -2, -8, -4, 8, -8,
    -- filter=21 channel=92
    0, -4, 4, 0, 3, -6, -5, -7, -8,
    -- filter=21 channel=93
    10, -1, 0, -8, -7, -5, 1, -9, 3,
    -- filter=21 channel=94
    -3, 6, 4, -7, 1, -3, 0, -7, -3,
    -- filter=21 channel=95
    6, 0, -7, 1, 0, -4, -5, 2, -4,
    -- filter=21 channel=96
    -3, 0, -2, 3, 0, 4, 3, -8, 1,
    -- filter=21 channel=97
    0, -8, -2, 7, 4, 3, 7, 0, -5,
    -- filter=21 channel=98
    7, -1, -4, 4, 9, -5, -11, -7, -10,
    -- filter=21 channel=99
    13, 8, 5, 4, -6, -5, -16, 0, -15,
    -- filter=21 channel=100
    2, -6, 0, 6, -6, -7, -5, 0, -2,
    -- filter=21 channel=101
    4, -9, 0, 2, 4, -2, 0, 3, 0,
    -- filter=21 channel=102
    3, 0, -1, -4, 5, -1, 6, -2, 7,
    -- filter=21 channel=103
    7, 8, -1, 12, -7, 10, -9, -13, -9,
    -- filter=21 channel=104
    16, 10, 8, 6, 3, -1, -4, -3, -3,
    -- filter=21 channel=105
    3, 0, 0, -3, 5, 0, 3, 14, 11,
    -- filter=21 channel=106
    -3, 5, -3, 2, -2, 3, -3, 7, 0,
    -- filter=21 channel=107
    -5, -6, 0, 1, 5, 5, 0, 4, 5,
    -- filter=21 channel=108
    -8, -6, -4, -3, 4, 1, 6, 0, 4,
    -- filter=21 channel=109
    13, -1, -6, -7, -2, -1, -19, -6, 0,
    -- filter=21 channel=110
    9, -4, 1, -1, -5, -2, -5, 0, -4,
    -- filter=21 channel=111
    1, 8, -2, -1, 0, -7, 0, -2, 0,
    -- filter=21 channel=112
    2, 1, -3, 7, -9, -5, 0, 0, 0,
    -- filter=21 channel=113
    7, 7, 2, 8, -1, 7, 2, 0, -7,
    -- filter=21 channel=114
    4, -11, -7, 4, -1, -5, -6, 10, 7,
    -- filter=21 channel=115
    -1, 6, 0, -4, -7, 0, 3, 0, 2,
    -- filter=21 channel=116
    7, 3, 3, 0, 4, -1, -13, 0, 0,
    -- filter=21 channel=117
    -6, 0, 5, 4, 0, 6, -4, 3, 3,
    -- filter=21 channel=118
    7, -3, -6, 3, 4, 5, -6, 0, 0,
    -- filter=21 channel=119
    -2, -6, 6, -2, -10, -10, 0, 2, -11,
    -- filter=21 channel=120
    0, 0, 3, -14, -1, 3, -4, 9, 0,
    -- filter=21 channel=121
    1, 2, 4, 1, -1, 0, -4, 0, -4,
    -- filter=21 channel=122
    0, 1, 12, 4, -8, 10, -15, -11, -10,
    -- filter=21 channel=123
    0, -4, -5, 6, 2, -1, 4, 0, -10,
    -- filter=21 channel=124
    0, 4, -5, -5, 8, -3, -4, 10, 2,
    -- filter=21 channel=125
    16, 4, -1, 5, 0, 3, -17, -9, -10,
    -- filter=21 channel=126
    4, -1, 0, 9, 0, 1, -7, -7, 1,
    -- filter=21 channel=127
    -2, 8, 2, 3, -6, -6, 4, -3, -8,
    -- filter=22 channel=0
    -3, 0, 4, -12, 1, -3, 1, 2, 0,
    -- filter=22 channel=1
    -4, 1, 8, -2, 0, -3, 9, 4, 7,
    -- filter=22 channel=2
    0, -1, -5, 4, 1, 1, 7, -1, 5,
    -- filter=22 channel=3
    0, 2, -2, -3, 5, 9, -6, 7, 8,
    -- filter=22 channel=4
    0, -14, -4, -1, -7, -4, 17, 4, 6,
    -- filter=22 channel=5
    -2, -5, -3, 4, 3, -4, 6, 12, 4,
    -- filter=22 channel=6
    -7, -2, -5, -2, 1, 0, -2, 2, -7,
    -- filter=22 channel=7
    -7, 3, -6, 1, -3, 4, -1, -6, 3,
    -- filter=22 channel=8
    -3, -1, 1, -1, 7, -5, -5, -3, -6,
    -- filter=22 channel=9
    -1, -1, 0, 1, -3, 1, -7, -8, -8,
    -- filter=22 channel=10
    5, 14, 7, -9, 4, 3, -8, -4, -1,
    -- filter=22 channel=11
    -3, 1, 3, -7, -2, -3, -6, -4, -8,
    -- filter=22 channel=12
    3, 3, -5, 2, 10, 0, 7, 0, -1,
    -- filter=22 channel=13
    0, 8, 6, -5, 10, 3, 0, -4, -6,
    -- filter=22 channel=14
    6, -1, -5, 5, 6, 5, 1, -4, -2,
    -- filter=22 channel=15
    -10, 3, 8, -16, 3, 7, 0, 1, -12,
    -- filter=22 channel=16
    8, 4, -1, 5, 5, 6, 4, 8, -5,
    -- filter=22 channel=17
    3, -6, 5, -6, -4, 7, 0, 4, -6,
    -- filter=22 channel=18
    -10, 3, 10, -18, 5, 1, -10, 1, -2,
    -- filter=22 channel=19
    -3, 6, 0, -6, 1, 5, 7, -5, 6,
    -- filter=22 channel=20
    -9, 9, 0, 0, 11, -3, 0, -3, -5,
    -- filter=22 channel=21
    8, 11, 4, 3, 6, 6, -1, -7, -3,
    -- filter=22 channel=22
    -1, 11, 3, -8, 6, 0, -4, -4, -9,
    -- filter=22 channel=23
    6, 19, 7, -6, 24, -4, -18, -2, -14,
    -- filter=22 channel=24
    -3, 0, -6, 1, -4, 7, -2, 5, -4,
    -- filter=22 channel=25
    -6, 13, 0, -17, -1, 3, 0, -11, 0,
    -- filter=22 channel=26
    6, 7, -9, 7, 9, -6, -1, 4, -3,
    -- filter=22 channel=27
    -3, 15, -2, -20, 11, -2, 0, -2, -10,
    -- filter=22 channel=28
    7, -1, -6, 5, 0, -4, 3, -1, 5,
    -- filter=22 channel=29
    -9, 8, 0, -4, -2, 3, -2, 0, 1,
    -- filter=22 channel=30
    -3, -1, -6, -12, 3, 2, 2, -7, -13,
    -- filter=22 channel=31
    0, 17, -8, -6, 12, 2, -9, -13, -19,
    -- filter=22 channel=32
    -16, 15, 4, -19, 12, 8, -7, 0, -12,
    -- filter=22 channel=33
    -7, 12, 11, -15, 8, 1, -16, 4, -3,
    -- filter=22 channel=34
    6, 15, 6, 6, 16, 7, -6, 7, -8,
    -- filter=22 channel=35
    1, -7, 5, -6, 0, -4, 0, 0, -1,
    -- filter=22 channel=36
    0, 1, 3, 5, -2, -1, 0, 1, 0,
    -- filter=22 channel=37
    -5, 7, 6, -4, 2, -3, 0, 14, 0,
    -- filter=22 channel=38
    -4, 0, 1, -9, 12, -5, 0, -3, -8,
    -- filter=22 channel=39
    -4, 9, -5, -3, -3, -6, 5, 0, 4,
    -- filter=22 channel=40
    5, 9, 6, -2, 10, 7, 2, -6, -1,
    -- filter=22 channel=41
    -10, 6, 13, -3, 4, 6, -10, 3, -1,
    -- filter=22 channel=42
    -7, -5, 4, -3, -6, 0, -5, -5, -4,
    -- filter=22 channel=43
    7, 4, -2, 0, 9, -1, -5, 2, 6,
    -- filter=22 channel=44
    -1, 3, 7, -3, 9, 1, 5, -3, 0,
    -- filter=22 channel=45
    0, 3, 5, 2, -2, 3, -4, -1, 6,
    -- filter=22 channel=46
    6, -4, -3, 6, 0, -4, 1, -2, -3,
    -- filter=22 channel=47
    2, 8, 8, -1, 11, 0, 3, -3, -3,
    -- filter=22 channel=48
    -12, -4, 0, -10, -3, 0, 2, 1, -14,
    -- filter=22 channel=49
    -16, 1, 4, -11, 2, 3, -1, 0, 1,
    -- filter=22 channel=50
    5, 7, 0, -12, 9, -1, -10, -2, -2,
    -- filter=22 channel=51
    2, 0, 0, 4, -6, 0, -6, -3, -4,
    -- filter=22 channel=52
    5, 17, 4, -1, 13, 4, 0, -4, 1,
    -- filter=22 channel=53
    -6, 5, 4, -8, -2, 0, 0, 3, -1,
    -- filter=22 channel=54
    0, 2, -4, 3, 3, -1, -2, 0, 2,
    -- filter=22 channel=55
    0, 10, 7, -17, 0, 9, -10, -8, -17,
    -- filter=22 channel=56
    10, 1, 8, -5, 9, -1, -8, -3, -4,
    -- filter=22 channel=57
    -6, -1, -1, 6, -2, -6, -4, -3, 4,
    -- filter=22 channel=58
    4, 0, -6, 5, 0, 1, 7, 3, 5,
    -- filter=22 channel=59
    -13, 10, -3, -7, 3, 4, -8, -8, -14,
    -- filter=22 channel=60
    -3, -6, 4, -1, -7, 2, -3, -4, 2,
    -- filter=22 channel=61
    -2, -2, -2, -3, 10, -5, 5, 0, -2,
    -- filter=22 channel=62
    5, 0, -1, 0, 0, 1, -7, -4, 7,
    -- filter=22 channel=63
    -1, -8, -4, -1, -3, -8, 6, 8, -6,
    -- filter=22 channel=64
    -3, -3, -4, -2, 6, -6, 5, -4, 5,
    -- filter=22 channel=65
    3, 6, -3, -6, 1, 1, 0, 0, 6,
    -- filter=22 channel=66
    -1, 18, 1, 1, 11, -5, 6, 0, -5,
    -- filter=22 channel=67
    0, -6, 2, 7, -5, -2, -7, 5, 5,
    -- filter=22 channel=68
    3, 5, -7, -7, 2, 3, 3, 3, 3,
    -- filter=22 channel=69
    0, -2, -4, -2, -5, -3, 4, -8, 7,
    -- filter=22 channel=70
    3, 13, 7, -18, 7, 1, -8, -9, -9,
    -- filter=22 channel=71
    0, 0, 4, -3, 3, 0, 0, 2, -2,
    -- filter=22 channel=72
    -9, 8, 1, -5, -2, 3, -5, -4, -17,
    -- filter=22 channel=73
    0, -1, 4, -14, 1, 4, -5, 5, -3,
    -- filter=22 channel=74
    8, 19, -2, -3, 7, -3, 3, 5, -10,
    -- filter=22 channel=75
    0, 12, 10, -12, -1, 7, -10, 11, 13,
    -- filter=22 channel=76
    5, 6, 7, -8, 5, 0, -8, 0, -1,
    -- filter=22 channel=77
    3, 6, -7, 5, -6, 0, -4, 0, 4,
    -- filter=22 channel=78
    4, 2, -7, 4, 9, 3, -5, -4, -5,
    -- filter=22 channel=79
    -13, 14, 9, -29, 7, 12, -1, -3, -15,
    -- filter=22 channel=80
    -8, 8, 2, -13, 2, 4, -8, -11, -9,
    -- filter=22 channel=81
    -4, -6, 6, 0, 3, 0, 6, -1, -3,
    -- filter=22 channel=82
    5, 0, 5, 5, -2, -5, -2, 0, -5,
    -- filter=22 channel=83
    -7, -6, -8, -4, 0, -5, -1, -2, -3,
    -- filter=22 channel=84
    -12, 1, 5, -12, 9, 4, -4, 3, -13,
    -- filter=22 channel=85
    1, 0, -3, 6, 0, -6, 0, -2, -2,
    -- filter=22 channel=86
    4, 3, -4, -9, 3, 5, -5, 9, 6,
    -- filter=22 channel=87
    6, 8, 4, 0, 11, 7, -3, 7, 3,
    -- filter=22 channel=88
    10, 9, 0, 8, 2, -9, 1, 2, -8,
    -- filter=22 channel=89
    -6, 17, 9, -20, 1, 12, -13, -8, -13,
    -- filter=22 channel=90
    17, 12, 6, 13, 10, 0, -4, -2, 1,
    -- filter=22 channel=91
    -15, 12, -2, -22, 10, -2, 5, -2, -13,
    -- filter=22 channel=92
    0, 11, 3, 8, 6, 8, -8, -4, -1,
    -- filter=22 channel=93
    -4, 8, -7, -8, 3, 2, 4, 0, -10,
    -- filter=22 channel=94
    -6, -7, -1, -1, -2, -3, 0, -4, -4,
    -- filter=22 channel=95
    0, 3, 4, -4, -2, 7, -2, 6, -7,
    -- filter=22 channel=96
    -3, 2, 3, -2, -7, -5, -3, -1, -3,
    -- filter=22 channel=97
    10, 3, 4, -5, 2, 5, 1, -2, 0,
    -- filter=22 channel=98
    -2, 15, -1, -27, 12, 9, -15, -3, -15,
    -- filter=22 channel=99
    11, 22, -7, -7, 11, -3, -19, -1, -19,
    -- filter=22 channel=100
    3, -4, 1, -1, 0, 4, -2, -6, -1,
    -- filter=22 channel=101
    0, -3, 0, -3, -6, -4, 6, 8, -2,
    -- filter=22 channel=102
    -5, -3, 4, 6, 4, -5, -5, -1, 1,
    -- filter=22 channel=103
    8, 10, 5, -3, 6, 1, -9, 1, 5,
    -- filter=22 channel=104
    -3, 2, -3, -7, 3, -7, 1, -11, -6,
    -- filter=22 channel=105
    2, 8, 2, -7, -3, 8, -7, -1, -5,
    -- filter=22 channel=106
    4, 1, 6, -2, -5, 1, 2, 0, 4,
    -- filter=22 channel=107
    6, 12, -4, -4, 5, 3, -6, -3, 1,
    -- filter=22 channel=108
    -4, 0, 3, -4, -4, 5, 4, -5, -1,
    -- filter=22 channel=109
    -5, 6, 0, -23, 10, 4, -9, 0, -9,
    -- filter=22 channel=110
    6, 7, 7, -9, 9, -7, -4, -5, -9,
    -- filter=22 channel=111
    5, -1, 6, -4, -7, 0, 0, -6, 1,
    -- filter=22 channel=112
    -3, 12, -5, -10, 4, 0, 0, -2, 1,
    -- filter=22 channel=113
    1, 5, 1, -11, 7, 0, -5, -1, -2,
    -- filter=22 channel=114
    -21, 14, 3, -26, 4, -3, -5, 1, -18,
    -- filter=22 channel=115
    -6, 4, 4, 4, -1, 4, 3, 5, 0,
    -- filter=22 channel=116
    -16, 9, -2, -7, 1, 0, -7, 0, -13,
    -- filter=22 channel=117
    3, -2, 2, 1, 0, 0, -4, 0, -5,
    -- filter=22 channel=118
    -5, -6, 0, 6, -7, -6, 4, 0, 4,
    -- filter=22 channel=119
    14, 6, 4, -3, 10, 1, -1, 8, -3,
    -- filter=22 channel=120
    -3, 18, 0, -21, 3, -5, 0, -11, -25,
    -- filter=22 channel=121
    -3, 9, 10, -5, 8, 2, -11, 3, 0,
    -- filter=22 channel=122
    6, 9, 10, 0, 13, -4, -5, 8, -9,
    -- filter=22 channel=123
    10, 10, 0, 4, 1, 3, -3, 5, -1,
    -- filter=22 channel=124
    1, 9, -5, 1, 0, -1, -5, 0, -5,
    -- filter=22 channel=125
    -10, 14, 4, -11, 3, 4, 0, -5, -12,
    -- filter=22 channel=126
    -12, 10, 7, -11, 3, 9, -10, 3, -2,
    -- filter=22 channel=127
    7, -4, 4, -4, 5, 7, 2, -6, 1,
    -- filter=23 channel=0
    -16, -2, 7, -13, 13, 10, 3, 14, 19,
    -- filter=23 channel=1
    -4, -11, 1, -10, 13, 13, 8, 4, 16,
    -- filter=23 channel=2
    -2, -5, 0, 0, -2, 1, 0, 1, -3,
    -- filter=23 channel=3
    9, 8, 4, -9, 6, 0, -5, 3, 10,
    -- filter=23 channel=4
    8, 8, 6, -10, -6, -2, -1, 2, -6,
    -- filter=23 channel=5
    -15, 8, 3, -3, 15, 21, 6, 19, 21,
    -- filter=23 channel=6
    -7, -2, -4, 11, 5, 5, 7, -3, 0,
    -- filter=23 channel=7
    2, 2, 5, -3, -3, 7, 3, 7, 4,
    -- filter=23 channel=8
    3, 4, -9, 0, 0, -3, 2, -9, -5,
    -- filter=23 channel=9
    -6, 6, 3, -5, -1, 13, -5, 8, 1,
    -- filter=23 channel=10
    13, 2, -4, -3, 5, 0, -4, -1, -9,
    -- filter=23 channel=11
    -4, -1, 11, 7, 4, -5, -7, -4, -4,
    -- filter=23 channel=12
    8, -5, -19, 7, -8, -14, 4, -6, -4,
    -- filter=23 channel=13
    4, -8, -2, -5, -1, -4, 2, -9, -12,
    -- filter=23 channel=14
    5, 3, -1, 1, -2, 1, -4, 1, 0,
    -- filter=23 channel=15
    3, 8, -9, 8, 16, -3, 1, -1, -13,
    -- filter=23 channel=16
    -19, -11, 2, -16, -6, -2, -10, -9, -6,
    -- filter=23 channel=17
    -1, 2, 0, 0, 0, -7, 0, 5, 3,
    -- filter=23 channel=18
    2, 17, -7, 9, 28, 2, 0, -3, -11,
    -- filter=23 channel=19
    3, 7, 7, 3, 0, 2, -4, -3, 4,
    -- filter=23 channel=20
    -5, -6, -8, 0, 4, -1, 1, -13, -13,
    -- filter=23 channel=21
    -12, -4, 2, -15, -12, 1, -12, -14, -4,
    -- filter=23 channel=22
    -4, 3, -14, 3, 9, 0, 2, 0, -7,
    -- filter=23 channel=23
    13, 9, -16, 6, 10, -7, -2, -5, -15,
    -- filter=23 channel=24
    4, -4, -4, -5, -1, 7, -1, -6, 4,
    -- filter=23 channel=25
    2, 13, 5, -7, 8, -5, 3, -1, -6,
    -- filter=23 channel=26
    -3, -1, 2, -8, -7, 12, -7, -4, 2,
    -- filter=23 channel=27
    2, 18, -4, -10, 36, -2, 2, -1, -19,
    -- filter=23 channel=28
    -3, -5, 5, 2, -3, 4, 4, -2, 0,
    -- filter=23 channel=29
    -3, 0, 7, 9, 3, 6, 8, -3, -1,
    -- filter=23 channel=30
    0, 7, 4, -5, 10, 13, -13, -3, 9,
    -- filter=23 channel=31
    -8, -7, -4, -16, -7, 2, -23, -18, -10,
    -- filter=23 channel=32
    2, 11, 0, 4, 21, 0, -4, 4, -3,
    -- filter=23 channel=33
    0, 7, -6, -1, 22, 6, 1, 12, 0,
    -- filter=23 channel=34
    -3, -10, -16, 6, -8, -30, -2, -7, -11,
    -- filter=23 channel=35
    -3, 0, -1, 5, -3, 5, -1, 5, 2,
    -- filter=23 channel=36
    0, -12, 0, 2, -12, -13, -2, -22, -12,
    -- filter=23 channel=37
    -21, -4, 3, -6, -4, 8, 1, 4, 11,
    -- filter=23 channel=38
    5, 6, 3, 2, 9, -4, 1, 3, -9,
    -- filter=23 channel=39
    -2, 0, 8, 1, -1, 5, -7, -2, 0,
    -- filter=23 channel=40
    -14, 0, -15, -4, -6, -4, -13, -12, -13,
    -- filter=23 channel=41
    4, -5, -15, 0, -21, -18, -7, -14, -6,
    -- filter=23 channel=42
    -3, -4, 7, -3, 1, 7, 0, 0, 2,
    -- filter=23 channel=43
    3, -3, -8, 6, 7, -4, 3, -1, 4,
    -- filter=23 channel=44
    -14, -9, -5, -12, 4, 8, -14, 4, -1,
    -- filter=23 channel=45
    -2, 0, 3, -10, -1, 1, -4, 1, 7,
    -- filter=23 channel=46
    -5, 0, -3, -4, 5, 3, 1, -2, -1,
    -- filter=23 channel=47
    -24, -9, 0, -16, -6, 17, -6, 0, 1,
    -- filter=23 channel=48
    0, 7, 11, -4, 0, 8, -7, -10, 5,
    -- filter=23 channel=49
    10, 15, 0, 4, 2, -8, 1, -5, -8,
    -- filter=23 channel=50
    -1, 7, 2, -5, 14, -5, -12, 7, 0,
    -- filter=23 channel=51
    1, 1, -5, 7, -3, 1, -5, -2, 0,
    -- filter=23 channel=52
    1, 0, -17, 3, 0, -15, -2, -7, -8,
    -- filter=23 channel=53
    -7, -3, 0, 1, 2, 1, -6, 0, 3,
    -- filter=23 channel=54
    5, -5, 4, -3, 5, 6, -2, -2, -2,
    -- filter=23 channel=55
    3, 7, -9, 6, 15, -15, -8, -5, -17,
    -- filter=23 channel=56
    11, 3, -14, 0, -2, -9, 3, -9, -6,
    -- filter=23 channel=57
    6, 0, -3, 0, 0, 0, 0, -3, -7,
    -- filter=23 channel=58
    1, -8, 5, 0, 3, 7, -2, 8, 19,
    -- filter=23 channel=59
    6, 4, 3, -7, 7, 10, -6, -11, 0,
    -- filter=23 channel=60
    4, 0, 6, 4, 0, 1, 0, 0, 5,
    -- filter=23 channel=61
    -7, 3, -2, -6, 0, -7, 0, -7, -9,
    -- filter=23 channel=62
    5, 3, -4, -4, 1, -1, 0, -6, -1,
    -- filter=23 channel=63
    -3, 2, 11, -6, -4, 13, 4, 7, 18,
    -- filter=23 channel=64
    -3, -4, -3, -8, -4, -5, -9, -7, -12,
    -- filter=23 channel=65
    -1, -4, 2, -4, 2, 0, 0, 0, -1,
    -- filter=23 channel=66
    0, -2, -16, 10, -2, -18, 5, -13, -3,
    -- filter=23 channel=67
    3, -6, -3, -6, -7, 0, -5, 0, -1,
    -- filter=23 channel=68
    -6, 0, -7, -7, -10, -6, -2, -6, -8,
    -- filter=23 channel=69
    -4, -1, 0, 5, 2, 0, -2, 6, -2,
    -- filter=23 channel=70
    10, 3, -12, 2, 5, -13, -2, -6, -19,
    -- filter=23 channel=71
    6, 1, 2, -11, -2, -5, -10, 0, -3,
    -- filter=23 channel=72
    -4, 3, 2, 2, 0, -5, -3, -5, -5,
    -- filter=23 channel=73
    3, 4, 4, 3, 10, -10, 6, -2, -6,
    -- filter=23 channel=74
    -4, 6, -22, 5, 1, -22, -10, -10, -19,
    -- filter=23 channel=75
    -1, -4, 3, -17, 9, 12, 0, 18, 22,
    -- filter=23 channel=76
    -8, -7, -2, 6, 0, -7, -2, -2, -7,
    -- filter=23 channel=77
    -6, -2, -7, 5, -2, 6, 6, 4, -4,
    -- filter=23 channel=78
    2, 2, 2, -2, -6, 7, 2, 6, 11,
    -- filter=23 channel=79
    2, 13, -9, 7, 29, 1, 0, 7, -9,
    -- filter=23 channel=80
    -2, 0, 9, -16, -7, 16, -6, -6, -5,
    -- filter=23 channel=81
    0, 7, -2, 1, -5, 0, -2, 4, 4,
    -- filter=23 channel=82
    3, 4, -5, -3, 5, 5, 3, 3, -5,
    -- filter=23 channel=83
    0, 10, 4, 0, -2, -1, -3, -1, 1,
    -- filter=23 channel=84
    -5, 4, -2, -2, 13, -10, 0, 3, -3,
    -- filter=23 channel=85
    -2, 7, -7, 0, 0, -5, -6, 4, 6,
    -- filter=23 channel=86
    -5, -8, -4, -4, 9, -1, -1, 1, 2,
    -- filter=23 channel=87
    2, -2, -13, 5, -1, -3, 4, 2, -7,
    -- filter=23 channel=88
    -4, 0, -7, -8, -13, -14, -13, -7, -13,
    -- filter=23 channel=89
    8, 12, -6, -3, -1, -5, 4, -17, -6,
    -- filter=23 channel=90
    -9, -19, -14, -6, -7, -12, -6, -16, -12,
    -- filter=23 channel=91
    4, 11, -12, 2, 18, -17, -4, -3, -12,
    -- filter=23 channel=92
    -3, -1, -14, 6, -8, -4, 5, 3, -8,
    -- filter=23 channel=93
    -7, -9, 12, -12, -4, 15, -4, -1, 10,
    -- filter=23 channel=94
    -5, 5, 4, 4, 2, 2, -6, 0, -2,
    -- filter=23 channel=95
    0, 0, -5, 3, -5, -6, 0, -5, -4,
    -- filter=23 channel=96
    -4, 5, -1, 0, -5, 1, -7, 3, 5,
    -- filter=23 channel=97
    -1, 1, -5, 0, 0, 1, -4, 4, 8,
    -- filter=23 channel=98
    10, 22, 10, -8, 20, 10, 4, -4, 0,
    -- filter=23 channel=99
    9, 1, 0, 8, 15, -7, -6, -4, -13,
    -- filter=23 channel=100
    8, 4, -11, 8, -1, -4, 4, 0, -9,
    -- filter=23 channel=101
    7, -7, 1, -10, 0, -8, -6, 2, 0,
    -- filter=23 channel=102
    -7, -2, 3, 2, -5, 0, 7, 4, 0,
    -- filter=23 channel=103
    -11, 0, 2, -23, 6, 11, -7, 3, 2,
    -- filter=23 channel=104
    0, 5, -4, -11, -1, 0, -7, -5, 0,
    -- filter=23 channel=105
    -7, 0, -6, 10, 6, -1, -1, -5, -2,
    -- filter=23 channel=106
    -7, -11, -3, -1, -4, -3, -1, -7, -7,
    -- filter=23 channel=107
    -5, -3, -12, 8, 0, -1, -3, -3, -7,
    -- filter=23 channel=108
    2, -2, 1, 8, -2, 6, 7, 11, 11,
    -- filter=23 channel=109
    0, 11, -9, 10, 32, -2, 8, 2, -20,
    -- filter=23 channel=110
    2, -7, -6, -6, -5, -3, 0, -9, 1,
    -- filter=23 channel=111
    5, 0, -5, 8, 1, 3, 5, 6, 0,
    -- filter=23 channel=112
    2, 4, -5, -6, 14, 1, 1, 7, -6,
    -- filter=23 channel=113
    2, 11, 1, 0, 9, 2, -4, 0, -8,
    -- filter=23 channel=114
    -17, 16, -5, 8, 29, 13, 12, 15, -3,
    -- filter=23 channel=115
    -4, 3, -2, 6, -4, 0, -5, -5, 3,
    -- filter=23 channel=116
    10, 18, 10, -2, 4, 6, -2, -7, -13,
    -- filter=23 channel=117
    2, -5, 4, 0, -9, -8, 1, -10, 0,
    -- filter=23 channel=118
    1, 6, -1, -7, 7, 1, -8, 0, 3,
    -- filter=23 channel=119
    0, -7, -16, 16, -4, -18, -6, -1, -13,
    -- filter=23 channel=120
    8, 17, -15, 9, 12, -17, -2, -2, -19,
    -- filter=23 channel=121
    8, -4, -10, 0, -9, -9, 3, 0, -1,
    -- filter=23 channel=122
    -35, -10, 2, -26, -7, 0, -29, -5, 2,
    -- filter=23 channel=123
    -3, 0, -7, 3, -5, -17, 1, -2, -14,
    -- filter=23 channel=124
    2, 2, -4, 9, -1, 4, 6, -8, -1,
    -- filter=23 channel=125
    -5, 13, 0, -1, 4, 3, -8, -7, -6,
    -- filter=23 channel=126
    -2, 4, -3, -3, 12, 7, 7, 2, 7,
    -- filter=23 channel=127
    3, -5, -1, -2, 2, 4, 5, -5, -9,
    -- filter=24 channel=0
    -2, 3, 3, 0, 14, 5, 8, 4, 2,
    -- filter=24 channel=1
    4, 0, -11, 8, -3, 4, 13, 13, 5,
    -- filter=24 channel=2
    0, 5, 0, 0, -3, -6, -4, 0, -2,
    -- filter=24 channel=3
    7, 2, 5, 3, 9, 0, -6, -6, -3,
    -- filter=24 channel=4
    4, -7, 1, 4, 3, 0, -2, 5, 5,
    -- filter=24 channel=5
    -2, 4, 0, 0, 4, 0, 5, 3, 6,
    -- filter=24 channel=6
    1, 0, -6, 5, 3, -5, -1, -5, 3,
    -- filter=24 channel=7
    -7, 1, 0, 2, -1, -2, -4, -5, -4,
    -- filter=24 channel=8
    -2, 2, 3, -5, 0, -2, 0, 0, -3,
    -- filter=24 channel=9
    7, 5, -4, -3, -9, 1, 0, -2, -3,
    -- filter=24 channel=10
    -1, -5, -2, 7, -1, -2, 5, 0, -10,
    -- filter=24 channel=11
    -8, 0, 6, -9, -8, 3, 4, -1, 0,
    -- filter=24 channel=12
    -7, -7, 4, 8, -8, -2, 8, 1, -8,
    -- filter=24 channel=13
    0, 4, 4, 4, -11, -3, 14, -7, -2,
    -- filter=24 channel=14
    -4, 5, -1, -3, 2, -4, -4, -3, -2,
    -- filter=24 channel=15
    -3, -7, 0, -2, -3, -8, 10, 0, -9,
    -- filter=24 channel=16
    1, 7, 1, 1, -1, 5, -2, -7, 7,
    -- filter=24 channel=17
    -1, 0, -6, 0, -4, -3, 0, 0, 4,
    -- filter=24 channel=18
    7, -10, -3, 6, -14, -4, 14, 0, -7,
    -- filter=24 channel=19
    0, -6, 0, 5, -5, -1, 0, 1, -3,
    -- filter=24 channel=20
    -1, -1, -1, -1, -3, 7, 2, -3, 0,
    -- filter=24 channel=21
    0, -2, -2, -1, -6, -6, 4, -10, 1,
    -- filter=24 channel=22
    4, 1, -6, 4, 1, -5, 5, -3, 6,
    -- filter=24 channel=23
    4, -7, 0, -16, -1, -1, -2, -14, -3,
    -- filter=24 channel=24
    -7, -5, 5, 0, 6, -1, -2, -6, -1,
    -- filter=24 channel=25
    8, 5, -3, 0, -10, -4, 6, -9, 2,
    -- filter=24 channel=26
    -7, 6, -5, -7, -1, 8, -4, -1, 2,
    -- filter=24 channel=27
    0, -3, 6, -2, -16, 4, 5, -16, -3,
    -- filter=24 channel=28
    2, -3, -5, -2, -4, -1, 1, -7, 2,
    -- filter=24 channel=29
    -10, 3, 9, 0, -8, -6, 4, -6, 4,
    -- filter=24 channel=30
    5, 0, 1, -4, -1, 6, 3, -7, 1,
    -- filter=24 channel=31
    8, 2, 4, -3, -14, -5, -1, -11, -7,
    -- filter=24 channel=32
    -5, 3, 3, -1, -3, 1, 5, -12, -5,
    -- filter=24 channel=33
    9, 7, 3, -3, -11, -5, 5, -1, 0,
    -- filter=24 channel=34
    -5, -4, -4, -7, 5, 1, -2, 0, -7,
    -- filter=24 channel=35
    0, 2, 6, -7, 1, -5, -1, 1, -1,
    -- filter=24 channel=36
    -4, -7, -1, -3, -1, -6, -6, -5, 4,
    -- filter=24 channel=37
    3, 0, 1, -2, 11, -2, 7, -1, 3,
    -- filter=24 channel=38
    0, 1, -1, 1, 0, 1, 0, -2, -8,
    -- filter=24 channel=39
    2, 4, -1, -1, 3, 0, 4, 4, -4,
    -- filter=24 channel=40
    -1, -6, 4, -4, -5, 0, 0, 0, -2,
    -- filter=24 channel=41
    13, -5, 1, 17, 0, -7, 24, 7, -16,
    -- filter=24 channel=42
    2, -3, -4, 4, -4, -3, 6, -1, -3,
    -- filter=24 channel=43
    -2, 6, 1, 5, 6, -5, 5, 5, -2,
    -- filter=24 channel=44
    9, 2, -4, 3, 4, 2, 0, -6, 8,
    -- filter=24 channel=45
    3, 0, 0, -6, 3, 6, -5, 3, 0,
    -- filter=24 channel=46
    1, 0, 3, -4, 0, -7, 0, 0, -4,
    -- filter=24 channel=47
    2, 5, -3, 3, -4, -1, 5, -6, 3,
    -- filter=24 channel=48
    4, -4, -4, 9, -6, -8, 10, 3, 2,
    -- filter=24 channel=49
    -4, -9, -2, -1, -2, -8, -1, 2, -8,
    -- filter=24 channel=50
    -2, -4, 9, -7, 0, 0, -1, -9, -2,
    -- filter=24 channel=51
    -1, 5, 0, 7, 3, -3, -3, 3, 7,
    -- filter=24 channel=52
    -2, -4, 7, -4, -5, 4, -3, 2, -4,
    -- filter=24 channel=53
    -4, -5, 1, -3, 2, 7, -6, -2, 3,
    -- filter=24 channel=54
    -7, 6, 6, -6, 4, 4, 6, -7, -2,
    -- filter=24 channel=55
    6, 1, 4, -7, -10, -4, -1, -13, -8,
    -- filter=24 channel=56
    0, 5, 3, 0, -6, -7, -4, 0, -6,
    -- filter=24 channel=57
    -2, -6, 0, 0, 6, 3, 3, -2, -2,
    -- filter=24 channel=58
    2, 0, 0, 0, 0, 5, -2, -3, 5,
    -- filter=24 channel=59
    6, 3, 0, 12, -11, 1, 13, -5, 1,
    -- filter=24 channel=60
    -7, 3, -4, -5, -3, -5, 6, 7, -6,
    -- filter=24 channel=61
    0, 0, 4, -1, -3, 4, 1, -4, -7,
    -- filter=24 channel=62
    -3, 6, 1, -2, 6, 2, -2, -7, 3,
    -- filter=24 channel=63
    -1, 1, 0, -7, 0, 4, 2, -2, 1,
    -- filter=24 channel=64
    -6, -4, 8, -3, -7, 7, 2, 1, 5,
    -- filter=24 channel=65
    7, 5, -6, -4, -5, -5, -3, 0, 2,
    -- filter=24 channel=66
    3, 2, 2, 1, -1, -1, 7, -1, -2,
    -- filter=24 channel=67
    -2, 5, 0, -4, 6, -4, 0, 0, -3,
    -- filter=24 channel=68
    1, 0, -2, 7, 5, 4, -5, 0, 0,
    -- filter=24 channel=69
    4, 5, 6, 0, 6, -6, 5, 4, -4,
    -- filter=24 channel=70
    4, 0, -4, -3, -6, 2, -5, -8, 3,
    -- filter=24 channel=71
    -3, 10, 1, -3, 9, 3, 0, -7, -5,
    -- filter=24 channel=72
    8, 0, 8, -4, -12, -2, 7, -6, -10,
    -- filter=24 channel=73
    -5, -6, -3, -3, -1, -5, 2, -6, 3,
    -- filter=24 channel=74
    -9, -5, -1, -14, -1, 0, -10, -6, -2,
    -- filter=24 channel=75
    10, 3, -4, 6, 4, 1, 10, 2, 0,
    -- filter=24 channel=76
    0, -8, 8, -4, -8, -7, 0, -1, -6,
    -- filter=24 channel=77
    0, -1, 1, 4, 2, -7, -5, 0, 4,
    -- filter=24 channel=78
    4, 0, -3, 4, 0, 5, -8, -8, -3,
    -- filter=24 channel=79
    2, 3, -3, 11, -3, -3, 9, -7, -11,
    -- filter=24 channel=80
    10, 3, -1, 1, -16, -8, 9, -15, -7,
    -- filter=24 channel=81
    0, -5, 7, 1, 0, 5, -4, 0, -3,
    -- filter=24 channel=82
    -5, -2, 6, 0, 1, -3, 0, 3, 5,
    -- filter=24 channel=83
    -2, -8, 1, -3, 0, -6, 0, 6, -3,
    -- filter=24 channel=84
    -4, -10, 4, -4, -10, 2, 4, -6, -8,
    -- filter=24 channel=85
    4, -7, 5, 2, 2, 0, -1, 5, 5,
    -- filter=24 channel=86
    -4, 1, -5, 0, 0, -5, 1, 3, -4,
    -- filter=24 channel=87
    -8, -6, -3, -4, 0, 4, 5, 3, -3,
    -- filter=24 channel=88
    -1, -4, 5, -4, -7, -4, -8, 2, 2,
    -- filter=24 channel=89
    6, 3, 4, 6, -10, -3, 4, -14, -9,
    -- filter=24 channel=90
    4, -6, 8, -5, 1, 0, -1, 0, -6,
    -- filter=24 channel=91
    -6, 3, -2, 0, -8, -8, 9, -1, -6,
    -- filter=24 channel=92
    -7, 1, 5, 4, 2, -6, 2, 0, -6,
    -- filter=24 channel=93
    -3, -3, -8, 4, -6, 2, 6, 0, 4,
    -- filter=24 channel=94
    -3, -1, 3, -2, -6, 2, 1, 0, 4,
    -- filter=24 channel=95
    -6, 0, 0, 4, -5, 5, -7, -6, -6,
    -- filter=24 channel=96
    -3, 0, 5, -2, 0, 2, 2, -5, -5,
    -- filter=24 channel=97
    0, 1, 10, 3, 0, 8, 1, 1, 2,
    -- filter=24 channel=98
    6, 1, 4, 9, -6, -4, 11, -12, -6,
    -- filter=24 channel=99
    0, -6, 4, -11, -13, 3, 0, -10, 1,
    -- filter=24 channel=100
    -5, 1, 3, -4, 5, 3, -2, -5, -9,
    -- filter=24 channel=101
    4, 2, 2, -5, 1, -7, 3, 2, 1,
    -- filter=24 channel=102
    -1, -7, -6, 6, 3, -4, -2, 0, -6,
    -- filter=24 channel=103
    6, 10, -2, 0, -2, 8, 2, -13, 5,
    -- filter=24 channel=104
    -2, 3, 1, -2, -12, 2, 1, -10, -9,
    -- filter=24 channel=105
    1, -1, -2, 1, 5, 7, 0, -2, 4,
    -- filter=24 channel=106
    4, -1, -3, -4, 2, -7, 0, -1, -5,
    -- filter=24 channel=107
    -8, 3, 4, -11, 4, 0, 4, 1, 6,
    -- filter=24 channel=108
    0, -2, -6, 1, 3, -4, 11, -2, -3,
    -- filter=24 channel=109
    5, -4, 2, 0, -3, -10, 7, -13, -1,
    -- filter=24 channel=110
    -6, 1, 1, -8, 1, -5, -3, -1, 0,
    -- filter=24 channel=111
    -4, 0, 3, -2, -4, 0, -2, 0, -1,
    -- filter=24 channel=112
    -5, -7, 2, -11, -7, -2, -8, -7, -1,
    -- filter=24 channel=113
    6, 2, -4, -1, 4, -6, 0, 0, -8,
    -- filter=24 channel=114
    2, -8, 0, 2, -7, -6, 12, -2, 1,
    -- filter=24 channel=115
    -1, -6, -6, -7, -6, 3, 1, 4, -5,
    -- filter=24 channel=116
    0, -3, 7, -4, -12, 3, 14, 1, -1,
    -- filter=24 channel=117
    4, -6, 5, -2, 0, -5, -2, 0, 0,
    -- filter=24 channel=118
    -5, -5, 3, 0, 0, 4, -2, 7, -1,
    -- filter=24 channel=119
    5, -7, 7, -6, 6, -6, -8, 3, -10,
    -- filter=24 channel=120
    2, -12, 6, -5, -7, 4, 0, -9, 3,
    -- filter=24 channel=121
    -4, 6, -7, 1, -3, 2, 4, -10, 3,
    -- filter=24 channel=122
    8, 12, 1, 4, -6, 0, -5, -12, 5,
    -- filter=24 channel=123
    -7, -7, 4, -8, -4, -7, 0, -2, 2,
    -- filter=24 channel=124
    -6, -2, 0, -8, 2, 7, -5, -2, 2,
    -- filter=24 channel=125
    5, 0, -5, -8, -3, -5, 9, -11, -9,
    -- filter=24 channel=126
    0, 9, 3, 11, -2, 2, 8, 3, 0,
    -- filter=24 channel=127
    -2, 2, 1, 6, 5, -4, 5, 2, -2,
    -- filter=25 channel=0
    7, 12, 1, 16, 22, 0, 0, -1, -9,
    -- filter=25 channel=1
    -10, 6, 0, 10, 13, 2, -12, -9, -21,
    -- filter=25 channel=2
    3, -3, 4, -7, -8, 6, 3, -4, 1,
    -- filter=25 channel=3
    13, 8, -9, 15, 6, 2, 12, 1, 0,
    -- filter=25 channel=4
    6, 2, 5, 3, 3, -4, -10, -1, -6,
    -- filter=25 channel=5
    3, 10, -4, 10, 20, 9, 3, 8, 0,
    -- filter=25 channel=6
    0, -1, 0, -7, -6, 0, 3, -3, 0,
    -- filter=25 channel=7
    3, -4, 3, 3, 2, -7, 0, 3, -5,
    -- filter=25 channel=8
    -4, -9, 3, -7, -8, 0, -8, -6, 5,
    -- filter=25 channel=9
    1, 1, 7, -3, 1, 3, -3, -3, -5,
    -- filter=25 channel=10
    2, 13, -1, -2, -2, 2, -3, -2, 9,
    -- filter=25 channel=11
    7, 3, 3, -10, -9, 6, -5, -1, 5,
    -- filter=25 channel=12
    -2, 0, -8, -6, -7, -4, 4, -6, 0,
    -- filter=25 channel=13
    17, 10, 1, 0, -6, -2, -13, -8, 2,
    -- filter=25 channel=14
    7, -6, 0, -4, -1, -3, -1, 4, 2,
    -- filter=25 channel=15
    25, 13, -9, 1, -8, 3, -16, -3, 4,
    -- filter=25 channel=16
    -8, 0, -7, -5, 3, -1, -1, 4, -11,
    -- filter=25 channel=17
    0, -4, 0, 1, 2, -6, 5, -6, 5,
    -- filter=25 channel=18
    31, 15, -7, -6, -8, 0, -15, -22, -5,
    -- filter=25 channel=19
    -3, -3, 7, 0, 2, -5, 6, 3, 5,
    -- filter=25 channel=20
    19, 9, -3, -3, -2, 1, 0, 3, 16,
    -- filter=25 channel=21
    -11, -3, 2, 6, 8, 0, 9, -3, 2,
    -- filter=25 channel=22
    0, 9, 0, 7, 1, -1, -4, -4, 1,
    -- filter=25 channel=23
    24, 4, -6, -3, -20, 8, -15, 7, 13,
    -- filter=25 channel=24
    3, 1, 5, -7, -6, 7, 0, 7, -6,
    -- filter=25 channel=25
    15, 6, -8, -5, -5, 4, -17, -13, -1,
    -- filter=25 channel=26
    -3, -3, -2, -7, 11, 3, 2, 0, -5,
    -- filter=25 channel=27
    22, 10, -5, -9, -3, -3, -11, -1, 13,
    -- filter=25 channel=28
    5, -1, 3, -6, 6, 0, 2, -6, -5,
    -- filter=25 channel=29
    24, 10, 2, -3, 0, -3, -4, 3, 3,
    -- filter=25 channel=30
    7, 2, 1, -10, 2, 6, 1, -3, 5,
    -- filter=25 channel=31
    -6, -7, 0, -1, -9, 4, 0, 1, 9,
    -- filter=25 channel=32
    28, 8, -8, -5, -14, 1, -19, -7, 0,
    -- filter=25 channel=33
    21, 13, -3, 0, 2, -4, -13, -3, 5,
    -- filter=25 channel=34
    0, -5, 1, -8, -2, -4, 0, -3, -3,
    -- filter=25 channel=35
    -3, 2, 0, 3, 0, 1, 2, -4, 2,
    -- filter=25 channel=36
    -12, -5, 3, -9, -4, 3, -8, -1, -3,
    -- filter=25 channel=37
    -9, 0, 7, 2, 11, -3, -2, 2, -13,
    -- filter=25 channel=38
    14, 7, 1, 1, -1, 2, 5, 7, 6,
    -- filter=25 channel=39
    11, 7, -2, -8, -5, 7, -2, 3, 9,
    -- filter=25 channel=40
    12, 3, -2, -3, -9, 0, -7, 2, 3,
    -- filter=25 channel=41
    -2, 12, -1, -4, -10, -13, -3, -23, -7,
    -- filter=25 channel=42
    -7, 5, 8, -3, 3, 6, -9, 6, 1,
    -- filter=25 channel=43
    13, 13, 1, 12, 3, 0, 2, -8, -2,
    -- filter=25 channel=44
    0, 0, -6, 4, 9, 0, -5, 3, 0,
    -- filter=25 channel=45
    -7, 2, 0, 6, 9, -4, 6, 6, 2,
    -- filter=25 channel=46
    -5, 9, 6, -3, -2, 1, 2, 4, 1,
    -- filter=25 channel=47
    -16, 0, 9, 0, 11, 4, -1, 0, -7,
    -- filter=25 channel=48
    -1, 4, 4, -8, 2, 0, -13, -9, -2,
    -- filter=25 channel=49
    6, 4, 1, -8, -6, 2, -18, -2, 1,
    -- filter=25 channel=50
    13, -4, -1, 0, 2, 6, 1, 0, 5,
    -- filter=25 channel=51
    1, -4, 3, -3, 0, 6, -7, -2, 3,
    -- filter=25 channel=52
    6, 1, 1, -1, -11, -2, 3, 0, 0,
    -- filter=25 channel=53
    15, 1, 5, 1, 2, -4, -9, -4, 4,
    -- filter=25 channel=54
    2, -4, -5, 0, -2, 3, 0, -5, -5,
    -- filter=25 channel=55
    26, 9, -3, -7, -17, -6, -19, -5, 8,
    -- filter=25 channel=56
    5, 3, 6, 3, -5, 0, -5, -6, -6,
    -- filter=25 channel=57
    4, -6, -3, -9, -3, -4, -4, -7, 1,
    -- filter=25 channel=58
    -10, 2, -3, 5, 10, 9, -6, 11, 0,
    -- filter=25 channel=59
    11, 9, 0, -1, -1, 5, -7, -9, 4,
    -- filter=25 channel=60
    -5, 0, 1, 0, 1, -3, 4, 0, -2,
    -- filter=25 channel=61
    -4, 2, -2, -5, -5, -9, 1, 1, 6,
    -- filter=25 channel=62
    0, -1, 7, -2, -2, -6, 6, 4, -3,
    -- filter=25 channel=63
    2, 7, 6, 2, 8, 1, 2, 1, -7,
    -- filter=25 channel=64
    -1, -4, 6, -8, 3, 3, 1, 4, 2,
    -- filter=25 channel=65
    0, -2, 0, -4, -2, 3, 2, 6, 4,
    -- filter=25 channel=66
    7, -2, -8, -5, -10, -9, -6, -15, -9,
    -- filter=25 channel=67
    -6, 0, -1, -3, -5, 0, 3, -7, 2,
    -- filter=25 channel=68
    1, -6, -5, -7, -6, 7, -9, -3, -6,
    -- filter=25 channel=69
    4, -5, -3, 7, -2, -3, -5, 4, -4,
    -- filter=25 channel=70
    13, 5, -1, -7, -4, -1, -12, -9, 0,
    -- filter=25 channel=71
    7, 6, -8, 0, -4, 4, 10, 0, -5,
    -- filter=25 channel=72
    -1, 1, 6, 0, 2, 0, -9, -2, 2,
    -- filter=25 channel=73
    7, -6, 3, -3, -8, 1, -6, -2, -1,
    -- filter=25 channel=74
    0, -15, -7, -10, -8, 5, -2, 2, 11,
    -- filter=25 channel=75
    9, 21, -10, 9, 16, -4, -2, -4, -18,
    -- filter=25 channel=76
    16, 1, -8, -8, -18, 0, -7, -9, 5,
    -- filter=25 channel=77
    -7, -2, 0, -5, 3, -6, 7, 0, 5,
    -- filter=25 channel=78
    -3, 4, -5, -6, 4, 0, -9, -5, -5,
    -- filter=25 channel=79
    38, 10, -17, 3, -15, -9, -12, -7, -4,
    -- filter=25 channel=80
    -4, 2, -2, 1, -4, 4, -2, -1, 4,
    -- filter=25 channel=81
    0, -5, 2, 3, -2, -2, 5, 3, -4,
    -- filter=25 channel=82
    -3, -2, 0, 2, 0, 7, 0, 1, 7,
    -- filter=25 channel=83
    -4, 3, 4, 0, 1, 6, -7, 4, -2,
    -- filter=25 channel=84
    16, 1, 1, -15, -9, -2, -13, -6, 0,
    -- filter=25 channel=85
    -1, 0, 5, -5, 0, 4, 0, 0, 0,
    -- filter=25 channel=86
    -4, -3, -3, 2, 3, 5, -4, -5, 1,
    -- filter=25 channel=87
    13, 3, 4, -2, -11, -5, -3, -5, -6,
    -- filter=25 channel=88
    -3, -14, 1, 0, -3, -2, -2, -2, -2,
    -- filter=25 channel=89
    26, 11, -8, -6, -11, 7, -9, -7, 9,
    -- filter=25 channel=90
    0, -11, 4, -3, -1, 1, 4, 0, 2,
    -- filter=25 channel=91
    16, -3, 0, -12, -4, -1, -21, -1, 0,
    -- filter=25 channel=92
    6, -6, -8, -4, 6, 3, -1, -6, -2,
    -- filter=25 channel=93
    -4, 0, 2, -2, 11, -4, -10, -7, -2,
    -- filter=25 channel=94
    -3, 3, 5, 0, -4, -4, 4, 5, 0,
    -- filter=25 channel=95
    1, -5, -3, -2, 2, -2, 4, 3, 0,
    -- filter=25 channel=96
    -1, 4, 0, -1, 0, 0, 1, -8, 6,
    -- filter=25 channel=97
    6, 8, 3, 2, 5, 1, 0, 2, -6,
    -- filter=25 channel=98
    24, 12, -13, 0, 2, -2, -14, 4, 6,
    -- filter=25 channel=99
    2, -6, 0, -4, -15, 4, -11, 6, 13,
    -- filter=25 channel=100
    -1, 5, 2, -7, -5, -5, 1, 1, 2,
    -- filter=25 channel=101
    -2, 4, 6, 1, -4, 4, 3, -5, 0,
    -- filter=25 channel=102
    -3, -3, -2, 1, -6, -4, 2, 7, -4,
    -- filter=25 channel=103
    -4, 7, 5, 14, 10, 5, 0, 4, -8,
    -- filter=25 channel=104
    -5, -8, 1, -6, -7, 1, -7, 5, 0,
    -- filter=25 channel=105
    18, 7, 0, 3, -4, -3, 0, -9, 0,
    -- filter=25 channel=106
    0, 0, -7, 3, -7, 0, 1, -7, -4,
    -- filter=25 channel=107
    9, -2, 1, 0, -11, 2, -15, -1, 4,
    -- filter=25 channel=108
    -3, 4, -5, 5, 4, 0, -6, -2, -10,
    -- filter=25 channel=109
    26, -1, 0, -10, -13, -3, -17, -2, 6,
    -- filter=25 channel=110
    5, -4, 6, -8, 0, 6, 5, 1, 2,
    -- filter=25 channel=111
    -3, 2, -6, -2, -3, -2, 1, -6, -2,
    -- filter=25 channel=112
    2, -5, 1, -6, 4, 0, 0, 5, 1,
    -- filter=25 channel=113
    6, 11, -2, 0, -2, 3, 4, -2, -4,
    -- filter=25 channel=114
    29, 11, -2, 0, 2, -7, -25, -11, 3,
    -- filter=25 channel=115
    0, 5, -2, -1, 0, 2, 1, -4, -3,
    -- filter=25 channel=116
    3, -3, 1, -12, -12, 4, -13, -9, 0,
    -- filter=25 channel=117
    0, 2, 1, -3, 1, -1, -8, -5, 1,
    -- filter=25 channel=118
    4, 5, 2, 5, -1, -7, -1, -4, 0,
    -- filter=25 channel=119
    5, -8, 3, -7, 1, -6, -3, -7, -1,
    -- filter=25 channel=120
    21, -13, -6, -17, -6, 12, -9, 7, 17,
    -- filter=25 channel=121
    11, 3, 5, 0, 1, -4, -3, -2, -3,
    -- filter=25 channel=122
    -14, -9, 12, -8, 12, -2, 4, -2, 1,
    -- filter=25 channel=123
    -4, 0, 0, 6, 4, 1, -7, -2, 2,
    -- filter=25 channel=124
    3, 3, -4, 0, -2, 6, 3, 2, 7,
    -- filter=25 channel=125
    7, -6, 2, -11, -1, 5, -5, 3, 6,
    -- filter=25 channel=126
    19, 21, -2, 4, 4, 0, 3, -8, -9,
    -- filter=25 channel=127
    -1, -3, 3, -8, 0, -1, -7, -5, -5,
    -- filter=26 channel=0
    3, 8, -21, 24, 31, -11, 7, 27, -18,
    -- filter=26 channel=1
    -6, 16, -9, 13, 39, 0, 6, 20, 1,
    -- filter=26 channel=2
    -2, 3, -7, 2, 0, -2, -1, -4, -6,
    -- filter=26 channel=3
    3, 7, 1, 1, 4, 1, 7, 2, 7,
    -- filter=26 channel=4
    -6, 7, -3, 4, 9, 7, 0, 12, 13,
    -- filter=26 channel=5
    -1, 10, -11, -1, 8, -12, -3, 10, -17,
    -- filter=26 channel=6
    -6, 0, -1, 12, 7, -4, -6, 5, -3,
    -- filter=26 channel=7
    -7, 6, -1, -7, -5, 0, -6, 0, -2,
    -- filter=26 channel=8
    -4, 6, 5, -2, 0, 2, 5, 2, 4,
    -- filter=26 channel=9
    -9, -5, -8, -10, -3, -10, -3, -3, 0,
    -- filter=26 channel=10
    -8, -5, 3, -16, -15, 2, -8, -19, -1,
    -- filter=26 channel=11
    -3, -1, 9, -7, -9, 7, -9, -16, 7,
    -- filter=26 channel=12
    -1, 1, -2, 6, 0, 3, 0, 5, 6,
    -- filter=26 channel=13
    2, 0, 12, -3, -8, 2, 3, -2, 7,
    -- filter=26 channel=14
    0, -7, -7, -6, 5, 6, -6, -4, -2,
    -- filter=26 channel=15
    -3, 2, -10, 19, 11, 1, 3, -6, -7,
    -- filter=26 channel=16
    -2, 4, 0, -12, -9, 3, -6, -8, -2,
    -- filter=26 channel=17
    3, -3, -1, 0, 1, 3, 4, 0, -5,
    -- filter=26 channel=18
    6, -4, -20, 22, 10, -6, 9, 9, -4,
    -- filter=26 channel=19
    -6, 2, 0, 0, 3, 4, -2, 6, -5,
    -- filter=26 channel=20
    -10, -10, -3, -4, -11, 6, -10, -21, 2,
    -- filter=26 channel=21
    0, -2, 17, -14, -16, 2, -6, -7, 0,
    -- filter=26 channel=22
    7, 6, -3, 7, 9, 0, 13, 11, -9,
    -- filter=26 channel=23
    4, -5, 2, 0, -6, 6, 0, 0, 12,
    -- filter=26 channel=24
    2, 4, 1, 0, -7, -7, -5, -5, -5,
    -- filter=26 channel=25
    -3, -1, -2, -6, 7, 4, 2, -2, -2,
    -- filter=26 channel=26
    0, -4, 4, -5, -10, 0, -1, -8, 4,
    -- filter=26 channel=27
    4, 4, -3, 3, 13, -9, 15, 12, 1,
    -- filter=26 channel=28
    -5, -4, -1, 5, -1, 0, -1, 3, 2,
    -- filter=26 channel=29
    -1, -19, 1, 0, -15, -4, -14, -11, 0,
    -- filter=26 channel=30
    -7, 10, -5, 5, 5, -3, 4, 14, -7,
    -- filter=26 channel=31
    -9, 4, 27, -36, -29, 16, -13, -16, 12,
    -- filter=26 channel=32
    6, -3, -14, 6, 12, -2, 4, 9, -6,
    -- filter=26 channel=33
    4, 8, -1, 7, 3, -6, 4, 9, -7,
    -- filter=26 channel=34
    -3, 0, 8, 9, 12, 2, 0, -1, -8,
    -- filter=26 channel=35
    -2, 0, 6, 3, 3, -3, 3, 5, 6,
    -- filter=26 channel=36
    2, -11, 10, -20, -9, 2, 0, -9, 12,
    -- filter=26 channel=37
    -8, 22, -7, 10, 23, -2, -2, 28, 4,
    -- filter=26 channel=38
    6, -1, -1, -1, 1, -4, 5, -3, 1,
    -- filter=26 channel=39
    -2, -2, 5, -6, -11, 6, -1, -6, -3,
    -- filter=26 channel=40
    5, 2, 9, 6, 1, 9, 2, 6, -1,
    -- filter=26 channel=41
    -6, -15, -10, -6, -3, 6, -3, -7, -3,
    -- filter=26 channel=42
    -9, 3, 0, 4, 1, 1, 0, 8, -8,
    -- filter=26 channel=43
    6, 0, 0, 15, 13, -3, 2, 9, -4,
    -- filter=26 channel=44
    -7, 11, 0, -1, 11, -4, -3, 13, 2,
    -- filter=26 channel=45
    1, 0, -2, 7, 13, 0, 13, 5, -2,
    -- filter=26 channel=46
    -2, 0, -8, 2, -1, 0, -4, -2, 6,
    -- filter=26 channel=47
    5, 4, 10, -15, -14, -4, 0, -5, 1,
    -- filter=26 channel=48
    -8, 0, 9, -7, -12, -7, -5, 2, 3,
    -- filter=26 channel=49
    5, 0, -10, 10, 8, 2, 1, -4, 3,
    -- filter=26 channel=50
    6, 2, 8, -4, 8, 4, 0, -2, -1,
    -- filter=26 channel=51
    -4, -1, -2, 6, -2, 5, -5, -5, 2,
    -- filter=26 channel=52
    3, 3, -4, 0, -3, 5, 4, 3, 9,
    -- filter=26 channel=53
    -8, 0, 6, -1, -5, 4, -3, -4, 0,
    -- filter=26 channel=54
    7, 6, -5, -2, 4, -2, -3, 3, 5,
    -- filter=26 channel=55
    3, -15, -1, 2, -13, 4, -11, -14, 5,
    -- filter=26 channel=56
    0, -5, 3, 8, 6, -4, 5, -5, 4,
    -- filter=26 channel=57
    4, 3, 5, 0, -4, -3, -6, -8, 7,
    -- filter=26 channel=58
    -2, -4, -10, 0, 5, -4, 3, 6, -8,
    -- filter=26 channel=59
    6, -6, 8, -11, -6, 3, 4, -9, -5,
    -- filter=26 channel=60
    -4, 0, -4, 5, -1, -4, -6, 1, -4,
    -- filter=26 channel=61
    -7, 5, 8, -7, -8, 7, -1, 0, 5,
    -- filter=26 channel=62
    0, -7, 4, 6, 5, 0, 6, -7, 0,
    -- filter=26 channel=63
    -8, -2, -2, -10, -12, -5, -11, -5, -1,
    -- filter=26 channel=64
    5, 0, 7, -3, -11, 10, -5, -8, 2,
    -- filter=26 channel=65
    2, 5, -3, 1, -1, -3, 2, -5, -5,
    -- filter=26 channel=66
    -2, 0, 0, -9, 4, 2, 5, -10, -1,
    -- filter=26 channel=67
    0, 0, -2, 2, -5, -4, -6, -2, 0,
    -- filter=26 channel=68
    -5, 0, 10, 5, 5, 7, -2, -4, 2,
    -- filter=26 channel=69
    0, -4, -5, -3, -5, 6, 1, 6, 5,
    -- filter=26 channel=70
    -2, 9, 1, 9, 19, 9, 5, 15, 0,
    -- filter=26 channel=71
    8, -5, 0, -6, -7, -5, 2, 1, 9,
    -- filter=26 channel=72
    0, -1, 18, -16, -21, 6, -17, -22, 11,
    -- filter=26 channel=73
    -6, 3, -5, -5, 7, 3, -2, -2, -6,
    -- filter=26 channel=74
    6, -2, 4, -9, 10, 1, 0, 4, -2,
    -- filter=26 channel=75
    -4, 13, -11, 1, 24, -6, 3, 18, -2,
    -- filter=26 channel=76
    -2, -10, 3, 1, -8, -5, -3, -19, 1,
    -- filter=26 channel=77
    -7, -2, 0, -1, -3, 0, -6, -5, 1,
    -- filter=26 channel=78
    -5, 5, 0, -7, -1, -10, -12, -7, -8,
    -- filter=26 channel=79
    11, -4, -17, 21, 13, -1, 16, 13, 1,
    -- filter=26 channel=80
    -11, 1, 12, -32, -17, 0, -8, -19, 0,
    -- filter=26 channel=81
    3, 4, 0, 6, 5, -2, 1, -7, 6,
    -- filter=26 channel=82
    2, 1, 0, 3, 4, -6, -1, 2, 3,
    -- filter=26 channel=83
    -3, 4, 3, -6, -3, -2, -4, 0, -6,
    -- filter=26 channel=84
    -6, -6, -8, 5, 7, -9, 5, -2, -3,
    -- filter=26 channel=85
    1, 6, 5, -3, -6, -6, -6, -2, -6,
    -- filter=26 channel=86
    0, 2, 0, 4, 9, 3, 0, 0, 0,
    -- filter=26 channel=87
    -5, -10, -6, 0, -5, 5, 0, -4, 7,
    -- filter=26 channel=88
    1, -8, 9, -17, -18, 7, -10, -14, 7,
    -- filter=26 channel=89
    1, -15, 7, -12, -18, 0, -9, -17, 8,
    -- filter=26 channel=90
    -5, -8, 14, -5, -6, 9, -2, -10, 9,
    -- filter=26 channel=91
    4, 1, -2, 4, 0, 5, 10, 2, -7,
    -- filter=26 channel=92
    0, 7, -2, 8, -2, 1, -6, 6, 5,
    -- filter=26 channel=93
    -8, 11, 1, -14, -1, 1, -12, 8, -2,
    -- filter=26 channel=94
    4, 1, 2, 3, 5, 7, -3, 5, 2,
    -- filter=26 channel=95
    -2, 0, -5, -4, 3, 0, -1, -7, 1,
    -- filter=26 channel=96
    -2, 6, 0, 3, 0, 7, -4, 5, -4,
    -- filter=26 channel=97
    -4, 1, 4, -1, 5, -3, -3, 3, 0,
    -- filter=26 channel=98
    -3, 3, 4, -17, -6, -3, -8, -8, -9,
    -- filter=26 channel=99
    -13, -7, 11, -27, -25, 8, -18, -21, 13,
    -- filter=26 channel=100
    -9, 4, -7, -6, 0, -4, -4, 4, 2,
    -- filter=26 channel=101
    -2, 5, -4, 4, -4, 3, 0, 7, 6,
    -- filter=26 channel=102
    5, 1, -6, -1, 7, -1, 0, -1, -2,
    -- filter=26 channel=103
    -3, 7, 12, -11, -4, 0, -15, -6, 2,
    -- filter=26 channel=104
    -3, 6, 5, -17, -26, 4, -12, -14, -1,
    -- filter=26 channel=105
    -8, -5, -10, -3, -2, 4, -9, -10, -7,
    -- filter=26 channel=106
    3, -6, 4, 6, 0, 9, -9, -8, 7,
    -- filter=26 channel=107
    12, -2, -15, 10, 8, -6, 10, 7, -10,
    -- filter=26 channel=108
    2, -8, -3, -2, 0, -2, -3, 1, -3,
    -- filter=26 channel=109
    6, -7, -17, -5, -5, -17, 2, 0, -14,
    -- filter=26 channel=110
    -2, -8, 12, -18, -19, -1, -14, -17, 10,
    -- filter=26 channel=111
    -5, 2, 0, 4, 3, 3, -1, 3, -4,
    -- filter=26 channel=112
    -6, 11, -13, 3, 1, 0, -1, 0, -6,
    -- filter=26 channel=113
    1, 8, 11, 0, 0, 1, -3, -8, 3,
    -- filter=26 channel=114
    -4, -4, -28, 34, 41, -27, 19, 27, -25,
    -- filter=26 channel=115
    1, -7, -6, -2, 5, -1, -3, 5, 5,
    -- filter=26 channel=116
    -3, -4, 3, -11, -8, 1, -13, -19, 0,
    -- filter=26 channel=117
    0, -2, 4, -2, 2, 7, -1, 0, 11,
    -- filter=26 channel=118
    -3, -7, -1, -5, 0, -2, -3, -5, -1,
    -- filter=26 channel=119
    0, -6, 3, -2, 13, 0, -2, -1, -5,
    -- filter=26 channel=120
    -1, -8, -12, 7, -6, -2, 5, -7, -5,
    -- filter=26 channel=121
    0, -9, 7, 0, -8, 7, -2, -7, 6,
    -- filter=26 channel=122
    -1, 5, 24, -32, -17, 11, -4, -19, 21,
    -- filter=26 channel=123
    6, -2, -3, 0, 8, 7, -3, -3, 2,
    -- filter=26 channel=124
    0, -2, 4, 1, 1, 5, -8, -8, 1,
    -- filter=26 channel=125
    5, 5, 8, -23, -12, -4, -3, -13, 6,
    -- filter=26 channel=126
    -2, -13, -9, 0, -9, -6, -1, -5, 3,
    -- filter=26 channel=127
    0, -7, -4, 1, 0, 0, -6, -2, -2,
    -- filter=27 channel=0
    3, -5, -2, 7, -6, -7, 8, 4, 9,
    -- filter=27 channel=1
    7, 4, -4, 10, 1, -3, 10, 9, 13,
    -- filter=27 channel=2
    0, -7, 5, 4, -3, 6, 2, 11, 1,
    -- filter=27 channel=3
    -8, 0, -6, -8, -2, 0, 7, 11, 9,
    -- filter=27 channel=4
    7, 0, 4, -6, 7, 13, 1, 19, 27,
    -- filter=27 channel=5
    -6, -8, -1, -1, -5, -2, 5, -6, 7,
    -- filter=27 channel=6
    7, 6, 7, 9, 3, -2, 5, 9, 0,
    -- filter=27 channel=7
    5, -5, 3, 3, 5, -7, 6, -5, 1,
    -- filter=27 channel=8
    0, 1, 2, 6, -5, 0, 6, 5, 7,
    -- filter=27 channel=9
    0, -11, -4, 0, -3, -10, -8, 6, -2,
    -- filter=27 channel=10
    -6, -8, -8, -8, -2, -3, -5, -6, -4,
    -- filter=27 channel=11
    6, 5, 0, 7, 8, -3, 9, 0, 1,
    -- filter=27 channel=12
    9, 8, -3, 4, 2, 7, 3, -3, 2,
    -- filter=27 channel=13
    -4, 1, -14, 0, 1, 0, -2, 8, 7,
    -- filter=27 channel=14
    -3, 5, 6, 0, 0, -7, -4, -5, -6,
    -- filter=27 channel=15
    -1, -3, -9, 6, -11, -4, 2, 7, -3,
    -- filter=27 channel=16
    8, 2, 8, -3, 3, 3, 5, 6, 3,
    -- filter=27 channel=17
    2, 0, 2, -4, 2, -4, 4, 2, -5,
    -- filter=27 channel=18
    3, -1, -16, -1, -10, -8, -2, 5, 9,
    -- filter=27 channel=19
    -4, 8, 0, 5, 4, -2, 5, -6, 4,
    -- filter=27 channel=20
    9, 11, -1, 6, 12, 1, 8, 11, -5,
    -- filter=27 channel=21
    -4, 4, -1, 5, 5, 11, 7, 9, 1,
    -- filter=27 channel=22
    -7, -6, -3, 5, -5, 0, -5, 10, 0,
    -- filter=27 channel=23
    2, -11, -11, -1, -12, -6, -5, 11, -8,
    -- filter=27 channel=24
    3, 6, -3, 5, 0, -5, -4, 6, 0,
    -- filter=27 channel=25
    -4, -16, -16, -11, -11, -5, -3, 7, 6,
    -- filter=27 channel=26
    -3, -3, -1, 8, -2, 6, -3, 0, 2,
    -- filter=27 channel=27
    -15, -22, -23, -11, -20, -6, -6, 0, 13,
    -- filter=27 channel=28
    0, 0, 3, 5, 3, -2, -1, 1, 2,
    -- filter=27 channel=29
    6, 4, -6, 6, 3, -4, 9, -5, 2,
    -- filter=27 channel=30
    -9, -3, -9, -4, -4, 0, 0, 1, 7,
    -- filter=27 channel=31
    -9, -11, -8, -1, -17, -3, -4, 8, -4,
    -- filter=27 channel=32
    3, -17, -7, -1, -11, -13, -5, 3, -3,
    -- filter=27 channel=33
    -12, -12, -18, -1, -15, -1, -4, -3, -5,
    -- filter=27 channel=34
    4, 5, 3, -3, 2, 14, -3, 3, 12,
    -- filter=27 channel=35
    -6, -2, 1, 1, -4, 2, -5, 5, 4,
    -- filter=27 channel=36
    7, 12, 13, 7, 3, 18, 9, 13, 12,
    -- filter=27 channel=37
    8, -4, 6, 0, 2, 1, 6, 16, 10,
    -- filter=27 channel=38
    1, 0, -12, -8, 0, -1, 3, 4, -7,
    -- filter=27 channel=39
    2, 3, 0, 3, 3, -4, 0, -2, 5,
    -- filter=27 channel=40
    6, 13, 7, 9, 8, 8, 12, 4, 1,
    -- filter=27 channel=41
    0, 10, -5, 10, 20, 6, -5, 3, 8,
    -- filter=27 channel=42
    2, 2, -1, 5, -3, -9, 0, -3, 2,
    -- filter=27 channel=43
    -4, 5, -8, 5, -7, -6, 7, -2, 6,
    -- filter=27 channel=44
    1, -15, -5, -12, -14, -1, 1, 0, 4,
    -- filter=27 channel=45
    9, 5, 8, 7, 8, 0, 10, 4, 0,
    -- filter=27 channel=46
    -5, 3, -6, 1, 7, -2, -2, -1, 5,
    -- filter=27 channel=47
    -9, -12, 4, 4, -10, -8, 1, 1, 10,
    -- filter=27 channel=48
    0, -19, -8, -10, -10, -2, -4, 6, 15,
    -- filter=27 channel=49
    0, -11, -8, 6, 4, -6, 7, 12, 8,
    -- filter=27 channel=50
    -11, -6, -7, -6, -5, 1, -9, 0, 0,
    -- filter=27 channel=51
    -4, -3, 0, -3, -3, 4, -5, -5, 1,
    -- filter=27 channel=52
    -1, 6, 10, 7, 6, 9, 10, 7, 10,
    -- filter=27 channel=53
    6, -1, 0, 0, 3, 2, -6, 3, 2,
    -- filter=27 channel=54
    -7, -4, -4, 2, -3, 6, -7, -1, -1,
    -- filter=27 channel=55
    0, -5, -14, -4, -2, -15, 1, 5, 0,
    -- filter=27 channel=56
    0, 2, 10, 3, -2, 2, -4, 0, 8,
    -- filter=27 channel=57
    -2, 5, 2, -6, 0, -2, 3, -1, 0,
    -- filter=27 channel=58
    8, 5, 0, -4, 0, -4, 4, 5, 0,
    -- filter=27 channel=59
    -2, -7, -2, 0, -4, 0, -9, 6, 4,
    -- filter=27 channel=60
    2, 1, -5, 5, -1, 4, -6, 6, 0,
    -- filter=27 channel=61
    3, 0, -2, 0, 6, 6, 3, -2, 0,
    -- filter=27 channel=62
    0, -5, 0, 6, -5, 0, -4, -1, 1,
    -- filter=27 channel=63
    9, -3, 0, 0, 0, 8, -4, 0, 4,
    -- filter=27 channel=64
    6, 11, 4, 5, 11, 1, 9, 0, 5,
    -- filter=27 channel=65
    6, -2, 1, 0, -3, 0, 3, -1, -6,
    -- filter=27 channel=66
    7, -1, -2, 8, 6, 9, 5, -6, -1,
    -- filter=27 channel=67
    3, -2, 4, -3, 7, 2, -6, -3, 0,
    -- filter=27 channel=68
    8, 0, -4, 5, -4, 4, 8, 1, 2,
    -- filter=27 channel=69
    -5, 4, 1, -4, 0, 2, -6, -5, 4,
    -- filter=27 channel=70
    1, -10, -9, -1, -4, -4, 0, 2, 5,
    -- filter=27 channel=71
    -2, 0, -4, -5, -1, 5, 9, 2, 0,
    -- filter=27 channel=72
    -11, -6, -5, 0, -15, -9, -1, 1, 3,
    -- filter=27 channel=73
    -1, -2, -4, -3, 0, -6, -5, 10, 6,
    -- filter=27 channel=74
    -8, -4, 1, -5, -2, 14, -3, 9, 14,
    -- filter=27 channel=75
    0, -2, -8, 5, -12, -10, -1, -1, 0,
    -- filter=27 channel=76
    12, 5, -2, 13, 6, -3, 12, 6, -4,
    -- filter=27 channel=77
    2, 2, 4, 9, 1, 5, 1, 0, 5,
    -- filter=27 channel=78
    -1, 1, 5, 4, 0, 0, -7, -6, 0,
    -- filter=27 channel=79
    -1, -18, -11, -1, -14, -15, 0, 2, 8,
    -- filter=27 channel=80
    -13, -17, -7, -12, -10, -12, -8, 0, -1,
    -- filter=27 channel=81
    -5, 0, -3, -6, -6, 0, -2, -6, 0,
    -- filter=27 channel=82
    -5, 1, 7, 5, -1, 2, 4, 4, -4,
    -- filter=27 channel=83
    -3, 0, -1, -9, 4, 0, 1, 2, 8,
    -- filter=27 channel=84
    3, 1, -8, -5, 6, 0, -3, 12, 3,
    -- filter=27 channel=85
    5, 0, -6, -1, 2, -5, 6, 1, -6,
    -- filter=27 channel=86
    5, -5, 7, 0, 0, 0, 4, 6, 4,
    -- filter=27 channel=87
    5, 0, 2, 1, 10, 12, 10, 4, -3,
    -- filter=27 channel=88
    5, 4, 17, 0, 1, 11, 3, 7, 3,
    -- filter=27 channel=89
    -9, -7, -10, -12, -10, -7, -11, -6, 1,
    -- filter=27 channel=90
    -1, 10, 7, 11, 12, 18, 8, 10, 0,
    -- filter=27 channel=91
    -11, -7, -8, -4, -10, 3, -7, 11, 10,
    -- filter=27 channel=92
    -5, 0, 6, -8, 7, 0, 2, -2, -2,
    -- filter=27 channel=93
    0, -12, -11, 0, -8, -6, 2, 6, 12,
    -- filter=27 channel=94
    -1, -6, 2, -4, 0, -3, 0, 3, -1,
    -- filter=27 channel=95
    1, -2, -4, -5, 4, 2, -6, -4, 4,
    -- filter=27 channel=96
    6, 6, -5, 3, -7, -4, -6, 4, 5,
    -- filter=27 channel=97
    5, 4, 4, -1, 2, -6, -3, -4, 0,
    -- filter=27 channel=98
    -11, -11, -12, -6, -13, -7, -6, -3, 4,
    -- filter=27 channel=99
    -3, -8, -5, -11, -11, -3, 0, 3, -4,
    -- filter=27 channel=100
    5, 0, 0, 2, 8, -1, 1, -3, 6,
    -- filter=27 channel=101
    4, 0, -6, 7, 10, 3, -2, 9, 7,
    -- filter=27 channel=102
    5, -5, -7, 0, 4, -2, -2, 5, 3,
    -- filter=27 channel=103
    4, -4, -9, -8, -13, -9, -3, 5, 0,
    -- filter=27 channel=104
    -11, -13, -1, -1, -2, -1, 2, 4, 7,
    -- filter=27 channel=105
    7, 12, 6, 3, 7, 0, 9, 8, -7,
    -- filter=27 channel=106
    11, 1, 0, 6, 11, 0, 5, 4, -3,
    -- filter=27 channel=107
    6, 8, 6, 16, 12, 0, 4, 10, 1,
    -- filter=27 channel=108
    -2, 7, 4, 1, 2, 4, -2, 2, 2,
    -- filter=27 channel=109
    -5, -17, -19, -3, -14, -1, -11, 3, 5,
    -- filter=27 channel=110
    -7, -9, 2, 4, -12, 0, -5, 5, -6,
    -- filter=27 channel=111
    -5, 3, 9, -1, 5, 4, 0, 3, 3,
    -- filter=27 channel=112
    2, -9, 1, -10, -9, 6, -9, 2, -5,
    -- filter=27 channel=113
    -6, -3, -5, 2, -10, -11, 0, -5, 2,
    -- filter=27 channel=114
    -3, -10, -14, 5, -12, -9, -6, 15, 13,
    -- filter=27 channel=115
    -3, -7, -2, -2, 4, 7, 5, 5, 5,
    -- filter=27 channel=116
    -11, -11, -11, -2, -11, -1, -9, 7, 5,
    -- filter=27 channel=117
    -5, -4, -8, 6, -1, -1, -6, 4, 1,
    -- filter=27 channel=118
    7, -1, -1, 6, 8, 0, -2, 5, 7,
    -- filter=27 channel=119
    -2, 8, 3, 2, 10, 6, -4, 11, 5,
    -- filter=27 channel=120
    -9, -19, -4, -9, -8, -3, -1, 16, 5,
    -- filter=27 channel=121
    -8, 1, -3, 2, -1, 1, -4, -6, 0,
    -- filter=27 channel=122
    -1, 0, 1, 2, -4, 4, 10, 11, 14,
    -- filter=27 channel=123
    0, -1, -4, -4, 8, -4, -5, -3, 7,
    -- filter=27 channel=124
    3, -2, -1, 6, 3, -6, 6, -3, -3,
    -- filter=27 channel=125
    -2, -15, -15, -10, -11, 4, -2, 0, 10,
    -- filter=27 channel=126
    -5, -7, -9, 2, -6, 0, 0, 1, -2,
    -- filter=27 channel=127
    5, -2, -4, -4, 8, 1, 0, -5, 1,
    -- filter=28 channel=0
    6, 11, -6, 0, -2, -4, 3, -4, 6,
    -- filter=28 channel=1
    14, -2, 1, -8, 7, 3, -5, -6, -2,
    -- filter=28 channel=2
    -4, -4, 0, -8, 6, 0, -7, -9, 1,
    -- filter=28 channel=3
    -13, -9, 1, -1, -14, -12, -10, 1, -6,
    -- filter=28 channel=4
    -8, -7, -12, -16, 0, -1, -5, -13, -1,
    -- filter=28 channel=5
    4, -1, 6, 0, -11, -5, 4, -6, 3,
    -- filter=28 channel=6
    -5, 8, 0, 7, 2, 1, -3, 0, 0,
    -- filter=28 channel=7
    3, -1, -1, 7, 5, -3, -2, -7, -5,
    -- filter=28 channel=8
    2, -10, 0, 2, -4, -13, -6, -1, -9,
    -- filter=28 channel=9
    4, 4, -4, 5, 0, 4, -4, -7, 0,
    -- filter=28 channel=10
    0, -4, -7, 2, 2, -11, 7, -3, -3,
    -- filter=28 channel=11
    -1, -2, -1, 8, 17, 2, -10, 13, 9,
    -- filter=28 channel=12
    6, -4, -3, -10, 1, -20, -4, 2, -5,
    -- filter=28 channel=13
    -2, -7, -4, -2, 19, -11, -5, 1, -4,
    -- filter=28 channel=14
    5, 0, -5, -4, 5, -4, 0, 2, 4,
    -- filter=28 channel=15
    -12, -7, -17, 12, 11, -7, -11, 16, -1,
    -- filter=28 channel=16
    5, -9, 3, -2, 0, 2, -5, 0, -3,
    -- filter=28 channel=17
    3, -6, -1, -2, -6, 7, -3, 4, 2,
    -- filter=28 channel=18
    -1, 2, -28, 6, 36, -11, -4, 22, 0,
    -- filter=28 channel=19
    -5, 6, -2, -2, 4, 0, 2, 3, -5,
    -- filter=28 channel=20
    -15, -7, -8, 8, 21, -8, -2, 14, 2,
    -- filter=28 channel=21
    12, 4, 17, 0, -2, 4, 3, 0, 5,
    -- filter=28 channel=22
    0, -3, -5, 10, 3, -2, -6, 13, -4,
    -- filter=28 channel=23
    -12, -13, -11, 19, 6, -17, 6, 15, -9,
    -- filter=28 channel=24
    4, -1, -1, -2, 2, 7, -4, 0, 2,
    -- filter=28 channel=25
    4, -9, -8, 3, 23, 3, -5, 5, 2,
    -- filter=28 channel=26
    4, 11, 2, -9, 4, 0, -6, -8, -2,
    -- filter=28 channel=27
    2, -7, -15, 8, 18, -11, -8, 7, 5,
    -- filter=28 channel=28
    -6, 0, -1, -2, -5, -3, 4, 0, -3,
    -- filter=28 channel=29
    -8, 3, -2, -1, 26, 0, -7, 18, 9,
    -- filter=28 channel=30
    -2, 1, 6, 0, 12, 6, 0, -8, 5,
    -- filter=28 channel=31
    -3, -20, 12, 4, 0, -3, -5, 3, -3,
    -- filter=28 channel=32
    3, -14, -18, 2, 30, -7, -14, 9, -3,
    -- filter=28 channel=33
    -2, -12, -19, 4, 15, -8, 2, 17, 3,
    -- filter=28 channel=34
    -8, -7, -2, 14, -16, -16, 0, 5, -14,
    -- filter=28 channel=35
    0, 5, 2, -1, -4, -2, 0, -1, 2,
    -- filter=28 channel=36
    -3, -5, 3, -2, -2, 5, -5, -10, -7,
    -- filter=28 channel=37
    1, -6, -3, 2, -10, -2, -5, -9, 7,
    -- filter=28 channel=38
    0, -5, -11, 10, 0, -4, -4, 11, 7,
    -- filter=28 channel=39
    -8, 1, -2, 0, 2, -3, -9, -3, 0,
    -- filter=28 channel=40
    -7, -3, -1, -6, 3, -1, 1, 7, -8,
    -- filter=28 channel=41
    17, 0, -13, -3, 5, 3, -2, 1, -6,
    -- filter=28 channel=42
    4, -3, 4, 4, -2, 4, 0, 3, 9,
    -- filter=28 channel=43
    -14, 0, 0, 0, -5, -5, 0, 6, -7,
    -- filter=28 channel=44
    8, -9, 11, 8, -11, -4, 3, -1, -2,
    -- filter=28 channel=45
    -6, -3, 10, -1, 1, -3, -5, 3, 2,
    -- filter=28 channel=46
    -1, 7, 2, 0, -1, -1, 4, -5, 4,
    -- filter=28 channel=47
    11, -2, 5, -5, -7, -1, 0, -6, 10,
    -- filter=28 channel=48
    10, -5, -1, 0, 9, 12, -5, -12, 13,
    -- filter=28 channel=49
    5, -6, -7, 8, 26, -6, -13, 2, 2,
    -- filter=28 channel=50
    3, -8, -8, 8, 2, -8, -2, 5, 9,
    -- filter=28 channel=51
    2, 3, 7, 6, 6, -4, -1, -2, 1,
    -- filter=28 channel=52
    -10, -13, -14, -2, -10, -13, -3, 7, 0,
    -- filter=28 channel=53
    -10, -8, -3, 6, 14, 0, -1, 10, -3,
    -- filter=28 channel=54
    0, 0, -7, 0, 2, 2, 0, 5, 3,
    -- filter=28 channel=55
    -8, -15, -22, 8, 12, -14, -5, 14, -2,
    -- filter=28 channel=56
    -5, -8, -1, 9, -4, -2, -2, 5, -14,
    -- filter=28 channel=57
    0, 7, -9, 1, 0, 8, -6, -9, 5,
    -- filter=28 channel=58
    3, 2, 8, 4, 2, -9, 1, -7, 2,
    -- filter=28 channel=59
    5, -3, -4, -7, 21, 5, -5, -5, 7,
    -- filter=28 channel=60
    -4, -5, 5, 3, 2, -5, 0, 0, 4,
    -- filter=28 channel=61
    -1, -7, 2, -8, -5, -6, 0, -7, -5,
    -- filter=28 channel=62
    3, 2, -8, -6, -4, -8, -1, 4, 4,
    -- filter=28 channel=63
    8, 0, 10, -7, 0, 4, -1, -6, 2,
    -- filter=28 channel=64
    -4, -8, -2, -5, -7, 1, -2, 5, 0,
    -- filter=28 channel=65
    0, 3, -7, 7, 0, 0, 2, 0, 6,
    -- filter=28 channel=66
    1, -4, -10, 2, 5, -12, -1, 0, -9,
    -- filter=28 channel=67
    -2, 5, 3, 5, 1, -6, 0, -6, 3,
    -- filter=28 channel=68
    -8, -5, -5, -1, -2, 7, 0, 3, -5,
    -- filter=28 channel=69
    1, 4, 6, 0, 6, -7, 5, 2, 4,
    -- filter=28 channel=70
    -11, -12, -17, 13, 3, -15, 3, 13, 0,
    -- filter=28 channel=71
    -2, -6, 5, 0, -10, -8, 0, 1, 4,
    -- filter=28 channel=72
    3, -5, 3, -2, 1, 3, -4, 3, 4,
    -- filter=28 channel=73
    -6, -5, -8, 1, 13, 4, 0, -3, 1,
    -- filter=28 channel=74
    4, -13, -5, 14, -3, -18, 0, 9, -18,
    -- filter=28 channel=75
    -8, -3, -8, 1, -1, -16, -7, 7, 11,
    -- filter=28 channel=76
    -12, -7, -12, -3, 21, -10, 0, 13, -6,
    -- filter=28 channel=77
    7, -7, -6, 0, 2, -3, -2, 1, 6,
    -- filter=28 channel=78
    -2, 3, -4, -3, -5, 0, 11, -3, 1,
    -- filter=28 channel=79
    4, -7, -29, 9, 39, -19, -9, 25, -6,
    -- filter=28 channel=80
    6, 3, 6, -7, 9, 0, -10, -1, 7,
    -- filter=28 channel=81
    5, 0, 5, 5, 0, 6, 4, -2, -1,
    -- filter=28 channel=82
    -2, -2, 1, -1, -4, -5, 6, 0, -5,
    -- filter=28 channel=83
    9, 0, 4, -6, 5, 14, -8, -8, 7,
    -- filter=28 channel=84
    4, -10, -9, 0, 11, -5, -1, 1, -4,
    -- filter=28 channel=85
    -4, 3, -5, -2, 1, 0, 1, -3, -5,
    -- filter=28 channel=86
    5, -10, -1, 3, 2, -15, -2, -1, -4,
    -- filter=28 channel=87
    -4, -6, -4, 7, 7, -6, -8, 2, -4,
    -- filter=28 channel=88
    4, -5, 7, -7, 0, 2, -1, -4, -7,
    -- filter=28 channel=89
    2, -10, -5, 1, 23, -1, -5, 12, 4,
    -- filter=28 channel=90
    -3, -8, 0, -1, -20, -6, 2, 7, 0,
    -- filter=28 channel=91
    4, -2, -11, 8, 29, 2, -11, 8, -6,
    -- filter=28 channel=92
    -5, -3, -2, -2, -4, 0, 1, 5, 1,
    -- filter=28 channel=93
    19, -8, -2, -2, -4, 12, -1, -18, 7,
    -- filter=28 channel=94
    -3, 1, 2, 6, 5, 3, -1, 1, -1,
    -- filter=28 channel=95
    3, -8, -3, 1, -4, -9, 7, 0, -3,
    -- filter=28 channel=96
    -2, 0, 0, 4, 0, -5, 1, 8, 4,
    -- filter=28 channel=97
    -1, -10, 0, 1, -10, -4, -4, -2, 0,
    -- filter=28 channel=98
    8, -14, -5, 1, 9, -13, -1, 10, -1,
    -- filter=28 channel=99
    -5, -20, -11, 17, -2, -14, 1, 12, -10,
    -- filter=28 channel=100
    -2, 0, 0, 2, -9, -3, 4, 4, -5,
    -- filter=28 channel=101
    -1, -3, -8, -10, -3, 4, -6, -3, -5,
    -- filter=28 channel=102
    1, -3, 1, -6, 4, 0, -6, -4, -3,
    -- filter=28 channel=103
    -5, -7, 8, 2, -5, -1, 5, 2, 7,
    -- filter=28 channel=104
    4, -6, 6, -6, 9, 11, 2, -7, -2,
    -- filter=28 channel=105
    -4, 2, -5, 6, 6, -2, 7, 14, -3,
    -- filter=28 channel=106
    4, -5, -5, -8, 4, 1, 1, 0, 1,
    -- filter=28 channel=107
    -5, 0, -14, 12, 10, -7, 5, 16, -5,
    -- filter=28 channel=108
    2, -3, -5, 1, 6, 5, 3, -2, 2,
    -- filter=28 channel=109
    8, -2, -18, 11, 21, -2, -14, 8, 4,
    -- filter=28 channel=110
    -3, -9, 2, 7, -8, -4, 0, -4, -7,
    -- filter=28 channel=111
    2, 2, 0, 0, 0, 5, 6, -1, 0,
    -- filter=28 channel=112
    -2, -6, -12, 0, 1, -16, 4, 11, 0,
    -- filter=28 channel=113
    -7, -17, -4, -1, -4, -16, -3, 14, 3,
    -- filter=28 channel=114
    4, 1, -16, 10, 28, -11, -6, 9, 1,
    -- filter=28 channel=115
    -1, 0, 1, -5, 5, -2, 8, 7, 0,
    -- filter=28 channel=116
    3, -5, -13, 6, 22, 7, -9, 1, 11,
    -- filter=28 channel=117
    2, -4, -2, 3, 0, 4, -4, 3, 1,
    -- filter=28 channel=118
    -4, 5, -4, -6, 0, -7, -1, -2, -1,
    -- filter=28 channel=119
    2, -1, -9, 3, -4, -22, 8, 0, -16,
    -- filter=28 channel=120
    -10, -9, -28, 26, 10, -11, -2, 13, -3,
    -- filter=28 channel=121
    7, -10, -10, 4, -3, -1, -6, 0, 0,
    -- filter=28 channel=122
    7, -5, 21, -2, -7, 0, -3, -6, 7,
    -- filter=28 channel=123
    5, -1, 0, -1, 0, 2, -1, -1, -10,
    -- filter=28 channel=124
    2, -1, -1, 7, 9, -10, 2, 3, 6,
    -- filter=28 channel=125
    11, -13, -13, 6, 7, -3, 0, 1, 9,
    -- filter=28 channel=126
    -9, -13, -7, 5, 13, -7, 4, 4, 8,
    -- filter=28 channel=127
    5, -3, -6, 7, -6, 0, 4, -8, -5,
    -- filter=29 channel=0
    6, 9, 0, 7, 15, 1, 7, -9, -7,
    -- filter=29 channel=1
    11, 0, -3, 15, 6, -1, 4, -4, -3,
    -- filter=29 channel=2
    0, -4, -1, 1, -2, 5, -7, 5, 8,
    -- filter=29 channel=3
    -2, 11, 4, -14, -3, -7, -5, -8, 1,
    -- filter=29 channel=4
    -3, -11, 1, -11, 5, 7, -7, 9, 9,
    -- filter=29 channel=5
    -8, 8, 3, -2, 9, -3, -10, 3, -6,
    -- filter=29 channel=6
    8, -8, -3, -2, 6, 5, 1, -6, 6,
    -- filter=29 channel=7
    6, 1, 3, -4, 0, -4, 2, -4, -2,
    -- filter=29 channel=8
    -2, 5, 2, -6, 5, 4, 1, 5, 5,
    -- filter=29 channel=9
    5, 5, -7, 1, -6, -3, 4, 5, -4,
    -- filter=29 channel=10
    12, -4, 0, 14, -11, 4, 5, -6, 1,
    -- filter=29 channel=11
    6, 3, -4, -4, -2, 1, -1, 1, 13,
    -- filter=29 channel=12
    7, 7, 4, 19, -7, 5, 2, -1, 2,
    -- filter=29 channel=13
    14, -1, 0, 29, -23, -7, 13, -11, 1,
    -- filter=29 channel=14
    -3, -3, 0, 4, 4, 2, 1, 3, -4,
    -- filter=29 channel=15
    15, -3, -4, 6, -11, -14, 4, -7, -5,
    -- filter=29 channel=16
    -1, 6, 10, -8, -6, 5, 2, 2, -6,
    -- filter=29 channel=17
    -2, 5, 0, 1, 2, -4, -2, -6, 3,
    -- filter=29 channel=18
    33, -12, -22, 34, -15, -6, 15, -17, -6,
    -- filter=29 channel=19
    5, -1, -2, 2, 3, -2, -4, 4, 0,
    -- filter=29 channel=20
    6, -7, -4, -3, 0, 6, 3, -4, 7,
    -- filter=29 channel=21
    2, 9, 10, 0, 3, -6, 0, 10, -8,
    -- filter=29 channel=22
    -3, -4, 3, 6, -6, -9, -2, -9, -8,
    -- filter=29 channel=23
    2, -10, -10, -7, -27, -7, -14, -5, 2,
    -- filter=29 channel=24
    -2, -6, 0, 2, 0, -3, 4, 4, 0,
    -- filter=29 channel=25
    25, -1, -1, 17, -15, -2, 4, -4, -12,
    -- filter=29 channel=26
    -10, -3, -1, -8, 0, -1, -9, 5, 0,
    -- filter=29 channel=27
    12, -19, -6, 15, -23, -10, 0, 1, -6,
    -- filter=29 channel=28
    7, 6, 0, 2, 0, -5, 7, -1, -4,
    -- filter=29 channel=29
    13, 2, -13, 7, 0, 3, 5, 2, 4,
    -- filter=29 channel=30
    -2, 0, 1, 0, -1, 3, -4, 0, 5,
    -- filter=29 channel=31
    6, 0, -1, -11, -5, -4, -2, 16, 15,
    -- filter=29 channel=32
    27, -9, -8, 16, -24, -8, 7, -6, -10,
    -- filter=29 channel=33
    12, -8, -11, 14, -14, -5, -3, -16, -11,
    -- filter=29 channel=34
    7, 0, 5, 2, 12, -5, -1, -7, 0,
    -- filter=29 channel=35
    5, 4, 6, -4, 5, -3, 3, 1, 3,
    -- filter=29 channel=36
    11, 3, 7, -3, -3, 2, -3, 2, 6,
    -- filter=29 channel=37
    -7, 2, 12, -12, 6, 5, -9, 0, -1,
    -- filter=29 channel=38
    11, 0, 3, 6, -12, -5, 0, 0, 1,
    -- filter=29 channel=39
    -3, 2, -3, 1, -5, 0, 3, -3, 0,
    -- filter=29 channel=40
    7, -8, -6, 0, -7, 3, 0, -1, 0,
    -- filter=29 channel=41
    30, 5, 5, 48, -6, -7, 31, -11, -16,
    -- filter=29 channel=42
    6, -2, -6, -5, 7, -4, -3, 9, 2,
    -- filter=29 channel=43
    5, 12, -5, -4, -10, 0, -8, -16, -3,
    -- filter=29 channel=44
    3, 5, 7, -8, 0, 0, -10, 8, -2,
    -- filter=29 channel=45
    -10, 6, -6, -5, 6, 3, -2, 4, 6,
    -- filter=29 channel=46
    0, 0, -2, 10, -3, -4, -2, -5, 4,
    -- filter=29 channel=47
    -1, -2, 7, -2, -5, -2, 0, 7, 0,
    -- filter=29 channel=48
    16, -8, -2, 3, -4, -1, -7, 3, 4,
    -- filter=29 channel=49
    1, -9, -8, 4, -9, -8, -6, 1, 4,
    -- filter=29 channel=50
    -1, -4, -5, 0, -14, -5, 8, 3, -5,
    -- filter=29 channel=51
    4, 6, 3, 6, -5, -5, 1, 0, 3,
    -- filter=29 channel=52
    -2, -3, -2, -9, 3, -2, -10, -1, 7,
    -- filter=29 channel=53
    -3, 4, -5, 7, -3, 5, 5, 1, 6,
    -- filter=29 channel=54
    2, 1, 0, 1, 3, -4, 5, 5, 0,
    -- filter=29 channel=55
    22, -13, -15, 22, -17, -9, 11, -18, 2,
    -- filter=29 channel=56
    0, 7, 1, -2, 7, -2, 4, 0, 10,
    -- filter=29 channel=57
    3, -9, -1, 9, -9, -6, 8, -7, -4,
    -- filter=29 channel=58
    -3, 2, 3, -5, 17, 2, -10, 9, -3,
    -- filter=29 channel=59
    22, -5, 3, 14, -20, -13, 13, 0, 0,
    -- filter=29 channel=60
    -5, -6, 5, -6, -2, -1, 5, 3, -2,
    -- filter=29 channel=61
    5, 7, -1, 0, 2, 2, 3, 3, 1,
    -- filter=29 channel=62
    7, -4, -6, -7, 1, 1, 5, -7, -1,
    -- filter=29 channel=63
    -10, 11, 9, -1, 9, 7, -10, 0, 6,
    -- filter=29 channel=64
    -3, 8, -1, -3, -4, -1, 6, -2, 9,
    -- filter=29 channel=65
    1, -4, -6, 6, -3, -7, 1, -1, 4,
    -- filter=29 channel=66
    5, -2, 10, 25, -16, 6, 4, -11, 1,
    -- filter=29 channel=67
    -1, 0, -4, 0, 0, 6, 2, 4, -1,
    -- filter=29 channel=68
    2, -1, 0, -1, 4, -4, 3, 2, 5,
    -- filter=29 channel=69
    2, 6, 7, 9, 3, -1, 3, -5, 1,
    -- filter=29 channel=70
    6, -8, -6, -4, -6, -6, -7, -9, 1,
    -- filter=29 channel=71
    1, -2, -2, -8, 2, -7, -7, -10, 1,
    -- filter=29 channel=72
    17, 0, -2, 7, -12, -4, 0, 6, 1,
    -- filter=29 channel=73
    10, -3, -2, 0, -14, 1, -3, -7, 1,
    -- filter=29 channel=74
    6, -7, 2, -9, -2, -5, -15, 3, 0,
    -- filter=29 channel=75
    4, 15, 5, 19, 4, -1, 1, -14, -11,
    -- filter=29 channel=76
    15, 0, -4, 15, -13, -8, 5, -3, -1,
    -- filter=29 channel=77
    -3, -7, 6, 6, 3, -3, -4, -4, 4,
    -- filter=29 channel=78
    -2, 3, 5, -12, 4, 4, -10, -4, 3,
    -- filter=29 channel=79
    35, -4, -15, 39, -28, -9, 11, -16, -11,
    -- filter=29 channel=80
    22, -4, 0, 19, -8, 0, 7, 3, 5,
    -- filter=29 channel=81
    -4, 0, 1, -3, 0, 5, 3, -7, 6,
    -- filter=29 channel=82
    3, -6, 0, -3, -5, -7, -2, -3, -2,
    -- filter=29 channel=83
    5, -3, -8, -1, -3, -2, 3, 3, 3,
    -- filter=29 channel=84
    9, -18, -3, 2, -2, -2, 3, -3, 3,
    -- filter=29 channel=85
    6, 1, 6, -1, -4, -2, 3, 4, 0,
    -- filter=29 channel=86
    0, -5, 5, 4, 6, 7, -7, -8, -4,
    -- filter=29 channel=87
    -1, -8, 6, -3, -3, -2, 5, 0, 4,
    -- filter=29 channel=88
    -2, 4, 8, -3, 0, 11, -2, 3, 9,
    -- filter=29 channel=89
    29, -6, 0, 27, -25, -2, 12, -4, 1,
    -- filter=29 channel=90
    -7, 5, 7, -12, 0, -3, -5, -2, 8,
    -- filter=29 channel=91
    7, -18, 0, -4, -15, -10, 6, -6, 6,
    -- filter=29 channel=92
    -5, 4, -3, -2, -5, 0, -3, -4, -4,
    -- filter=29 channel=93
    7, 6, 7, -11, 1, -7, -4, 0, 2,
    -- filter=29 channel=94
    -6, -2, -4, 4, 4, 5, 5, 1, 1,
    -- filter=29 channel=95
    -4, 2, 3, -6, 3, 2, 1, 0, -3,
    -- filter=29 channel=96
    4, -4, -1, 2, 5, -6, 8, 2, -1,
    -- filter=29 channel=97
    -5, 8, 7, 0, 2, 0, -1, -8, 0,
    -- filter=29 channel=98
    20, 5, -6, 20, -15, -6, 1, -7, 0,
    -- filter=29 channel=99
    11, -11, -9, 1, -11, -5, -8, 6, 8,
    -- filter=29 channel=100
    0, 10, -3, -1, 1, -2, 8, -8, -2,
    -- filter=29 channel=101
    -1, -4, 0, -13, -6, 0, -12, 1, 0,
    -- filter=29 channel=102
    -6, 0, 7, 0, 4, 2, 1, 5, -6,
    -- filter=29 channel=103
    -1, 1, 1, -11, -1, -9, 3, 6, -10,
    -- filter=29 channel=104
    9, 0, -2, 10, -9, -5, 4, 2, 2,
    -- filter=29 channel=105
    -1, -4, 3, 1, -4, -7, -5, -10, -3,
    -- filter=29 channel=106
    11, 4, -8, 5, 1, 1, 9, 0, -2,
    -- filter=29 channel=107
    0, -6, -8, -1, 1, 6, -8, -5, 0,
    -- filter=29 channel=108
    6, 3, 6, 12, 3, 2, 1, 1, 0,
    -- filter=29 channel=109
    31, -16, -11, 20, -24, -12, 0, -8, 2,
    -- filter=29 channel=110
    -1, 1, -1, 7, -6, 0, 0, 7, 0,
    -- filter=29 channel=111
    1, 1, -5, 14, -4, -6, 5, 3, 4,
    -- filter=29 channel=112
    -9, 0, 0, -6, -6, -1, -9, -11, 0,
    -- filter=29 channel=113
    16, 2, 3, 2, -5, -10, 2, -12, -7,
    -- filter=29 channel=114
    29, -8, -5, 27, -13, 0, 1, 1, 0,
    -- filter=29 channel=115
    -1, -5, 0, -1, 1, -6, 7, 5, 3,
    -- filter=29 channel=116
    27, -4, 1, 14, -7, -10, 11, 0, 0,
    -- filter=29 channel=117
    8, -2, 2, 9, -3, -2, -6, -2, 5,
    -- filter=29 channel=118
    -3, 4, 1, 3, 1, 1, -3, 2, -1,
    -- filter=29 channel=119
    6, -3, 5, 4, 11, -3, 7, -6, 5,
    -- filter=29 channel=120
    16, -23, 0, -12, -21, -5, -5, -2, 8,
    -- filter=29 channel=121
    13, 2, 0, 16, -10, -4, 7, -9, 3,
    -- filter=29 channel=122
    -2, -3, 8, -16, -7, -3, -16, 6, -7,
    -- filter=29 channel=123
    1, 3, 5, -8, 4, -6, -7, 0, 6,
    -- filter=29 channel=124
    0, -4, 0, 5, -7, -2, 2, -6, 1,
    -- filter=29 channel=125
    10, 3, 5, 3, -12, -7, 9, 1, 3,
    -- filter=29 channel=126
    26, 12, -10, 32, -10, 0, 12, -14, -7,
    -- filter=29 channel=127
    11, 4, -6, 14, -8, 3, 4, -4, 1,
    -- filter=30 channel=0
    0, 14, 16, 0, 10, 0, -14, -19, -5,
    -- filter=30 channel=1
    6, 8, 15, 1, 2, -12, -4, -9, -18,
    -- filter=30 channel=2
    -5, 13, 0, -1, -8, 1, 4, -6, 0,
    -- filter=30 channel=3
    5, 19, 30, -8, 30, 15, -4, -11, 2,
    -- filter=30 channel=4
    4, 25, 13, 6, -8, 13, -9, 5, 7,
    -- filter=30 channel=5
    7, 12, 11, 12, 15, 10, -17, -20, -11,
    -- filter=30 channel=6
    1, 3, -1, 4, 0, -6, 6, -1, 7,
    -- filter=30 channel=7
    1, -3, 4, -5, -6, 6, -6, -4, 1,
    -- filter=30 channel=8
    7, 8, 5, 0, -6, -3, -11, -4, -1,
    -- filter=30 channel=9
    3, 7, 0, 4, -9, -4, -2, -4, -6,
    -- filter=30 channel=10
    -4, 13, 8, 0, 13, 3, 2, -17, -12,
    -- filter=30 channel=11
    -5, 2, 0, -2, -5, -2, 3, -1, 1,
    -- filter=30 channel=12
    -5, -3, -2, 6, -4, -2, 0, -11, 4,
    -- filter=30 channel=13
    1, 0, 24, -1, -6, -7, 8, -15, -11,
    -- filter=30 channel=14
    4, -6, -2, -7, 6, -5, 2, -6, -5,
    -- filter=30 channel=15
    -2, 3, 13, -9, 7, 4, 1, -4, -9,
    -- filter=30 channel=16
    -1, 0, 12, 7, 9, -1, -8, -11, -6,
    -- filter=30 channel=17
    3, 1, -1, -1, 6, -6, -6, 0, -6,
    -- filter=30 channel=18
    -14, 7, 30, -4, 2, -15, 4, -12, -18,
    -- filter=30 channel=19
    -6, -1, 0, -6, -3, 1, 5, -2, 7,
    -- filter=30 channel=20
    -9, -4, 5, -10, 0, 1, 8, -4, 10,
    -- filter=30 channel=21
    6, 11, 0, -2, 3, 1, -1, -3, -2,
    -- filter=30 channel=22
    0, 3, 1, -6, 4, 10, 0, 0, 1,
    -- filter=30 channel=23
    -2, 14, 21, -10, 10, 4, 5, -26, -6,
    -- filter=30 channel=24
    1, -6, 3, -6, 4, 5, -1, -1, -5,
    -- filter=30 channel=25
    4, 19, 14, 3, -11, -14, 4, -11, -13,
    -- filter=30 channel=26
    1, 5, -1, 2, -8, -5, -6, 0, 3,
    -- filter=30 channel=27
    0, 35, 18, 0, -3, -17, 3, -27, -9,
    -- filter=30 channel=28
    -5, -4, 2, 3, -6, -6, 0, -2, 2,
    -- filter=30 channel=29
    -7, 4, 9, 0, -5, 3, 15, 0, 4,
    -- filter=30 channel=30
    6, 20, 2, -6, -6, -14, -5, -19, -3,
    -- filter=30 channel=31
    2, 21, 7, -13, -8, 3, -10, -27, -11,
    -- filter=30 channel=32
    -4, 21, 15, -7, -8, -11, -4, -9, -5,
    -- filter=30 channel=33
    -6, 16, 13, 5, 21, 3, 4, -26, -21,
    -- filter=30 channel=34
    -9, 17, -5, 5, -1, -2, -2, -12, -3,
    -- filter=30 channel=35
    -6, 1, 5, -5, -1, 5, 1, 4, -5,
    -- filter=30 channel=36
    -6, -3, 2, 2, -18, -5, 4, -1, 0,
    -- filter=30 channel=37
    1, 13, 9, 6, -7, -9, -8, -15, 2,
    -- filter=30 channel=38
    -3, 9, 8, -4, 6, -6, -3, -5, -12,
    -- filter=30 channel=39
    -7, 2, -4, -5, -5, -4, 8, 4, 12,
    -- filter=30 channel=40
    -4, -8, 1, -7, 0, -3, 4, -8, -3,
    -- filter=30 channel=41
    -4, 2, 6, -12, 3, -2, 8, 19, -15,
    -- filter=30 channel=42
    4, 8, -1, 3, 0, -2, -2, -10, -8,
    -- filter=30 channel=43
    -1, 12, 16, -8, 14, 16, -8, -1, -2,
    -- filter=30 channel=44
    11, 22, 2, 0, -4, -1, -11, -12, -6,
    -- filter=30 channel=45
    1, 0, -2, -5, -7, 2, -4, -5, -3,
    -- filter=30 channel=46
    -4, -5, 4, -3, 7, -6, -2, 0, 0,
    -- filter=30 channel=47
    5, 14, 3, 0, 1, 5, -9, -10, -11,
    -- filter=30 channel=48
    5, 28, 17, -2, -20, -25, -4, -19, -1,
    -- filter=30 channel=49
    -8, 10, 10, -8, -17, -11, -1, -5, 0,
    -- filter=30 channel=50
    -7, 16, 5, -7, -5, 0, 3, -16, -6,
    -- filter=30 channel=51
    0, -6, -3, -4, 6, -3, -4, 5, -3,
    -- filter=30 channel=52
    3, 7, 3, 0, 0, 3, 3, 2, 3,
    -- filter=30 channel=53
    0, -6, -1, -5, -9, 0, 10, -9, 7,
    -- filter=30 channel=54
    0, 0, 7, 5, -7, 0, -5, 0, 1,
    -- filter=30 channel=55
    1, 1, 20, -1, -1, -11, 12, -17, -7,
    -- filter=30 channel=56
    -1, 7, -4, -5, 0, -2, -3, 5, 5,
    -- filter=30 channel=57
    0, -2, 8, -8, 0, -5, -6, 4, 3,
    -- filter=30 channel=58
    -4, -5, -1, -6, -3, 2, -1, -5, -1,
    -- filter=30 channel=59
    -1, 9, 19, -3, -7, -9, -4, -6, -8,
    -- filter=30 channel=60
    -2, -5, -2, 0, -3, -1, 3, 2, -2,
    -- filter=30 channel=61
    3, 10, 1, -7, -4, -10, 0, -5, 2,
    -- filter=30 channel=62
    7, -4, 5, 4, -4, -5, 3, 4, 1,
    -- filter=30 channel=63
    -6, -4, 4, 7, -3, -8, -3, 0, -4,
    -- filter=30 channel=64
    -3, 0, -6, 0, 2, 8, 1, 8, 8,
    -- filter=30 channel=65
    -5, -2, -4, 1, 0, 4, 0, 6, -3,
    -- filter=30 channel=66
    -4, -1, 0, 6, -4, -11, 2, 4, -4,
    -- filter=30 channel=67
    -5, -3, -1, -7, -3, 6, -4, 0, 1,
    -- filter=30 channel=68
    -5, 4, 5, -7, -7, -5, 0, 6, 9,
    -- filter=30 channel=69
    1, -2, -5, -2, 1, -1, 6, -5, -4,
    -- filter=30 channel=70
    0, 20, 6, 1, -3, -10, -7, -16, -11,
    -- filter=30 channel=71
    6, 10, 2, 0, 7, 9, 3, -9, -7,
    -- filter=30 channel=72
    0, 5, 7, -8, 3, 1, 2, -15, -1,
    -- filter=30 channel=73
    5, 6, 9, -2, 0, -16, 0, -4, 3,
    -- filter=30 channel=74
    7, 21, -2, 3, -12, -2, -5, -18, 2,
    -- filter=30 channel=75
    14, 18, 21, 6, 17, 14, -17, -29, -26,
    -- filter=30 channel=76
    -10, -11, -1, 2, 0, -2, 9, 5, -2,
    -- filter=30 channel=77
    1, 3, 1, 4, 3, 0, 6, -2, 3,
    -- filter=30 channel=78
    9, 7, 0, 5, 0, 6, 0, -4, -5,
    -- filter=30 channel=79
    -13, 14, 27, 3, 3, -3, 10, -21, -24,
    -- filter=30 channel=80
    -7, 15, 18, -4, -7, -7, -7, -26, -11,
    -- filter=30 channel=81
    1, -5, -7, -4, -4, 6, 2, -3, 5,
    -- filter=30 channel=82
    5, 3, 3, 6, -4, 1, -2, -10, 2,
    -- filter=30 channel=83
    -1, 8, -4, -5, -16, -3, -8, -3, -2,
    -- filter=30 channel=84
    -4, 11, 7, 0, -10, -16, 3, -6, -5,
    -- filter=30 channel=85
    7, -4, 6, 5, 2, -4, 1, -6, 0,
    -- filter=30 channel=86
    3, 13, -6, 2, -5, 1, 0, -8, -3,
    -- filter=30 channel=87
    6, -1, 8, 2, -9, 1, 8, 3, 1,
    -- filter=30 channel=88
    -3, 11, -2, 1, -1, 3, -1, -4, 9,
    -- filter=30 channel=89
    -8, 0, 17, 0, 7, -2, 4, -16, -10,
    -- filter=30 channel=90
    4, 10, 0, -3, -3, 9, 0, -7, 0,
    -- filter=30 channel=91
    0, 18, 7, -8, -25, -19, -3, -17, -8,
    -- filter=30 channel=92
    -5, 3, -4, 0, 8, -1, -5, -2, -5,
    -- filter=30 channel=93
    11, 16, 10, 5, -7, -14, -5, -8, -5,
    -- filter=30 channel=94
    -2, -1, 4, -1, -6, 6, -5, -5, -7,
    -- filter=30 channel=95
    4, 0, 6, -5, 8, 4, 0, 6, 2,
    -- filter=30 channel=96
    3, -4, 5, -4, -7, 8, 7, 2, -7,
    -- filter=30 channel=97
    6, 8, 4, 0, 13, 17, -6, -12, -8,
    -- filter=30 channel=98
    -6, 14, 20, 2, 16, -10, 6, -14, -7,
    -- filter=30 channel=99
    -1, 21, 11, -3, -9, -13, 2, -28, -9,
    -- filter=30 channel=100
    4, -3, -2, -4, 0, -9, -6, 0, -8,
    -- filter=30 channel=101
    7, 16, 8, -2, -6, 8, -6, 7, 12,
    -- filter=30 channel=102
    -6, -2, -3, 5, -1, -1, -7, -6, -3,
    -- filter=30 channel=103
    0, 19, 12, 2, 11, 0, -4, -12, -10,
    -- filter=30 channel=104
    6, 21, 5, 0, -5, -3, -5, -6, -8,
    -- filter=30 channel=105
    -1, 0, 12, -1, -4, 2, 8, 0, 2,
    -- filter=30 channel=106
    -3, -7, 1, -2, 5, -5, 10, 2, -4,
    -- filter=30 channel=107
    1, 5, -1, -1, 6, 0, -2, 0, 2,
    -- filter=30 channel=108
    -5, 6, 8, 1, 6, -4, 1, -5, -1,
    -- filter=30 channel=109
    -5, 27, 11, -3, -11, -25, -2, -25, -12,
    -- filter=30 channel=110
    0, 10, 6, -1, 6, 6, 4, -15, -6,
    -- filter=30 channel=111
    5, 5, 6, 0, 7, 1, 8, 3, -3,
    -- filter=30 channel=112
    0, 15, 0, 0, -4, 0, -4, -16, 0,
    -- filter=30 channel=113
    -2, 15, 17, 1, 18, 13, -5, -14, -11,
    -- filter=30 channel=114
    -8, 27, 14, -4, -2, -22, -4, -24, -1,
    -- filter=30 channel=115
    2, -3, -5, -6, -5, -4, 4, 1, 2,
    -- filter=30 channel=116
    0, 22, 8, -1, -10, -14, -2, -9, -9,
    -- filter=30 channel=117
    -5, 5, 3, 0, -1, -8, -4, -10, -5,
    -- filter=30 channel=118
    1, -2, -2, 3, 4, -4, 1, -3, -6,
    -- filter=30 channel=119
    -2, 2, -11, 2, -14, 0, -8, -2, -1,
    -- filter=30 channel=120
    7, 36, 9, 6, -26, -19, -1, -29, -3,
    -- filter=30 channel=121
    4, 5, 14, -5, 11, 7, 1, 2, -11,
    -- filter=30 channel=122
    12, 22, 7, 6, -2, 0, -4, -20, 3,
    -- filter=30 channel=123
    -1, 8, 5, -3, 6, 6, 2, 0, -4,
    -- filter=30 channel=124
    -4, 1, 10, 6, 5, 1, 9, 4, -3,
    -- filter=30 channel=125
    1, 22, 18, 0, -9, -20, -5, -11, -5,
    -- filter=30 channel=126
    -3, 7, 11, 3, 16, 1, -6, -4, -21,
    -- filter=30 channel=127
    -1, -1, 0, -7, 3, -8, -1, 2, -4,
    -- filter=31 channel=0
    -6, -9, 4, -13, 14, 16, -5, 7, 15,
    -- filter=31 channel=1
    -7, -10, 1, -12, 5, 19, -13, -5, 13,
    -- filter=31 channel=2
    5, 7, -5, 2, 1, -5, -2, 1, -9,
    -- filter=31 channel=3
    -5, -16, -12, 1, -10, 5, 6, -4, -3,
    -- filter=31 channel=4
    0, -11, -4, -2, -8, -4, -8, -22, -7,
    -- filter=31 channel=5
    -5, -9, -7, 13, 5, 2, 0, 0, 7,
    -- filter=31 channel=6
    -8, 10, 7, -1, 10, 3, -1, 5, -2,
    -- filter=31 channel=7
    5, 6, -2, -4, -1, 0, 5, 6, 6,
    -- filter=31 channel=8
    -4, 3, 3, -6, -5, -5, 0, -1, -1,
    -- filter=31 channel=9
    6, 0, 8, 4, 1, 3, 8, -6, 5,
    -- filter=31 channel=10
    0, 4, -6, 3, 6, -3, 2, -2, -7,
    -- filter=31 channel=11
    7, 0, 0, 3, 8, -1, 5, 4, 3,
    -- filter=31 channel=12
    -5, 2, -6, -11, 3, -1, 0, 3, 4,
    -- filter=31 channel=13
    -10, -6, -10, -16, 14, 3, -15, 4, 0,
    -- filter=31 channel=14
    6, -5, -6, 7, 0, 6, -3, 1, -5,
    -- filter=31 channel=15
    -12, 4, 5, -3, 18, 3, -12, 15, 0,
    -- filter=31 channel=16
    3, -8, -2, 7, 6, -2, -1, -2, 3,
    -- filter=31 channel=17
    -1, 0, 6, -4, 4, 1, 6, 4, -1,
    -- filter=31 channel=18
    -17, 1, 6, -22, 21, 16, -10, 14, 6,
    -- filter=31 channel=19
    7, -2, 2, 5, -3, 1, 7, 5, 1,
    -- filter=31 channel=20
    -10, 9, 1, 2, 7, -6, 4, 11, -10,
    -- filter=31 channel=21
    13, -4, -4, 20, -8, 0, 10, -11, -11,
    -- filter=31 channel=22
    -1, -2, 4, -9, 9, 11, -11, 0, 5,
    -- filter=31 channel=23
    -17, -4, 6, -6, 4, -6, -5, 14, -4,
    -- filter=31 channel=24
    0, -4, 7, 3, -6, 6, 6, 6, -2,
    -- filter=31 channel=25
    0, -6, 9, -10, 12, 5, -12, 7, -4,
    -- filter=31 channel=26
    2, 2, 3, 11, -5, -11, 7, -6, -1,
    -- filter=31 channel=27
    -2, -3, -1, -7, 24, 13, -16, 9, -1,
    -- filter=31 channel=28
    4, -5, -5, 2, -4, 0, 2, 0, -6,
    -- filter=31 channel=29
    5, 11, 1, 3, 9, -13, 5, 14, -1,
    -- filter=31 channel=30
    -5, -3, 3, 0, 8, 9, 2, -5, 3,
    -- filter=31 channel=31
    15, 0, -2, 12, -6, -7, 9, -9, -10,
    -- filter=31 channel=32
    -15, 0, 2, -18, 21, 4, -5, 5, 5,
    -- filter=31 channel=33
    -18, -6, -2, -7, 17, 10, -7, 17, 3,
    -- filter=31 channel=34
    -9, 5, 5, -4, 5, 0, -13, 0, -1,
    -- filter=31 channel=35
    6, -5, 4, 0, 4, 5, 0, 5, 4,
    -- filter=31 channel=36
    7, 4, -3, 8, 4, -12, -5, -11, -11,
    -- filter=31 channel=37
    -9, -5, -2, 5, -2, 0, -7, -6, 6,
    -- filter=31 channel=38
    4, 1, 2, 1, 7, -5, -5, 0, 3,
    -- filter=31 channel=39
    -1, 1, 6, -3, -1, -10, 2, 0, -5,
    -- filter=31 channel=40
    -5, 0, -2, 2, -2, -8, -5, 12, -3,
    -- filter=31 channel=41
    -30, -2, -7, -35, 10, -2, -25, 5, -3,
    -- filter=31 channel=42
    7, -2, -1, 3, 6, 7, 0, -2, 5,
    -- filter=31 channel=43
    -9, -12, -6, -1, -5, 10, -2, 13, 3,
    -- filter=31 channel=44
    -1, 5, -3, 12, 9, 0, 0, 0, 0,
    -- filter=31 channel=45
    -5, 4, -6, -1, -6, 8, 1, 9, 5,
    -- filter=31 channel=46
    0, 4, -5, 0, -2, 6, -2, -5, 6,
    -- filter=31 channel=47
    0, -8, 3, 18, 1, 8, 8, -12, 3,
    -- filter=31 channel=48
    13, 9, 2, -3, 4, 1, -5, -14, -5,
    -- filter=31 channel=49
    -4, 3, 4, -2, 3, 5, -1, 5, 2,
    -- filter=31 channel=50
    -2, 2, 2, 1, 0, 7, 0, -7, -2,
    -- filter=31 channel=51
    -6, 5, 3, -4, 3, -5, 1, -2, 6,
    -- filter=31 channel=52
    -2, 3, -1, -5, 0, 2, -7, -6, 2,
    -- filter=31 channel=53
    0, 3, 3, -7, 7, -1, -2, -4, -7,
    -- filter=31 channel=54
    -1, -2, -6, -5, -5, -7, -7, -2, -5,
    -- filter=31 channel=55
    -12, 1, 4, -9, 5, 1, -8, 13, -4,
    -- filter=31 channel=56
    0, -2, -7, 1, -2, -7, -12, 0, -6,
    -- filter=31 channel=57
    -2, -2, 2, -1, -8, 0, -9, -10, -2,
    -- filter=31 channel=58
    6, 2, -10, 3, 0, 1, 2, 1, 1,
    -- filter=31 channel=59
    -1, 5, 0, 0, 13, 11, -8, -7, -6,
    -- filter=31 channel=60
    5, 1, -7, -6, 3, -3, 3, 5, -5,
    -- filter=31 channel=61
    -5, 3, -1, -6, 1, 4, -2, -1, -3,
    -- filter=31 channel=62
    0, -2, -9, 0, 3, 3, -3, -6, 4,
    -- filter=31 channel=63
    0, -7, 5, 5, 1, 5, 9, -3, 4,
    -- filter=31 channel=64
    9, 7, -4, 0, -2, -10, -3, 1, -10,
    -- filter=31 channel=65
    -3, 5, 6, -5, -5, -3, -6, 3, -6,
    -- filter=31 channel=66
    -9, 7, -12, -10, 2, 1, 0, -3, -6,
    -- filter=31 channel=67
    -2, -6, 3, 2, 2, 6, -6, 5, -8,
    -- filter=31 channel=68
    -5, 4, -2, 0, 0, -6, 0, 0, -7,
    -- filter=31 channel=69
    -7, 0, -6, 1, -2, 7, 2, -4, -4,
    -- filter=31 channel=70
    -13, -4, -4, -11, 0, 7, -17, 0, -6,
    -- filter=31 channel=71
    2, -11, -4, -1, -5, -3, -5, -6, 5,
    -- filter=31 channel=72
    4, 5, 6, 2, 9, 0, -5, -5, -2,
    -- filter=31 channel=73
    -9, 3, 0, -1, 10, 6, -7, 7, -5,
    -- filter=31 channel=74
    -3, 5, -5, 0, 7, -4, -4, 3, 1,
    -- filter=31 channel=75
    -14, -11, 3, -12, 9, 10, -4, 2, 11,
    -- filter=31 channel=76
    0, 9, 0, 2, 9, -12, 3, 4, -5,
    -- filter=31 channel=77
    -2, -5, -6, -6, -2, 2, 7, -1, 0,
    -- filter=31 channel=78
    3, -2, -6, 12, -1, 0, 7, 0, -5,
    -- filter=31 channel=79
    -26, 4, 5, -27, 24, 6, -20, 21, 9,
    -- filter=31 channel=80
    6, -2, 4, 15, 14, 6, -1, -12, -4,
    -- filter=31 channel=81
    4, 5, -2, -5, 2, 6, 4, -6, 1,
    -- filter=31 channel=82
    4, 4, -3, 6, 0, -4, 7, -5, -5,
    -- filter=31 channel=83
    7, 8, -4, 5, 2, -6, -2, 0, -5,
    -- filter=31 channel=84
    -4, 8, -4, -2, 4, 5, -12, 0, -5,
    -- filter=31 channel=85
    0, -5, 6, 5, -7, 6, 3, -4, -4,
    -- filter=31 channel=86
    -8, 3, -8, -8, 5, 0, -5, 0, -1,
    -- filter=31 channel=87
    -11, 1, 0, -10, 4, 1, -8, 5, 4,
    -- filter=31 channel=88
    13, 11, 1, -1, 1, -13, 3, -2, -7,
    -- filter=31 channel=89
    -11, -5, 4, -5, 2, -6, -14, 3, -4,
    -- filter=31 channel=90
    6, -6, -1, 7, -11, -7, -5, -12, -12,
    -- filter=31 channel=91
    0, 10, 6, -6, 15, -1, -12, -2, -3,
    -- filter=31 channel=92
    0, -5, -7, 1, -8, -5, -2, -6, -4,
    -- filter=31 channel=93
    2, 5, 2, 1, -4, 2, 0, -5, 5,
    -- filter=31 channel=94
    3, -3, 2, -5, -2, -5, 2, -6, 3,
    -- filter=31 channel=95
    -1, -4, -7, -7, 0, -3, 5, -3, -2,
    -- filter=31 channel=96
    -7, -4, -1, -9, 6, 1, -9, -3, 2,
    -- filter=31 channel=97
    -6, -6, -3, -2, -11, -1, -6, -1, 0,
    -- filter=31 channel=98
    0, 3, -1, -5, 21, 7, -1, 7, 6,
    -- filter=31 channel=99
    4, 0, 9, 5, 2, -10, -8, 2, -16,
    -- filter=31 channel=100
    -1, 0, 2, 2, 0, -7, 2, 0, -4,
    -- filter=31 channel=101
    -7, -7, -4, -10, -6, -6, -10, -9, -4,
    -- filter=31 channel=102
    2, -3, -7, -1, 2, 3, 6, 2, 6,
    -- filter=31 channel=103
    1, 0, 5, 17, -7, 3, 8, 4, 3,
    -- filter=31 channel=104
    19, -1, 6, 17, 4, -1, 10, -14, -11,
    -- filter=31 channel=105
    3, 4, 3, -2, 3, 1, 2, -2, 2,
    -- filter=31 channel=106
    -5, -4, 3, 3, 4, -3, 0, 3, 1,
    -- filter=31 channel=107
    -11, 2, 11, -11, 1, 5, -2, 0, -2,
    -- filter=31 channel=108
    -5, -8, 4, -6, 7, 0, -8, -6, 5,
    -- filter=31 channel=109
    -5, 11, 13, -11, 26, 2, -8, -3, -7,
    -- filter=31 channel=110
    6, -5, -2, 0, 4, -12, -1, -7, 0,
    -- filter=31 channel=111
    1, 4, -5, -8, -4, 0, -7, 3, 7,
    -- filter=31 channel=112
    -1, -2, -2, 0, 0, 7, 0, 2, 5,
    -- filter=31 channel=113
    -11, 1, -1, 3, -3, 8, -6, 10, -6,
    -- filter=31 channel=114
    -16, 2, 14, -25, 30, 22, -8, 18, 3,
    -- filter=31 channel=115
    -2, -5, 1, 1, -3, -3, 0, -2, -6,
    -- filter=31 channel=116
    4, 5, 2, 0, 4, 0, -5, 3, -6,
    -- filter=31 channel=117
    0, -5, 5, 0, -6, 3, 0, -5, 0,
    -- filter=31 channel=118
    5, 4, 7, 1, 2, -4, -1, 0, 0,
    -- filter=31 channel=119
    -13, 0, -2, 0, -12, -5, -11, 2, -11,
    -- filter=31 channel=120
    2, 16, 3, -9, 11, -5, -8, 5, -2,
    -- filter=31 channel=121
    -2, -4, -4, -10, 3, 4, -7, 2, 6,
    -- filter=31 channel=122
    11, -8, -13, 27, -5, -11, 6, -11, -10,
    -- filter=31 channel=123
    -13, -4, 4, -6, 0, 1, -8, -4, -6,
    -- filter=31 channel=124
    1, -5, 4, -6, -3, -5, 2, 2, -5,
    -- filter=31 channel=125
    7, 5, 8, 8, 4, -4, -2, 0, 0,
    -- filter=31 channel=126
    -16, -12, -1, -13, 4, 11, -11, 6, 3,
    -- filter=31 channel=127
    0, -4, 4, 0, 0, 3, -3, -3, -1,
    -- filter=32 channel=0
    -4, -4, -2, 1, -6, -11, -3, -2, 4,
    -- filter=32 channel=1
    3, -2, 2, -4, -2, -2, 9, 0, 7,
    -- filter=32 channel=2
    0, 0, 0, -4, 3, -2, 8, 0, -1,
    -- filter=32 channel=3
    -7, 1, 18, 4, 12, 3, 0, 0, 12,
    -- filter=32 channel=4
    0, 3, 3, 3, 4, 21, 10, 25, 13,
    -- filter=32 channel=5
    5, 3, -2, -3, 0, -9, -8, 1, -6,
    -- filter=32 channel=6
    0, -2, 2, 2, -8, -6, -1, 6, 5,
    -- filter=32 channel=7
    -4, -4, 0, 4, 0, -7, 1, -1, -6,
    -- filter=32 channel=8
    -1, 1, 0, 0, -3, 9, -4, 13, 4,
    -- filter=32 channel=9
    0, 8, -6, -3, -7, -3, -8, -3, 0,
    -- filter=32 channel=10
    7, 4, 2, -4, -2, -8, -5, -2, 11,
    -- filter=32 channel=11
    -3, -1, 1, -6, -10, -7, -8, 6, 7,
    -- filter=32 channel=12
    -1, 0, 4, -4, 0, -8, 5, 0, 0,
    -- filter=32 channel=13
    -6, 1, 9, 0, -7, -19, -7, 7, 12,
    -- filter=32 channel=14
    -4, -6, 4, 5, 5, -2, 0, -3, 3,
    -- filter=32 channel=15
    -6, -2, 2, -2, -2, -6, -6, -1, 5,
    -- filter=32 channel=16
    -2, 8, 9, 0, 3, -6, -1, 2, -5,
    -- filter=32 channel=17
    1, -2, 6, -5, -4, -3, 1, 1, 4,
    -- filter=32 channel=18
    7, 7, 8, 9, 0, -13, -9, 4, 13,
    -- filter=32 channel=19
    6, -2, 4, -3, 1, -1, 7, 3, -7,
    -- filter=32 channel=20
    -1, -5, -10, -6, 1, -4, 0, 6, 0,
    -- filter=32 channel=21
    1, 11, -2, -1, -11, -10, 5, -4, -5,
    -- filter=32 channel=22
    -3, 5, 5, -1, 6, -2, -4, -6, 7,
    -- filter=32 channel=23
    3, 14, 10, -1, -15, -17, -12, 1, 10,
    -- filter=32 channel=24
    -4, -4, -7, 5, -3, -6, -5, 7, 4,
    -- filter=32 channel=25
    8, 6, 3, -4, -15, -24, 3, 3, 17,
    -- filter=32 channel=26
    9, 7, -1, -5, 0, 5, 0, 4, -3,
    -- filter=32 channel=27
    4, 19, 4, -13, -18, -22, 1, 11, 23,
    -- filter=32 channel=28
    -6, 6, 7, 7, 5, 3, 6, 3, -4,
    -- filter=32 channel=29
    6, 1, -2, -5, -7, -10, 5, 9, 6,
    -- filter=32 channel=30
    11, 12, -5, -9, -15, -13, -3, 2, 10,
    -- filter=32 channel=31
    7, 13, 8, -4, -18, -19, -7, 1, 13,
    -- filter=32 channel=32
    0, 0, 3, -2, -12, -9, -4, 3, 16,
    -- filter=32 channel=33
    0, 2, 11, 8, -1, -10, 0, -3, 0,
    -- filter=32 channel=34
    -2, 3, -9, 2, -12, -5, -3, 10, 11,
    -- filter=32 channel=35
    -4, 0, 4, -1, 0, -3, 1, 0, 4,
    -- filter=32 channel=36
    8, 6, -6, -8, -6, -8, 1, 10, 3,
    -- filter=32 channel=37
    3, 6, -9, 2, -2, -2, 5, 0, 3,
    -- filter=32 channel=38
    4, 6, 10, 0, -4, -11, -3, 6, 9,
    -- filter=32 channel=39
    -5, 6, -6, 3, 1, 0, 1, 7, 5,
    -- filter=32 channel=40
    4, 7, 0, 0, 6, 5, -7, 2, 0,
    -- filter=32 channel=41
    7, -18, 4, 7, -7, -7, -8, -11, 9,
    -- filter=32 channel=42
    -3, 0, -5, -6, -8, 2, 0, -2, 8,
    -- filter=32 channel=43
    -5, 3, 3, 11, 4, -7, 1, 3, 7,
    -- filter=32 channel=44
    3, 2, -5, 2, -3, -9, 0, 8, 0,
    -- filter=32 channel=45
    0, 7, -2, -7, 6, 1, -4, 7, 3,
    -- filter=32 channel=46
    4, 3, 0, 2, 2, -4, 7, -2, 0,
    -- filter=32 channel=47
    3, 15, 0, 6, -10, -16, -10, -2, 0,
    -- filter=32 channel=48
    2, 8, 1, -12, -13, -17, -4, 10, 8,
    -- filter=32 channel=49
    8, 8, 1, -4, -3, 1, 5, 16, 6,
    -- filter=32 channel=50
    2, 12, 7, 2, -11, -6, -6, 8, 12,
    -- filter=32 channel=51
    2, 5, 0, -4, -5, -1, 0, 0, -5,
    -- filter=32 channel=52
    -2, 0, 2, -5, -6, -3, 3, 7, -4,
    -- filter=32 channel=53
    -4, 3, -7, -1, -7, -8, 0, -1, 5,
    -- filter=32 channel=54
    -3, 6, -3, 7, 3, 6, -1, 7, -1,
    -- filter=32 channel=55
    0, 8, 0, -5, -6, -4, -11, -7, 11,
    -- filter=32 channel=56
    -1, -3, 2, -9, -8, 9, 6, -3, 7,
    -- filter=32 channel=57
    7, 4, 0, -2, 4, 2, -2, 6, 9,
    -- filter=32 channel=58
    -5, 3, 1, 6, -5, -1, -4, 3, -5,
    -- filter=32 channel=59
    9, 9, 1, -1, -3, -21, -10, -9, 7,
    -- filter=32 channel=60
    -6, -6, 2, 1, -4, -1, 0, 3, -3,
    -- filter=32 channel=61
    7, -3, -3, -3, -10, 6, 1, 0, -8,
    -- filter=32 channel=62
    4, 3, 4, 6, -3, -2, 4, -4, 0,
    -- filter=32 channel=63
    1, 0, 0, 2, 1, -1, -7, -4, -3,
    -- filter=32 channel=64
    -5, -3, -6, 0, 0, -3, 0, 0, -5,
    -- filter=32 channel=65
    4, -6, 0, -5, 0, -3, 5, -7, 0,
    -- filter=32 channel=66
    0, -6, 8, -2, -6, -13, 0, -6, 4,
    -- filter=32 channel=67
    -7, 3, 3, -3, -4, -3, 3, -4, -6,
    -- filter=32 channel=68
    8, -5, -1, 2, 3, 1, -4, 6, -3,
    -- filter=32 channel=69
    2, 0, 6, 2, 3, 0, -4, -1, 5,
    -- filter=32 channel=70
    -1, 4, -1, -4, -5, 2, -8, 4, 14,
    -- filter=32 channel=71
    -4, -4, 5, 4, 12, 4, -3, 4, 6,
    -- filter=32 channel=72
    2, 13, 6, -5, -10, -21, -14, -7, 7,
    -- filter=32 channel=73
    7, 2, -4, 0, -12, -4, -5, 0, 9,
    -- filter=32 channel=74
    5, 8, -12, -4, -18, 3, -7, 5, 3,
    -- filter=32 channel=75
    -6, 2, 18, 1, 6, -10, -8, -12, 0,
    -- filter=32 channel=76
    -2, -1, 4, 2, 3, -3, -1, 5, 0,
    -- filter=32 channel=77
    -3, 1, 7, 0, -3, 4, 0, -2, 0,
    -- filter=32 channel=78
    -1, -1, -1, -7, -10, -6, -6, 3, 5,
    -- filter=32 channel=79
    -6, 13, 11, 1, -11, -17, -9, -1, 7,
    -- filter=32 channel=80
    10, 15, 5, -9, -8, -23, -12, -8, 1,
    -- filter=32 channel=81
    1, 3, -3, 7, 0, -5, -4, -5, -2,
    -- filter=32 channel=82
    0, -1, 6, -5, -1, -2, 2, -4, 0,
    -- filter=32 channel=83
    2, 2, -8, -9, -8, 3, 6, 6, 7,
    -- filter=32 channel=84
    5, -1, 0, -6, -4, -5, 0, 6, 0,
    -- filter=32 channel=85
    -4, -5, -6, 0, -3, -6, -6, -3, 0,
    -- filter=32 channel=86
    -4, 0, 1, -3, -7, -6, 6, 0, -6,
    -- filter=32 channel=87
    6, -2, -6, 1, 0, -4, -2, 1, 5,
    -- filter=32 channel=88
    4, 0, -1, 0, -3, -6, -6, -1, 10,
    -- filter=32 channel=89
    -3, 12, 13, 6, 1, -14, -5, 1, 17,
    -- filter=32 channel=90
    5, -1, 5, 3, -1, 6, -6, -6, 2,
    -- filter=32 channel=91
    -1, 10, -4, -11, -19, -7, 6, 11, 13,
    -- filter=32 channel=92
    -3, -2, -6, 6, -4, 2, -1, 4, 6,
    -- filter=32 channel=93
    5, 14, -5, -10, -4, 0, 7, 6, 10,
    -- filter=32 channel=94
    -5, 5, -1, -1, -2, -5, 0, -2, 2,
    -- filter=32 channel=95
    2, 7, 3, 5, -1, 6, -6, 4, 4,
    -- filter=32 channel=96
    -4, 1, 0, 0, 0, 0, 6, -7, 0,
    -- filter=32 channel=97
    -5, -5, 5, 4, 15, 6, 0, -4, 7,
    -- filter=32 channel=98
    6, 7, 12, -8, -15, -14, -2, 0, 17,
    -- filter=32 channel=99
    4, 5, 6, 1, -17, -13, -11, 0, 9,
    -- filter=32 channel=100
    3, -8, -3, 4, 0, 2, -8, 0, 4,
    -- filter=32 channel=101
    0, 3, 1, 0, 7, 15, 0, 8, 11,
    -- filter=32 channel=102
    -4, -7, -5, -5, -6, 6, 4, -5, 5,
    -- filter=32 channel=103
    -4, 12, 6, 1, 2, -13, -8, -2, 2,
    -- filter=32 channel=104
    7, 12, 0, -3, -14, -9, -2, 0, -5,
    -- filter=32 channel=105
    -2, -3, -1, 0, -6, -1, 0, -4, 3,
    -- filter=32 channel=106
    0, -2, -2, 6, -3, -2, -7, 3, 5,
    -- filter=32 channel=107
    2, 1, -4, -2, 5, 1, 2, 0, 9,
    -- filter=32 channel=108
    6, -8, 4, -3, 2, -1, -7, -5, 3,
    -- filter=32 channel=109
    3, 2, -1, -5, -21, -21, -5, 8, 13,
    -- filter=32 channel=110
    6, 8, -1, 3, 2, -8, 0, 2, -1,
    -- filter=32 channel=111
    2, -5, -3, -3, 5, 6, 1, -3, 5,
    -- filter=32 channel=112
    -4, 5, 2, 3, -2, -1, -5, 8, 10,
    -- filter=32 channel=113
    4, 3, 7, -2, -1, -9, -6, 0, 0,
    -- filter=32 channel=114
    7, 17, -3, -1, -14, -19, 7, 8, 5,
    -- filter=32 channel=115
    4, 4, -7, -5, -2, 2, -6, -1, 5,
    -- filter=32 channel=116
    1, 7, -4, -12, -15, -20, -6, 4, 12,
    -- filter=32 channel=117
    -1, 9, 1, -3, -5, -8, 2, 6, 2,
    -- filter=32 channel=118
    0, 4, -1, 0, 0, 3, -1, -1, 4,
    -- filter=32 channel=119
    0, 1, -3, -4, -15, 0, 4, -3, -3,
    -- filter=32 channel=120
    2, 6, -3, -7, -29, -5, 3, 10, 11,
    -- filter=32 channel=121
    0, -4, 6, -3, 3, 0, 3, -7, 2,
    -- filter=32 channel=122
    5, 8, 1, 6, -10, -7, -1, 1, 10,
    -- filter=32 channel=123
    5, 5, -6, -4, -7, 7, -1, 5, 7,
    -- filter=32 channel=124
    -7, 7, -3, 8, 6, -4, 3, 5, -5,
    -- filter=32 channel=125
    4, 15, -9, -10, -22, -20, -13, -3, 8,
    -- filter=32 channel=126
    -2, 0, 10, 2, 5, -13, 0, 0, 5,
    -- filter=32 channel=127
    0, -7, 6, 0, 2, -9, 1, 4, 5,
    -- filter=33 channel=0
    -5, 2, 14, -7, 11, 3, -8, 6, 5,
    -- filter=33 channel=1
    -3, 10, 5, -6, 3, 10, -5, 13, 0,
    -- filter=33 channel=2
    -3, 0, 4, 7, -2, 4, -5, -3, 1,
    -- filter=33 channel=3
    2, 7, 1, 5, -6, 6, 12, 9, 6,
    -- filter=33 channel=4
    2, 2, -2, -2, 2, -6, 1, -1, -3,
    -- filter=33 channel=5
    0, 2, 5, -2, 1, 2, 2, 10, 6,
    -- filter=33 channel=6
    -4, -2, 4, -4, -1, 0, -4, 9, 1,
    -- filter=33 channel=7
    5, 6, 3, -3, -2, 1, 6, 4, -5,
    -- filter=33 channel=8
    0, 4, -1, 7, -7, -7, 6, 1, 0,
    -- filter=33 channel=9
    6, 1, -5, -6, -5, -2, -5, -8, -5,
    -- filter=33 channel=10
    -4, -8, -10, 5, 0, -3, 5, 4, -13,
    -- filter=33 channel=11
    -2, 4, -8, -3, 9, 0, -1, -4, 1,
    -- filter=33 channel=12
    -4, 2, -3, 3, 1, 5, 3, 0, -3,
    -- filter=33 channel=13
    5, 6, -9, 9, 13, -3, 2, 2, -14,
    -- filter=33 channel=14
    -3, 0, 5, 5, 0, 4, 0, 2, 5,
    -- filter=33 channel=15
    5, -5, 0, 2, -1, -17, 1, 9, -20,
    -- filter=33 channel=16
    0, -5, 1, 0, -4, 1, -5, -4, -1,
    -- filter=33 channel=17
    4, 6, 2, -4, -3, 1, -4, 3, -5,
    -- filter=33 channel=18
    2, 1, 5, -6, 13, -7, -3, 3, -15,
    -- filter=33 channel=19
    4, -6, 2, -5, 6, 4, 2, -1, 4,
    -- filter=33 channel=20
    10, -6, 0, 3, 0, -7, 9, 5, 0,
    -- filter=33 channel=21
    6, -8, -5, -4, -1, -5, 3, -5, -5,
    -- filter=33 channel=22
    2, -3, -5, 0, 3, -5, 7, -1, 1,
    -- filter=33 channel=23
    5, -13, -5, 11, -10, -17, 17, -3, -31,
    -- filter=33 channel=24
    5, 3, -5, 0, 0, 0, 4, -1, 0,
    -- filter=33 channel=25
    7, -3, -12, 7, 0, -18, -2, -4, -20,
    -- filter=33 channel=26
    -4, 4, 1, 5, 3, 8, -1, 4, 3,
    -- filter=33 channel=27
    -1, -13, -12, 11, -17, -36, 5, -16, -29,
    -- filter=33 channel=28
    -1, 2, -4, 3, 1, -6, 1, 6, -6,
    -- filter=33 channel=29
    3, -4, -3, 0, 12, -10, 8, 2, -7,
    -- filter=33 channel=30
    -2, -2, -2, -6, -4, -10, -5, -6, -15,
    -- filter=33 channel=31
    6, -7, -16, 16, -10, -24, 11, -6, -15,
    -- filter=33 channel=32
    -3, 1, -8, 8, 10, -16, 8, 1, -15,
    -- filter=33 channel=33
    -8, -7, 1, -3, -6, -9, -1, 0, -22,
    -- filter=33 channel=34
    -5, -4, 1, 2, -4, 0, -1, 3, -6,
    -- filter=33 channel=35
    3, -4, -6, 0, 5, 0, 1, 4, 5,
    -- filter=33 channel=36
    1, 1, 2, 8, 6, -6, 8, -7, -6,
    -- filter=33 channel=37
    3, 7, 2, -1, -6, 0, -3, -3, -4,
    -- filter=33 channel=38
    5, -4, -7, 1, -5, -6, -2, -8, -15,
    -- filter=33 channel=39
    0, 5, 0, 6, 3, 3, 0, -3, -4,
    -- filter=33 channel=40
    0, -2, 3, -1, 7, -10, 5, 7, -2,
    -- filter=33 channel=41
    4, 15, 12, 12, 28, 22, 7, 19, 17,
    -- filter=33 channel=42
    3, -1, -4, 3, 0, -9, 0, 4, -5,
    -- filter=33 channel=43
    -6, 2, 14, 6, 7, 9, 8, 9, 6,
    -- filter=33 channel=44
    4, 0, 1, -6, -1, -13, -6, -8, -9,
    -- filter=33 channel=45
    1, 4, 1, 6, -5, -3, 4, 2, 8,
    -- filter=33 channel=46
    4, 2, 3, -2, 3, -1, 0, 6, 4,
    -- filter=33 channel=47
    -5, -1, -13, -1, -8, -12, -4, -5, -9,
    -- filter=33 channel=48
    0, -10, -6, -3, -4, -18, 3, -12, -14,
    -- filter=33 channel=49
    0, -3, -9, 8, 7, -6, 2, 4, -10,
    -- filter=33 channel=50
    5, -4, -7, -3, -10, -17, -2, -13, -23,
    -- filter=33 channel=51
    4, -6, -7, -3, 6, -5, -6, -1, -7,
    -- filter=33 channel=52
    4, 3, -6, -2, -3, -4, 7, -2, 2,
    -- filter=33 channel=53
    3, -2, -4, -4, 5, -11, 0, -4, -12,
    -- filter=33 channel=54
    3, 1, 0, -1, 3, 6, 6, -6, 5,
    -- filter=33 channel=55
    1, 0, 0, -1, 3, -11, 7, 5, -10,
    -- filter=33 channel=56
    0, 2, 4, 1, 0, -7, 6, 6, -7,
    -- filter=33 channel=57
    4, 9, 1, 2, 0, 6, 0, 9, 1,
    -- filter=33 channel=58
    3, 0, 10, 3, -2, 10, -2, 5, 11,
    -- filter=33 channel=59
    6, 2, -18, 9, 2, -23, 7, -1, -13,
    -- filter=33 channel=60
    0, 0, 4, 6, -1, 5, -2, -4, 2,
    -- filter=33 channel=61
    -2, 2, -2, -5, -5, -4, 1, 3, -5,
    -- filter=33 channel=62
    -6, -4, 3, 0, 2, 0, 2, 7, -7,
    -- filter=33 channel=63
    -4, 0, -2, 4, 5, 13, 5, 1, 12,
    -- filter=33 channel=64
    6, -6, -7, -4, 8, 0, 6, 5, -6,
    -- filter=33 channel=65
    0, 1, 0, 0, -2, 2, 3, -1, 6,
    -- filter=33 channel=66
    3, -1, 2, 8, 5, 11, 2, 6, 10,
    -- filter=33 channel=67
    -6, -7, 1, -3, 2, 0, 0, 7, 2,
    -- filter=33 channel=68
    4, -4, 0, 7, 0, 2, -1, 4, -4,
    -- filter=33 channel=69
    -3, -3, 0, 4, 0, -2, 1, 1, 7,
    -- filter=33 channel=70
    5, -8, -10, 9, -4, -27, -5, -16, -14,
    -- filter=33 channel=71
    -8, -1, 8, -6, -5, -4, -2, 5, -4,
    -- filter=33 channel=72
    7, 1, -11, 6, 4, -13, 9, -2, -14,
    -- filter=33 channel=73
    -3, -1, -1, -2, 1, -17, 4, -9, -5,
    -- filter=33 channel=74
    -5, -6, 0, 8, -6, -9, 0, -9, -16,
    -- filter=33 channel=75
    -12, -3, 11, 0, 14, 7, 5, 16, 4,
    -- filter=33 channel=76
    9, 6, 2, 1, 15, 1, 2, 15, 5,
    -- filter=33 channel=77
    0, -4, 0, -6, 5, 1, 0, 2, 2,
    -- filter=33 channel=78
    -7, 2, -6, 6, 0, 5, 1, -4, 0,
    -- filter=33 channel=79
    5, 0, -4, 0, 11, -8, 5, 15, -16,
    -- filter=33 channel=80
    9, 0, -17, 0, -3, -16, 6, -7, -24,
    -- filter=33 channel=81
    5, 1, 1, -7, -3, 6, -4, -2, 6,
    -- filter=33 channel=82
    6, -6, -3, 4, 1, 4, 7, -4, -1,
    -- filter=33 channel=83
    4, -9, -9, 6, 3, -10, -4, 1, -9,
    -- filter=33 channel=84
    0, -1, -2, 8, 5, -1, 4, -1, -2,
    -- filter=33 channel=85
    7, 6, -5, 0, -3, 3, -7, 2, -6,
    -- filter=33 channel=86
    -3, 2, 4, 7, -1, 5, 5, 1, -1,
    -- filter=33 channel=87
    0, -4, -4, 8, -5, 1, 3, 2, 5,
    -- filter=33 channel=88
    6, 6, 0, -2, 0, -5, 4, 1, -6,
    -- filter=33 channel=89
    -2, -4, 0, -2, 0, -21, 9, 9, -18,
    -- filter=33 channel=90
    0, -8, -3, 0, -6, 0, 8, -8, 3,
    -- filter=33 channel=91
    7, -10, -14, 2, -8, -24, 4, -1, -17,
    -- filter=33 channel=92
    -7, -2, 6, -6, 0, -3, 1, -2, 5,
    -- filter=33 channel=93
    3, 6, 0, -4, -4, -8, -8, -2, -12,
    -- filter=33 channel=94
    -1, 5, 0, 7, -1, -5, -2, 4, 7,
    -- filter=33 channel=95
    -3, 5, -2, 0, 7, 0, 5, -3, -7,
    -- filter=33 channel=96
    -6, 0, 1, -6, 0, 3, -2, 4, 2,
    -- filter=33 channel=97
    1, 3, 2, -4, -4, -5, 0, 7, 5,
    -- filter=33 channel=98
    -7, -5, -8, 8, -6, -23, 9, -5, -23,
    -- filter=33 channel=99
    8, -8, -13, 16, -13, -12, 9, -10, -26,
    -- filter=33 channel=100
    -1, -3, -3, 6, -1, 0, 7, 3, -1,
    -- filter=33 channel=101
    6, -5, 0, 7, 0, -9, -1, -4, 7,
    -- filter=33 channel=102
    4, 0, 6, 0, 0, 2, 4, 3, -5,
    -- filter=33 channel=103
    -13, -14, -4, -9, -3, -15, 1, -9, -11,
    -- filter=33 channel=104
    8, -9, -12, 13, -8, -16, -5, -10, -20,
    -- filter=33 channel=105
    6, -2, 3, -2, 0, 6, 11, 4, 1,
    -- filter=33 channel=106
    -2, 5, 6, -3, 3, 5, 3, 5, 1,
    -- filter=33 channel=107
    1, 1, 4, 11, -3, 4, 2, 7, 0,
    -- filter=33 channel=108
    2, 0, 12, -1, 16, 16, 3, 8, 1,
    -- filter=33 channel=109
    6, -3, -13, 11, -1, -20, 2, -12, -30,
    -- filter=33 channel=110
    5, -2, 2, 10, -4, 1, 5, -7, -2,
    -- filter=33 channel=111
    -4, 9, 1, 6, -2, 10, 2, 1, 7,
    -- filter=33 channel=112
    -2, -9, -10, -4, -7, -5, -2, -10, -4,
    -- filter=33 channel=113
    0, -5, 1, -1, 0, -8, 8, -6, -7,
    -- filter=33 channel=114
    1, 5, -3, -2, 12, -2, -4, 14, -1,
    -- filter=33 channel=115
    5, 1, 6, -1, 0, -3, 4, 0, 3,
    -- filter=33 channel=116
    5, -1, -15, 10, -5, -21, 0, 4, -13,
    -- filter=33 channel=117
    1, 1, -4, 0, 1, 1, 4, 0, -7,
    -- filter=33 channel=118
    5, 4, -5, 0, -1, -1, -3, -6, 5,
    -- filter=33 channel=119
    -8, -7, 3, 3, -8, -2, 4, -2, -4,
    -- filter=33 channel=120
    14, -6, -15, 9, -4, -22, 10, -7, -24,
    -- filter=33 channel=121
    0, 5, -6, 0, 6, 2, 1, 3, 2,
    -- filter=33 channel=122
    -3, -5, -13, 3, -8, -22, -1, -18, -18,
    -- filter=33 channel=123
    -3, -6, 5, 4, 2, 2, 5, -6, -2,
    -- filter=33 channel=124
    2, 6, 9, 7, -2, 0, 4, 0, -7,
    -- filter=33 channel=125
    9, -4, -6, 1, 5, -17, 0, -1, -25,
    -- filter=33 channel=126
    2, 4, 7, -6, 8, 7, 8, 15, 0,
    -- filter=33 channel=127
    0, 4, 0, 2, -3, 1, 4, 1, 0,
    -- filter=34 channel=0
    -5, -1, -10, 4, -7, -9, 1, 0, -1,
    -- filter=34 channel=1
    5, -12, -3, -4, -11, -8, 1, 3, -8,
    -- filter=34 channel=2
    -1, 1, 4, 6, 5, 3, -7, 4, 5,
    -- filter=34 channel=3
    -5, -3, -4, -10, -7, -5, 5, 1, 4,
    -- filter=34 channel=4
    6, -7, 0, -4, 0, 5, -7, -2, 2,
    -- filter=34 channel=5
    6, -2, -8, 3, 5, -1, 4, 6, -6,
    -- filter=34 channel=6
    1, 0, 0, -4, 0, -4, -2, -3, 5,
    -- filter=34 channel=7
    2, 0, -2, -5, 0, 1, -5, -2, 1,
    -- filter=34 channel=8
    0, 5, 0, 3, 0, -5, -7, 7, -4,
    -- filter=34 channel=9
    -4, 7, 2, 2, 4, -1, -1, 4, 7,
    -- filter=34 channel=10
    -1, 0, 7, 2, 5, -1, -4, 7, 0,
    -- filter=34 channel=11
    3, -7, -3, 6, -5, -4, -5, -4, 1,
    -- filter=34 channel=12
    5, -2, 0, 3, -6, 5, 6, 6, -4,
    -- filter=34 channel=13
    -2, -11, 0, 1, 0, -1, 0, -8, 3,
    -- filter=34 channel=14
    -2, 7, -6, -6, -5, 4, 0, -1, 4,
    -- filter=34 channel=15
    0, -4, 2, 0, -7, -9, 0, 1, -2,
    -- filter=34 channel=16
    -2, 3, -1, -1, 8, 0, 1, 0, 0,
    -- filter=34 channel=17
    -3, 3, 5, -1, -4, -2, 1, 1, -1,
    -- filter=34 channel=18
    -5, 0, -8, -6, -9, -9, -3, -11, -1,
    -- filter=34 channel=19
    1, 5, -1, -5, 0, 1, -2, 1, -2,
    -- filter=34 channel=20
    4, -6, 2, -2, -1, 3, -5, -1, -2,
    -- filter=34 channel=21
    2, 1, 6, -3, 3, 3, -2, 3, 1,
    -- filter=34 channel=22
    -9, -10, 0, 3, -10, -3, -1, -1, 1,
    -- filter=34 channel=23
    -13, -8, -8, -1, -13, 0, -2, -7, -3,
    -- filter=34 channel=24
    1, -5, -6, 1, 7, 6, -3, 0, 6,
    -- filter=34 channel=25
    -8, -2, -2, -3, 4, 4, -4, -6, 9,
    -- filter=34 channel=26
    2, 0, -3, -3, 10, 10, -6, 0, 5,
    -- filter=34 channel=27
    -12, -11, -10, 1, -8, -4, 4, -3, -2,
    -- filter=34 channel=28
    -5, -3, -5, 4, -5, 0, 0, 5, -2,
    -- filter=34 channel=29
    0, 0, -7, 2, 2, 5, 8, 0, -8,
    -- filter=34 channel=30
    5, 4, -3, 7, 6, 0, 4, -1, 4,
    -- filter=34 channel=31
    -5, 1, 4, -9, 8, -2, -2, -2, 11,
    -- filter=34 channel=32
    -6, -3, -1, -3, -1, -4, 4, -1, -8,
    -- filter=34 channel=33
    -1, -13, -5, -5, 0, -3, 3, -8, -6,
    -- filter=34 channel=34
    -3, 3, 7, -6, -6, -1, -3, 1, 0,
    -- filter=34 channel=35
    -2, 6, 6, 0, -3, -4, -1, 6, -1,
    -- filter=34 channel=36
    4, 2, -1, 5, 7, -3, 1, -9, 0,
    -- filter=34 channel=37
    -9, -2, -6, -3, -3, -5, -3, -2, 4,
    -- filter=34 channel=38
    -9, 4, -1, 3, -5, -6, 1, 4, -3,
    -- filter=34 channel=39
    -4, -6, 1, 0, 6, 3, 6, 3, 2,
    -- filter=34 channel=40
    -5, 0, -5, -3, -8, -7, -3, 1, 2,
    -- filter=34 channel=41
    -1, 10, -2, 0, 3, -2, 6, 3, 4,
    -- filter=34 channel=42
    -1, -4, -4, 5, 7, -4, -2, -3, 0,
    -- filter=34 channel=43
    -5, -8, -6, -6, 1, -1, -1, -4, 0,
    -- filter=34 channel=44
    -6, -1, 2, 3, 5, 1, 0, 8, 5,
    -- filter=34 channel=45
    -8, 3, -6, 1, 0, 0, -6, -6, -4,
    -- filter=34 channel=46
    -1, -4, 3, -4, 0, 0, -7, -1, 0,
    -- filter=34 channel=47
    -7, 0, -2, 7, 5, 5, 1, 5, 12,
    -- filter=34 channel=48
    3, -3, 2, -4, 11, 5, -3, 2, 5,
    -- filter=34 channel=49
    1, -3, 2, -3, -6, 4, 3, 1, -6,
    -- filter=34 channel=50
    -3, -1, -2, 2, 0, -6, -4, -4, -1,
    -- filter=34 channel=51
    5, -5, 5, -7, -4, -4, -2, 6, 3,
    -- filter=34 channel=52
    0, 4, 2, -6, 2, -1, 4, -7, -3,
    -- filter=34 channel=53
    -4, -7, 2, 0, -2, 3, 4, -4, -4,
    -- filter=34 channel=54
    -1, 3, -7, -3, -6, 0, -1, -3, -2,
    -- filter=34 channel=55
    -4, -11, -12, -3, -1, 0, -2, -8, -3,
    -- filter=34 channel=56
    3, 3, 1, 8, 0, -4, -5, -4, -1,
    -- filter=34 channel=57
    -4, 7, 7, -6, 4, -3, -5, 0, 2,
    -- filter=34 channel=58
    -5, 1, 5, 5, -3, -7, -6, 8, 1,
    -- filter=34 channel=59
    0, 1, -7, 1, -2, -5, 3, -3, 1,
    -- filter=34 channel=60
    6, 0, 1, -4, -3, 0, -6, 6, 5,
    -- filter=34 channel=61
    3, -4, 7, 1, 7, 6, -4, 7, 0,
    -- filter=34 channel=62
    -2, 6, 4, -7, 0, 5, -2, 4, -3,
    -- filter=34 channel=63
    -3, 9, 6, 5, 3, 3, -3, 5, 1,
    -- filter=34 channel=64
    -7, -1, 0, 1, 3, 1, 3, -7, -3,
    -- filter=34 channel=65
    -6, 5, -4, 3, 2, -5, -2, -6, 2,
    -- filter=34 channel=66
    4, -3, -6, 10, -7, 6, 4, 1, -3,
    -- filter=34 channel=67
    1, -5, 5, 4, 4, 5, -4, 0, -2,
    -- filter=34 channel=68
    0, 6, 0, -3, -5, -2, -5, -5, 1,
    -- filter=34 channel=69
    5, 0, 6, 0, 1, 2, -4, -1, 1,
    -- filter=34 channel=70
    -9, -8, 3, -10, -13, 0, -8, 0, 0,
    -- filter=34 channel=71
    3, -8, 6, -2, 5, 4, -1, 5, -6,
    -- filter=34 channel=72
    -1, -7, -8, -5, 9, -2, -4, -6, -2,
    -- filter=34 channel=73
    -9, 1, -1, 5, -2, 4, -4, 3, -5,
    -- filter=34 channel=74
    -1, -1, 4, 4, 2, -1, -8, 1, 1,
    -- filter=34 channel=75
    -1, -5, 0, -6, -1, -5, 4, -3, 0,
    -- filter=34 channel=76
    -5, -5, 4, 3, 0, -4, -6, -5, 3,
    -- filter=34 channel=77
    0, -2, -1, -5, 0, 7, 5, -2, 1,
    -- filter=34 channel=78
    -2, 4, 1, 1, 3, 0, -6, 4, 0,
    -- filter=34 channel=79
    -6, -2, -10, -3, -19, -15, 4, -8, -7,
    -- filter=34 channel=80
    4, 8, -7, 3, 11, 5, 4, 12, 10,
    -- filter=34 channel=81
    2, 1, -3, 7, 6, 0, 4, 6, 4,
    -- filter=34 channel=82
    6, 5, 0, -2, 2, 0, -4, 4, 3,
    -- filter=34 channel=83
    7, -2, 6, -6, 2, -3, -8, 3, 6,
    -- filter=34 channel=84
    -8, 0, 2, 1, 3, 1, 2, 0, 1,
    -- filter=34 channel=85
    -2, -2, -3, -6, -1, 6, -1, -2, -3,
    -- filter=34 channel=86
    4, 2, 4, -7, -5, 0, -7, -3, 0,
    -- filter=34 channel=87
    5, -1, -2, -2, -3, -3, 0, 0, 0,
    -- filter=34 channel=88
    -10, -2, -4, -1, 8, -3, -7, -3, 3,
    -- filter=34 channel=89
    -10, -6, -1, -1, -9, -4, -2, -9, 1,
    -- filter=34 channel=90
    -2, 0, 2, -9, 2, 0, -10, 6, 3,
    -- filter=34 channel=91
    0, 0, -8, -10, -6, -4, -9, 3, -6,
    -- filter=34 channel=92
    0, -1, -2, 0, 3, -7, 0, 0, -3,
    -- filter=34 channel=93
    4, 3, -5, 3, 6, 11, 0, 4, 12,
    -- filter=34 channel=94
    5, -1, 0, 6, -7, 1, -3, 0, -5,
    -- filter=34 channel=95
    -2, 0, 0, -2, 0, 4, 8, 5, -4,
    -- filter=34 channel=96
    0, -3, -7, 6, -7, -3, -7, 4, -5,
    -- filter=34 channel=97
    5, 5, 3, 3, -5, -8, 0, -4, 2,
    -- filter=34 channel=98
    0, -3, -7, 4, 0, -4, 3, 8, 2,
    -- filter=34 channel=99
    -1, 3, 4, 1, -3, 5, 2, 0, 0,
    -- filter=34 channel=100
    -4, 6, 7, -5, 8, 4, -6, 1, -3,
    -- filter=34 channel=101
    -2, 1, 1, 0, -3, 3, 4, 6, 0,
    -- filter=34 channel=102
    4, 4, 6, -5, 5, -6, -4, -2, 4,
    -- filter=34 channel=103
    4, -1, -5, -3, 10, 10, 1, 8, 11,
    -- filter=34 channel=104
    1, 7, 6, 0, 6, 10, -3, 6, 3,
    -- filter=34 channel=105
    -2, -2, 3, 5, 7, 0, 7, 0, 1,
    -- filter=34 channel=106
    -4, 0, 5, -3, 6, -1, -7, -7, -1,
    -- filter=34 channel=107
    -2, -6, 0, -6, -5, -10, -8, -8, -3,
    -- filter=34 channel=108
    -3, -6, -6, -5, 7, 1, -5, 0, 7,
    -- filter=34 channel=109
    1, 0, -1, -4, -2, 5, 5, -2, 5,
    -- filter=34 channel=110
    -7, -1, 1, 0, 7, 6, -6, 5, 6,
    -- filter=34 channel=111
    -2, 1, 4, 6, 0, -6, 0, -5, 5,
    -- filter=34 channel=112
    -6, 0, 1, -5, -4, 3, 0, -4, -3,
    -- filter=34 channel=113
    -6, 1, -8, -1, 3, 0, -4, 3, 1,
    -- filter=34 channel=114
    1, -9, -17, -6, -8, -16, 1, -2, -11,
    -- filter=34 channel=115
    1, 0, 7, -1, -3, 3, 1, -3, -1,
    -- filter=34 channel=116
    3, -4, -6, 5, 2, 0, -1, 4, 7,
    -- filter=34 channel=117
    1, -4, 4, -6, 0, -6, 3, 1, -7,
    -- filter=34 channel=118
    0, 1, -2, 4, -5, -1, -4, 0, -6,
    -- filter=34 channel=119
    3, -1, 4, 0, -3, -2, 0, 3, 5,
    -- filter=34 channel=120
    -2, -3, -6, -3, -10, -1, 0, -7, -4,
    -- filter=34 channel=121
    -6, 0, -6, 1, 4, 5, -5, -3, -5,
    -- filter=34 channel=122
    -1, 13, -4, -4, 12, 17, -7, 1, 14,
    -- filter=34 channel=123
    3, 2, 2, 0, 6, 2, 0, -2, 0,
    -- filter=34 channel=124
    0, 0, -5, -1, 0, -5, 1, -4, 2,
    -- filter=34 channel=125
    -2, 2, 0, 4, 4, -1, 2, 7, 8,
    -- filter=34 channel=126
    0, -7, -8, 5, 3, -3, 5, 0, -3,
    -- filter=34 channel=127
    -1, 0, 0, 7, 2, 7, 2, -5, -1,
    -- filter=35 channel=0
    8, 7, 7, 1, -1, 2, 6, 3, 2,
    -- filter=35 channel=1
    0, -2, 3, 0, -3, 3, -5, -5, -4,
    -- filter=35 channel=2
    -4, 0, -4, 2, 4, 5, 4, -3, 2,
    -- filter=35 channel=3
    2, -1, 0, -7, 3, -3, -3, -2, -4,
    -- filter=35 channel=4
    -1, 0, -6, 6, -1, 4, 0, 0, 3,
    -- filter=35 channel=5
    -3, -3, -4, 6, 5, -5, -2, 6, -4,
    -- filter=35 channel=6
    -7, 1, 6, -4, 5, 2, -2, -6, -2,
    -- filter=35 channel=7
    -6, -6, 0, -2, 1, -7, -1, -6, -1,
    -- filter=35 channel=8
    0, 3, -2, 4, 0, 4, 6, 1, 4,
    -- filter=35 channel=9
    -1, -1, 0, 2, -6, -2, -1, 2, -3,
    -- filter=35 channel=10
    2, -3, -2, 3, 4, -2, -7, 0, -2,
    -- filter=35 channel=11
    0, 1, -5, 2, -2, -4, -1, -7, 8,
    -- filter=35 channel=12
    -3, -2, 0, -5, 2, 6, 1, 2, 6,
    -- filter=35 channel=13
    6, 5, 0, -5, -7, 5, 3, -5, 0,
    -- filter=35 channel=14
    -2, 0, 6, 1, 4, -3, 4, -7, 3,
    -- filter=35 channel=15
    3, 7, 7, -5, -4, 1, 3, -5, -2,
    -- filter=35 channel=16
    7, -5, -1, 3, 5, -2, -5, 0, 5,
    -- filter=35 channel=17
    -4, -4, -4, -1, -2, -3, -5, -4, -3,
    -- filter=35 channel=18
    -4, -5, -6, -3, -9, -4, -5, -4, 3,
    -- filter=35 channel=19
    0, 4, -6, -2, -6, 5, 6, 2, 4,
    -- filter=35 channel=20
    0, 5, 0, 6, 3, 0, -3, -6, 1,
    -- filter=35 channel=21
    -2, -1, -5, 0, 2, -5, 3, -3, 4,
    -- filter=35 channel=22
    -5, 1, 1, -5, -1, 1, 6, -4, 3,
    -- filter=35 channel=23
    -5, -2, -2, -1, 4, -3, -5, 0, 1,
    -- filter=35 channel=24
    -4, -2, -2, 4, 3, -2, 5, -3, -4,
    -- filter=35 channel=25
    0, 0, -5, 0, 4, -7, 5, 4, -5,
    -- filter=35 channel=26
    -5, 5, 1, 0, -6, 0, 3, 0, 6,
    -- filter=35 channel=27
    -3, 0, -2, -6, -3, -1, -1, -3, 0,
    -- filter=35 channel=28
    6, 6, 2, -3, 3, 5, -3, -7, 0,
    -- filter=35 channel=29
    0, -2, -4, 3, 6, 7, 0, 3, 5,
    -- filter=35 channel=30
    0, 3, -2, 0, -3, 2, -7, 0, 5,
    -- filter=35 channel=31
    7, 0, 3, 0, -2, 1, 3, 6, -7,
    -- filter=35 channel=32
    0, 3, 5, 0, 3, 2, 2, -1, -6,
    -- filter=35 channel=33
    4, 1, -3, -3, 2, -2, 2, 0, -5,
    -- filter=35 channel=34
    -3, -1, 3, -3, 0, 0, -4, 5, -3,
    -- filter=35 channel=35
    -1, 0, -5, 1, -5, -6, 0, -3, 2,
    -- filter=35 channel=36
    0, 8, 3, -5, 8, 7, 5, 3, -5,
    -- filter=35 channel=37
    -2, 0, 6, 0, 1, 0, -1, 2, 3,
    -- filter=35 channel=38
    -5, 7, 0, -5, -7, 2, 4, 4, 0,
    -- filter=35 channel=39
    -4, 3, -4, -6, 5, 7, -3, 1, 0,
    -- filter=35 channel=40
    5, -1, 9, -2, -2, 5, 4, 0, 5,
    -- filter=35 channel=41
    -5, 7, 5, -1, 3, 3, 2, -7, 7,
    -- filter=35 channel=42
    4, 7, 2, -7, 5, 3, 5, 1, 0,
    -- filter=35 channel=43
    1, 5, -2, 0, 0, 1, -6, -7, 5,
    -- filter=35 channel=44
    4, -1, -3, -5, 0, -3, 0, 1, 2,
    -- filter=35 channel=45
    1, 5, 6, -5, 8, 7, -1, 6, -4,
    -- filter=35 channel=46
    -6, -2, 7, 7, 0, 4, 4, 0, 5,
    -- filter=35 channel=47
    1, -7, -1, 0, -4, -6, 0, 4, -1,
    -- filter=35 channel=48
    0, -3, -6, -7, -6, -1, 2, 4, -2,
    -- filter=35 channel=49
    5, 5, 1, 3, 3, 1, -3, -2, 0,
    -- filter=35 channel=50
    7, 6, -5, -2, 6, -4, 1, 5, -6,
    -- filter=35 channel=51
    -1, 4, 1, 0, 3, 6, -6, 1, 5,
    -- filter=35 channel=52
    0, 3, 6, -4, 7, 3, 6, -2, 3,
    -- filter=35 channel=53
    6, 0, -7, 0, 5, 6, 6, -1, 0,
    -- filter=35 channel=54
    -6, 5, 6, 0, 4, -1, -3, -4, 3,
    -- filter=35 channel=55
    4, 0, -2, 3, -1, 3, 2, -3, 0,
    -- filter=35 channel=56
    1, -7, 3, 4, -4, -3, 2, 3, 0,
    -- filter=35 channel=57
    -1, -7, -3, -7, 4, 8, -2, -2, -1,
    -- filter=35 channel=58
    2, 2, 0, -6, 5, -4, -2, -2, 4,
    -- filter=35 channel=59
    -5, 0, 5, -4, 0, 1, -4, 2, 2,
    -- filter=35 channel=60
    6, -4, -1, 2, -3, 3, -4, -1, 4,
    -- filter=35 channel=61
    5, -2, 2, 4, 1, -4, 0, 7, 0,
    -- filter=35 channel=62
    3, 2, -5, -7, 5, -1, 5, -5, -6,
    -- filter=35 channel=63
    2, -4, 5, 3, -6, -5, -5, 4, 4,
    -- filter=35 channel=64
    3, 2, 0, 5, -5, 1, 0, -4, 0,
    -- filter=35 channel=65
    -6, 3, -5, -4, -5, -3, 3, -5, -4,
    -- filter=35 channel=66
    -1, 5, 6, -2, 6, -6, 1, 0, -1,
    -- filter=35 channel=67
    -6, 0, -7, 7, 5, -4, -1, 0, -6,
    -- filter=35 channel=68
    -5, 4, 5, -4, 3, 0, -3, -4, -4,
    -- filter=35 channel=69
    1, -5, 3, 1, -6, 2, 4, -1, 4,
    -- filter=35 channel=70
    1, 4, -3, 0, 3, -5, 3, 4, -1,
    -- filter=35 channel=71
    3, 7, 7, -5, -3, 2, 0, 4, -3,
    -- filter=35 channel=72
    -7, 0, 2, 0, 3, 0, -1, -3, -5,
    -- filter=35 channel=73
    -2, -2, -3, -2, -3, -1, -6, 3, -3,
    -- filter=35 channel=74
    4, -1, 0, -4, -2, 0, 2, 4, 0,
    -- filter=35 channel=75
    0, 6, -5, 4, -3, 1, 4, 2, -4,
    -- filter=35 channel=76
    -1, -4, -5, 4, -4, 7, 7, 3, 2,
    -- filter=35 channel=77
    -4, 3, -4, -5, 0, 0, 0, -2, 3,
    -- filter=35 channel=78
    -5, -6, -2, 0, 4, -5, -7, -6, -5,
    -- filter=35 channel=79
    -1, 2, 4, 2, 0, 3, -6, -3, 0,
    -- filter=35 channel=80
    -1, -7, 5, 4, -7, -2, -4, 1, 6,
    -- filter=35 channel=81
    -1, 0, 2, -2, 3, 4, 2, 5, -3,
    -- filter=35 channel=82
    0, -5, 7, -6, -6, -5, -3, 0, 0,
    -- filter=35 channel=83
    -6, 6, 0, 4, -5, 6, -1, -5, 5,
    -- filter=35 channel=84
    -2, 6, 1, -1, 0, 6, -7, 2, -7,
    -- filter=35 channel=85
    4, -1, 0, -3, -3, 7, -3, -1, 0,
    -- filter=35 channel=86
    1, 4, 2, -4, 2, 7, -5, 5, -4,
    -- filter=35 channel=87
    5, 5, 2, 0, -3, 2, 0, 3, 1,
    -- filter=35 channel=88
    7, -2, 5, 4, 5, -2, -3, 6, 0,
    -- filter=35 channel=89
    0, -3, -7, -5, 4, 0, -5, -4, -2,
    -- filter=35 channel=90
    4, -3, -3, 4, 9, 2, 2, 0, 0,
    -- filter=35 channel=91
    -5, -6, 1, -2, 6, -3, 2, 3, 1,
    -- filter=35 channel=92
    -4, -2, 3, -6, 2, -4, -7, -3, -3,
    -- filter=35 channel=93
    3, 0, 4, -7, -3, -5, 5, -7, -7,
    -- filter=35 channel=94
    -6, 2, -1, 3, 6, 6, 0, -2, 6,
    -- filter=35 channel=95
    -4, -5, -5, 0, -3, -1, 5, 0, 0,
    -- filter=35 channel=96
    0, 0, 4, 3, -3, 5, 2, 0, 7,
    -- filter=35 channel=97
    6, -1, 4, -4, 5, -5, 4, -2, 1,
    -- filter=35 channel=98
    3, -4, -4, 0, 2, 2, 2, -7, -1,
    -- filter=35 channel=99
    0, -1, -5, 3, -1, 4, -1, -1, 0,
    -- filter=35 channel=100
    -1, 1, 0, -6, 3, 3, 3, 1, -7,
    -- filter=35 channel=101
    0, 2, -7, 2, 5, 2, -1, -4, -1,
    -- filter=35 channel=102
    2, 7, 7, -1, -4, 0, 1, 4, 6,
    -- filter=35 channel=103
    0, 6, 0, -5, -5, -6, -6, -7, 0,
    -- filter=35 channel=104
    -4, 2, 5, 2, 5, 5, 5, 2, 3,
    -- filter=35 channel=105
    -4, 6, 0, 0, -1, 1, 5, 0, 0,
    -- filter=35 channel=106
    -3, 1, -3, 3, -6, 7, -1, -6, 7,
    -- filter=35 channel=107
    5, -5, -1, 7, 6, 3, -7, -3, 0,
    -- filter=35 channel=108
    -4, 0, 5, 5, -2, 0, 4, 2, -6,
    -- filter=35 channel=109
    4, -6, 0, -9, -5, 3, -1, 0, 5,
    -- filter=35 channel=110
    -4, 3, 0, -7, -5, 6, 0, 1, 1,
    -- filter=35 channel=111
    -4, 0, 7, -6, -5, -1, 4, 1, -2,
    -- filter=35 channel=112
    -6, 6, 0, -2, -5, 6, 5, 4, -5,
    -- filter=35 channel=113
    0, 0, 2, 5, 6, -3, -6, -7, -7,
    -- filter=35 channel=114
    1, -4, 3, -6, 3, -6, -7, -1, 2,
    -- filter=35 channel=115
    7, 0, 2, -7, -2, -4, -6, 1, 7,
    -- filter=35 channel=116
    0, 4, -3, 4, -8, -6, 1, -7, -2,
    -- filter=35 channel=117
    -4, 1, -2, 6, -6, 5, -2, 4, -7,
    -- filter=35 channel=118
    3, -1, 1, -3, -5, -6, 3, 5, -4,
    -- filter=35 channel=119
    -3, 3, 1, -5, 0, -3, 4, 3, 0,
    -- filter=35 channel=120
    -1, 2, 0, 1, 6, 4, 1, -2, -3,
    -- filter=35 channel=121
    -3, 7, 0, -3, -4, 2, 4, -2, -2,
    -- filter=35 channel=122
    -6, 1, -6, 3, -1, -6, -4, -3, -2,
    -- filter=35 channel=123
    0, 7, 0, -2, 6, 4, 2, 4, -2,
    -- filter=35 channel=124
    -3, -6, 5, 4, 0, -6, 4, 5, 5,
    -- filter=35 channel=125
    -4, 4, 5, 0, 4, -2, 0, 2, -4,
    -- filter=35 channel=126
    -7, 0, 4, -6, -6, -7, 0, -7, 5,
    -- filter=35 channel=127
    1, 2, 3, 1, -7, 0, 6, -1, 1,
    -- filter=36 channel=0
    6, -5, -4, -1, 0, -4, -11, 5, -12,
    -- filter=36 channel=1
    -1, 4, -11, -13, 17, 5, -5, 8, 8,
    -- filter=36 channel=2
    -5, 5, 3, -8, 4, -5, 3, -8, 8,
    -- filter=36 channel=3
    -5, -17, 7, 0, -12, 2, -7, -5, -6,
    -- filter=36 channel=4
    -15, -6, -11, -14, 0, 0, -9, -7, 13,
    -- filter=36 channel=5
    -7, -5, 2, -10, -2, -4, -5, 6, -10,
    -- filter=36 channel=6
    3, 10, 2, 2, 13, -10, -1, 0, 0,
    -- filter=36 channel=7
    0, 7, 0, -7, 2, 5, 5, -4, 0,
    -- filter=36 channel=8
    3, 5, 8, -1, -3, 3, -8, -2, -1,
    -- filter=36 channel=9
    0, -8, 4, 0, 0, 0, -7, -6, 5,
    -- filter=36 channel=10
    0, -8, 2, -2, 12, 0, -10, 4, -1,
    -- filter=36 channel=11
    -4, 2, -9, 0, 11, -13, -1, 0, -6,
    -- filter=36 channel=12
    -1, 9, -2, -1, 12, 7, 12, 9, -2,
    -- filter=36 channel=13
    -2, 4, -2, -8, 25, -4, -8, 6, -6,
    -- filter=36 channel=14
    6, 7, -2, -2, 3, -1, 2, -6, -4,
    -- filter=36 channel=15
    3, 8, -4, 4, 9, -23, 0, 14, -8,
    -- filter=36 channel=16
    6, -2, 9, -3, 0, 7, 3, -5, 5,
    -- filter=36 channel=17
    -6, 3, 2, -6, 3, -2, -2, -5, 0,
    -- filter=36 channel=18
    5, 3, -11, -7, 27, -30, -8, 9, -9,
    -- filter=36 channel=19
    -5, 4, -3, 0, 5, -6, 2, -3, 2,
    -- filter=36 channel=20
    -5, 11, -14, 5, 19, -21, -8, 13, -9,
    -- filter=36 channel=21
    5, -5, 2, -6, -6, 3, 0, -8, 8,
    -- filter=36 channel=22
    3, 0, 0, -5, 8, -6, -4, 11, -7,
    -- filter=36 channel=23
    -7, -5, 3, 21, 5, -9, -4, 11, -15,
    -- filter=36 channel=24
    5, 3, -5, 4, -6, -2, -4, -3, -5,
    -- filter=36 channel=25
    0, 7, -1, -13, 20, -8, -14, 3, 7,
    -- filter=36 channel=26
    4, -2, 6, -2, -1, 2, 1, -6, 1,
    -- filter=36 channel=27
    5, -5, -3, 2, 12, -16, -18, 9, 3,
    -- filter=36 channel=28
    5, -1, 0, -2, 2, -5, -6, -5, 1,
    -- filter=36 channel=29
    -5, 9, -13, 7, 15, -18, -3, 13, -4,
    -- filter=36 channel=30
    3, 0, 0, 0, 3, -11, -5, -1, 5,
    -- filter=36 channel=31
    6, -14, 0, 0, -1, -10, -19, -3, 0,
    -- filter=36 channel=32
    0, 0, -8, -6, 31, -17, -12, 5, -5,
    -- filter=36 channel=33
    2, -1, -5, 0, 9, -18, -6, 11, -15,
    -- filter=36 channel=34
    -7, 1, 24, 17, 9, 22, -8, 19, 6,
    -- filter=36 channel=35
    -5, -4, 2, 5, -5, -3, 2, 2, -2,
    -- filter=36 channel=36
    5, 0, 3, 2, -2, 8, 0, 6, 5,
    -- filter=36 channel=37
    0, 7, 5, -8, 7, 2, 0, -4, -5,
    -- filter=36 channel=38
    0, -7, -3, 0, 2, -9, 0, 7, 0,
    -- filter=36 channel=39
    -6, 4, 0, 7, 3, -7, -3, 3, -11,
    -- filter=36 channel=40
    -7, -5, -4, 4, 0, -1, -2, -1, -10,
    -- filter=36 channel=41
    1, 26, 4, -12, 35, 25, 0, 4, 27,
    -- filter=36 channel=42
    6, 4, -7, -1, -9, -4, -2, -8, -8,
    -- filter=36 channel=43
    -11, 0, -4, 1, 6, 4, -5, 5, -15,
    -- filter=36 channel=44
    7, 3, 10, 4, 3, 3, -1, -8, 6,
    -- filter=36 channel=45
    2, -9, -12, 2, -10, -13, 0, -2, -6,
    -- filter=36 channel=46
    -6, 5, -2, 2, 6, 10, 1, 5, 4,
    -- filter=36 channel=47
    5, 0, 1, -8, 8, 3, -4, -2, 4,
    -- filter=36 channel=48
    -2, -1, 8, -10, 6, -12, -8, -9, 6,
    -- filter=36 channel=49
    -7, -4, -9, 2, 7, -16, -9, 0, -6,
    -- filter=36 channel=50
    8, -12, -1, -3, 0, -10, -8, -2, 2,
    -- filter=36 channel=51
    -1, -6, 0, -3, -1, 3, -4, -3, -6,
    -- filter=36 channel=52
    0, 0, 13, 10, 11, 7, -1, 14, -3,
    -- filter=36 channel=53
    -4, -2, -3, 2, 5, -2, -7, 6, 3,
    -- filter=36 channel=54
    -5, 5, -4, 0, -5, -2, -5, -7, -1,
    -- filter=36 channel=55
    0, 4, -11, 4, 19, -19, -2, 9, -1,
    -- filter=36 channel=56
    -8, 8, 5, 9, 12, 9, 0, 9, 1,
    -- filter=36 channel=57
    1, 11, -4, 0, 1, 11, 4, -1, 2,
    -- filter=36 channel=58
    1, 4, 5, 2, -1, 5, 2, -5, 0,
    -- filter=36 channel=59
    -3, 0, 0, -2, 10, -8, 0, 1, -2,
    -- filter=36 channel=60
    6, -4, -4, -5, -6, 8, -3, -1, 7,
    -- filter=36 channel=61
    3, 0, 0, -3, 3, 0, 3, 0, 4,
    -- filter=36 channel=62
    0, -6, 3, -2, -7, 3, 3, 4, 3,
    -- filter=36 channel=63
    1, 6, 1, -7, 4, -1, 4, -6, -1,
    -- filter=36 channel=64
    -6, 6, -6, -3, 8, 4, -4, 1, 7,
    -- filter=36 channel=65
    6, -3, 3, 6, 5, 1, -6, 7, 2,
    -- filter=36 channel=66
    0, 14, 7, 6, 32, 6, 7, 17, 9,
    -- filter=36 channel=67
    5, -6, -6, 6, 2, 5, -6, 4, 3,
    -- filter=36 channel=68
    0, 6, -9, 0, 5, 0, 0, -1, 0,
    -- filter=36 channel=69
    -5, -3, -2, 6, 2, -6, 0, 5, -3,
    -- filter=36 channel=70
    -2, 0, 2, 12, 9, -8, -7, 0, -8,
    -- filter=36 channel=71
    -6, -4, -6, 5, -11, -5, -3, -7, -5,
    -- filter=36 channel=72
    10, 3, -5, -7, 4, -14, -7, 2, 3,
    -- filter=36 channel=73
    -1, 1, -8, -6, 6, -15, -7, 2, 0,
    -- filter=36 channel=74
    -6, -2, 18, 2, -1, 0, -11, 16, -6,
    -- filter=36 channel=75
    -6, -12, -6, -12, 10, 3, 1, 0, 0,
    -- filter=36 channel=76
    0, 5, -15, 7, 16, -21, -3, 13, -9,
    -- filter=36 channel=77
    -2, 0, -1, 3, 0, -5, 7, -5, 6,
    -- filter=36 channel=78
    -3, 2, 9, 1, -8, -1, -4, 0, -6,
    -- filter=36 channel=79
    -2, 0, -18, 0, 37, -31, -4, 14, -7,
    -- filter=36 channel=80
    3, -5, 1, -8, 12, -12, -3, -2, 1,
    -- filter=36 channel=81
    4, 1, -4, 2, -1, 4, -1, 5, 5,
    -- filter=36 channel=82
    -6, 5, 4, -2, -6, -8, 0, 1, -5,
    -- filter=36 channel=83
    0, -6, -4, 4, -4, -7, -2, -8, -2,
    -- filter=36 channel=84
    -3, 7, -13, 2, 10, -8, -10, 14, -3,
    -- filter=36 channel=85
    -4, 1, -5, -4, 0, -3, -6, 0, 5,
    -- filter=36 channel=86
    -1, 3, 11, -1, 10, 8, 2, 7, 1,
    -- filter=36 channel=87
    -1, 7, 0, 7, 10, -7, 4, 7, 5,
    -- filter=36 channel=88
    -6, 0, 0, 1, -7, 4, -1, -5, 9,
    -- filter=36 channel=89
    0, 4, -14, 1, 19, -9, -5, 2, -1,
    -- filter=36 channel=90
    0, 0, 17, 5, -2, 3, -1, 6, -1,
    -- filter=36 channel=91
    -4, 5, -10, 2, 8, -11, -12, 5, -3,
    -- filter=36 channel=92
    1, -2, 12, 9, 2, 6, 0, 5, 7,
    -- filter=36 channel=93
    0, -5, -2, -7, 4, 1, 2, -11, 9,
    -- filter=36 channel=94
    -1, -4, 1, -1, 0, -3, -5, 1, -4,
    -- filter=36 channel=95
    -2, -6, 2, 7, 0, 0, 1, -1, -5,
    -- filter=36 channel=96
    1, -6, 0, -6, 6, -2, -2, 1, -3,
    -- filter=36 channel=97
    -2, -3, 5, -3, 0, -3, 0, -2, -4,
    -- filter=36 channel=98
    -4, -5, -1, -5, 9, -19, -1, -1, -7,
    -- filter=36 channel=99
    -1, 4, 11, 2, 7, -6, -14, 11, -3,
    -- filter=36 channel=100
    2, 4, 4, 6, 7, 12, 6, 14, 1,
    -- filter=36 channel=101
    -10, -7, -2, -4, 0, 5, -13, 0, 9,
    -- filter=36 channel=102
    6, -2, 0, -3, -2, 4, 4, 5, -6,
    -- filter=36 channel=103
    4, -3, 2, 3, -6, -6, 3, -8, -9,
    -- filter=36 channel=104
    -3, 2, 5, -8, 1, -10, -10, -4, -1,
    -- filter=36 channel=105
    -4, 9, -11, 8, 9, -7, -5, 11, -4,
    -- filter=36 channel=106
    0, 6, -3, -1, 8, -3, -1, 5, -1,
    -- filter=36 channel=107
    -6, 9, 2, 0, 6, -13, 2, 11, -12,
    -- filter=36 channel=108
    7, 4, 0, -7, 2, -1, -3, 1, 5,
    -- filter=36 channel=109
    2, 8, -7, -1, 22, -13, -8, 4, 2,
    -- filter=36 channel=110
    -5, -4, 5, 2, 2, 0, -4, 0, 6,
    -- filter=36 channel=111
    -5, 2, -5, -7, 10, 2, 3, 0, 2,
    -- filter=36 channel=112
    -5, -9, 11, -1, 0, -7, -9, 4, -11,
    -- filter=36 channel=113
    4, -11, 6, 9, 5, 3, -2, 6, -1,
    -- filter=36 channel=114
    0, 3, -23, -9, 27, -35, -16, 10, -12,
    -- filter=36 channel=115
    3, 0, -5, -4, -4, -2, -6, -3, 6,
    -- filter=36 channel=116
    -1, 11, 0, -2, 11, -7, -14, 4, 9,
    -- filter=36 channel=117
    -3, 1, 4, 3, 5, 1, 6, 0, 4,
    -- filter=36 channel=118
    5, -1, -7, 1, 5, 7, -2, 0, -3,
    -- filter=36 channel=119
    -7, 15, 20, 0, 11, 11, -1, 22, -3,
    -- filter=36 channel=120
    -8, -1, 4, 11, 0, -10, -13, 12, -6,
    -- filter=36 channel=121
    0, 8, 9, -13, 5, 6, -5, 4, 9,
    -- filter=36 channel=122
    6, -5, 11, 0, 9, 10, 7, -4, 14,
    -- filter=36 channel=123
    -7, 0, 4, 10, 12, 16, -9, 5, 1,
    -- filter=36 channel=124
    2, 5, -3, 9, 3, -13, 0, 7, -12,
    -- filter=36 channel=125
    1, 1, 0, -8, 4, -17, -11, 0, 4,
    -- filter=36 channel=126
    -4, -2, -3, -13, 18, -11, -10, 3, -2,
    -- filter=36 channel=127
    5, 8, -2, -1, 6, 7, 3, 9, 0,
    -- filter=37 channel=0
    9, 6, 5, 11, 11, 4, 8, 2, -1,
    -- filter=37 channel=1
    12, 4, 0, 12, 9, 0, 8, 15, 5,
    -- filter=37 channel=2
    1, -4, 1, 5, 0, -2, 3, -5, -4,
    -- filter=37 channel=3
    8, 10, 1, -4, 4, -4, -5, 5, -7,
    -- filter=37 channel=4
    7, 8, 5, -2, 1, -4, 7, 4, 1,
    -- filter=37 channel=5
    -2, 3, 10, 0, 0, 3, 5, 2, 7,
    -- filter=37 channel=6
    2, 14, 14, 4, 8, 12, -2, 5, 1,
    -- filter=37 channel=7
    1, 5, -1, -2, 2, -6, 4, -5, -6,
    -- filter=37 channel=8
    2, -8, 4, -2, -5, -3, 3, 0, 3,
    -- filter=37 channel=9
    0, -9, -3, -2, -2, 0, 5, -2, -7,
    -- filter=37 channel=10
    0, -3, -10, 8, -11, -14, 7, -5, -10,
    -- filter=37 channel=11
    -1, 10, 9, 2, 6, 15, -9, -3, 13,
    -- filter=37 channel=12
    1, 5, 0, 11, -3, -8, 12, -8, -5,
    -- filter=37 channel=13
    2, 1, -14, -3, 2, -10, 6, -7, -4,
    -- filter=37 channel=14
    -4, 4, 0, 5, -7, 5, -1, 3, -3,
    -- filter=37 channel=15
    0, 4, 5, -5, -2, 1, -4, -8, -5,
    -- filter=37 channel=16
    2, 4, 0, -2, -6, 3, 2, -6, 1,
    -- filter=37 channel=17
    -5, -7, 5, 5, 6, -6, -3, -2, -4,
    -- filter=37 channel=18
    3, 9, 1, 4, 11, -10, -4, 1, -12,
    -- filter=37 channel=19
    6, 2, 3, -4, -3, 3, 0, 0, 1,
    -- filter=37 channel=20
    1, 10, 18, 2, 16, 30, 0, 3, 17,
    -- filter=37 channel=21
    2, -7, -11, 1, -6, 3, 0, 0, 0,
    -- filter=37 channel=22
    8, -6, 0, 3, -5, 1, -1, 6, -9,
    -- filter=37 channel=23
    -10, -15, -10, 3, -20, -11, 3, -15, -17,
    -- filter=37 channel=24
    0, -5, 2, -5, 0, -2, 0, -2, 6,
    -- filter=37 channel=25
    5, -14, -14, 2, -16, -25, -1, -11, -16,
    -- filter=37 channel=26
    -1, -7, -3, 3, 7, -1, 3, 2, 10,
    -- filter=37 channel=27
    -1, -20, -26, -8, -20, -27, -4, -18, -28,
    -- filter=37 channel=28
    6, -3, -3, 1, 0, -2, 4, 4, -1,
    -- filter=37 channel=29
    8, 17, 18, 2, 21, 21, -3, 13, 17,
    -- filter=37 channel=30
    7, -6, -12, -6, 0, -2, 2, -1, -10,
    -- filter=37 channel=31
    -5, -12, -21, -1, -8, -18, 0, -7, -12,
    -- filter=37 channel=32
    6, -6, -7, -7, -12, -6, -1, -7, -8,
    -- filter=37 channel=33
    4, -11, -10, -6, -9, -18, -5, -15, -19,
    -- filter=37 channel=34
    2, -9, -2, 7, -12, -13, 10, -10, -4,
    -- filter=37 channel=35
    6, -1, 3, 5, -2, -5, 0, 3, -7,
    -- filter=37 channel=36
    4, 5, -4, 5, 0, 0, 5, 5, 1,
    -- filter=37 channel=37
    -3, 7, 0, 2, -3, 2, 8, 5, 3,
    -- filter=37 channel=38
    0, -1, 1, 4, -12, -8, -2, -8, -7,
    -- filter=37 channel=39
    1, 0, 16, 0, 12, 8, 4, 0, 10,
    -- filter=37 channel=40
    3, 4, 3, -3, -2, 4, 3, 0, 0,
    -- filter=37 channel=41
    19, 4, -7, 15, 10, -11, 14, 11, -7,
    -- filter=37 channel=42
    3, 0, 0, -9, -1, 0, -5, 5, 1,
    -- filter=37 channel=43
    3, 3, 7, 4, 6, 0, 8, 4, 10,
    -- filter=37 channel=44
    0, 0, -12, 3, -8, -12, -3, 1, -3,
    -- filter=37 channel=45
    1, 0, 6, 0, 3, 5, 0, 3, 9,
    -- filter=37 channel=46
    1, -3, 2, 7, -2, -6, 5, 0, 4,
    -- filter=37 channel=47
    -5, -13, -13, 5, -12, -3, 4, -5, -9,
    -- filter=37 channel=48
    2, -12, -22, 0, -7, -19, -1, -10, -17,
    -- filter=37 channel=49
    7, 3, -4, 0, 4, -4, -1, 1, -4,
    -- filter=37 channel=50
    2, -18, -12, -3, -20, -16, -5, -5, -17,
    -- filter=37 channel=51
    0, 8, -4, -3, 7, 0, 0, 0, 0,
    -- filter=37 channel=52
    4, -1, 3, 6, 4, -3, -4, -5, -6,
    -- filter=37 channel=53
    -1, -1, 1, 5, 9, 2, 0, -5, 9,
    -- filter=37 channel=54
    -6, -1, -7, 6, -4, -1, -2, -2, 5,
    -- filter=37 channel=55
    1, -10, 0, 2, -1, 0, -12, 0, -10,
    -- filter=37 channel=56
    2, -2, -5, -5, 2, -7, 3, 4, -6,
    -- filter=37 channel=57
    7, 4, -2, 0, -3, 0, -1, 7, 1,
    -- filter=37 channel=58
    2, 12, 7, 2, 7, -1, 7, 7, 3,
    -- filter=37 channel=59
    5, -6, -20, 4, -14, -21, 0, -7, -11,
    -- filter=37 channel=60
    2, 4, 1, -1, 4, 7, 3, -2, 2,
    -- filter=37 channel=61
    -4, 8, 4, 2, 1, 0, -1, 0, 5,
    -- filter=37 channel=62
    2, -4, -6, -3, 6, -2, -5, 3, 5,
    -- filter=37 channel=63
    -2, 5, 9, 8, 2, 4, -3, 7, 8,
    -- filter=37 channel=64
    -4, 5, 6, 7, 1, 6, -3, -3, -1,
    -- filter=37 channel=65
    -2, -2, 4, 1, -6, 0, 5, 2, -6,
    -- filter=37 channel=66
    8, 2, -7, 11, 3, -13, 0, 1, 2,
    -- filter=37 channel=67
    -4, 6, 1, -3, 4, -2, 0, 4, -3,
    -- filter=37 channel=68
    5, 0, -3, 5, 6, 8, -3, 6, 4,
    -- filter=37 channel=69
    5, 6, 1, 0, -3, -1, -4, 8, -3,
    -- filter=37 channel=70
    0, -19, -17, -1, -16, -13, -5, -11, -19,
    -- filter=37 channel=71
    -2, 0, 5, -5, -5, -2, -5, -2, -2,
    -- filter=37 channel=72
    -5, -12, -8, 6, -8, -7, -7, -6, -3,
    -- filter=37 channel=73
    -6, 0, -3, 3, -7, 1, -2, -1, -2,
    -- filter=37 channel=74
    -1, -11, -12, 7, -10, -3, 7, -7, -5,
    -- filter=37 channel=75
    4, 14, 6, 10, 6, -10, 0, 0, 2,
    -- filter=37 channel=76
    3, 4, 17, 12, 20, 19, 1, 3, 18,
    -- filter=37 channel=77
    4, 1, -3, 4, -4, 0, 6, -3, 7,
    -- filter=37 channel=78
    -6, -7, -1, 4, 2, -1, -1, 0, 5,
    -- filter=37 channel=79
    8, -5, -6, 8, 0, -13, 0, -5, -16,
    -- filter=37 channel=80
    4, -16, -15, 4, -12, -11, 5, -2, -17,
    -- filter=37 channel=81
    -5, 1, -3, -3, -3, -1, 5, 1, 6,
    -- filter=37 channel=82
    1, -5, -3, 0, 4, -2, -2, 4, -3,
    -- filter=37 channel=83
    -7, -9, -10, 0, 3, -5, -7, 0, -10,
    -- filter=37 channel=84
    8, 4, 4, 4, 0, -7, -9, -7, -8,
    -- filter=37 channel=85
    6, -6, -7, -6, 4, 2, 0, -6, -2,
    -- filter=37 channel=86
    1, -2, -5, 10, 0, -1, 5, -7, -3,
    -- filter=37 channel=87
    -3, 5, 2, 5, 10, 10, -1, 1, 7,
    -- filter=37 channel=88
    12, 6, 1, 10, -2, 0, -1, 7, 10,
    -- filter=37 channel=89
    1, -5, -11, -8, -10, -8, 1, -9, -9,
    -- filter=37 channel=90
    7, 0, 0, 8, -8, 0, 3, 1, -2,
    -- filter=37 channel=91
    2, -3, -5, 0, -10, -16, -10, -13, -6,
    -- filter=37 channel=92
    0, 2, -4, -2, -8, 1, 4, -7, 4,
    -- filter=37 channel=93
    -3, -9, -8, 2, -5, 1, 8, 5, -5,
    -- filter=37 channel=94
    -1, 4, 0, 3, 2, -2, 1, 6, 2,
    -- filter=37 channel=95
    5, 5, 2, 2, 0, -5, -7, 2, -6,
    -- filter=37 channel=96
    0, 4, -3, 0, -7, -3, -4, 4, -5,
    -- filter=37 channel=97
    6, -4, 8, -6, -2, -7, 5, -2, 5,
    -- filter=37 channel=98
    -5, -12, -14, -8, -7, -8, -7, -7, -14,
    -- filter=37 channel=99
    -4, -6, -17, 7, -17, -12, 3, -12, -6,
    -- filter=37 channel=100
    -5, -4, -4, 2, -6, 2, 7, -4, -6,
    -- filter=37 channel=101
    0, -3, 0, -1, -5, 0, -3, 0, 3,
    -- filter=37 channel=102
    0, 2, -1, -3, 0, 2, -2, 6, 4,
    -- filter=37 channel=103
    -4, -3, -2, -1, -11, -3, -6, -10, -6,
    -- filter=37 channel=104
    1, -7, -7, -2, -14, 0, -6, 0, -8,
    -- filter=37 channel=105
    -1, 11, 21, 8, 5, 21, -4, 13, 9,
    -- filter=37 channel=106
    3, 0, 0, 10, 7, 13, 0, 2, 8,
    -- filter=37 channel=107
    11, 4, 16, 4, 13, 14, 0, 9, 9,
    -- filter=37 channel=108
    10, 3, 1, 0, 5, -1, 4, 12, 5,
    -- filter=37 channel=109
    -4, -8, -19, 0, -11, -22, -7, -15, -11,
    -- filter=37 channel=110
    -8, -4, -2, -3, 0, 3, -5, -4, 2,
    -- filter=37 channel=111
    -2, -2, -3, -1, 10, 2, 6, 0, 6,
    -- filter=37 channel=112
    0, -9, -7, -1, -17, -2, 0, -4, -5,
    -- filter=37 channel=113
    0, -2, -11, 4, -3, -6, -5, -7, -8,
    -- filter=37 channel=114
    10, 10, 3, 6, 0, 1, 0, 9, -3,
    -- filter=37 channel=115
    -3, -1, 0, -5, -7, 5, -1, -6, -1,
    -- filter=37 channel=116
    3, -8, -14, -10, -13, -10, -4, -10, -7,
    -- filter=37 channel=117
    -5, 1, -10, 0, -9, -6, 6, -5, -9,
    -- filter=37 channel=118
    2, 7, 4, 5, 3, 8, -6, 0, 0,
    -- filter=37 channel=119
    5, -4, -11, -3, -11, -1, -6, -3, -3,
    -- filter=37 channel=120
    0, -4, -10, -4, -18, -12, -10, -21, -8,
    -- filter=37 channel=121
    -5, -7, -8, -3, 1, -5, -5, -7, -12,
    -- filter=37 channel=122
    -3, -19, -14, 10, -10, -13, 5, -12, 0,
    -- filter=37 channel=123
    1, 0, -6, -4, -6, -6, 6, -2, -7,
    -- filter=37 channel=124
    7, 9, 8, -2, 7, 14, 5, 0, 14,
    -- filter=37 channel=125
    5, -5, -13, -5, -3, -10, -3, -7, -10,
    -- filter=37 channel=126
    8, 3, -6, 6, 1, -3, 7, 2, -4,
    -- filter=37 channel=127
    1, -5, 0, -3, 9, 3, 7, 5, -4,
    -- filter=38 channel=0
    3, 10, 2, 0, 17, 17, -9, -9, -7,
    -- filter=38 channel=1
    1, 10, 13, 0, 23, 11, -17, -1, 5,
    -- filter=38 channel=2
    -1, 0, 0, 1, 6, 2, 0, 7, 7,
    -- filter=38 channel=3
    3, 16, 12, 2, 1, 7, 7, 9, 2,
    -- filter=38 channel=4
    2, 12, 0, -1, 3, 0, 0, 10, 9,
    -- filter=38 channel=5
    -1, -4, 0, -1, 10, 9, -10, -6, -7,
    -- filter=38 channel=6
    -3, -4, 0, -2, -1, 8, -4, 2, -9,
    -- filter=38 channel=7
    5, -2, 0, -1, -3, 5, -2, 5, 2,
    -- filter=38 channel=8
    -5, -5, -2, 1, 4, 3, 4, -2, 1,
    -- filter=38 channel=9
    -4, 6, 3, -5, -7, -11, -4, 9, -6,
    -- filter=38 channel=10
    -2, -7, -3, 0, -1, -9, 8, -3, -8,
    -- filter=38 channel=11
    -5, -7, -7, 1, -8, -3, -4, -2, -4,
    -- filter=38 channel=12
    0, -3, -4, 0, 0, 5, -7, 6, 5,
    -- filter=38 channel=13
    1, -1, 11, -7, 2, -8, -4, 12, 3,
    -- filter=38 channel=14
    -5, 0, 0, -4, 1, 1, 5, -4, 2,
    -- filter=38 channel=15
    2, 5, 8, 0, 2, -9, -5, -3, -8,
    -- filter=38 channel=16
    3, -6, -2, 0, -1, -5, 0, 2, -4,
    -- filter=38 channel=17
    1, -6, -1, 6, 0, 2, 6, 6, 1,
    -- filter=38 channel=18
    1, 6, 3, -8, 15, -13, -6, 0, -9,
    -- filter=38 channel=19
    5, -6, -4, 6, -5, 0, 2, -5, -6,
    -- filter=38 channel=20
    -6, 0, -7, -3, 0, 4, 0, 3, -11,
    -- filter=38 channel=21
    -1, 0, -7, -6, -13, -16, 2, 13, 3,
    -- filter=38 channel=22
    6, 2, 0, -4, 6, 2, -7, -6, -4,
    -- filter=38 channel=23
    2, -5, 12, 5, -11, 4, 6, 10, -9,
    -- filter=38 channel=24
    -4, -2, -5, -3, 4, 0, 5, 1, 4,
    -- filter=38 channel=25
    -1, 5, -1, -10, 5, -11, 1, 15, 6,
    -- filter=38 channel=26
    -1, 2, -8, -1, 2, -1, 3, 4, 8,
    -- filter=38 channel=27
    -3, 9, 10, 2, -9, -20, 4, 15, 4,
    -- filter=38 channel=28
    6, -3, 2, 3, -6, 4, 2, -1, -1,
    -- filter=38 channel=29
    -2, -5, -4, 0, -2, 3, -6, -6, -1,
    -- filter=38 channel=30
    2, 7, 3, 4, 4, -2, 2, 1, 0,
    -- filter=38 channel=31
    -5, -1, -3, 7, -25, -13, 20, 22, 5,
    -- filter=38 channel=32
    0, 10, -2, -1, 11, -1, 0, 3, -5,
    -- filter=38 channel=33
    -1, -2, 6, 2, 0, 0, -12, 6, -4,
    -- filter=38 channel=34
    0, 7, 2, -5, -9, 15, -2, 6, 6,
    -- filter=38 channel=35
    6, 6, -6, 3, -3, 0, 3, 5, 6,
    -- filter=38 channel=36
    3, -9, -6, 0, 0, -11, 8, 7, 11,
    -- filter=38 channel=37
    4, 4, 12, -2, 11, 6, -3, -2, 7,
    -- filter=38 channel=38
    -6, -4, -3, -1, -9, -8, 2, 0, -5,
    -- filter=38 channel=39
    -7, -7, 3, -2, 1, -7, -3, 2, -9,
    -- filter=38 channel=40
    1, 7, 6, 2, 2, 0, 4, -3, 2,
    -- filter=38 channel=41
    -4, -2, 4, -10, 14, 6, 3, 8, 14,
    -- filter=38 channel=42
    -3, 7, 6, -4, -1, -3, -3, 1, 6,
    -- filter=38 channel=43
    -5, 8, 10, -5, -5, 1, 0, 5, 3,
    -- filter=38 channel=44
    -1, 7, -1, 7, -6, 2, 7, 7, 0,
    -- filter=38 channel=45
    3, -5, 2, 1, 9, -3, -1, -2, 3,
    -- filter=38 channel=46
    5, 2, 7, 5, -1, -3, 3, 2, 1,
    -- filter=38 channel=47
    1, 0, 4, -3, -5, -8, 12, 11, 0,
    -- filter=38 channel=48
    -2, 1, 4, 2, -1, -14, 4, 13, 9,
    -- filter=38 channel=49
    3, 3, 3, 4, -2, -3, -6, 2, 4,
    -- filter=38 channel=50
    -3, 0, 7, 5, -1, -13, -2, 2, 3,
    -- filter=38 channel=51
    0, 0, -2, 7, -3, 2, 6, 1, 7,
    -- filter=38 channel=52
    4, 0, -1, -6, -5, 7, -5, 6, 7,
    -- filter=38 channel=53
    -7, 2, 5, -1, 0, -2, 0, 7, -2,
    -- filter=38 channel=54
    3, -3, -1, 7, -3, 0, -6, 7, -7,
    -- filter=38 channel=55
    -11, -5, -6, -6, -9, -15, 7, 10, -9,
    -- filter=38 channel=56
    -1, 5, 4, 2, 1, 2, 8, 0, 2,
    -- filter=38 channel=57
    -7, -5, -3, 7, 7, 8, 0, 2, 4,
    -- filter=38 channel=58
    0, -7, 6, -4, 0, 5, -9, 2, 3,
    -- filter=38 channel=59
    0, 3, 1, -6, -5, -18, 9, 14, -4,
    -- filter=38 channel=60
    3, -6, -3, 3, 5, 6, 2, 3, 0,
    -- filter=38 channel=61
    -6, 0, -5, -3, -3, 6, -6, -1, -5,
    -- filter=38 channel=62
    0, 4, 7, 4, 5, -4, 4, 5, 0,
    -- filter=38 channel=63
    -7, -7, -2, 0, -4, -1, 3, -7, 0,
    -- filter=38 channel=64
    -5, -3, 0, 7, -7, -2, 8, 0, 0,
    -- filter=38 channel=65
    -5, 7, 6, -6, -6, 3, -2, 6, 5,
    -- filter=38 channel=66
    -8, 2, 7, -7, 1, -7, -7, 0, 3,
    -- filter=38 channel=67
    -4, 0, 0, -3, 4, 2, 4, -5, -5,
    -- filter=38 channel=68
    0, 2, 4, -3, 0, -3, -1, 7, 0,
    -- filter=38 channel=69
    0, -5, 4, 3, 3, -7, 4, 5, 7,
    -- filter=38 channel=70
    0, 4, 8, 0, -1, -7, -1, 8, 1,
    -- filter=38 channel=71
    3, 0, -2, -3, -4, 1, -1, -3, 0,
    -- filter=38 channel=72
    -6, -1, -4, -8, -16, -16, 0, 9, 0,
    -- filter=38 channel=73
    3, 5, 5, 0, 7, 0, -6, -1, -3,
    -- filter=38 channel=74
    3, -2, -5, 6, -10, 4, -2, 4, -4,
    -- filter=38 channel=75
    0, 8, 18, -13, 11, 12, -12, -3, 1,
    -- filter=38 channel=76
    -3, 3, -2, 1, -8, -11, -7, -6, -7,
    -- filter=38 channel=77
    -3, 6, -2, 2, 1, 5, 4, 7, -1,
    -- filter=38 channel=78
    5, 0, 7, -4, -9, 2, -1, 2, -5,
    -- filter=38 channel=79
    1, 7, 12, -6, 10, -13, -1, 0, 1,
    -- filter=38 channel=80
    -4, -5, 5, -3, -16, -21, 3, 13, -1,
    -- filter=38 channel=81
    4, 4, -4, 5, 4, 0, 5, 2, -1,
    -- filter=38 channel=82
    3, 5, 6, -7, -6, 1, 0, 5, -9,
    -- filter=38 channel=83
    -5, -7, -7, 5, -6, -7, 4, 0, 0,
    -- filter=38 channel=84
    2, -6, 2, 3, 11, -5, -7, 10, -4,
    -- filter=38 channel=85
    -5, 0, -4, 1, 6, 3, -3, 0, 0,
    -- filter=38 channel=86
    1, -4, 5, 2, 7, 2, -10, -7, -4,
    -- filter=38 channel=87
    -4, -5, -3, -1, 2, 1, 1, 8, 6,
    -- filter=38 channel=88
    2, -3, -6, -4, -1, 4, 7, 3, 0,
    -- filter=38 channel=89
    2, 0, 2, -11, -10, -20, -2, 6, -5,
    -- filter=38 channel=90
    0, -3, 2, 1, -10, -2, 13, 2, 6,
    -- filter=38 channel=91
    5, 4, 6, -3, 1, -15, 0, 4, -1,
    -- filter=38 channel=92
    -3, -3, -1, -1, -6, 5, 8, 9, 4,
    -- filter=38 channel=93
    0, -2, 2, 2, -1, -9, 5, 6, 9,
    -- filter=38 channel=94
    3, -5, -3, -7, 4, -3, 0, -2, 0,
    -- filter=38 channel=95
    3, -4, 3, 5, 0, 0, -5, -5, -6,
    -- filter=38 channel=96
    -5, -2, -1, 6, 8, -4, 0, 3, -6,
    -- filter=38 channel=97
    4, 7, 7, 6, 5, 0, 6, -3, -4,
    -- filter=38 channel=98
    -8, 6, 4, -13, -3, -20, -6, 7, -6,
    -- filter=38 channel=99
    -12, 0, -3, 6, -24, -8, 14, 13, 2,
    -- filter=38 channel=100
    4, -1, 5, 2, 2, 2, 8, 3, 7,
    -- filter=38 channel=101
    6, -2, 9, -3, 8, 1, 8, -1, 4,
    -- filter=38 channel=102
    -6, -2, -5, 5, 0, 6, -5, 0, 0,
    -- filter=38 channel=103
    -1, 0, 0, -2, 1, -13, 5, 10, 1,
    -- filter=38 channel=104
    -5, -4, -1, 5, -6, -24, 12, 1, -4,
    -- filter=38 channel=105
    -8, -1, 7, 4, 0, -2, 6, -2, 1,
    -- filter=38 channel=106
    -6, -3, -4, -3, 4, -4, 6, 2, 6,
    -- filter=38 channel=107
    7, 7, 3, 6, 8, 0, 1, -8, 3,
    -- filter=38 channel=108
    1, -3, -1, -6, 10, -3, 0, 1, 7,
    -- filter=38 channel=109
    -8, -6, 0, -7, 3, -16, 0, -1, 7,
    -- filter=38 channel=110
    -9, 0, 5, 2, -2, -8, 4, 5, -2,
    -- filter=38 channel=111
    2, -4, -3, 5, 8, 2, -3, -1, -4,
    -- filter=38 channel=112
    -7, 4, -4, -4, -2, -3, 1, 3, -9,
    -- filter=38 channel=113
    -2, 3, 1, -7, -3, -7, -4, -2, -2,
    -- filter=38 channel=114
    1, 1, 5, -3, 18, 2, -12, -3, -5,
    -- filter=38 channel=115
    -1, -3, -5, -4, 5, 5, 4, 7, -3,
    -- filter=38 channel=116
    1, -2, -1, 4, -9, -12, 8, 9, 4,
    -- filter=38 channel=117
    5, 0, 7, -6, -6, -5, -4, -1, 1,
    -- filter=38 channel=118
    0, -3, -2, -5, -3, -5, -1, 3, -4,
    -- filter=38 channel=119
    -3, -8, -7, -1, -3, 0, -2, 5, 1,
    -- filter=38 channel=120
    -10, 0, 4, 0, -14, -10, -3, 0, 5,
    -- filter=38 channel=121
    0, -4, 1, -10, -5, -5, 0, 0, 0,
    -- filter=38 channel=122
    -6, -3, -1, 9, -11, -14, 11, 16, 9,
    -- filter=38 channel=123
    4, 2, 3, 7, 4, 3, -3, 8, 7,
    -- filter=38 channel=124
    -4, 2, 8, -6, -1, -2, 3, -4, -7,
    -- filter=38 channel=125
    0, -1, 3, -4, -14, -20, -2, 7, -2,
    -- filter=38 channel=126
    -3, 1, -3, -11, 9, -8, -7, 0, -7,
    -- filter=38 channel=127
    2, 5, -7, 2, 0, -1, -3, 1, 0,
    -- filter=39 channel=0
    5, -4, -6, 0, -8, 0, -6, 0, 0,
    -- filter=39 channel=1
    6, 2, -2, 6, -9, 1, -5, 10, 0,
    -- filter=39 channel=2
    0, 0, 0, 2, 5, -2, 2, 2, 1,
    -- filter=39 channel=3
    0, 17, -3, 1, -1, -3, -12, 0, 2,
    -- filter=39 channel=4
    -1, 0, 12, 1, 13, -1, 14, -11, -7,
    -- filter=39 channel=5
    6, -7, 1, -5, -5, 5, -8, -2, 4,
    -- filter=39 channel=6
    -5, -1, -1, -6, -2, -2, 5, 1, -8,
    -- filter=39 channel=7
    1, 6, -5, 6, -6, 2, -3, 1, -1,
    -- filter=39 channel=8
    -7, -5, 4, -4, 14, -4, 2, -8, 4,
    -- filter=39 channel=9
    4, -1, 1, 0, 0, 5, 6, 4, -5,
    -- filter=39 channel=10
    4, -1, 5, -4, 0, 5, -8, 14, 2,
    -- filter=39 channel=11
    -8, 5, 5, 0, 5, 1, 3, -5, 2,
    -- filter=39 channel=12
    9, -1, -3, 5, 2, -2, -1, 4, -1,
    -- filter=39 channel=13
    2, 3, -6, 1, -8, -5, 2, 5, -9,
    -- filter=39 channel=14
    0, -5, 4, -2, 1, 0, 4, 1, 1,
    -- filter=39 channel=15
    -7, -2, 6, -5, 0, 10, 1, 5, -10,
    -- filter=39 channel=16
    9, 8, 2, 2, 2, -7, -5, 7, -8,
    -- filter=39 channel=17
    2, -5, -6, 2, -7, -6, -3, -7, -4,
    -- filter=39 channel=18
    3, 0, 0, -13, -5, 11, -1, 18, -11,
    -- filter=39 channel=19
    2, 5, 2, -5, 4, 5, 0, 1, 6,
    -- filter=39 channel=20
    -3, 5, -4, 0, 11, 6, -3, 6, -13,
    -- filter=39 channel=21
    1, -9, -7, 5, -7, 0, -6, 5, -4,
    -- filter=39 channel=22
    -2, -2, -6, -1, 8, 2, 4, -8, 4,
    -- filter=39 channel=23
    2, -3, 7, -8, 12, 5, 0, 6, -12,
    -- filter=39 channel=24
    0, 0, -2, 3, -4, 4, -1, -5, -5,
    -- filter=39 channel=25
    15, -3, -4, -12, -5, 8, -7, 11, -8,
    -- filter=39 channel=26
    -4, -1, 3, 2, 7, -5, 8, 2, -1,
    -- filter=39 channel=27
    9, -4, 11, -27, 9, 9, 1, 9, -11,
    -- filter=39 channel=28
    0, -3, -6, -5, 0, 2, 3, 7, 5,
    -- filter=39 channel=29
    2, -1, 0, -7, 11, -1, -5, 6, -13,
    -- filter=39 channel=30
    1, -8, -2, -11, 4, 10, 5, 7, -6,
    -- filter=39 channel=31
    1, -7, -7, -18, 6, -4, -3, 2, -8,
    -- filter=39 channel=32
    13, -7, 1, -13, 10, 6, 3, 14, -16,
    -- filter=39 channel=33
    11, 6, -5, 0, -9, -2, -3, 2, 0,
    -- filter=39 channel=34
    -4, 3, 0, -7, 14, -2, 5, -13, 2,
    -- filter=39 channel=35
    -4, 3, -1, -2, 3, -3, -2, 6, -3,
    -- filter=39 channel=36
    2, -7, -2, -2, 12, 4, 0, -3, 4,
    -- filter=39 channel=37
    9, -3, 0, 0, 4, -9, 0, 6, 1,
    -- filter=39 channel=38
    10, -7, -2, 0, 3, 8, -5, 12, -8,
    -- filter=39 channel=39
    -3, 4, 0, -2, 8, 0, -3, 0, -9,
    -- filter=39 channel=40
    -3, 5, -1, 2, -3, 0, 1, 5, 2,
    -- filter=39 channel=41
    -8, 15, -9, 11, -1, -7, 2, 2, -15,
    -- filter=39 channel=42
    6, -7, 0, -5, -7, -4, 1, -6, 4,
    -- filter=39 channel=43
    6, 1, 0, -1, -7, -6, -8, 8, 2,
    -- filter=39 channel=44
    5, 2, 3, -12, -4, 7, 2, -2, 2,
    -- filter=39 channel=45
    2, -6, -5, 3, 3, -4, 5, 0, 1,
    -- filter=39 channel=46
    -4, 1, 3, 2, 2, -2, 0, -6, -4,
    -- filter=39 channel=47
    18, 1, -3, 3, -15, 7, -9, 10, 5,
    -- filter=39 channel=48
    1, -18, -8, -18, 9, 7, 0, 0, -1,
    -- filter=39 channel=49
    -11, 2, 6, -8, 8, 3, 13, 0, -4,
    -- filter=39 channel=50
    -1, -9, 6, -7, -1, 0, 2, -3, 4,
    -- filter=39 channel=51
    3, -1, -3, -3, -6, 5, 0, 6, 0,
    -- filter=39 channel=52
    -1, 3, -6, -7, 16, -8, 2, 1, -10,
    -- filter=39 channel=53
    4, -6, 7, -6, 3, -3, 5, 8, 2,
    -- filter=39 channel=54
    -6, 2, 3, -7, 4, 5, -1, 7, 4,
    -- filter=39 channel=55
    -1, 0, -2, -12, 2, 1, -6, 8, -1,
    -- filter=39 channel=56
    0, 7, -1, -6, 8, -9, 12, 0, 0,
    -- filter=39 channel=57
    5, -7, -5, -1, -3, -7, -3, -5, -8,
    -- filter=39 channel=58
    3, 7, -3, 0, -1, 1, -1, -7, -3,
    -- filter=39 channel=59
    2, 0, -2, -4, 0, 5, -6, 14, -3,
    -- filter=39 channel=60
    4, -3, -2, -5, 6, -1, -2, 0, 6,
    -- filter=39 channel=61
    -3, -3, -3, 5, 1, -3, 1, 3, 2,
    -- filter=39 channel=62
    0, 2, -6, -3, -7, 4, 3, 7, 1,
    -- filter=39 channel=63
    0, -4, -1, -4, 0, 5, 0, -5, 5,
    -- filter=39 channel=64
    -9, -3, 0, 5, 3, 4, 4, -1, 1,
    -- filter=39 channel=65
    2, 0, 0, -6, 5, -7, -1, 1, -4,
    -- filter=39 channel=66
    0, -6, -5, 5, -5, 2, 0, 12, -14,
    -- filter=39 channel=67
    2, -4, -3, 7, -1, -5, -1, 1, 4,
    -- filter=39 channel=68
    -5, 1, -2, 2, 3, 0, -3, -5, -2,
    -- filter=39 channel=69
    0, 6, -3, 5, -8, 0, 4, 5, -5,
    -- filter=39 channel=70
    -7, 1, 3, -10, 7, 0, 4, -6, 2,
    -- filter=39 channel=71
    8, 9, 3, 10, 0, -5, -3, -3, 8,
    -- filter=39 channel=72
    2, -4, -4, -12, -5, 0, -8, 7, -2,
    -- filter=39 channel=73
    0, -1, 1, -18, 12, -1, 1, 14, -6,
    -- filter=39 channel=74
    -1, -9, 6, -17, 14, -13, 19, 0, -1,
    -- filter=39 channel=75
    5, 4, -2, 6, -16, -1, -9, -1, 2,
    -- filter=39 channel=76
    -6, 10, -3, 4, 1, -4, 0, 9, 0,
    -- filter=39 channel=77
    5, 1, 2, -6, 3, 5, 4, 1, 4,
    -- filter=39 channel=78
    0, -1, 2, -6, -2, 7, 0, -3, -6,
    -- filter=39 channel=79
    1, 8, -4, -16, 0, 10, -7, 13, -12,
    -- filter=39 channel=80
    21, -9, 0, -11, -15, 8, -10, 7, 2,
    -- filter=39 channel=81
    3, -6, -1, 1, 1, 2, 4, 5, -3,
    -- filter=39 channel=82
    0, 5, 0, 7, 0, -5, -5, 2, -2,
    -- filter=39 channel=83
    -6, -6, -4, -9, 2, -4, 0, -3, -1,
    -- filter=39 channel=84
    3, -8, 4, -12, 14, 5, 14, -4, -10,
    -- filter=39 channel=85
    0, -5, -6, 0, -3, 1, -3, -5, 3,
    -- filter=39 channel=86
    6, -7, 3, -8, 2, -3, 4, 2, -12,
    -- filter=39 channel=87
    -6, 8, 1, -1, 15, -6, 12, 2, -6,
    -- filter=39 channel=88
    0, 1, -3, -8, 9, -3, 2, -2, -7,
    -- filter=39 channel=89
    4, 7, -2, -6, -3, 11, -8, 16, -9,
    -- filter=39 channel=90
    -7, -3, 5, 2, 6, 2, 5, 0, 5,
    -- filter=39 channel=91
    -5, -15, -2, -14, 18, 5, 17, -3, -9,
    -- filter=39 channel=92
    1, 8, 2, -7, 1, -8, 2, -1, 2,
    -- filter=39 channel=93
    7, 0, -5, -8, -5, -5, 10, -5, 0,
    -- filter=39 channel=94
    0, 0, -3, 3, 5, -5, 0, -1, -4,
    -- filter=39 channel=95
    7, 0, -1, -3, -4, -3, -1, -2, -5,
    -- filter=39 channel=96
    4, 2, -5, 4, -4, 0, -1, 6, -1,
    -- filter=39 channel=97
    4, 11, -6, -1, -1, -3, -10, -5, 7,
    -- filter=39 channel=98
    15, -4, -8, -12, 3, 7, -4, 14, -2,
    -- filter=39 channel=99
    10, -1, -5, -18, 8, -2, 4, 10, -14,
    -- filter=39 channel=100
    -8, 2, 4, 5, 2, 6, 2, -5, 0,
    -- filter=39 channel=101
    -8, -7, -1, -10, 18, -1, 13, -1, -3,
    -- filter=39 channel=102
    -4, -1, 3, 2, 6, -6, -5, 6, -4,
    -- filter=39 channel=103
    10, -5, 0, 7, -15, -2, -1, 5, 8,
    -- filter=39 channel=104
    13, 0, -7, -6, 0, 6, 0, 2, -3,
    -- filter=39 channel=105
    -5, -3, 0, 0, 9, 4, -5, 4, -1,
    -- filter=39 channel=106
    -7, -2, -6, -6, 6, 6, 2, 3, -5,
    -- filter=39 channel=107
    -4, 6, 1, -6, 17, 0, 5, 3, -8,
    -- filter=39 channel=108
    3, 4, 0, 0, -3, 4, -1, 1, -3,
    -- filter=39 channel=109
    13, -13, -1, -20, 13, 11, 12, 12, -5,
    -- filter=39 channel=110
    -3, 4, 1, 6, 5, 2, -6, 5, -6,
    -- filter=39 channel=111
    -4, 1, 0, 0, -1, -4, -8, -5, -5,
    -- filter=39 channel=112
    -7, 1, -2, -11, 8, 4, 9, 2, 2,
    -- filter=39 channel=113
    2, -1, -7, -2, -12, -5, -1, 8, -4,
    -- filter=39 channel=114
    12, -5, -6, -23, 9, 9, -2, 14, -13,
    -- filter=39 channel=115
    -6, -6, -4, 0, -2, -4, 0, 0, 5,
    -- filter=39 channel=116
    12, -3, -6, -15, 0, 10, 3, 2, -9,
    -- filter=39 channel=117
    2, -2, -8, 1, -4, -3, 5, 6, -7,
    -- filter=39 channel=118
    -2, 4, -3, -1, -3, -3, 0, 2, -3,
    -- filter=39 channel=119
    -15, -3, 2, 0, 15, -3, 18, -17, 4,
    -- filter=39 channel=120
    -7, -13, 5, -26, 28, 2, 26, 8, -12,
    -- filter=39 channel=121
    10, 10, -9, 2, -10, 7, -10, 15, -1,
    -- filter=39 channel=122
    15, 1, -2, 8, -7, -10, 0, 0, -6,
    -- filter=39 channel=123
    2, -5, 6, -2, -5, 3, -4, -8, 0,
    -- filter=39 channel=124
    5, 0, 2, 4, 4, -3, 3, -5, -9,
    -- filter=39 channel=125
    13, -16, 5, -20, 9, 2, 7, 11, -10,
    -- filter=39 channel=126
    12, 12, 2, 3, -8, -4, -10, 8, 0,
    -- filter=39 channel=127
    6, 6, 0, -4, -3, 3, 5, -2, -7,
    -- filter=40 channel=0
    8, 8, 2, 1, 3, -9, 6, -7, -12,
    -- filter=40 channel=1
    9, 11, -1, 13, -12, -1, 5, -10, -8,
    -- filter=40 channel=2
    -3, -5, 0, -5, -5, 2, 4, 1, 4,
    -- filter=40 channel=3
    3, 1, -9, 2, -6, 1, 9, 11, -4,
    -- filter=40 channel=4
    2, -1, -3, 5, 1, 0, 8, 0, 4,
    -- filter=40 channel=5
    17, 5, 0, 5, -1, -6, 2, -3, -7,
    -- filter=40 channel=6
    3, 3, 0, 4, -1, 5, -4, 3, 0,
    -- filter=40 channel=7
    0, -4, -3, -5, 3, -3, -5, -1, -5,
    -- filter=40 channel=8
    0, 0, 3, 5, 2, 3, -4, 0, -5,
    -- filter=40 channel=9
    3, -5, 4, 0, -8, 6, 4, 7, 0,
    -- filter=40 channel=10
    -3, -6, 0, -1, -5, 3, -3, -3, 7,
    -- filter=40 channel=11
    -1, -12, 7, -7, -3, 9, -6, -3, 0,
    -- filter=40 channel=12
    -4, -2, 9, 6, -7, 5, 1, -2, -1,
    -- filter=40 channel=13
    -5, -11, 0, -1, -10, 0, 6, 6, -2,
    -- filter=40 channel=14
    3, -3, 2, -3, -7, 3, 1, -1, 0,
    -- filter=40 channel=15
    -13, -11, 7, -3, 6, 7, 3, 6, 5,
    -- filter=40 channel=16
    9, -6, -3, -5, 1, -6, -7, 1, 3,
    -- filter=40 channel=17
    0, -4, 0, 4, -6, -7, 2, 0, -4,
    -- filter=40 channel=18
    -9, -14, 7, -7, -4, 17, 0, 0, 3,
    -- filter=40 channel=19
    -6, 6, -3, -1, 1, 6, -3, -4, -6,
    -- filter=40 channel=20
    -18, -16, -1, -10, 1, 3, -1, 3, 4,
    -- filter=40 channel=21
    3, -2, -6, -5, -14, -9, 0, -10, -9,
    -- filter=40 channel=22
    -6, -4, 4, -6, 2, -3, -3, 0, 3,
    -- filter=40 channel=23
    -7, -9, 7, -19, 12, 3, -3, 8, 2,
    -- filter=40 channel=24
    4, 5, 2, -1, -2, -3, 5, 2, -2,
    -- filter=40 channel=25
    -2, -3, 4, 1, -9, 7, -6, -1, 8,
    -- filter=40 channel=26
    2, 10, -7, 7, -3, -9, -1, 0, -3,
    -- filter=40 channel=27
    -12, -11, 4, -19, -1, 18, 1, 10, 5,
    -- filter=40 channel=28
    -1, 5, 0, -6, 2, -4, 2, 3, 1,
    -- filter=40 channel=29
    -3, -3, 0, -6, 5, 16, -6, 9, 3,
    -- filter=40 channel=30
    0, -3, -2, -1, -5, 7, -4, -4, -2,
    -- filter=40 channel=31
    -2, -5, -6, -12, 0, 4, -6, -6, -7,
    -- filter=40 channel=32
    -10, -13, 9, -4, 0, 20, 6, 6, 3,
    -- filter=40 channel=33
    -4, -2, 0, -7, -4, 8, 4, 12, -2,
    -- filter=40 channel=34
    -10, 0, -1, -3, 14, -3, 9, 0, -5,
    -- filter=40 channel=35
    0, -1, -2, 0, -2, 0, 7, -7, 3,
    -- filter=40 channel=36
    -7, -6, -1, 2, -1, -5, 2, -5, 0,
    -- filter=40 channel=37
    5, 0, 5, 1, -1, -13, 4, -5, -9,
    -- filter=40 channel=38
    -4, 0, 0, -9, 3, 9, -5, 2, 4,
    -- filter=40 channel=39
    -4, -1, 5, -7, 4, -1, -8, 6, -4,
    -- filter=40 channel=40
    -5, -10, -9, -2, -12, -5, -11, 5, -7,
    -- filter=40 channel=41
    7, -3, -5, 14, -9, 6, 6, -13, 0,
    -- filter=40 channel=42
    0, 5, 3, 2, 5, 1, -5, -3, 2,
    -- filter=40 channel=43
    0, 0, -7, -7, -5, 3, 1, 8, 2,
    -- filter=40 channel=44
    -1, -5, 4, 5, -3, -1, -1, -3, -10,
    -- filter=40 channel=45
    -1, -8, -8, -1, -1, -6, -7, 0, 4,
    -- filter=40 channel=46
    -5, -4, -2, 3, 6, -6, -6, 5, -4,
    -- filter=40 channel=47
    2, 0, -3, 6, -13, -3, 4, -13, -5,
    -- filter=40 channel=48
    7, -8, 5, 0, -6, -7, 2, 7, 1,
    -- filter=40 channel=49
    0, -6, 10, -7, 1, 5, -7, 6, -5,
    -- filter=40 channel=50
    -6, -1, 6, -8, 7, 5, 6, -4, -2,
    -- filter=40 channel=51
    6, 1, 6, 6, -3, 0, -1, 0, 4,
    -- filter=40 channel=52
    -3, -8, 4, -2, -4, -7, 1, 4, -6,
    -- filter=40 channel=53
    2, 0, 1, -6, 0, -1, -3, 6, 2,
    -- filter=40 channel=54
    0, 2, 0, 0, 0, 5, -6, -6, 7,
    -- filter=40 channel=55
    -1, -12, 4, -10, -6, 9, 2, 9, 10,
    -- filter=40 channel=56
    4, 5, 6, -5, 3, -5, 1, 0, -7,
    -- filter=40 channel=57
    7, 1, -6, -3, -5, -3, -4, -1, 0,
    -- filter=40 channel=58
    8, 11, 0, 9, -5, 1, 1, -1, -1,
    -- filter=40 channel=59
    1, -7, -6, 4, -12, 13, 5, 0, 5,
    -- filter=40 channel=60
    -3, 6, 1, -4, -4, 0, 3, -6, -7,
    -- filter=40 channel=61
    1, -3, 0, 0, -3, 2, -1, -7, 2,
    -- filter=40 channel=62
    -6, -4, 1, -3, 5, -6, 7, 3, 5,
    -- filter=40 channel=63
    10, 4, 0, 0, 0, 5, -1, -2, 3,
    -- filter=40 channel=64
    -2, -1, -5, 3, 1, -2, 0, -5, 4,
    -- filter=40 channel=65
    -7, -7, -2, 0, 0, 4, -3, 0, -2,
    -- filter=40 channel=66
    9, 3, 4, 0, -4, -1, -3, 1, 2,
    -- filter=40 channel=67
    3, 3, -6, 2, 0, 2, 4, -7, 0,
    -- filter=40 channel=68
    0, 3, -2, -2, 2, 2, 5, -8, 3,
    -- filter=40 channel=69
    7, -6, -2, 8, -7, 1, 5, -2, 5,
    -- filter=40 channel=70
    -10, -10, 0, -13, 2, 1, 5, 0, -2,
    -- filter=40 channel=71
    -6, 0, -10, 0, -7, -6, -4, 6, 1,
    -- filter=40 channel=72
    -6, -9, 3, -11, 2, 0, -6, 7, 8,
    -- filter=40 channel=73
    -5, -3, 10, -4, 11, 15, 7, 9, -5,
    -- filter=40 channel=74
    -2, 0, 13, 0, 0, 4, 5, -5, -2,
    -- filter=40 channel=75
    17, 2, -12, 1, -10, -2, 1, -2, 0,
    -- filter=40 channel=76
    -6, -9, -1, -16, 1, 5, -3, -5, 1,
    -- filter=40 channel=77
    -3, -3, 0, 1, 5, 7, 6, 3, -6,
    -- filter=40 channel=78
    4, 6, 4, 0, -5, 2, -2, -5, -4,
    -- filter=40 channel=79
    -11, -14, 10, -8, -1, 20, -6, 4, 5,
    -- filter=40 channel=80
    8, -13, -3, -1, -5, 2, -2, 0, 5,
    -- filter=40 channel=81
    2, 4, -1, -3, 3, 0, -3, 6, 7,
    -- filter=40 channel=82
    -5, 0, -1, -1, -6, -3, 5, 5, -5,
    -- filter=40 channel=83
    5, 2, 6, 1, 0, -8, 4, 6, -3,
    -- filter=40 channel=84
    -9, -4, 4, -8, 0, 9, -3, 4, 4,
    -- filter=40 channel=85
    0, 1, 3, 3, 6, 6, 3, 2, 3,
    -- filter=40 channel=86
    6, -4, -1, -4, 6, 2, 1, 1, 3,
    -- filter=40 channel=87
    -11, -7, -3, -10, 0, 6, -6, 1, -1,
    -- filter=40 channel=88
    -1, -3, -3, -1, -6, 1, -10, 2, -6,
    -- filter=40 channel=89
    -4, -14, 4, 2, -3, 21, 0, 14, 10,
    -- filter=40 channel=90
    -10, -2, 0, -1, -8, -10, -3, -11, -1,
    -- filter=40 channel=91
    -8, -4, 0, -2, -1, 10, -7, 5, -6,
    -- filter=40 channel=92
    -9, 2, -5, 3, -5, 8, 7, -6, 0,
    -- filter=40 channel=93
    7, 3, 3, 8, -3, -7, -1, 0, 0,
    -- filter=40 channel=94
    -1, 1, -3, 0, 0, 3, -3, -6, -2,
    -- filter=40 channel=95
    -3, 2, 1, -2, -1, -2, 4, -3, 7,
    -- filter=40 channel=96
    6, -5, 0, -1, -7, -3, -2, 3, 6,
    -- filter=40 channel=97
    2, -5, -9, -6, 1, -5, -5, 4, -6,
    -- filter=40 channel=98
    6, -2, 6, -9, -7, 21, -1, 4, 10,
    -- filter=40 channel=99
    -8, -17, 8, -8, 4, 5, -7, 0, 5,
    -- filter=40 channel=100
    5, 0, -6, -4, 0, 0, 0, 0, 5,
    -- filter=40 channel=101
    3, -4, 5, 6, 5, -5, 3, -1, -1,
    -- filter=40 channel=102
    -6, -5, -1, -1, 2, -7, 4, 4, 7,
    -- filter=40 channel=103
    10, 4, -12, 2, -16, -6, -4, -6, -2,
    -- filter=40 channel=104
    0, -8, -6, 1, -5, 6, 1, 0, -7,
    -- filter=40 channel=105
    -3, -12, 0, 0, 4, 7, 3, 0, 4,
    -- filter=40 channel=106
    -1, 1, -6, -3, -6, 3, 3, 0, 0,
    -- filter=40 channel=107
    -7, 0, 0, -3, 0, -3, -10, -1, 3,
    -- filter=40 channel=108
    3, 0, 6, 10, 5, 0, 5, -4, 0,
    -- filter=40 channel=109
    -5, -15, 6, -8, 4, 15, -1, 9, -2,
    -- filter=40 channel=110
    -3, -1, 0, 3, -6, 3, -2, -5, -1,
    -- filter=40 channel=111
    -5, -5, -4, 3, 6, -2, 5, -7, 1,
    -- filter=40 channel=112
    5, 4, 9, 1, 2, -3, 6, 6, -5,
    -- filter=40 channel=113
    -1, -14, 1, 2, -6, -2, 7, 9, 5,
    -- filter=40 channel=114
    2, -13, 11, -10, 3, 17, 4, -1, -2,
    -- filter=40 channel=115
    0, -5, 0, 6, -6, -6, 0, 5, -5,
    -- filter=40 channel=116
    0, 0, 8, 3, 1, 11, 6, 2, 1,
    -- filter=40 channel=117
    0, 1, 0, -8, -4, -4, 4, -6, 5,
    -- filter=40 channel=118
    -5, -7, 1, -2, 3, -7, -6, -5, -4,
    -- filter=40 channel=119
    -4, 9, 10, 3, 4, 8, -2, -12, -3,
    -- filter=40 channel=120
    -13, -15, 14, -8, 23, 10, 7, 8, -6,
    -- filter=40 channel=121
    5, -1, 0, -4, -7, 6, 0, -6, 2,
    -- filter=40 channel=122
    7, -4, -21, 5, -8, -18, -2, -17, -18,
    -- filter=40 channel=123
    -3, 4, -4, -8, -6, -7, -1, -3, -4,
    -- filter=40 channel=124
    -8, 2, 7, -9, 0, -3, 3, -4, 0,
    -- filter=40 channel=125
    -6, -15, 0, 2, 0, 6, 3, 0, 8,
    -- filter=40 channel=126
    9, -12, 3, -5, 0, 12, 0, 0, 6,
    -- filter=40 channel=127
    0, -4, 0, -1, 5, 8, -5, -6, 1,
    -- filter=41 channel=0
    -6, 5, -4, 1, 4, 2, -5, 4, 1,
    -- filter=41 channel=1
    4, 0, -7, 2, -2, -5, -5, -1, 0,
    -- filter=41 channel=2
    -6, -2, -6, -5, -5, 7, 0, -2, -6,
    -- filter=41 channel=3
    0, 1, -4, -5, -1, 0, 0, 3, 4,
    -- filter=41 channel=4
    -2, -5, -2, 2, 5, -4, -1, -5, 5,
    -- filter=41 channel=5
    -2, -1, -5, 4, 4, -7, 6, 0, 0,
    -- filter=41 channel=6
    -6, -5, 0, 0, -6, -5, 1, 4, -1,
    -- filter=41 channel=7
    0, 6, 0, -3, 3, -4, -4, -5, -4,
    -- filter=41 channel=8
    -1, 0, -2, -6, 7, 4, 1, 4, 6,
    -- filter=41 channel=9
    1, -5, -4, 5, -4, 4, -2, -1, -1,
    -- filter=41 channel=10
    -5, -2, 0, -2, 0, -4, -2, -1, -6,
    -- filter=41 channel=11
    3, 1, 6, 5, 7, 3, -3, 0, 4,
    -- filter=41 channel=12
    5, -2, 0, 0, 0, -4, -2, 5, -5,
    -- filter=41 channel=13
    -2, -4, 0, -4, 4, 7, -4, 5, -5,
    -- filter=41 channel=14
    0, 1, 5, -7, 7, -6, -1, -1, -1,
    -- filter=41 channel=15
    -5, -2, 0, 3, -7, 0, -4, -3, 2,
    -- filter=41 channel=16
    -5, 7, 6, -4, 5, 1, 5, -2, 5,
    -- filter=41 channel=17
    2, -5, 2, 2, 5, 4, -4, -1, -2,
    -- filter=41 channel=18
    0, 0, 2, 3, 6, -6, -6, 3, -7,
    -- filter=41 channel=19
    4, 3, 2, -5, -2, -4, 1, 7, -5,
    -- filter=41 channel=20
    -4, -5, -4, 4, 3, -2, -4, -7, -1,
    -- filter=41 channel=21
    0, 0, -3, -5, -5, -2, 0, 6, -5,
    -- filter=41 channel=22
    4, -3, 0, 0, -7, -4, 0, -7, -3,
    -- filter=41 channel=23
    -4, 3, 5, 3, 0, 6, 0, 0, 4,
    -- filter=41 channel=24
    -1, -5, 2, -4, 7, -4, -6, -5, 7,
    -- filter=41 channel=25
    -7, -1, -2, -4, 4, -2, 1, -4, 4,
    -- filter=41 channel=26
    1, 0, -1, -3, -4, -5, -4, 3, -3,
    -- filter=41 channel=27
    -2, 7, -6, 0, 4, 2, -7, -4, -5,
    -- filter=41 channel=28
    -3, -3, 7, 1, -4, 7, -2, -1, -2,
    -- filter=41 channel=29
    3, -2, 3, -2, 4, -5, 3, 2, -3,
    -- filter=41 channel=30
    -1, 0, -4, -4, 4, 0, -2, 6, 1,
    -- filter=41 channel=31
    0, -3, -7, -4, -7, -2, -3, -2, 1,
    -- filter=41 channel=32
    3, 2, 6, 1, -6, 2, -5, -6, 2,
    -- filter=41 channel=33
    -1, -6, -7, -1, -5, -6, 2, -6, -4,
    -- filter=41 channel=34
    2, 5, 5, -1, 6, -3, 1, -2, -3,
    -- filter=41 channel=35
    4, -2, 0, -7, -1, 5, 2, 0, 0,
    -- filter=41 channel=36
    3, 0, 6, 2, 0, 5, 3, -6, -2,
    -- filter=41 channel=37
    2, 0, -3, 0, -2, 0, 7, 8, -1,
    -- filter=41 channel=38
    0, 4, 7, 3, -7, 1, -1, 6, -2,
    -- filter=41 channel=39
    -5, -2, 4, -5, 1, 0, 2, -1, 3,
    -- filter=41 channel=40
    -6, 2, 0, -2, -7, 0, -4, 6, 0,
    -- filter=41 channel=41
    1, -2, -4, 4, 0, 0, -3, -8, -4,
    -- filter=41 channel=42
    0, -7, 3, -2, -4, -3, 4, 0, 3,
    -- filter=41 channel=43
    -2, -6, 0, 5, 1, 0, 3, -6, 1,
    -- filter=41 channel=44
    -3, 4, -3, 5, -6, 0, 5, 1, -4,
    -- filter=41 channel=45
    1, -7, -4, -6, 1, 2, 3, 7, 1,
    -- filter=41 channel=46
    1, 0, 4, 3, 0, -5, -1, 1, -2,
    -- filter=41 channel=47
    7, -4, -2, -1, -2, 6, 0, 2, 4,
    -- filter=41 channel=48
    -5, 0, -7, -6, 4, 4, 2, 3, -1,
    -- filter=41 channel=49
    4, 2, -2, 3, -2, -2, 3, 2, 7,
    -- filter=41 channel=50
    5, -1, 1, 3, 5, 0, 3, 1, -6,
    -- filter=41 channel=51
    -4, 2, -1, -1, 0, 7, -5, -5, -1,
    -- filter=41 channel=52
    3, 3, -5, 4, 3, 3, -6, -5, 2,
    -- filter=41 channel=53
    2, 2, -7, -2, 0, -4, -3, 1, -1,
    -- filter=41 channel=54
    1, 5, -1, 5, 0, 2, 6, 3, 2,
    -- filter=41 channel=55
    3, 0, -3, -3, -2, -5, 2, 3, -4,
    -- filter=41 channel=56
    5, -3, 1, 7, -2, 5, 4, -6, -3,
    -- filter=41 channel=57
    1, 4, 7, 6, -4, -7, 0, 0, 0,
    -- filter=41 channel=58
    -3, 6, -7, 1, -4, 2, 0, 1, 2,
    -- filter=41 channel=59
    0, 1, -3, -1, 2, -2, -6, -4, 6,
    -- filter=41 channel=60
    -3, 4, 6, -6, 4, -2, -2, 4, 0,
    -- filter=41 channel=61
    0, 4, 6, 2, -2, -2, -7, 4, -5,
    -- filter=41 channel=62
    -6, -2, 7, -4, -2, -1, 4, -3, 1,
    -- filter=41 channel=63
    3, -1, 3, -1, -4, 4, 5, 4, 0,
    -- filter=41 channel=64
    0, 6, 0, 2, -3, 0, -1, -7, -3,
    -- filter=41 channel=65
    -4, -7, 2, 3, 3, 2, -1, 4, -1,
    -- filter=41 channel=66
    1, -1, 4, 1, -2, 6, -1, -2, -3,
    -- filter=41 channel=67
    -1, 2, -1, -2, -4, -5, 0, -5, 0,
    -- filter=41 channel=68
    0, 0, 2, -4, 3, -4, 2, -3, 0,
    -- filter=41 channel=69
    -5, -1, 1, -5, 2, -3, 4, -1, 2,
    -- filter=41 channel=70
    6, 4, 2, -7, -2, -7, 1, 0, -1,
    -- filter=41 channel=71
    -7, -3, 3, 4, 0, 1, 0, -6, 7,
    -- filter=41 channel=72
    0, 1, 4, -6, 5, -2, -1, -4, -5,
    -- filter=41 channel=73
    2, 7, -1, -6, 5, -4, -6, 2, 4,
    -- filter=41 channel=74
    0, 0, -4, -4, -5, 0, 0, 7, 0,
    -- filter=41 channel=75
    2, -2, 3, 1, -2, 1, 7, -1, -4,
    -- filter=41 channel=76
    -7, 2, -1, -8, 0, 3, -3, -1, 6,
    -- filter=41 channel=77
    -2, -2, 2, -2, 3, 0, 4, 7, 3,
    -- filter=41 channel=78
    -5, 0, 1, -2, 0, -7, 0, 3, -3,
    -- filter=41 channel=79
    1, 1, 4, 2, 0, -7, -7, 0, -4,
    -- filter=41 channel=80
    -2, -1, -4, -1, -2, -6, -3, 5, -2,
    -- filter=41 channel=81
    -6, -3, 0, -7, 6, -2, 4, 0, -3,
    -- filter=41 channel=82
    5, -5, -1, -7, 6, -3, 0, -3, 1,
    -- filter=41 channel=83
    -6, -3, -4, -1, -4, 0, -6, 5, 0,
    -- filter=41 channel=84
    -2, 3, -2, -5, -3, 1, 5, 3, 7,
    -- filter=41 channel=85
    2, 4, -3, 6, -1, 1, 6, -3, -6,
    -- filter=41 channel=86
    0, 7, -5, 4, -4, -7, 3, 3, 4,
    -- filter=41 channel=87
    2, -5, 2, 1, -2, 6, 5, -7, -5,
    -- filter=41 channel=88
    2, 5, 0, -2, 3, 6, 7, -3, 4,
    -- filter=41 channel=89
    -2, 1, -4, 2, -3, -4, -3, -3, 0,
    -- filter=41 channel=90
    4, 4, -4, -4, -1, -5, 0, -4, 1,
    -- filter=41 channel=91
    -7, -6, 0, -1, 5, -3, -2, 1, -2,
    -- filter=41 channel=92
    0, -4, 2, -2, 6, -6, 6, -5, 3,
    -- filter=41 channel=93
    -2, -2, 3, 4, 3, -4, -2, -2, 6,
    -- filter=41 channel=94
    -2, -6, -5, 0, -2, -3, 0, 5, -3,
    -- filter=41 channel=95
    4, -5, 1, 4, 0, 1, 4, 5, 2,
    -- filter=41 channel=96
    -6, -1, -3, 5, -3, 0, 3, 3, -2,
    -- filter=41 channel=97
    -1, 1, 6, 7, -6, 6, 1, -2, -2,
    -- filter=41 channel=98
    3, 0, -7, -7, 1, -7, -2, 1, 3,
    -- filter=41 channel=99
    0, 0, 3, 1, 0, 2, -5, -3, -3,
    -- filter=41 channel=100
    -4, 2, 0, -7, -4, 6, -3, 3, 5,
    -- filter=41 channel=101
    -1, 2, -3, 5, 5, -2, -4, 3, 0,
    -- filter=41 channel=102
    -3, 6, -5, 4, -1, -1, -1, -2, 3,
    -- filter=41 channel=103
    5, -4, 0, 2, -5, -6, 1, -5, 0,
    -- filter=41 channel=104
    -4, 5, 5, 3, -2, 4, 0, 1, -2,
    -- filter=41 channel=105
    -2, 2, 4, 3, 2, -7, 1, 1, -2,
    -- filter=41 channel=106
    6, 0, 1, -6, 0, -5, 2, 4, 5,
    -- filter=41 channel=107
    -4, -2, 0, -7, 3, -5, 7, 5, -2,
    -- filter=41 channel=108
    -3, 0, -6, -1, -3, 3, 4, 0, 4,
    -- filter=41 channel=109
    -5, -3, -2, 6, -5, 4, 5, -4, 1,
    -- filter=41 channel=110
    6, -6, -3, 2, -2, 6, -6, 4, -3,
    -- filter=41 channel=111
    -5, 0, 6, 7, 0, 1, 0, -3, 3,
    -- filter=41 channel=112
    -1, -1, -4, 2, 5, -4, -4, 3, 4,
    -- filter=41 channel=113
    -1, -3, 3, 3, -6, 0, 5, -3, 2,
    -- filter=41 channel=114
    5, -2, -3, -7, -1, 4, 0, 6, 4,
    -- filter=41 channel=115
    4, -5, 0, 0, 3, -6, -6, 3, 3,
    -- filter=41 channel=116
    -4, 5, 1, 4, -6, 2, 0, 3, 4,
    -- filter=41 channel=117
    -5, -7, -1, 5, -5, -5, -5, 4, 7,
    -- filter=41 channel=118
    3, 3, -6, 2, -4, 3, -3, 6, -6,
    -- filter=41 channel=119
    1, 5, 6, 4, 4, 2, 0, -6, 4,
    -- filter=41 channel=120
    -5, 0, 4, -1, 0, 0, -4, -6, 0,
    -- filter=41 channel=121
    -4, 3, 1, 0, 2, -1, -4, -2, 5,
    -- filter=41 channel=122
    -6, 0, 6, 2, -4, 5, 1, -1, 0,
    -- filter=41 channel=123
    -4, 4, -4, -3, 5, 5, -1, 7, 3,
    -- filter=41 channel=124
    -3, -2, 1, -4, 1, -5, 3, 4, 0,
    -- filter=41 channel=125
    0, -1, 1, -4, 2, -3, -4, 3, -2,
    -- filter=41 channel=126
    -6, 3, 0, 5, 6, 0, 2, 7, 4,
    -- filter=41 channel=127
    0, -6, 2, 0, -3, -5, 2, -5, 0,
    -- filter=42 channel=0
    2, 0, 1, -3, -4, 4, 9, 9, 3,
    -- filter=42 channel=1
    -5, -6, -11, -8, -6, -7, 5, 5, -3,
    -- filter=42 channel=2
    3, -4, 6, -3, 4, -3, 2, 4, 2,
    -- filter=42 channel=3
    2, 4, 3, -8, -1, 10, 1, 1, 3,
    -- filter=42 channel=4
    -15, -6, 0, -18, -5, -2, -2, -9, -13,
    -- filter=42 channel=5
    -8, -13, -1, -5, -2, -6, 11, 3, -7,
    -- filter=42 channel=6
    -6, -3, 5, -9, -7, -3, 0, -3, 2,
    -- filter=42 channel=7
    6, 2, 2, 0, -7, -5, -2, 7, 0,
    -- filter=42 channel=8
    0, -6, 5, -1, -1, -5, -11, -6, -8,
    -- filter=42 channel=9
    10, -4, 0, 13, 0, -8, 11, 0, -8,
    -- filter=42 channel=10
    8, 9, 3, 9, -1, 0, -4, -4, 0,
    -- filter=42 channel=11
    3, 4, 12, 3, -6, 4, -7, -6, -8,
    -- filter=42 channel=12
    -9, 0, -5, -12, -5, -7, -5, 3, -7,
    -- filter=42 channel=13
    8, 6, -1, 0, 6, 0, 1, 1, -11,
    -- filter=42 channel=14
    5, -5, 2, -2, -5, 5, 5, -4, 6,
    -- filter=42 channel=15
    -2, 8, 0, 0, -12, -8, 2, -2, -6,
    -- filter=42 channel=16
    -5, -9, -9, -1, -4, -8, 0, 0, 2,
    -- filter=42 channel=17
    -4, 1, -2, -6, -3, 1, -5, 0, -5,
    -- filter=42 channel=18
    4, 5, 9, -3, -3, -5, -2, -8, -12,
    -- filter=42 channel=19
    6, -1, 3, -2, 5, 2, -6, -1, 5,
    -- filter=42 channel=20
    -10, 1, 12, -6, -5, -3, -14, -14, -5,
    -- filter=42 channel=21
    13, 8, -14, 8, 11, -12, 0, 0, -9,
    -- filter=42 channel=22
    -5, -3, 7, -3, -5, 0, -8, -3, 2,
    -- filter=42 channel=23
    12, 10, 3, -6, -22, -10, -6, -15, -9,
    -- filter=42 channel=24
    6, 0, 5, 0, 4, -6, -7, 0, -5,
    -- filter=42 channel=25
    2, 9, -8, 5, 10, -4, 12, 6, -14,
    -- filter=42 channel=26
    -3, -8, -13, 0, -3, -7, 2, -2, 1,
    -- filter=42 channel=27
    11, 2, -1, 17, -13, -9, 18, -11, -13,
    -- filter=42 channel=28
    -6, -1, 6, -3, 3, -7, 0, -3, 7,
    -- filter=42 channel=29
    -8, -6, 14, -12, -6, -8, -9, -13, -1,
    -- filter=42 channel=30
    -3, -5, -4, 4, -8, -3, 4, 3, 0,
    -- filter=42 channel=31
    18, 0, -3, 33, 0, -7, 5, -9, -14,
    -- filter=42 channel=32
    -1, 12, 4, -4, -8, -10, 1, -1, -8,
    -- filter=42 channel=33
    14, 9, 0, 10, -3, -2, 14, 5, -3,
    -- filter=42 channel=34
    0, -15, -8, -14, -23, -7, -12, -18, -7,
    -- filter=42 channel=35
    0, -2, -1, 3, -4, -6, 3, 0, 3,
    -- filter=42 channel=36
    -1, 1, 0, 4, -4, -10, -7, -5, -10,
    -- filter=42 channel=37
    4, -4, -6, 5, -7, 2, 2, 0, -7,
    -- filter=42 channel=38
    1, 7, 1, 4, 4, -7, 5, -5, -6,
    -- filter=42 channel=39
    -8, 0, 2, 0, -4, 5, -1, 0, 6,
    -- filter=42 channel=40
    1, 8, 1, -7, -8, -3, -6, -4, -5,
    -- filter=42 channel=41
    -5, 3, -7, -19, 0, -11, 1, 5, -3,
    -- filter=42 channel=42
    0, -1, -1, 7, 8, -3, 14, 3, 5,
    -- filter=42 channel=43
    -8, 4, 8, -9, -5, -2, -3, -7, 7,
    -- filter=42 channel=44
    13, -8, -13, 9, -4, -12, 14, -7, 0,
    -- filter=42 channel=45
    1, -5, -4, -4, -4, -2, -3, -2, -3,
    -- filter=42 channel=46
    0, -2, -6, -1, -3, -6, -1, -6, -5,
    -- filter=42 channel=47
    14, -7, -9, 16, 16, -9, 14, 11, -5,
    -- filter=42 channel=48
    9, -1, -8, 24, 13, -7, 16, 7, -9,
    -- filter=42 channel=49
    1, -2, 0, 2, -4, 2, 7, 0, -1,
    -- filter=42 channel=50
    15, 6, -2, 18, 4, -6, 12, -7, -3,
    -- filter=42 channel=51
    -6, 0, 5, -1, -2, 3, 6, 5, 5,
    -- filter=42 channel=52
    -4, -4, 0, -13, -17, -8, -6, -13, 0,
    -- filter=42 channel=53
    -1, -3, 5, 3, -4, -2, 3, 0, -5,
    -- filter=42 channel=54
    -6, 4, 0, 2, -3, 5, -5, 3, 0,
    -- filter=42 channel=55
    6, 4, 7, 5, -5, -5, -8, -5, -11,
    -- filter=42 channel=56
    -3, -7, -9, -9, -2, -5, -3, -5, 0,
    -- filter=42 channel=57
    0, -5, 0, 4, 2, 0, 4, 2, 3,
    -- filter=42 channel=58
    0, -2, -4, -1, -6, -9, 6, 0, -6,
    -- filter=42 channel=59
    8, 7, -7, 24, 14, -13, 12, -2, -9,
    -- filter=42 channel=60
    0, 3, -1, -2, -3, 4, 0, -5, 0,
    -- filter=42 channel=61
    0, -8, 4, -1, 0, 1, -10, -8, -4,
    -- filter=42 channel=62
    6, -1, 1, -6, -5, 2, 0, 0, 2,
    -- filter=42 channel=63
    -11, -10, -11, -1, -11, -10, 0, -6, -5,
    -- filter=42 channel=64
    -5, 4, -1, -7, 0, -4, -2, -9, 2,
    -- filter=42 channel=65
    4, 4, 1, -3, 1, -6, 4, 1, 6,
    -- filter=42 channel=66
    -12, 3, -4, -16, -5, -7, -9, -4, 0,
    -- filter=42 channel=67
    0, 4, 6, -3, -5, -3, 1, -6, 0,
    -- filter=42 channel=68
    -5, -1, 2, 6, -5, 5, 5, -6, 6,
    -- filter=42 channel=69
    -3, -2, -5, -4, -3, 4, 4, 7, 3,
    -- filter=42 channel=70
    9, -4, -9, 10, -11, -4, 3, -9, -10,
    -- filter=42 channel=71
    -2, -4, 9, 1, 2, -5, -4, -4, 0,
    -- filter=42 channel=72
    18, 12, 4, 23, 0, -10, 12, -7, -13,
    -- filter=42 channel=73
    9, 2, 3, -5, -13, -6, 5, -4, -4,
    -- filter=42 channel=74
    5, -11, -12, 8, -16, -10, 0, -16, -8,
    -- filter=42 channel=75
    -1, 1, -3, 3, -5, 3, 6, 8, 5,
    -- filter=42 channel=76
    4, 6, 10, -14, -14, 0, 0, -4, 7,
    -- filter=42 channel=77
    2, 1, 2, -4, 6, -2, -5, -5, 2,
    -- filter=42 channel=78
    -4, -4, 4, 6, 3, 0, 4, -7, -7,
    -- filter=42 channel=79
    2, 5, 1, -3, -5, -10, 10, -4, -8,
    -- filter=42 channel=80
    23, 14, 0, 37, 10, -14, 16, 8, -9,
    -- filter=42 channel=81
    -5, 2, 1, -1, 6, 6, 0, -5, -4,
    -- filter=42 channel=82
    0, 5, -4, 2, 2, 5, -5, -1, -2,
    -- filter=42 channel=83
    11, 7, -9, 4, 0, -6, 9, 0, -11,
    -- filter=42 channel=84
    -6, 7, 4, -1, -15, -2, -3, -6, -13,
    -- filter=42 channel=85
    4, 3, 7, 3, 7, 1, -4, 0, 6,
    -- filter=42 channel=86
    1, -10, 1, -10, -6, -2, 0, -10, -3,
    -- filter=42 channel=87
    -2, -5, 4, -15, -9, -7, -5, -6, 1,
    -- filter=42 channel=88
    -3, -1, -5, 6, -12, -2, -9, -12, -5,
    -- filter=42 channel=89
    14, 19, 0, 7, 9, -16, 4, 8, -13,
    -- filter=42 channel=90
    -8, -7, 6, 0, -15, 0, -11, -19, -9,
    -- filter=42 channel=91
    13, 8, 2, 0, -1, -12, 5, -7, -15,
    -- filter=42 channel=92
    0, 2, 6, -8, -6, 4, 0, -7, 0,
    -- filter=42 channel=93
    8, 0, -5, 11, -9, -9, 11, 1, -3,
    -- filter=42 channel=94
    0, -5, -1, -6, 5, -5, 0, -2, -7,
    -- filter=42 channel=95
    -6, 0, 4, -6, 5, 0, -3, -6, 1,
    -- filter=42 channel=96
    9, 9, -6, 3, 0, 7, 0, 1, 2,
    -- filter=42 channel=97
    0, 0, 10, 3, 7, 0, -1, 2, 0,
    -- filter=42 channel=98
    22, 3, 4, 16, 14, -11, 18, 10, 0,
    -- filter=42 channel=99
    20, 5, 0, 16, -11, -9, 1, -18, -23,
    -- filter=42 channel=100
    -1, -1, -9, -7, 1, -5, -1, -7, 0,
    -- filter=42 channel=101
    -8, 4, 8, -4, -10, 4, -9, 4, -8,
    -- filter=42 channel=102
    -4, 4, -1, -3, 5, -5, -6, -1, 0,
    -- filter=42 channel=103
    9, 0, -10, 23, 14, 0, 7, 7, -7,
    -- filter=42 channel=104
    14, 8, -7, 29, 12, -2, 9, 3, -7,
    -- filter=42 channel=105
    4, -3, 2, -6, 0, -3, -10, -7, -1,
    -- filter=42 channel=106
    -2, 7, 2, -7, 3, 4, -9, 3, 4,
    -- filter=42 channel=107
    -7, -5, 5, -17, -15, -7, -15, -12, 5,
    -- filter=42 channel=108
    0, 0, 4, -1, -3, -7, -6, -1, 3,
    -- filter=42 channel=109
    12, 7, -1, 7, -5, -12, 12, -6, -14,
    -- filter=42 channel=110
    9, 10, 3, 9, 0, -11, 0, -13, -8,
    -- filter=42 channel=111
    4, -7, -7, -2, -7, 2, 0, 5, 6,
    -- filter=42 channel=112
    10, -10, -2, 1, -2, -6, 10, -9, -7,
    -- filter=42 channel=113
    16, 9, 5, 4, 2, -5, 5, 0, -9,
    -- filter=42 channel=114
    6, 7, 5, 0, -18, -12, 5, -15, -8,
    -- filter=42 channel=115
    -6, 2, -1, 5, 4, -1, -5, -2, 2,
    -- filter=42 channel=116
    15, 0, -1, 7, -5, -15, 12, 7, -10,
    -- filter=42 channel=117
    3, 3, -6, -4, 0, 5, 7, 4, 5,
    -- filter=42 channel=118
    6, 5, 5, -5, 5, -3, 0, 0, -3,
    -- filter=42 channel=119
    -3, -8, -11, -12, -21, -14, -5, -14, -5,
    -- filter=42 channel=120
    11, 0, -3, 5, -19, -13, 0, -12, -19,
    -- filter=42 channel=121
    4, 0, 7, 3, 6, 2, -6, 3, 2,
    -- filter=42 channel=122
    11, -2, -17, 20, 5, -9, 11, -2, -16,
    -- filter=42 channel=123
    -9, 0, 3, -9, -10, -10, -5, -9, 4,
    -- filter=42 channel=124
    -5, 2, 0, 0, -11, 3, -2, -1, -1,
    -- filter=42 channel=125
    13, 9, 2, 17, 8, -4, 15, -9, -10,
    -- filter=42 channel=126
    12, 4, 9, 0, 10, 2, 0, 0, -8,
    -- filter=42 channel=127
    -3, -4, -3, -8, -5, -1, -5, 0, 5,
    -- filter=43 channel=0
    7, -5, -13, 10, -5, -12, 9, -4, -3,
    -- filter=43 channel=1
    1, -2, -10, 3, 0, -6, 7, -3, -16,
    -- filter=43 channel=2
    7, -6, 1, -5, -4, -7, -3, 2, -3,
    -- filter=43 channel=3
    -2, -11, 3, -18, -4, -11, 3, 0, -5,
    -- filter=43 channel=4
    -2, -13, 0, -16, -15, -18, -6, -20, -5,
    -- filter=43 channel=5
    0, 0, 0, -7, -1, 2, 5, 1, -3,
    -- filter=43 channel=6
    5, 6, -8, 15, 8, -3, 3, 9, 0,
    -- filter=43 channel=7
    -6, 1, -1, 2, -2, -3, -2, 0, 1,
    -- filter=43 channel=8
    3, -6, 0, 10, -14, -9, 2, -10, -7,
    -- filter=43 channel=9
    -7, -4, 5, -6, 9, 8, -3, 7, -5,
    -- filter=43 channel=10
    -5, 1, 5, 0, 2, 6, 5, 5, -10,
    -- filter=43 channel=11
    -8, 6, -3, -4, 8, 4, -1, 5, 13,
    -- filter=43 channel=12
    0, 3, -13, 2, 4, -17, -3, -5, -1,
    -- filter=43 channel=13
    2, 4, -5, 1, 0, -16, -1, -5, -12,
    -- filter=43 channel=14
    0, 2, 0, -5, -3, 6, 0, 7, -3,
    -- filter=43 channel=15
    7, 1, -18, 15, 5, -14, 5, -3, -15,
    -- filter=43 channel=16
    -3, -7, 6, -9, 2, 10, -2, -2, 4,
    -- filter=43 channel=17
    -1, 0, -3, -4, -7, -1, -7, -2, -3,
    -- filter=43 channel=18
    6, 16, -6, 18, 18, -26, 9, 6, -15,
    -- filter=43 channel=19
    0, -6, -3, 0, -2, -2, 4, -1, 4,
    -- filter=43 channel=20
    0, 7, -6, -2, 7, 2, 0, 3, 1,
    -- filter=43 channel=21
    -13, -1, 24, -10, 1, 20, -4, 0, 15,
    -- filter=43 channel=22
    4, 3, -8, 0, 4, -4, 5, -7, -7,
    -- filter=43 channel=23
    6, 0, -16, 7, -6, -9, 2, -2, -15,
    -- filter=43 channel=24
    -4, 5, 7, 4, 0, -5, 3, -1, 1,
    -- filter=43 channel=25
    -1, 3, 8, 5, 13, -3, 2, -7, -3,
    -- filter=43 channel=26
    -2, 4, 13, -2, 1, 4, 0, -3, 1,
    -- filter=43 channel=27
    12, 20, -17, 16, 5, -11, 4, -5, -12,
    -- filter=43 channel=28
    -2, -4, 1, 3, 5, -2, -3, -6, -6,
    -- filter=43 channel=29
    -5, 11, -1, 10, 24, 5, 5, 13, 13,
    -- filter=43 channel=30
    -2, 11, 0, -1, 0, 3, -5, 1, -2,
    -- filter=43 channel=31
    -16, 0, 15, -6, -9, 10, -12, -15, 11,
    -- filter=43 channel=32
    6, 6, -18, 1, 11, -23, 5, 4, -11,
    -- filter=43 channel=33
    7, 9, 3, 8, 18, -12, 10, 1, -18,
    -- filter=43 channel=34
    5, -16, -25, 12, -15, -22, 5, -18, -27,
    -- filter=43 channel=35
    1, 7, -4, 4, -3, -3, 3, 2, -6,
    -- filter=43 channel=36
    -4, 0, 0, -9, -5, 0, -12, -11, 7,
    -- filter=43 channel=37
    1, 9, 0, -1, -7, 2, 0, -10, -7,
    -- filter=43 channel=38
    -1, 6, 8, -4, 5, -1, -8, -3, 1,
    -- filter=43 channel=39
    -9, 7, 8, 6, 1, -3, -1, 2, 11,
    -- filter=43 channel=40
    -6, 2, -9, 4, -3, 3, 0, 0, -5,
    -- filter=43 channel=41
    14, -2, -13, 10, 8, -41, 12, -10, -23,
    -- filter=43 channel=42
    -1, 9, -2, -2, -2, 2, -2, -3, 0,
    -- filter=43 channel=43
    10, 0, -11, 9, 0, -6, 5, 1, -8,
    -- filter=43 channel=44
    1, 1, -4, 0, -6, -6, 1, -1, -5,
    -- filter=43 channel=45
    -6, 3, 0, -3, 1, 0, 6, 9, -1,
    -- filter=43 channel=46
    -4, -1, -5, 0, -4, -6, 3, -3, -2,
    -- filter=43 channel=47
    -9, 0, 17, -15, 2, 13, 1, 6, 5,
    -- filter=43 channel=48
    4, 4, 7, 1, 4, 6, -15, -4, -5,
    -- filter=43 channel=49
    4, 14, -2, 14, 1, -15, 5, -4, -4,
    -- filter=43 channel=50
    5, 2, 5, 0, 0, 5, 2, 6, -3,
    -- filter=43 channel=51
    6, 1, 4, 4, -2, 2, 6, 0, -4,
    -- filter=43 channel=52
    4, 1, -14, 9, -13, -15, -5, -15, -6,
    -- filter=43 channel=53
    -3, 5, -5, 0, 5, -3, -5, 10, 1,
    -- filter=43 channel=54
    2, -6, -6, -6, -3, -7, 3, 1, 2,
    -- filter=43 channel=55
    1, 1, -4, 5, 12, -8, 4, 9, -6,
    -- filter=43 channel=56
    13, -11, -10, 14, -6, -1, 0, 1, -18,
    -- filter=43 channel=57
    1, -7, 0, 0, -11, -13, 0, -2, -3,
    -- filter=43 channel=58
    2, -4, -2, -6, -3, 7, 2, -1, 5,
    -- filter=43 channel=59
    2, 10, 2, 2, 6, 6, -8, -2, 2,
    -- filter=43 channel=60
    -5, -6, -3, 3, -2, -7, -3, -3, -1,
    -- filter=43 channel=61
    -9, -5, 0, -2, -11, -1, 0, 1, 3,
    -- filter=43 channel=62
    0, -2, 5, -5, 0, -1, -3, -4, -5,
    -- filter=43 channel=63
    3, 0, 4, -2, 2, 9, -4, 3, 8,
    -- filter=43 channel=64
    -3, -10, 3, -7, 0, -4, -9, 0, 0,
    -- filter=43 channel=65
    -4, 6, -4, -1, -1, 4, -4, 1, 7,
    -- filter=43 channel=66
    9, 0, -12, 2, 3, -13, 9, 1, -13,
    -- filter=43 channel=67
    -1, -7, 2, 6, -3, -8, 2, -4, -8,
    -- filter=43 channel=68
    -2, -2, -5, -1, -2, 4, -1, 5, 8,
    -- filter=43 channel=69
    -6, 4, 7, 6, 1, 0, 0, 0, 4,
    -- filter=43 channel=70
    10, 6, -11, 20, -11, -12, 7, -6, -15,
    -- filter=43 channel=71
    0, 2, -5, -1, -2, -5, 2, 1, -2,
    -- filter=43 channel=72
    0, 12, 5, -3, 8, 14, -7, 1, 6,
    -- filter=43 channel=73
    0, 4, -1, 15, 3, -6, -4, -11, -6,
    -- filter=43 channel=74
    7, -5, -19, 10, -8, -22, -6, -14, -17,
    -- filter=43 channel=75
    0, -4, -6, 4, 1, -7, 10, -3, -10,
    -- filter=43 channel=76
    -3, 5, -6, 4, 8, 0, -7, 6, 8,
    -- filter=43 channel=77
    -7, 7, 6, -6, 2, -4, 5, 1, -1,
    -- filter=43 channel=78
    -4, -4, -2, 3, -9, -1, -1, -7, -2,
    -- filter=43 channel=79
    4, 18, -13, 20, 24, -28, 13, 3, -24,
    -- filter=43 channel=80
    -3, 11, 22, -12, 16, 16, -10, 3, 15,
    -- filter=43 channel=81
    2, 6, 7, 4, 1, 1, 1, 3, 2,
    -- filter=43 channel=82
    3, -3, -2, -2, -3, -2, 1, -1, 1,
    -- filter=43 channel=83
    -5, 0, 8, -2, 0, -2, -1, -6, 0,
    -- filter=43 channel=84
    9, 7, -10, 1, 2, -11, -7, 2, -17,
    -- filter=43 channel=85
    0, 7, 0, -4, 1, 0, -7, 0, -6,
    -- filter=43 channel=86
    8, 2, -13, 3, -9, -7, 8, 0, -7,
    -- filter=43 channel=87
    4, -9, -17, 0, -1, -14, 0, -4, -3,
    -- filter=43 channel=88
    -4, -8, 1, -10, -11, 0, -8, -5, 0,
    -- filter=43 channel=89
    0, 4, 3, 6, 18, 3, 4, 1, -3,
    -- filter=43 channel=90
    -5, -12, -11, -8, -15, -6, -9, -17, 0,
    -- filter=43 channel=91
    5, 15, -8, 5, 4, -10, -1, 0, -17,
    -- filter=43 channel=92
    -3, -6, -13, -3, -14, -13, -2, -10, -11,
    -- filter=43 channel=93
    8, 7, 17, 5, -7, 9, -6, -12, 5,
    -- filter=43 channel=94
    -3, 6, 4, 0, -4, 6, -1, 1, -5,
    -- filter=43 channel=95
    3, -4, 2, 2, 0, 2, 6, -4, 0,
    -- filter=43 channel=96
    2, 2, 0, 7, 5, 1, 1, -1, 0,
    -- filter=43 channel=97
    -8, -8, 1, -10, 0, 0, 5, 0, -10,
    -- filter=43 channel=98
    2, 11, 8, 8, 18, 3, -1, -6, 0,
    -- filter=43 channel=99
    -8, 4, -10, 9, -10, 3, -4, -13, -5,
    -- filter=43 channel=100
    0, -5, -14, 1, -9, -12, 8, 0, -6,
    -- filter=43 channel=101
    3, -12, -8, -10, -6, -6, -10, -14, -8,
    -- filter=43 channel=102
    3, -5, -6, 5, 0, 5, 3, -1, -4,
    -- filter=43 channel=103
    -10, 2, 11, -11, 8, 12, 5, -2, 12,
    -- filter=43 channel=104
    -5, 6, 20, -9, 5, 15, -5, -4, 10,
    -- filter=43 channel=105
    -11, -2, 0, 12, 8, 4, 0, 13, 3,
    -- filter=43 channel=106
    6, -1, -2, 6, 0, -5, -3, 5, 4,
    -- filter=43 channel=107
    -1, 7, -17, 18, 6, -19, 5, 5, -8,
    -- filter=43 channel=108
    -6, 0, 2, 7, 7, -14, -1, 0, 0,
    -- filter=43 channel=109
    10, 10, -9, 14, 6, -8, -6, -4, -20,
    -- filter=43 channel=110
    -7, 1, -1, 3, -7, 0, -3, 0, -1,
    -- filter=43 channel=111
    9, -7, 5, 8, -7, 2, -4, 5, -7,
    -- filter=43 channel=112
    -2, -3, -1, 0, -5, -12, 7, -8, -9,
    -- filter=43 channel=113
    1, 5, -5, 3, 10, -4, 6, -1, -15,
    -- filter=43 channel=114
    11, 7, -19, 19, 16, -19, 17, 9, -13,
    -- filter=43 channel=115
    2, 7, 5, 5, -1, 3, -2, 7, -5,
    -- filter=43 channel=116
    5, 13, 8, 6, 11, -5, -3, 2, 5,
    -- filter=43 channel=117
    -6, -1, 2, -5, 2, -6, 0, -1, -1,
    -- filter=43 channel=118
    2, -3, -2, -4, 5, -1, 0, 0, -1,
    -- filter=43 channel=119
    10, -15, -14, 9, -17, -22, 9, -5, -17,
    -- filter=43 channel=120
    9, 17, -17, 26, -2, -17, -3, -12, -19,
    -- filter=43 channel=121
    3, -5, -4, -3, 6, -2, 6, 2, -5,
    -- filter=43 channel=122
    -6, -2, 25, -6, 4, 21, -15, -10, 6,
    -- filter=43 channel=123
    8, -8, -6, 0, -9, -13, -9, -1, -9,
    -- filter=43 channel=124
    3, 5, -1, 7, 10, -8, 6, -1, -2,
    -- filter=43 channel=125
    -10, 3, 9, -3, 0, 1, -5, 4, 0,
    -- filter=43 channel=126
    3, 1, -3, 4, 21, -9, 18, 11, -4,
    -- filter=43 channel=127
    4, -7, -5, 4, -5, 0, 2, 1, -3,
    -- filter=44 channel=0
    -5, 4, -3, 13, 0, -7, 14, 9, 0,
    -- filter=44 channel=1
    3, -6, -4, 11, -3, -8, 6, 8, -4,
    -- filter=44 channel=2
    -3, 1, 6, 4, 9, 6, -5, -8, -6,
    -- filter=44 channel=3
    -4, -1, -4, -4, -6, -1, 6, 11, 11,
    -- filter=44 channel=4
    7, -1, -1, -5, -8, -4, -2, 1, -1,
    -- filter=44 channel=5
    6, -1, 5, 7, -1, 4, 15, 21, 12,
    -- filter=44 channel=6
    0, 9, 1, -4, 0, 6, 5, 2, 2,
    -- filter=44 channel=7
    -6, 5, -6, 0, 0, -2, 0, -6, 0,
    -- filter=44 channel=8
    1, 7, -4, 1, 2, -9, 2, -6, -9,
    -- filter=44 channel=9
    -5, -9, -5, 5, -4, 6, 8, 0, -3,
    -- filter=44 channel=10
    -2, -2, 3, 2, -3, 6, 12, 4, -4,
    -- filter=44 channel=11
    -13, 11, 8, -6, 4, 14, -1, -5, -4,
    -- filter=44 channel=12
    8, -8, -3, 0, -2, 0, 5, -4, -4,
    -- filter=44 channel=13
    2, -13, 4, 13, 2, 2, -2, -7, -7,
    -- filter=44 channel=14
    6, -5, -1, 3, -7, 0, 1, 0, 1,
    -- filter=44 channel=15
    -11, -6, 1, 5, 8, 8, -6, 0, 0,
    -- filter=44 channel=16
    -9, -16, -9, 0, -8, -5, 1, 1, 6,
    -- filter=44 channel=17
    2, 7, 3, -7, 7, -3, -6, -2, 0,
    -- filter=44 channel=18
    -3, -3, 9, 8, 11, 19, -6, -4, -2,
    -- filter=44 channel=19
    3, 6, -5, -1, 0, 0, -3, -4, 6,
    -- filter=44 channel=20
    -9, 1, 11, -3, 13, 11, -20, -9, -8,
    -- filter=44 channel=21
    -4, -24, -9, -8, -7, 0, 1, -5, 8,
    -- filter=44 channel=22
    -3, 0, 1, -4, 0, -7, -1, 5, -2,
    -- filter=44 channel=23
    -13, -9, -6, -3, 14, -1, 6, -7, -13,
    -- filter=44 channel=24
    0, 4, -4, 6, 6, 3, -4, 6, 4,
    -- filter=44 channel=25
    -2, -15, 6, 11, 6, 7, 4, -8, 4,
    -- filter=44 channel=26
    -1, -2, -5, 1, 4, 5, 0, 7, 8,
    -- filter=44 channel=27
    3, -3, 0, 12, 16, 10, 9, -7, -17,
    -- filter=44 channel=28
    -4, -3, 0, 0, 1, -4, 3, -6, -6,
    -- filter=44 channel=29
    -2, 15, 20, -6, 13, 18, -6, 0, -2,
    -- filter=44 channel=30
    1, -5, -2, 7, 2, -2, 8, -1, 4,
    -- filter=44 channel=31
    -8, -12, -11, 3, -7, 6, 5, 2, 5,
    -- filter=44 channel=32
    2, -10, 12, 4, 16, 18, -4, 0, 2,
    -- filter=44 channel=33
    -5, -6, 0, -1, 3, 1, 15, 3, -6,
    -- filter=44 channel=34
    -4, 8, -12, 6, 4, -21, 2, -5, -16,
    -- filter=44 channel=35
    -2, 5, 0, -1, 1, -1, 4, 6, 2,
    -- filter=44 channel=36
    -3, 1, 3, 8, -2, -4, -10, -9, -4,
    -- filter=44 channel=37
    -5, -11, -16, 12, -1, -10, 14, -1, 0,
    -- filter=44 channel=38
    0, -10, 3, 7, 8, 11, 8, -2, 4,
    -- filter=44 channel=39
    -8, 9, 0, 0, 3, 12, -2, -2, 4,
    -- filter=44 channel=40
    -15, -1, -9, -12, 0, -3, -11, -14, -11,
    -- filter=44 channel=41
    2, -7, -11, 11, -5, -6, -7, -16, -7,
    -- filter=44 channel=42
    -8, -6, 6, -2, -6, 3, -4, 9, 6,
    -- filter=44 channel=43
    -11, -6, -2, 4, 1, 6, 8, 9, 7,
    -- filter=44 channel=44
    0, -10, -13, 2, -8, -2, 5, -5, -2,
    -- filter=44 channel=45
    -10, -2, 1, -3, -7, -4, -6, 7, 7,
    -- filter=44 channel=46
    5, -1, -9, 4, 4, -4, -1, 4, -9,
    -- filter=44 channel=47
    -11, -26, -18, -14, -21, -13, -4, 6, 12,
    -- filter=44 channel=48
    -4, -19, -4, -1, 0, -5, 1, -3, -7,
    -- filter=44 channel=49
    -3, 1, 15, -3, 16, 10, -11, -7, -13,
    -- filter=44 channel=50
    0, -12, -1, 0, -4, 7, 1, -7, -1,
    -- filter=44 channel=51
    0, 1, 6, 3, 4, 5, 4, 3, 5,
    -- filter=44 channel=52
    -3, 3, -5, 9, 7, 2, 0, -11, 0,
    -- filter=44 channel=53
    -7, 10, 0, -4, 6, 6, -7, -3, 3,
    -- filter=44 channel=54
    0, 0, 2, -5, 1, -2, 3, -7, 7,
    -- filter=44 channel=55
    -3, 2, 0, 2, 8, 15, -4, -6, -17,
    -- filter=44 channel=56
    3, 6, -10, 3, -1, 2, -4, -10, -9,
    -- filter=44 channel=57
    -2, 7, -5, 0, -4, -8, 4, -1, 1,
    -- filter=44 channel=58
    6, 0, 1, -1, 7, 3, 12, 5, 6,
    -- filter=44 channel=59
    1, -14, 1, 5, -2, 0, 0, -2, -5,
    -- filter=44 channel=60
    -2, -1, 5, 1, 3, -5, 2, -4, 0,
    -- filter=44 channel=61
    6, 2, 0, 2, 3, 1, 3, -7, -1,
    -- filter=44 channel=62
    -5, 3, -5, -1, 3, -1, 3, 3, 1,
    -- filter=44 channel=63
    0, 2, -2, 0, 4, -2, 5, 10, 14,
    -- filter=44 channel=64
    0, 8, -7, 3, 5, -1, 1, -9, -7,
    -- filter=44 channel=65
    -3, 5, 7, 3, 4, 0, -2, -1, 4,
    -- filter=44 channel=66
    12, -1, -5, 5, 2, 3, 4, 0, -8,
    -- filter=44 channel=67
    -2, -5, 1, 0, 2, 4, 5, 5, -3,
    -- filter=44 channel=68
    -3, 6, -2, -5, -7, 6, -2, -5, -7,
    -- filter=44 channel=69
    -4, -6, -5, 8, 0, -3, 3, 4, 7,
    -- filter=44 channel=70
    -5, -5, -6, 3, 9, -1, -7, -3, -13,
    -- filter=44 channel=71
    -9, -10, -7, -7, -10, -7, 4, 2, -4,
    -- filter=44 channel=72
    5, 0, 1, 13, -2, 13, 9, -2, -6,
    -- filter=44 channel=73
    -3, 10, 0, 7, 6, 5, 2, -10, -12,
    -- filter=44 channel=74
    3, -3, -12, 7, 7, -6, -10, -18, -4,
    -- filter=44 channel=75
    0, 0, -9, 9, -2, -11, 23, 17, 20,
    -- filter=44 channel=76
    -14, 0, 10, -7, 5, 15, -13, -8, -2,
    -- filter=44 channel=77
    -2, -5, 6, 2, -1, -1, 2, -1, -6,
    -- filter=44 channel=78
    -1, 0, 5, -2, 0, 8, 5, 0, 7,
    -- filter=44 channel=79
    -9, -12, -2, 13, 21, 16, 0, -8, -16,
    -- filter=44 channel=80
    -6, -16, -10, 5, -7, 8, 12, -3, 9,
    -- filter=44 channel=81
    3, 4, 6, 6, 0, 0, 3, 6, 2,
    -- filter=44 channel=82
    -10, 0, -2, 0, 4, -6, 6, 1, 2,
    -- filter=44 channel=83
    -7, -1, -2, 0, -5, 1, 2, -3, -7,
    -- filter=44 channel=84
    3, 2, 11, 2, 8, 8, -6, -7, -11,
    -- filter=44 channel=85
    5, 4, 6, -6, 0, -6, -1, 5, 2,
    -- filter=44 channel=86
    12, 9, -8, 5, -2, -1, 3, 6, 1,
    -- filter=44 channel=87
    4, 3, 2, 8, 1, -6, -10, -2, -5,
    -- filter=44 channel=88
    -2, -3, -7, -6, -2, -6, -2, -11, -1,
    -- filter=44 channel=89
    -1, -4, 2, 9, 13, 16, 10, -3, -7,
    -- filter=44 channel=90
    -3, -7, -14, 0, -11, -10, -5, -6, -11,
    -- filter=44 channel=91
    3, -2, -1, 7, 7, 4, -9, -12, -19,
    -- filter=44 channel=92
    0, 3, -8, 4, 3, 2, 6, 0, -9,
    -- filter=44 channel=93
    -9, -9, -8, 1, -8, -9, 7, 0, -1,
    -- filter=44 channel=94
    -6, -1, -3, -2, 6, -3, 4, 3, 4,
    -- filter=44 channel=95
    6, -2, 0, -5, -6, 7, -5, 5, -6,
    -- filter=44 channel=96
    -6, -5, 1, -7, -6, 5, 3, 5, -1,
    -- filter=44 channel=97
    -6, -6, 1, -12, -11, -5, -2, -1, 1,
    -- filter=44 channel=98
    4, 0, 8, 7, -1, 16, 13, 4, -1,
    -- filter=44 channel=99
    -4, 8, -1, 2, 16, 1, 3, -7, -4,
    -- filter=44 channel=100
    9, 3, -3, 6, 0, -5, 8, -8, -1,
    -- filter=44 channel=101
    -3, 4, 7, -3, -2, -6, 2, -12, -8,
    -- filter=44 channel=102
    -4, 7, -3, 1, -5, 1, 2, -2, 2,
    -- filter=44 channel=103
    -12, -19, -6, -17, -21, 0, 1, 10, 17,
    -- filter=44 channel=104
    -9, -16, 0, 6, -2, -2, -3, -7, 2,
    -- filter=44 channel=105
    0, 6, 10, -3, 4, 7, -11, -6, -9,
    -- filter=44 channel=106
    -10, 1, -4, 0, 0, 0, -5, -10, -8,
    -- filter=44 channel=107
    -4, 1, 3, -5, 8, 6, -3, -11, -6,
    -- filter=44 channel=108
    -4, -2, -5, -3, 8, -3, 3, 12, -4,
    -- filter=44 channel=109
    4, 2, 2, 18, 20, 14, 0, -9, -16,
    -- filter=44 channel=110
    5, -3, 0, 8, 7, -1, 7, 1, 2,
    -- filter=44 channel=111
    3, 7, 0, 0, -4, -5, -4, -1, -1,
    -- filter=44 channel=112
    4, 3, -5, -1, 8, -9, 4, -5, 3,
    -- filter=44 channel=113
    1, -11, -9, 2, 5, 1, 5, 0, 0,
    -- filter=44 channel=114
    -7, 8, 16, 3, 30, 20, -1, -2, -3,
    -- filter=44 channel=115
    0, 7, 1, 3, -5, 4, -2, -2, 0,
    -- filter=44 channel=116
    -1, 7, 10, 9, 9, 12, 2, -3, -5,
    -- filter=44 channel=117
    -6, 0, 0, -2, 1, 3, -4, -8, 0,
    -- filter=44 channel=118
    3, 4, 0, 0, -1, 6, -2, 6, -7,
    -- filter=44 channel=119
    2, 0, -15, 2, 3, -12, -1, -13, -17,
    -- filter=44 channel=120
    1, 12, 9, 2, 19, 9, -4, -19, -22,
    -- filter=44 channel=121
    0, -10, -4, 1, -7, 3, 0, -1, 2,
    -- filter=44 channel=122
    -20, -39, -34, -13, -28, -21, -8, -7, 4,
    -- filter=44 channel=123
    -8, -6, -2, 0, -1, -11, 0, -8, 0,
    -- filter=44 channel=124
    -3, -1, -2, -4, 5, 1, 0, -2, 2,
    -- filter=44 channel=125
    0, -5, 0, 14, 6, 5, 0, -2, 0,
    -- filter=44 channel=126
    -9, -11, -8, 0, -5, 5, 1, 12, 14,
    -- filter=44 channel=127
    0, 1, -3, 8, -2, 0, -1, 0, -6,
    -- filter=45 channel=0
    5, -3, -2, -2, 4, -4, 1, -2, -7,
    -- filter=45 channel=1
    5, 6, -3, -2, 0, -3, 7, -3, 2,
    -- filter=45 channel=2
    0, -6, -5, 0, 3, -1, 1, -4, 4,
    -- filter=45 channel=3
    0, 3, 3, 6, -1, 4, 7, -3, -4,
    -- filter=45 channel=4
    -3, -7, 5, 1, 0, -3, -1, 5, 1,
    -- filter=45 channel=5
    4, -3, -4, 0, -3, 2, -4, 5, -5,
    -- filter=45 channel=6
    3, 6, 7, -3, -4, 3, 0, 5, 3,
    -- filter=45 channel=7
    0, 4, -6, 2, 0, -6, 1, -1, -2,
    -- filter=45 channel=8
    -6, 4, 7, -1, -3, -1, 1, 0, 2,
    -- filter=45 channel=9
    5, 4, -3, -7, 0, -1, 5, 0, 0,
    -- filter=45 channel=10
    -2, 0, 2, 7, -6, 0, -6, 0, 4,
    -- filter=45 channel=11
    -6, -3, -2, -6, 2, -2, -2, -1, 4,
    -- filter=45 channel=12
    -1, -2, 0, 2, 4, -4, 5, 3, -5,
    -- filter=45 channel=13
    -2, 2, -4, 9, -2, 0, 0, -8, 0,
    -- filter=45 channel=14
    4, -3, -2, 0, 7, -6, -4, 0, -5,
    -- filter=45 channel=15
    3, 2, -2, 4, -1, 5, -2, 0, -5,
    -- filter=45 channel=16
    5, 3, 4, 0, 0, 0, -4, -5, 2,
    -- filter=45 channel=17
    2, 6, -6, 4, 4, -4, 1, -5, 6,
    -- filter=45 channel=18
    7, 1, -6, 5, 5, -6, -4, -5, -7,
    -- filter=45 channel=19
    -5, 0, 3, 0, 5, -5, -5, -1, -3,
    -- filter=45 channel=20
    0, 2, 7, -2, -5, 5, 2, -4, 0,
    -- filter=45 channel=21
    8, 3, 6, 0, -4, 0, -3, 4, 4,
    -- filter=45 channel=22
    -4, 5, 4, -5, 0, 6, 2, -4, -5,
    -- filter=45 channel=23
    -3, 0, -3, -1, 0, -6, -6, -4, 0,
    -- filter=45 channel=24
    -7, 3, 5, 0, -4, 3, 1, 1, -7,
    -- filter=45 channel=25
    0, 0, -1, -5, -1, -7, -1, -4, -7,
    -- filter=45 channel=26
    0, -5, 7, 7, -1, 2, 7, 0, 0,
    -- filter=45 channel=27
    6, -7, 6, -6, -6, -7, -9, -7, 0,
    -- filter=45 channel=28
    -5, 0, 0, 2, -3, -3, -2, 0, 7,
    -- filter=45 channel=29
    -4, 7, 5, 3, 2, -5, 2, -5, -1,
    -- filter=45 channel=30
    -1, -1, -1, -7, 0, 0, -6, 2, 1,
    -- filter=45 channel=31
    2, 0, 2, -3, -5, 0, -7, -1, 2,
    -- filter=45 channel=32
    1, -4, 1, -5, -7, 3, -5, -3, 0,
    -- filter=45 channel=33
    1, 0, 1, 5, -5, 0, -8, -6, 6,
    -- filter=45 channel=34
    3, 1, -4, -1, -4, 2, -4, 3, 3,
    -- filter=45 channel=35
    4, 4, 1, -6, 2, -5, 4, 1, 0,
    -- filter=45 channel=36
    -4, 0, 0, 6, 5, 4, 5, -2, 0,
    -- filter=45 channel=37
    4, 3, 7, 1, 0, 6, -3, 3, 4,
    -- filter=45 channel=38
    -4, -4, 0, 0, 0, 0, -5, -8, -6,
    -- filter=45 channel=39
    -1, -1, 2, -1, -6, -2, 3, 4, 7,
    -- filter=45 channel=40
    5, 0, 0, -4, 7, 3, 5, 4, 4,
    -- filter=45 channel=41
    7, -3, 3, 8, -2, -5, 0, -3, 4,
    -- filter=45 channel=42
    4, 3, -6, -6, 4, 5, 7, 3, 6,
    -- filter=45 channel=43
    3, -4, -6, 0, 4, -7, 0, -1, 7,
    -- filter=45 channel=44
    7, -8, -5, -2, -6, 1, 1, -5, -1,
    -- filter=45 channel=45
    5, -3, -3, 3, 1, 5, 0, 0, 0,
    -- filter=45 channel=46
    0, -5, -5, -2, -6, 3, 0, -4, -3,
    -- filter=45 channel=47
    2, 4, -1, 6, -6, -5, -5, -3, -5,
    -- filter=45 channel=48
    6, -3, 5, -2, 3, 3, 4, 1, -1,
    -- filter=45 channel=49
    0, -5, -7, -2, -1, -2, 4, 0, 4,
    -- filter=45 channel=50
    -6, -4, -3, -5, 0, 3, -3, 2, 5,
    -- filter=45 channel=51
    -3, -6, 1, 2, -1, 2, 0, 2, -5,
    -- filter=45 channel=52
    1, -4, 6, -4, -6, 1, -2, -3, -6,
    -- filter=45 channel=53
    2, -4, 4, -6, -3, 3, -5, 1, 0,
    -- filter=45 channel=54
    3, 3, 5, -3, 0, 0, 0, -7, -1,
    -- filter=45 channel=55
    2, -6, -4, -4, -4, -8, -5, -8, -6,
    -- filter=45 channel=56
    4, 0, -3, 5, -7, 2, 3, -3, 6,
    -- filter=45 channel=57
    2, 0, 4, -1, 0, 0, -4, -3, 1,
    -- filter=45 channel=58
    1, -1, -3, -4, -6, 0, 6, 4, -4,
    -- filter=45 channel=59
    7, 0, 1, -6, 2, -1, 0, -7, -6,
    -- filter=45 channel=60
    0, -6, 0, 1, -4, 1, 4, 3, -2,
    -- filter=45 channel=61
    -7, 3, 4, -2, 1, -3, 0, 2, 0,
    -- filter=45 channel=62
    -6, -6, 7, -1, -3, 1, 7, -4, 0,
    -- filter=45 channel=63
    0, 6, 7, 5, -1, 0, 4, -4, 7,
    -- filter=45 channel=64
    -2, -3, 4, 0, -1, 6, 6, -7, -1,
    -- filter=45 channel=65
    3, -7, 4, -5, -4, 0, 3, 0, 0,
    -- filter=45 channel=66
    -3, 4, -4, 6, 3, -9, -4, 4, 2,
    -- filter=45 channel=67
    -3, 0, -6, 0, -5, 1, -3, 0, 1,
    -- filter=45 channel=68
    -6, 2, 0, -6, -6, 0, 0, 1, 1,
    -- filter=45 channel=69
    -2, -2, -4, 2, 5, 3, 7, 0, 3,
    -- filter=45 channel=70
    2, 0, 6, 1, -8, -6, -6, 3, 5,
    -- filter=45 channel=71
    7, 3, 1, 6, -2, -4, 4, -4, 7,
    -- filter=45 channel=72
    5, -7, 5, 0, 2, -4, -6, 0, -3,
    -- filter=45 channel=73
    4, -1, 3, 5, -2, 4, -1, 0, 3,
    -- filter=45 channel=74
    -1, 0, -1, -3, -2, -2, -7, -5, 4,
    -- filter=45 channel=75
    6, -2, -3, 9, -4, 0, 6, 3, 4,
    -- filter=45 channel=76
    0, 8, -6, 3, -2, -5, -2, 4, -4,
    -- filter=45 channel=77
    3, 5, -1, 6, -6, 4, -7, 0, 0,
    -- filter=45 channel=78
    4, 3, 3, 4, -6, -3, 1, 2, -4,
    -- filter=45 channel=79
    10, -2, -5, 5, 1, -10, -3, 4, -2,
    -- filter=45 channel=80
    4, -7, -8, -3, -5, -6, 2, 2, 3,
    -- filter=45 channel=81
    4, 3, -1, -2, 4, -6, 4, -6, -1,
    -- filter=45 channel=82
    2, -2, 0, -4, 2, -3, 0, 3, 0,
    -- filter=45 channel=83
    -6, -2, 0, -1, 3, 1, 2, -1, 1,
    -- filter=45 channel=84
    7, 3, -4, 2, -7, -1, 1, 2, 5,
    -- filter=45 channel=85
    0, 6, -2, -4, 6, -4, 3, -1, 2,
    -- filter=45 channel=86
    5, -7, 0, -6, -1, 5, 4, 1, -6,
    -- filter=45 channel=87
    2, 2, 0, 5, -4, 3, -4, -5, -6,
    -- filter=45 channel=88
    -1, -3, 2, -6, -5, 6, 4, 8, -5,
    -- filter=45 channel=89
    3, 6, 0, 7, 3, 4, 4, -4, 1,
    -- filter=45 channel=90
    0, -5, -2, 1, 7, 2, 6, 0, 7,
    -- filter=45 channel=91
    -5, 3, 3, 4, -2, 0, 0, -7, -4,
    -- filter=45 channel=92
    -3, -4, -3, -4, -1, 3, 7, 3, 3,
    -- filter=45 channel=93
    0, 2, -2, -7, 1, -3, 0, 0, -2,
    -- filter=45 channel=94
    -5, -3, 1, 0, 4, -5, 0, 4, 0,
    -- filter=45 channel=95
    6, 1, 0, 5, -4, -6, -1, -5, 4,
    -- filter=45 channel=96
    7, 2, 0, 0, -1, 0, -2, 0, 0,
    -- filter=45 channel=97
    2, 7, 0, 2, 6, 6, -1, 3, -2,
    -- filter=45 channel=98
    1, -1, 3, -6, -3, 5, -2, 0, 2,
    -- filter=45 channel=99
    1, -1, -6, -5, -9, -6, -3, -4, -3,
    -- filter=45 channel=100
    -2, 4, 3, -6, 0, 0, -5, -3, -3,
    -- filter=45 channel=101
    1, -3, 7, -5, -2, 6, 5, -1, 0,
    -- filter=45 channel=102
    -4, -4, 6, -4, -7, 4, -6, -1, 0,
    -- filter=45 channel=103
    4, 4, -5, 8, 4, -5, -1, -7, 1,
    -- filter=45 channel=104
    7, 1, 0, 5, 3, 2, -3, 3, -3,
    -- filter=45 channel=105
    6, -4, -3, -7, -3, 8, 4, -5, -2,
    -- filter=45 channel=106
    6, -4, 5, -1, 6, 4, 0, -5, -1,
    -- filter=45 channel=107
    2, -4, 1, -4, 0, 2, -4, 2, 4,
    -- filter=45 channel=108
    -5, -4, -4, 0, -1, 0, 0, -1, -6,
    -- filter=45 channel=109
    -3, -1, 0, 0, 0, -2, -4, 0, -4,
    -- filter=45 channel=110
    -1, -5, 6, 0, 0, 5, 3, -3, -1,
    -- filter=45 channel=111
    0, 0, -1, -3, 1, -4, 2, -6, -3,
    -- filter=45 channel=112
    3, 1, -2, 1, -1, 5, 3, -7, -2,
    -- filter=45 channel=113
    0, 5, 1, 2, -1, 4, -5, -1, 3,
    -- filter=45 channel=114
    4, -1, 0, 6, -6, -6, 2, -3, 2,
    -- filter=45 channel=115
    -7, 0, 3, -5, -3, 2, 1, 7, -3,
    -- filter=45 channel=116
    -1, -2, -9, 2, 0, -8, 3, -3, -7,
    -- filter=45 channel=117
    7, 4, -5, 5, -7, -4, 6, -4, 0,
    -- filter=45 channel=118
    -3, 3, 2, 1, -5, 0, 5, -5, -1,
    -- filter=45 channel=119
    -1, -3, 4, 6, -1, 3, 6, 5, 6,
    -- filter=45 channel=120
    7, -2, 4, -3, -3, 0, -6, 3, -3,
    -- filter=45 channel=121
    -3, -2, -8, -4, 3, -7, -4, 4, -3,
    -- filter=45 channel=122
    4, -3, -6, -4, 1, -7, 2, 0, 3,
    -- filter=45 channel=123
    -6, 6, -1, 3, -3, 3, 0, 2, -5,
    -- filter=45 channel=124
    -6, 0, -4, 0, 4, -3, 0, 2, 5,
    -- filter=45 channel=125
    7, 0, -3, 1, 1, -7, 0, 2, 5,
    -- filter=45 channel=126
    8, 4, -1, 0, 5, -2, 8, -7, -3,
    -- filter=45 channel=127
    5, 0, 2, 7, 4, 0, -2, -3, -2,
    -- filter=46 channel=0
    -3, 0, -7, 0, 2, 1, 6, -6, -6,
    -- filter=46 channel=1
    0, -1, -7, 6, -1, 4, -6, 0, 0,
    -- filter=46 channel=2
    -3, 0, 6, -4, 0, -3, -5, 5, 5,
    -- filter=46 channel=3
    5, -7, 6, 7, -4, 6, 6, -4, -7,
    -- filter=46 channel=4
    -6, -3, 1, 2, -4, -5, -1, 0, 3,
    -- filter=46 channel=5
    -4, 1, 4, -5, 2, -6, -4, -2, 0,
    -- filter=46 channel=6
    -4, 6, 1, 5, -1, -4, -1, 4, -2,
    -- filter=46 channel=7
    -7, -1, -5, 0, -4, 6, 2, -2, -1,
    -- filter=46 channel=8
    -3, -5, 3, -3, -6, 2, 2, 5, -4,
    -- filter=46 channel=9
    0, 0, 6, 7, 1, 6, 2, 7, -6,
    -- filter=46 channel=10
    -7, -1, -2, 6, 3, -3, 7, 0, 1,
    -- filter=46 channel=11
    -5, 3, -5, 1, -6, -7, 1, 6, 4,
    -- filter=46 channel=12
    -1, 3, 3, -5, 4, 5, 2, -2, 0,
    -- filter=46 channel=13
    -5, -7, 2, 1, -2, -4, -2, -2, 6,
    -- filter=46 channel=14
    -7, 4, -6, -7, 2, -3, -7, 6, -1,
    -- filter=46 channel=15
    -2, 4, -6, 7, 6, 2, 0, 6, 4,
    -- filter=46 channel=16
    -3, -3, 5, -5, -4, -3, 0, -3, 2,
    -- filter=46 channel=17
    3, 0, -4, -4, 0, 5, 6, 6, 2,
    -- filter=46 channel=18
    3, 0, 6, 1, 4, -2, 2, -1, 4,
    -- filter=46 channel=19
    -4, -5, 5, -4, 1, 0, -2, -4, -4,
    -- filter=46 channel=20
    3, 5, -6, 0, -5, 7, 6, -5, -2,
    -- filter=46 channel=21
    -5, -4, 6, -7, -1, -4, -2, -1, 4,
    -- filter=46 channel=22
    -4, -3, -5, 0, 3, -5, -2, -5, -2,
    -- filter=46 channel=23
    -1, 0, 0, 0, 5, -2, 2, -6, -1,
    -- filter=46 channel=24
    0, 0, -2, -3, 1, 2, 1, -6, -3,
    -- filter=46 channel=25
    3, 1, -2, -6, -5, 5, -1, -4, -3,
    -- filter=46 channel=26
    4, 3, -4, 3, 0, 1, 4, -4, 0,
    -- filter=46 channel=27
    -7, 6, -3, 0, -3, -1, 2, -1, -1,
    -- filter=46 channel=28
    -2, 2, 2, 4, -2, 2, -3, 2, -5,
    -- filter=46 channel=29
    -7, 4, 2, -5, 4, -1, -7, -2, -3,
    -- filter=46 channel=30
    1, -4, 0, 0, -2, 4, 3, -3, -3,
    -- filter=46 channel=31
    1, -4, -2, -3, -2, 3, 6, -5, 3,
    -- filter=46 channel=32
    -7, 0, 6, 3, 5, -5, -6, -4, -7,
    -- filter=46 channel=33
    2, -7, 5, -1, 3, 7, 0, -2, 4,
    -- filter=46 channel=34
    5, -3, 6, 1, 2, -6, 0, -1, -1,
    -- filter=46 channel=35
    -5, -3, -6, -1, -5, 3, 4, 4, 6,
    -- filter=46 channel=36
    4, -1, 3, -3, -6, 5, -2, 3, 6,
    -- filter=46 channel=37
    -5, -4, 4, -1, 1, -4, -4, -3, -1,
    -- filter=46 channel=38
    1, -1, -3, 0, -5, 5, -2, 0, -2,
    -- filter=46 channel=39
    -5, 1, 4, -3, -2, -1, 2, -1, 2,
    -- filter=46 channel=40
    4, 2, -2, -5, 5, 0, 6, -3, 7,
    -- filter=46 channel=41
    -1, -1, -6, 0, 4, -6, 0, -4, 0,
    -- filter=46 channel=42
    4, 0, 3, -1, 6, -1, 0, 0, 1,
    -- filter=46 channel=43
    -4, 2, 2, -6, -1, 2, 1, 4, 5,
    -- filter=46 channel=44
    0, 1, -4, 2, 7, -5, -3, -4, 5,
    -- filter=46 channel=45
    7, 7, 6, 1, -2, 0, 5, 0, 0,
    -- filter=46 channel=46
    -4, -7, 5, -1, -3, -5, 3, 6, -6,
    -- filter=46 channel=47
    -4, -6, 0, 1, -6, 2, -6, -1, 2,
    -- filter=46 channel=48
    2, 0, 0, 2, -3, -4, 4, 0, 7,
    -- filter=46 channel=49
    2, -5, 0, 0, 1, -5, -4, 3, -5,
    -- filter=46 channel=50
    -7, -4, -7, 3, 0, 2, 4, 4, 5,
    -- filter=46 channel=51
    -1, -4, 5, 2, 5, 4, 4, 6, -2,
    -- filter=46 channel=52
    3, 4, 6, -5, 5, -5, -3, 4, -2,
    -- filter=46 channel=53
    -2, -1, -3, 3, 7, 5, 5, -7, 4,
    -- filter=46 channel=54
    2, 4, -1, 1, 6, -4, -5, 0, 5,
    -- filter=46 channel=55
    -5, 6, 4, 0, -5, 4, -7, -4, 0,
    -- filter=46 channel=56
    7, -2, -1, -6, 1, -2, 6, 7, 0,
    -- filter=46 channel=57
    5, -2, -4, -6, -1, -3, 2, 1, 0,
    -- filter=46 channel=58
    2, -2, 5, 5, 2, 4, 0, 0, -1,
    -- filter=46 channel=59
    -1, -1, -4, 3, -5, 0, 0, 3, 1,
    -- filter=46 channel=60
    0, 0, 2, 6, 7, 5, -5, 0, 6,
    -- filter=46 channel=61
    -1, -2, -3, -6, 1, -7, -7, 5, 4,
    -- filter=46 channel=62
    -4, 4, 1, 0, -5, -7, 5, 7, 1,
    -- filter=46 channel=63
    1, 4, 2, 3, 0, -4, 2, -7, 2,
    -- filter=46 channel=64
    2, 4, 2, 4, 4, -1, -2, 5, 3,
    -- filter=46 channel=65
    -1, 1, -3, 2, 1, -3, 0, -6, 1,
    -- filter=46 channel=66
    -1, -4, -6, -4, -1, 5, 4, 3, -2,
    -- filter=46 channel=67
    -7, 2, 2, -6, 1, -1, -6, -2, -6,
    -- filter=46 channel=68
    3, -6, -2, 0, -5, 3, 0, 0, 3,
    -- filter=46 channel=69
    -5, -3, 3, -3, 0, -3, 1, 7, 0,
    -- filter=46 channel=70
    4, 0, 2, 1, 0, -4, -5, 1, -4,
    -- filter=46 channel=71
    -1, 1, 5, 3, 2, 0, 6, -7, 3,
    -- filter=46 channel=72
    -6, -1, 0, 7, 0, -1, 6, 6, 0,
    -- filter=46 channel=73
    -2, -1, -4, -4, 3, -4, -3, -1, 3,
    -- filter=46 channel=74
    6, -1, -7, 4, -7, -5, 4, -1, 4,
    -- filter=46 channel=75
    0, 3, 4, -3, -4, 3, 0, 6, -2,
    -- filter=46 channel=76
    -6, 5, 0, 2, -6, -4, 0, -2, 1,
    -- filter=46 channel=77
    -5, 5, 2, 0, -6, 0, -7, 2, -1,
    -- filter=46 channel=78
    -4, 5, -6, 4, 2, 5, 0, -2, 2,
    -- filter=46 channel=79
    -5, -3, -2, 3, 3, 2, 4, 4, 2,
    -- filter=46 channel=80
    2, 4, 0, -6, 4, -3, -3, 3, 6,
    -- filter=46 channel=81
    0, -3, -4, 0, -1, -3, 3, -7, 1,
    -- filter=46 channel=82
    4, 2, 1, -2, 1, 4, -3, -4, 6,
    -- filter=46 channel=83
    1, 4, 4, -2, 2, -1, 1, -5, -1,
    -- filter=46 channel=84
    5, 7, -1, -5, -5, 5, -4, 5, -6,
    -- filter=46 channel=85
    5, -3, 5, -2, 7, -6, 0, -3, 1,
    -- filter=46 channel=86
    -5, -5, 0, 0, 6, 0, -2, 4, -2,
    -- filter=46 channel=87
    1, 3, 4, 5, -2, 3, -4, -4, 3,
    -- filter=46 channel=88
    -3, 1, 0, 0, 0, -6, -3, 4, 3,
    -- filter=46 channel=89
    -4, -6, -4, 0, -4, 5, 0, -3, -5,
    -- filter=46 channel=90
    0, -5, 3, -1, -5, -7, 0, 4, 1,
    -- filter=46 channel=91
    2, 3, 6, -1, -2, -5, 0, -6, 1,
    -- filter=46 channel=92
    3, -4, 6, 5, -1, 3, 5, 3, -6,
    -- filter=46 channel=93
    5, -3, -4, -1, -4, -3, 6, -1, 0,
    -- filter=46 channel=94
    0, -4, 5, -1, -2, -1, 0, 4, -1,
    -- filter=46 channel=95
    2, 4, -3, -4, 3, -7, 6, -5, 4,
    -- filter=46 channel=96
    2, -7, -1, -3, 1, -5, 1, 4, -4,
    -- filter=46 channel=97
    0, 4, 2, -6, 0, -2, -1, 6, 5,
    -- filter=46 channel=98
    2, 4, -1, 1, 3, 3, 1, 6, 6,
    -- filter=46 channel=99
    6, -5, -4, -6, -4, 3, -2, 3, -6,
    -- filter=46 channel=100
    4, 0, -3, -7, -4, -6, 7, 4, 2,
    -- filter=46 channel=101
    5, 6, -6, 1, 2, 3, 6, -7, -2,
    -- filter=46 channel=102
    -1, -6, -3, 0, -3, 3, -1, 5, -3,
    -- filter=46 channel=103
    -1, -2, -6, 3, -5, 4, 5, 0, -2,
    -- filter=46 channel=104
    -5, 3, 5, -3, 3, 2, 0, 1, -1,
    -- filter=46 channel=105
    -3, -5, 0, 4, 0, -2, 0, -1, 0,
    -- filter=46 channel=106
    2, -1, -6, -4, -3, 5, 3, 1, -3,
    -- filter=46 channel=107
    2, 3, 0, -6, 3, -1, -5, 4, -7,
    -- filter=46 channel=108
    -4, 5, 0, 0, 0, -2, -5, 5, 4,
    -- filter=46 channel=109
    -3, -3, -2, 5, -5, -7, -2, -6, -2,
    -- filter=46 channel=110
    2, 0, 0, -6, -4, 3, -7, 1, -5,
    -- filter=46 channel=111
    -6, -3, -1, 0, -2, -5, 0, -5, -7,
    -- filter=46 channel=112
    -6, 2, -7, 0, -2, -7, -5, 1, -2,
    -- filter=46 channel=113
    0, 4, -5, -1, 5, 4, -1, 6, 2,
    -- filter=46 channel=114
    -5, -1, 0, 4, -3, -4, -1, -1, 4,
    -- filter=46 channel=115
    -7, -2, -7, 3, 0, 0, 4, 1, 0,
    -- filter=46 channel=116
    4, 3, 0, 5, 4, -1, 5, -4, 5,
    -- filter=46 channel=117
    0, 3, 6, -3, 1, 0, 2, -4, -3,
    -- filter=46 channel=118
    -2, 1, 0, 4, 1, -2, 0, 1, 5,
    -- filter=46 channel=119
    7, 7, -4, 4, -2, 0, 7, 6, 2,
    -- filter=46 channel=120
    -5, 4, 2, -7, -7, 6, -4, -4, -7,
    -- filter=46 channel=121
    -2, -4, -6, 3, 3, -4, 7, 5, 0,
    -- filter=46 channel=122
    0, -1, -4, -6, 2, -5, 1, 6, 4,
    -- filter=46 channel=123
    5, 0, -6, 4, 7, -2, -3, -2, 6,
    -- filter=46 channel=124
    4, 0, -5, -2, 0, -5, -2, 2, -4,
    -- filter=46 channel=125
    -3, -2, 5, -1, -7, -4, -3, 0, -4,
    -- filter=46 channel=126
    6, 7, 2, 5, 1, 0, -3, 2, 3,
    -- filter=46 channel=127
    2, 7, 5, 3, 2, 2, -5, -5, 0,
    -- filter=47 channel=0
    1, -2, -19, 17, 5, -12, 5, 7, -1,
    -- filter=47 channel=1
    9, -13, -13, 22, 0, -20, 10, -7, -5,
    -- filter=47 channel=2
    1, -1, 5, 2, -6, 4, 0, 1, 6,
    -- filter=47 channel=3
    0, 0, -9, 3, -15, -3, -4, -7, -9,
    -- filter=47 channel=4
    11, -9, -3, 2, -11, -15, 1, 2, 0,
    -- filter=47 channel=5
    1, -19, -23, 22, -9, -23, 12, 0, -3,
    -- filter=47 channel=6
    -2, 7, 0, -4, -1, 5, -9, -4, 2,
    -- filter=47 channel=7
    -7, 1, -5, -6, 7, -4, 0, 2, 7,
    -- filter=47 channel=8
    1, 1, 0, 4, -2, -12, -3, -1, 0,
    -- filter=47 channel=9
    3, 3, -4, 3, 0, -11, -1, 0, -3,
    -- filter=47 channel=10
    6, 0, -7, 5, -5, -6, 2, -2, -13,
    -- filter=47 channel=11
    -5, 2, 7, -18, 3, 15, -4, -8, 8,
    -- filter=47 channel=12
    4, 5, -4, 3, 3, -7, 1, 0, 1,
    -- filter=47 channel=13
    -2, 12, -4, -3, 0, 0, -8, -1, 6,
    -- filter=47 channel=14
    6, 3, -4, 5, 2, 6, -1, -5, -7,
    -- filter=47 channel=15
    -7, -5, 1, -11, 5, 17, -7, -6, 6,
    -- filter=47 channel=16
    11, -3, -18, 24, 3, -18, 12, -1, -20,
    -- filter=47 channel=17
    2, 0, -3, 6, -4, 2, -6, 7, 4,
    -- filter=47 channel=18
    8, -2, 14, -9, -1, 25, -10, 0, 23,
    -- filter=47 channel=19
    -4, 3, -3, -2, -2, 0, -1, -3, 0,
    -- filter=47 channel=20
    -8, 10, 13, -34, 3, 27, -19, -6, 5,
    -- filter=47 channel=21
    15, -2, -19, 21, 4, -24, 18, -1, -8,
    -- filter=47 channel=22
    1, 0, -4, -1, 4, 4, 0, 1, 0,
    -- filter=47 channel=23
    -8, -4, 2, -12, 0, 1, -13, -4, -9,
    -- filter=47 channel=24
    -2, 1, 6, 7, 4, -1, 0, 2, -5,
    -- filter=47 channel=25
    16, -3, -5, 5, -5, -8, 5, 8, 3,
    -- filter=47 channel=26
    4, -3, -10, 13, 8, -4, 1, -1, -8,
    -- filter=47 channel=27
    9, -8, -5, 2, 6, -2, -1, 0, 7,
    -- filter=47 channel=28
    1, -4, 3, 0, -2, 5, 4, 5, 3,
    -- filter=47 channel=29
    -9, -7, 18, -20, -4, 18, -17, -8, 6,
    -- filter=47 channel=30
    3, -10, -6, 15, -5, -4, 13, 1, 0,
    -- filter=47 channel=31
    14, -4, -5, 16, 3, -18, 11, 5, -14,
    -- filter=47 channel=32
    4, 4, 1, -11, 11, 9, 0, 1, 3,
    -- filter=47 channel=33
    8, -5, -7, 7, 1, -10, -4, 10, -4,
    -- filter=47 channel=34
    2, 5, 3, 12, -5, 0, 4, -1, 0,
    -- filter=47 channel=35
    -7, 5, -5, 1, 4, 3, -2, 3, 4,
    -- filter=47 channel=36
    9, 6, 0, 3, 3, -5, 8, 5, 0,
    -- filter=47 channel=37
    2, -12, -28, 23, -6, -29, 12, 6, -18,
    -- filter=47 channel=38
    0, 0, 4, 5, 1, -3, -2, -4, 0,
    -- filter=47 channel=39
    -11, 10, 8, -8, -1, 11, 1, 3, 12,
    -- filter=47 channel=40
    -2, 5, 1, -8, 2, 9, -3, -1, 6,
    -- filter=47 channel=41
    27, 16, 4, 26, 0, 1, 18, 3, -3,
    -- filter=47 channel=42
    -2, 5, -8, 1, 3, -7, 0, 10, 1,
    -- filter=47 channel=43
    -3, -1, 4, -3, -10, 4, -5, -8, -1,
    -- filter=47 channel=44
    3, -14, -18, 20, 5, -24, 13, 4, -16,
    -- filter=47 channel=45
    -8, -1, 6, 5, 6, 8, 0, 3, 5,
    -- filter=47 channel=46
    -2, 3, 2, 0, -3, -6, -4, 4, 1,
    -- filter=47 channel=47
    18, -6, -22, 28, 1, -34, 10, 0, -18,
    -- filter=47 channel=48
    18, -11, -14, 21, 5, -29, 17, 5, -7,
    -- filter=47 channel=49
    -6, -7, 0, -13, 8, 13, 0, 6, 4,
    -- filter=47 channel=50
    -2, -11, -2, 8, 1, -11, 4, -3, -3,
    -- filter=47 channel=51
    -2, 0, 6, -3, 2, 3, -1, -6, 3,
    -- filter=47 channel=52
    4, 2, 2, 0, -8, -7, -1, -9, 1,
    -- filter=47 channel=53
    -10, 7, 4, -11, 0, 9, 0, 0, 5,
    -- filter=47 channel=54
    -4, 4, 1, 4, 7, 5, 6, 5, 1,
    -- filter=47 channel=55
    -9, -3, 5, -11, 1, 20, -8, 3, 7,
    -- filter=47 channel=56
    2, -1, -8, 0, 4, -3, 10, -6, -5,
    -- filter=47 channel=57
    7, 0, -1, -1, -2, -5, 7, -2, 0,
    -- filter=47 channel=58
    7, -9, -9, 4, -1, -3, -4, 3, -8,
    -- filter=47 channel=59
    18, 7, -8, 5, -3, -6, 12, -1, 0,
    -- filter=47 channel=60
    -4, -2, 0, 6, 0, -3, -3, -3, -2,
    -- filter=47 channel=61
    0, -5, 0, -5, -1, -4, 7, -2, 4,
    -- filter=47 channel=62
    -1, 1, -3, -7, 1, -5, -2, -2, 0,
    -- filter=47 channel=63
    -2, -2, -5, 15, -2, -8, 0, 0, 0,
    -- filter=47 channel=64
    -3, -1, -5, -3, 7, -4, 7, 5, -3,
    -- filter=47 channel=65
    6, 4, 0, -4, 3, 5, -6, 7, 0,
    -- filter=47 channel=66
    3, 13, 5, 1, 2, 0, 8, -2, 0,
    -- filter=47 channel=67
    -6, 2, 3, -2, -4, -5, -1, 0, -3,
    -- filter=47 channel=68
    1, 5, 0, 0, 0, 2, 0, -4, 9,
    -- filter=47 channel=69
    -6, 6, -6, 2, 0, 0, 0, 3, 5,
    -- filter=47 channel=70
    0, -4, 4, -11, 7, 6, -7, 2, 3,
    -- filter=47 channel=71
    -5, 0, 5, 3, -3, -6, -6, 3, -10,
    -- filter=47 channel=72
    6, 7, 0, 9, -5, -14, 7, 2, -7,
    -- filter=47 channel=73
    3, 5, 0, -6, -1, 8, -5, 0, 7,
    -- filter=47 channel=74
    11, -8, -4, 0, 0, -11, 4, -2, -4,
    -- filter=47 channel=75
    20, -6, -28, 25, 6, -14, 1, -4, -3,
    -- filter=47 channel=76
    -11, 1, 23, -23, 0, 18, -8, 0, 9,
    -- filter=47 channel=77
    6, 3, -5, 4, -5, -1, 6, 0, -1,
    -- filter=47 channel=78
    10, 3, -9, 8, 7, -10, 2, -3, -9,
    -- filter=47 channel=79
    1, 0, 14, -7, 7, 21, -11, 0, 10,
    -- filter=47 channel=80
    18, -5, -10, 27, 2, -29, 15, 11, -15,
    -- filter=47 channel=81
    -4, 5, 5, 3, 6, -3, -5, 1, -2,
    -- filter=47 channel=82
    -6, 5, 5, -6, 0, -7, 3, 0, -6,
    -- filter=47 channel=83
    10, -6, 1, -2, -8, -6, 6, 7, 0,
    -- filter=47 channel=84
    4, 4, 4, -16, 7, 3, -4, -3, 11,
    -- filter=47 channel=85
    5, -7, 2, 4, 0, 3, 4, 5, 3,
    -- filter=47 channel=86
    8, -1, 1, 0, 2, -1, 10, 5, 0,
    -- filter=47 channel=87
    1, 1, 0, -15, 7, 8, 0, 4, 7,
    -- filter=47 channel=88
    1, 1, 3, 1, 7, -5, 3, -5, -1,
    -- filter=47 channel=89
    4, 2, 1, -8, 5, -6, -4, 1, 1,
    -- filter=47 channel=90
    2, 4, 0, 5, 3, -5, 3, -1, -7,
    -- filter=47 channel=91
    0, 0, 6, -17, 5, 3, 0, 8, 2,
    -- filter=47 channel=92
    -4, -7, 7, 2, -1, 1, 9, 0, -2,
    -- filter=47 channel=93
    11, -12, -26, 26, 0, -33, 17, 0, -15,
    -- filter=47 channel=94
    2, -2, 1, -1, 3, -1, -2, -5, 2,
    -- filter=47 channel=95
    7, 2, -1, 6, 6, -6, 3, -1, -2,
    -- filter=47 channel=96
    0, -6, 7, -4, 3, 0, -1, 1, 7,
    -- filter=47 channel=97
    3, -4, -2, 5, 0, -10, 2, -7, -4,
    -- filter=47 channel=98
    9, 5, -8, 12, -1, -20, 4, 6, -1,
    -- filter=47 channel=99
    1, 3, -4, -2, -4, -19, 2, 0, -7,
    -- filter=47 channel=100
    -2, -1, 0, 0, -1, 7, -3, -5, 0,
    -- filter=47 channel=101
    -4, 3, 5, -3, -10, -1, -3, -10, 1,
    -- filter=47 channel=102
    -7, -3, 0, 1, -4, 6, -6, 3, -1,
    -- filter=47 channel=103
    17, -8, -22, 28, 0, -28, 9, 0, -16,
    -- filter=47 channel=104
    10, -3, -18, 16, 4, -23, 10, 8, -8,
    -- filter=47 channel=105
    -10, -6, 14, -19, 3, 9, -5, 0, 0,
    -- filter=47 channel=106
    9, 0, 5, -8, -5, 11, 6, 0, 9,
    -- filter=47 channel=107
    -1, 0, 3, -19, 6, 13, -14, 2, 8,
    -- filter=47 channel=108
    6, 5, -2, 8, 4, -6, 1, -6, 5,
    -- filter=47 channel=109
    1, 1, 1, -1, -6, -6, 0, 0, 3,
    -- filter=47 channel=110
    0, 6, -3, -3, -1, -5, 7, 0, -9,
    -- filter=47 channel=111
    0, 2, 0, 6, -8, 0, 2, -4, 0,
    -- filter=47 channel=112
    10, -6, -2, 11, 0, -16, 4, -5, 3,
    -- filter=47 channel=113
    3, -1, -1, 3, -5, -15, 12, 0, 1,
    -- filter=47 channel=114
    7, -8, 10, -8, 4, 14, -3, 7, 19,
    -- filter=47 channel=115
    0, 0, -6, -7, 2, -2, -5, 3, 4,
    -- filter=47 channel=116
    9, 0, -4, 2, 5, -5, 7, 6, -2,
    -- filter=47 channel=117
    2, 0, 5, 3, 0, -2, 3, 0, 0,
    -- filter=47 channel=118
    6, 0, 3, 6, 0, 2, -2, -2, 4,
    -- filter=47 channel=119
    6, 0, 0, 3, 1, 2, 6, -9, -8,
    -- filter=47 channel=120
    -10, -8, 0, -20, -2, -9, -2, -4, 5,
    -- filter=47 channel=121
    5, 2, -7, 2, -6, -9, 7, 0, -11,
    -- filter=47 channel=122
    18, -15, -30, 40, 5, -44, 26, 6, -33,
    -- filter=47 channel=123
    8, -6, -1, 0, 0, -1, 0, 4, -9,
    -- filter=47 channel=124
    -3, 2, 2, -18, 2, 10, -9, 0, -3,
    -- filter=47 channel=125
    4, -3, -3, 10, 5, -10, 4, 12, 4,
    -- filter=47 channel=126
    1, -1, 4, 0, 4, 2, -7, -9, -8,
    -- filter=47 channel=127
    4, 7, 0, 0, -6, 0, -2, -2, 1,
    -- filter=48 channel=0
    1, -3, -15, -1, 5, -12, -1, 6, -4,
    -- filter=48 channel=1
    3, 7, -10, 0, 6, -6, 1, -3, -8,
    -- filter=48 channel=2
    -1, -5, 5, 6, 3, -6, 1, -3, -2,
    -- filter=48 channel=3
    0, -5, 0, -3, -9, -1, -2, -10, 0,
    -- filter=48 channel=4
    1, -1, 3, 4, -10, 3, -2, -5, 0,
    -- filter=48 channel=5
    0, 0, 3, 1, 5, -5, 4, 10, 8,
    -- filter=48 channel=6
    -1, -1, 0, 13, -5, -3, 7, 0, -9,
    -- filter=48 channel=7
    -6, 3, 7, 4, -2, 1, 1, -6, -2,
    -- filter=48 channel=8
    -1, -5, -1, 0, -4, 0, 4, -6, 2,
    -- filter=48 channel=9
    -1, 1, 7, -11, 1, -2, 3, 4, 1,
    -- filter=48 channel=10
    4, -4, -5, 0, -4, -5, 0, 0, -6,
    -- filter=48 channel=11
    4, 6, 1, 7, -2, 8, 3, -1, 3,
    -- filter=48 channel=12
    8, -1, -5, 3, 2, -10, 9, -5, 1,
    -- filter=48 channel=13
    3, -10, -8, 0, -9, 0, 8, 2, -2,
    -- filter=48 channel=14
    0, -2, -2, 1, -2, -4, -3, -6, 6,
    -- filter=48 channel=15
    7, -1, -4, 14, -4, 0, 9, -4, -5,
    -- filter=48 channel=16
    1, -6, -7, -4, -2, 0, -2, 0, 2,
    -- filter=48 channel=17
    7, -3, 4, 1, -3, -4, -6, 4, 7,
    -- filter=48 channel=18
    5, 3, -4, 15, 5, -13, 5, 4, -5,
    -- filter=48 channel=19
    5, -2, 0, 1, 0, 7, 1, 1, -2,
    -- filter=48 channel=20
    6, -6, 4, 17, 8, -4, 10, -4, -12,
    -- filter=48 channel=21
    -18, -4, -6, -20, -9, -2, -15, 0, 10,
    -- filter=48 channel=22
    3, 4, 3, 3, 3, -2, 7, -2, -3,
    -- filter=48 channel=23
    -1, -5, 14, 2, -1, 5, 1, -6, 3,
    -- filter=48 channel=24
    -5, 6, -7, -3, 1, 7, -7, -3, -5,
    -- filter=48 channel=25
    4, 2, 0, 4, 0, 0, -4, -7, -3,
    -- filter=48 channel=26
    -5, 1, -4, -7, -6, 2, -9, -7, -2,
    -- filter=48 channel=27
    6, -3, 5, 7, -5, -7, 4, -3, -2,
    -- filter=48 channel=28
    6, -5, 0, 5, 5, 2, 4, 0, 0,
    -- filter=48 channel=29
    0, -1, 7, 17, 8, -7, 1, -5, -14,
    -- filter=48 channel=30
    -2, 8, 4, 0, 1, -7, -1, -5, 4,
    -- filter=48 channel=31
    -14, -5, 8, -25, -7, 8, -20, -3, 13,
    -- filter=48 channel=32
    -1, 4, -6, 13, 3, -3, 2, 0, -5,
    -- filter=48 channel=33
    6, -1, 2, -7, 3, 3, -1, 0, -1,
    -- filter=48 channel=34
    6, -5, -4, 18, 3, 4, 6, -7, -3,
    -- filter=48 channel=35
    2, 3, 2, 1, 6, -1, -4, 7, -7,
    -- filter=48 channel=36
    2, 2, -2, 1, -1, 3, 5, -8, -1,
    -- filter=48 channel=37
    -7, 10, 0, -7, 8, -7, -3, -3, -1,
    -- filter=48 channel=38
    6, 3, -5, -2, 1, -2, 4, -2, -1,
    -- filter=48 channel=39
    -5, -1, -2, 2, -2, 5, 0, 2, -5,
    -- filter=48 channel=40
    4, -3, -4, 3, 0, -1, 0, -4, 0,
    -- filter=48 channel=41
    8, 1, -6, 17, -2, -13, 14, -8, -10,
    -- filter=48 channel=42
    -3, 3, -3, -8, -4, 1, -9, -7, -2,
    -- filter=48 channel=43
    7, 6, -1, 7, 4, 2, 3, 2, -7,
    -- filter=48 channel=44
    -1, -9, 1, -4, 2, -1, -11, -1, -6,
    -- filter=48 channel=45
    0, -4, 0, 5, 9, -2, -4, 0, 5,
    -- filter=48 channel=46
    7, 6, -2, -2, -4, 0, 9, -7, -1,
    -- filter=48 channel=47
    -17, -1, -9, -16, 1, 2, -10, -9, 5,
    -- filter=48 channel=48
    -10, -8, -5, -6, -4, -7, -8, -10, 5,
    -- filter=48 channel=49
    2, 0, 6, 11, 1, -8, 9, -1, -1,
    -- filter=48 channel=50
    0, 0, 5, -2, -6, 6, 0, 6, 7,
    -- filter=48 channel=51
    0, -1, -6, -1, -3, 3, -3, -7, 1,
    -- filter=48 channel=52
    -2, -8, -4, 4, -6, 3, 6, -9, -4,
    -- filter=48 channel=53
    5, 4, 1, 9, -2, 6, 5, 4, 3,
    -- filter=48 channel=54
    2, 2, 4, 0, 7, 2, -5, -4, 6,
    -- filter=48 channel=55
    8, -9, 1, 15, 4, -4, 5, -5, -5,
    -- filter=48 channel=56
    4, -3, 0, 7, 4, 0, -2, -5, -5,
    -- filter=48 channel=57
    -4, 0, -1, 6, 1, -4, 8, -4, -7,
    -- filter=48 channel=58
    7, -1, -5, -4, 0, 6, 0, 8, 8,
    -- filter=48 channel=59
    -6, 0, 2, -5, -10, 0, -2, -10, -6,
    -- filter=48 channel=60
    -2, -7, 5, 0, 3, 4, 4, -7, 0,
    -- filter=48 channel=61
    5, -3, -6, 5, -5, -8, -5, -2, 2,
    -- filter=48 channel=62
    -6, 5, -7, -4, -6, -2, 1, -1, 0,
    -- filter=48 channel=63
    -1, 6, -1, -3, 3, 1, -3, 1, -2,
    -- filter=48 channel=64
    -6, 0, 2, 6, -8, 0, -8, -3, -3,
    -- filter=48 channel=65
    3, 0, -1, 6, 6, 1, -2, -4, 6,
    -- filter=48 channel=66
    -3, -9, -9, -1, -10, -3, 9, -1, -12,
    -- filter=48 channel=67
    5, 6, 0, -6, 3, -2, -5, -3, -5,
    -- filter=48 channel=68
    -6, 5, 7, -1, -3, -3, 5, -3, 0,
    -- filter=48 channel=69
    -4, -3, -7, 6, -8, 7, -5, 4, 2,
    -- filter=48 channel=70
    -3, -1, 7, 7, -1, -5, 0, -2, -2,
    -- filter=48 channel=71
    2, 5, -2, -7, -6, -2, -2, -7, 1,
    -- filter=48 channel=72
    -5, -1, 0, -9, 0, 7, -1, 1, 0,
    -- filter=48 channel=73
    2, -6, -5, -1, 3, -1, 4, -6, 2,
    -- filter=48 channel=74
    3, -4, 7, -4, -7, 3, 6, -3, -6,
    -- filter=48 channel=75
    4, -2, -14, -1, 3, -3, 1, -5, 0,
    -- filter=48 channel=76
    1, -5, 0, 8, 1, 1, 5, -5, -8,
    -- filter=48 channel=77
    -4, 3, 4, -6, -7, 6, -1, 4, 5,
    -- filter=48 channel=78
    -8, -4, 5, 2, -4, 0, 1, -4, -4,
    -- filter=48 channel=79
    9, 0, -12, 7, 6, -4, 17, 7, -14,
    -- filter=48 channel=80
    -14, -9, 9, -14, 0, 8, -14, -3, 0,
    -- filter=48 channel=81
    -3, 1, 1, 1, 2, -6, -5, 7, -1,
    -- filter=48 channel=82
    -5, 3, -4, 2, 6, -4, 4, -6, -1,
    -- filter=48 channel=83
    -2, 1, 7, -2, 0, 9, 0, 4, 2,
    -- filter=48 channel=84
    -2, -1, -7, 1, -3, 0, 10, 3, -2,
    -- filter=48 channel=85
    1, -1, -1, 1, -2, 3, -4, 0, -2,
    -- filter=48 channel=86
    5, 4, -4, 0, 1, -5, 8, 1, -7,
    -- filter=48 channel=87
    1, -6, -2, 7, 0, 3, 5, -10, -10,
    -- filter=48 channel=88
    -4, 2, 8, -1, -5, 6, 0, -2, 0,
    -- filter=48 channel=89
    -3, 0, -3, 2, -9, -6, 6, -4, -4,
    -- filter=48 channel=90
    5, -11, 8, -3, -6, 0, -5, -8, 4,
    -- filter=48 channel=91
    -4, -5, 6, 8, -5, -6, 10, 0, -6,
    -- filter=48 channel=92
    8, -2, -2, -4, 1, -1, -3, 2, 5,
    -- filter=48 channel=93
    -9, 0, -8, -4, -9, 4, 1, -4, -4,
    -- filter=48 channel=94
    3, 5, 2, -2, 0, -1, -6, 3, 2,
    -- filter=48 channel=95
    -7, 4, 6, -3, -6, -5, -5, -1, -6,
    -- filter=48 channel=96
    -1, 5, 0, 4, 0, -4, 3, 5, -2,
    -- filter=48 channel=97
    2, 2, 9, -6, 2, 7, -2, 2, 5,
    -- filter=48 channel=98
    -8, 3, -8, -8, -9, -1, -4, 2, -3,
    -- filter=48 channel=99
    -6, -4, 0, 0, 3, 7, 1, -9, 0,
    -- filter=48 channel=100
    5, 4, 6, 8, 1, 1, -2, 6, 0,
    -- filter=48 channel=101
    1, 5, 2, 0, 2, -6, -5, -1, -1,
    -- filter=48 channel=102
    -5, -3, -2, -3, -4, -2, -4, 0, -6,
    -- filter=48 channel=103
    -9, -1, 5, -5, -4, 6, -15, -8, -5,
    -- filter=48 channel=104
    -3, -9, 2, -15, 0, 10, -14, 1, 5,
    -- filter=48 channel=105
    2, 0, 4, 7, 9, 2, 8, -6, -5,
    -- filter=48 channel=106
    6, -2, -2, 9, 0, 3, 5, -4, -8,
    -- filter=48 channel=107
    3, 3, 5, 16, 3, 0, 11, 4, 0,
    -- filter=48 channel=108
    -2, -6, -6, -1, 3, 1, 7, -4, 3,
    -- filter=48 channel=109
    -1, 2, -3, -2, -10, -8, 4, 5, -3,
    -- filter=48 channel=110
    -2, -8, 4, 1, 1, 6, 1, -1, 2,
    -- filter=48 channel=111
    0, 5, -6, 11, -7, 0, 5, -2, -2,
    -- filter=48 channel=112
    7, 1, -5, -1, -7, -4, -1, -2, 2,
    -- filter=48 channel=113
    0, -3, 6, -3, 5, 2, -8, -8, 1,
    -- filter=48 channel=114
    14, 3, -9, 21, 11, -5, 19, 7, -15,
    -- filter=48 channel=115
    -2, -4, 3, 7, -5, 3, -2, 3, -2,
    -- filter=48 channel=116
    2, 1, 7, -4, -2, -2, 7, 1, 5,
    -- filter=48 channel=117
    -3, -3, -2, 3, 0, 6, -3, 2, 2,
    -- filter=48 channel=118
    -4, 6, -5, -2, -3, -4, -5, -2, 0,
    -- filter=48 channel=119
    11, -9, 5, 10, -3, 0, 10, 4, 3,
    -- filter=48 channel=120
    0, 2, 4, 12, -8, 0, 6, 3, 0,
    -- filter=48 channel=121
    6, -9, 0, 3, -3, -4, 0, -11, -8,
    -- filter=48 channel=122
    -16, -15, -5, -20, -12, 5, -11, 0, 0,
    -- filter=48 channel=123
    5, -4, 9, 5, -3, 7, -3, -4, 4,
    -- filter=48 channel=124
    6, -3, 0, 9, -3, -5, -5, -3, -5,
    -- filter=48 channel=125
    0, 3, -1, -11, -8, 2, -3, -5, 7,
    -- filter=48 channel=126
    12, -6, -5, 8, 0, -8, 1, 3, -5,
    -- filter=48 channel=127
    -2, 2, -1, -1, -6, -7, 8, -5, -4,
    -- filter=49 channel=0
    1, 4, -6, 7, -4, -4, -3, 0, 4,
    -- filter=49 channel=1
    3, 0, 6, -1, -3, -2, 1, 2, -1,
    -- filter=49 channel=2
    3, 5, 2, 0, -5, -6, 4, 5, -2,
    -- filter=49 channel=3
    4, 2, -3, 5, 7, -4, 5, -3, 3,
    -- filter=49 channel=4
    0, 0, 7, -2, 3, -6, -3, 3, 7,
    -- filter=49 channel=5
    -1, -4, 3, 0, 3, -4, -1, -1, -7,
    -- filter=49 channel=6
    -2, -1, 1, -3, -1, 7, 3, 4, 0,
    -- filter=49 channel=7
    0, -4, -7, -6, -1, 5, 1, 2, -1,
    -- filter=49 channel=8
    -2, 0, 1, -6, 0, -3, 2, 1, -4,
    -- filter=49 channel=9
    0, 0, 0, -5, -4, 5, 2, 5, -1,
    -- filter=49 channel=10
    -7, 3, 3, 5, -5, 5, -1, -5, 3,
    -- filter=49 channel=11
    -7, 2, -1, -4, -3, 4, 2, 7, 4,
    -- filter=49 channel=12
    5, 0, 6, 5, -3, -1, 1, 5, 6,
    -- filter=49 channel=13
    3, 0, 6, 4, 2, 1, 0, -5, 3,
    -- filter=49 channel=14
    -5, 5, 0, 4, 2, 1, -6, 6, -6,
    -- filter=49 channel=15
    0, 2, -1, 6, -2, -1, -6, 2, -2,
    -- filter=49 channel=16
    0, -1, -2, -4, 1, 2, 2, -7, -1,
    -- filter=49 channel=17
    -4, 0, 2, 4, 6, 6, -1, 6, 4,
    -- filter=49 channel=18
    -6, -2, 1, 2, 6, 4, 5, -1, 4,
    -- filter=49 channel=19
    -1, -3, 0, 5, 0, -6, -1, -5, 0,
    -- filter=49 channel=20
    1, -5, -7, 3, -4, -1, -7, 4, 4,
    -- filter=49 channel=21
    5, 6, -2, -1, -5, 3, -1, -4, 4,
    -- filter=49 channel=22
    3, -7, -3, -6, -7, -6, 3, 1, 3,
    -- filter=49 channel=23
    1, -6, -1, 6, -3, -4, -2, 0, -7,
    -- filter=49 channel=24
    5, -7, -4, -2, -5, -3, 6, 3, 0,
    -- filter=49 channel=25
    -5, -1, -1, 5, -5, 4, 1, 2, 4,
    -- filter=49 channel=26
    1, 5, -2, 1, 5, -6, 2, 0, -1,
    -- filter=49 channel=27
    -6, -2, -4, -6, -5, 0, -6, -5, 3,
    -- filter=49 channel=28
    -7, 1, -3, -4, 1, -6, -2, 4, 3,
    -- filter=49 channel=29
    0, 3, 0, -1, 1, -3, 0, 0, -1,
    -- filter=49 channel=30
    -2, 0, -4, -5, 0, 4, 3, -6, 7,
    -- filter=49 channel=31
    0, 6, 4, -4, -5, -2, 5, 6, 0,
    -- filter=49 channel=32
    -3, 5, 0, -7, -5, 0, 0, 2, 6,
    -- filter=49 channel=33
    3, -5, -4, 2, 5, -6, 4, 7, -1,
    -- filter=49 channel=34
    4, 3, -5, 5, 0, -6, -6, 6, -6,
    -- filter=49 channel=35
    -6, -4, 5, 2, 0, -1, 4, -6, 0,
    -- filter=49 channel=36
    0, 2, -1, -2, -2, 2, -7, -1, -4,
    -- filter=49 channel=37
    0, -1, -5, 3, -5, 5, -3, 0, -6,
    -- filter=49 channel=38
    1, -4, -3, -5, -7, 0, -7, 4, 1,
    -- filter=49 channel=39
    6, -7, 6, -3, 7, -1, -4, 0, -2,
    -- filter=49 channel=40
    -7, -4, -7, -5, -5, 3, -2, 1, -4,
    -- filter=49 channel=41
    6, -2, -5, 5, -5, 6, 2, 4, -4,
    -- filter=49 channel=42
    4, -5, -4, 5, -3, 1, 5, 3, -1,
    -- filter=49 channel=43
    -5, 5, -4, -4, 6, 5, -2, 0, 3,
    -- filter=49 channel=44
    0, -1, 0, 0, 4, -5, 5, -7, 0,
    -- filter=49 channel=45
    0, 3, 1, -5, 0, 6, 1, -3, 0,
    -- filter=49 channel=46
    1, 0, 3, -3, 2, -3, -3, 0, 6,
    -- filter=49 channel=47
    1, 0, 4, 5, -5, 0, -5, 4, -1,
    -- filter=49 channel=48
    6, -5, 0, 1, -3, -2, 4, -3, -7,
    -- filter=49 channel=49
    -7, 6, -5, -3, 5, -5, -4, -3, 2,
    -- filter=49 channel=50
    -3, -1, -5, 4, -3, 6, 2, 1, 0,
    -- filter=49 channel=51
    -5, -3, 3, 6, 3, 5, 3, -5, -4,
    -- filter=49 channel=52
    -1, -6, -3, -2, -6, -1, 5, 4, -5,
    -- filter=49 channel=53
    -2, -3, -3, 1, 1, -6, -3, -4, 3,
    -- filter=49 channel=54
    6, -5, -4, -2, 3, 2, 5, 2, 6,
    -- filter=49 channel=55
    1, -4, 3, 3, 1, -1, -7, -3, 4,
    -- filter=49 channel=56
    0, 0, 5, -4, -6, 5, -4, 0, 2,
    -- filter=49 channel=57
    -1, -5, 4, -3, 5, -4, -4, 1, -4,
    -- filter=49 channel=58
    0, 6, 6, -5, -4, 1, -5, -5, 2,
    -- filter=49 channel=59
    0, 6, -4, 4, 0, 0, -4, -2, 1,
    -- filter=49 channel=60
    -2, -5, 2, -6, -1, -3, 6, 5, -7,
    -- filter=49 channel=61
    4, 1, 0, -2, 4, 4, -5, 5, 6,
    -- filter=49 channel=62
    -3, 7, 5, 0, 0, -5, -4, -1, -2,
    -- filter=49 channel=63
    2, 0, 3, 4, -3, -7, 2, 5, -1,
    -- filter=49 channel=64
    3, 6, 3, -2, 0, 6, 0, -5, 3,
    -- filter=49 channel=65
    -1, -1, -6, -6, 0, 3, -2, -6, 5,
    -- filter=49 channel=66
    -7, 0, 5, -7, -4, -6, -6, 3, 5,
    -- filter=49 channel=67
    2, 7, 4, 2, 0, -5, -5, 3, -3,
    -- filter=49 channel=68
    -6, 5, -7, -3, -1, -3, 5, -2, 0,
    -- filter=49 channel=69
    -1, -4, -5, 1, 6, -2, -1, 5, 2,
    -- filter=49 channel=70
    -4, -6, -1, -5, -7, 2, 4, 1, 2,
    -- filter=49 channel=71
    -1, -2, 2, -6, 0, -3, 3, -7, -5,
    -- filter=49 channel=72
    -2, -2, -2, -5, -5, -2, 3, -4, -6,
    -- filter=49 channel=73
    0, -5, 3, 0, -1, -6, 0, 0, -5,
    -- filter=49 channel=74
    7, 0, -4, 2, 6, 4, 3, -6, 4,
    -- filter=49 channel=75
    6, -2, 5, 5, -6, -6, -1, 6, -1,
    -- filter=49 channel=76
    0, -3, -6, 3, 0, 0, 3, 3, -2,
    -- filter=49 channel=77
    1, -1, -3, -7, -6, 4, -6, 0, -3,
    -- filter=49 channel=78
    5, -1, -5, 1, 2, 0, -4, 5, 3,
    -- filter=49 channel=79
    -1, 1, -4, -3, -3, 2, -2, 5, -5,
    -- filter=49 channel=80
    5, 5, -4, -7, -2, 2, 4, 6, 5,
    -- filter=49 channel=81
    0, 2, 1, 3, 7, 0, -7, 4, 0,
    -- filter=49 channel=82
    4, 3, 2, 0, -6, 0, 0, 2, -2,
    -- filter=49 channel=83
    -2, 0, 5, 0, 3, -1, 6, 7, -2,
    -- filter=49 channel=84
    1, -3, 0, 6, -6, 6, 1, -2, 5,
    -- filter=49 channel=85
    -2, 7, 0, -6, 5, -2, -7, 3, 6,
    -- filter=49 channel=86
    -5, 0, 5, -1, 5, -3, 4, -6, 0,
    -- filter=49 channel=87
    0, 4, -4, -7, -1, 1, -5, -2, -4,
    -- filter=49 channel=88
    3, 4, 4, -1, 7, 0, 4, 0, 0,
    -- filter=49 channel=89
    2, 0, 2, 4, -1, 6, -6, -7, 5,
    -- filter=49 channel=90
    1, -2, -5, 2, -6, -4, -2, -4, 5,
    -- filter=49 channel=91
    0, 1, -2, 2, -7, 0, 6, 7, 4,
    -- filter=49 channel=92
    3, 0, -1, 2, -5, -5, -5, 2, -3,
    -- filter=49 channel=93
    1, -1, 2, -7, 6, -6, 0, 2, -6,
    -- filter=49 channel=94
    -3, -3, 0, 7, -2, 6, -3, -1, -2,
    -- filter=49 channel=95
    2, -4, -1, 1, 5, 5, -4, -5, -1,
    -- filter=49 channel=96
    6, -4, 2, 3, 7, -7, -1, 3, -5,
    -- filter=49 channel=97
    2, 2, -3, -3, -6, -7, -5, 5, 6,
    -- filter=49 channel=98
    -4, -1, -4, 3, -1, 0, -4, -3, -6,
    -- filter=49 channel=99
    2, -2, -6, -4, 1, -4, 2, -1, -2,
    -- filter=49 channel=100
    -7, -3, -2, 6, 4, 7, 4, 0, 4,
    -- filter=49 channel=101
    4, -6, 6, 0, -3, -5, -6, -3, -4,
    -- filter=49 channel=102
    6, -6, -2, 3, 5, 2, 5, -1, 2,
    -- filter=49 channel=103
    6, -6, 4, 0, 6, -3, 3, 1, 4,
    -- filter=49 channel=104
    -3, -4, -3, 2, 6, 0, -3, 1, -1,
    -- filter=49 channel=105
    -6, -2, -5, 1, 0, -5, -3, 2, -5,
    -- filter=49 channel=106
    -4, -4, -7, 4, 1, -3, 2, 0, 0,
    -- filter=49 channel=107
    -4, 0, 0, 2, -6, -3, -3, -6, 6,
    -- filter=49 channel=108
    5, 4, -2, 4, 5, 6, 0, -2, 7,
    -- filter=49 channel=109
    -2, -5, 4, 5, -6, 6, -6, -5, 5,
    -- filter=49 channel=110
    -5, -1, 2, 4, -6, -5, 1, 4, 0,
    -- filter=49 channel=111
    -2, -1, 4, -3, -3, 3, -1, -4, -2,
    -- filter=49 channel=112
    -5, -5, -1, 6, 2, 3, -5, -1, 2,
    -- filter=49 channel=113
    -6, -1, -6, -7, 6, 0, 7, -1, 6,
    -- filter=49 channel=114
    5, 4, 6, 0, 5, -4, 7, -7, 4,
    -- filter=49 channel=115
    -4, 1, -5, -6, -3, -4, -7, -5, 7,
    -- filter=49 channel=116
    0, -1, 4, 0, 0, -6, -3, -1, 2,
    -- filter=49 channel=117
    -3, -1, 0, -4, 2, -5, 0, 2, 0,
    -- filter=49 channel=118
    6, 5, 0, -6, -5, -1, -3, 0, 4,
    -- filter=49 channel=119
    -4, -1, 4, 0, -4, 0, 2, -3, 0,
    -- filter=49 channel=120
    -4, -7, 1, 5, -7, 1, -2, -6, 1,
    -- filter=49 channel=121
    -2, -1, 0, -6, 3, -4, -2, -5, -1,
    -- filter=49 channel=122
    -5, -7, -4, -6, -7, 4, 5, -4, -6,
    -- filter=49 channel=123
    -1, -1, 6, -6, 2, 2, 3, -7, 4,
    -- filter=49 channel=124
    5, 6, 1, 6, -5, -5, 4, -4, 0,
    -- filter=49 channel=125
    6, 5, -3, 0, 3, 4, -7, 0, -7,
    -- filter=49 channel=126
    -6, -4, -5, -2, -2, 3, 0, -1, 0,
    -- filter=49 channel=127
    -4, -2, -3, 2, -4, 3, 0, 2, -6,
    -- filter=50 channel=0
    0, -28, -21, 8, 3, -14, 5, 27, 12,
    -- filter=50 channel=1
    -12, -16, -23, 2, 1, -6, 13, 13, -5,
    -- filter=50 channel=2
    1, 1, 3, 2, 0, 4, 7, 4, 2,
    -- filter=50 channel=3
    5, 4, -4, 15, 16, 0, 4, 8, 11,
    -- filter=50 channel=4
    3, 4, 0, 7, 17, 15, 11, 5, 1,
    -- filter=50 channel=5
    -16, -20, -8, 16, 11, -4, 17, 38, 8,
    -- filter=50 channel=6
    0, 4, 0, -2, 4, 11, 0, -3, -6,
    -- filter=50 channel=7
    2, 6, 0, -4, -3, -5, -6, 2, 1,
    -- filter=50 channel=8
    4, -3, 8, 2, -4, -6, -7, -5, -8,
    -- filter=50 channel=9
    1, -9, -1, 0, 10, 8, 0, -1, 1,
    -- filter=50 channel=10
    11, 3, 1, 6, 3, 8, -13, -14, 6,
    -- filter=50 channel=11
    10, 10, -4, 0, 3, 17, -11, -12, -7,
    -- filter=50 channel=12
    -2, 4, -4, -5, -4, -5, -4, -5, -9,
    -- filter=50 channel=13
    7, -1, 5, 0, 5, 16, -14, -27, -15,
    -- filter=50 channel=14
    1, 1, 0, 6, -2, -3, 0, -5, -4,
    -- filter=50 channel=15
    6, 7, 2, -9, 17, 11, -15, -29, -11,
    -- filter=50 channel=16
    -3, -13, -14, 0, 5, -1, 4, 16, -2,
    -- filter=50 channel=17
    0, 1, 4, -4, 2, 0, 0, -2, -2,
    -- filter=50 channel=18
    7, 2, -4, 5, 6, 26, -15, -23, -4,
    -- filter=50 channel=19
    -6, 5, 5, 5, -4, 4, 2, 0, -4,
    -- filter=50 channel=20
    18, 24, 11, -8, 15, 18, -21, -33, -10,
    -- filter=50 channel=21
    -9, 0, -5, -6, 1, -9, 3, 3, 9,
    -- filter=50 channel=22
    -1, -6, 0, 6, 11, 4, 1, -7, 6,
    -- filter=50 channel=23
    8, -4, -15, 2, 28, 3, -27, -27, 6,
    -- filter=50 channel=24
    6, 3, -7, 6, 1, -3, 6, 4, -4,
    -- filter=50 channel=25
    -9, -3, -7, -6, 8, 18, 0, -18, -5,
    -- filter=50 channel=26
    -6, -3, -3, 8, 7, 2, 11, 11, 8,
    -- filter=50 channel=27
    7, -5, -6, -5, 25, 7, -10, -24, -3,
    -- filter=50 channel=28
    0, 4, 0, 6, -6, 6, -4, 3, 1,
    -- filter=50 channel=29
    12, 14, 10, -11, 13, 18, -16, -12, -5,
    -- filter=50 channel=30
    -5, -10, -8, 6, 10, 0, 10, 5, -7,
    -- filter=50 channel=31
    9, -3, -7, 10, 18, 3, -11, -12, 7,
    -- filter=50 channel=32
    3, 10, -7, -7, 15, 17, -2, -30, 0,
    -- filter=50 channel=33
    0, -8, -15, 1, 15, 6, -5, -13, 1,
    -- filter=50 channel=34
    5, 4, 0, 1, 4, 1, -9, -5, -2,
    -- filter=50 channel=35
    -1, 4, -3, -6, 6, 6, -1, 0, 1,
    -- filter=50 channel=36
    0, 8, 2, -1, 0, -2, -1, -5, -10,
    -- filter=50 channel=37
    -15, -27, -18, 5, 8, -4, 15, 14, 4,
    -- filter=50 channel=38
    0, -6, -8, 0, 13, -2, 0, -8, -5,
    -- filter=50 channel=39
    -1, 13, -4, 0, 8, 14, -6, -8, 1,
    -- filter=50 channel=40
    -3, 7, -8, -10, -6, -5, -20, -13, -9,
    -- filter=50 channel=41
    9, 11, 2, -2, -6, 15, -5, -13, -25,
    -- filter=50 channel=42
    0, -1, -2, -5, 5, -6, 2, 1, 11,
    -- filter=50 channel=43
    0, 5, -6, 3, 0, 5, -4, -1, 3,
    -- filter=50 channel=44
    -13, -11, -13, 0, 0, 0, 10, 15, 6,
    -- filter=50 channel=45
    1, -4, -7, 3, -3, -6, 1, 1, 5,
    -- filter=50 channel=46
    -3, -6, 5, -2, -5, 4, 0, 4, -10,
    -- filter=50 channel=47
    -16, -19, -17, 12, 6, -7, 11, 28, 11,
    -- filter=50 channel=48
    -11, -12, -7, 0, 1, 10, 13, -2, -13,
    -- filter=50 channel=49
    6, 10, 0, -2, 11, 17, 6, -6, -5,
    -- filter=50 channel=50
    3, -10, -6, 1, 2, 2, 5, -11, 0,
    -- filter=50 channel=51
    1, 4, -2, -3, 0, -5, -7, 0, 5,
    -- filter=50 channel=52
    8, 7, 8, -5, 3, -5, -15, -10, -3,
    -- filter=50 channel=53
    -1, 2, 1, -8, 14, 13, -12, -7, -2,
    -- filter=50 channel=54
    1, -3, 0, -4, -6, 6, -1, 0, 0,
    -- filter=50 channel=55
    16, 13, 5, -2, 5, 16, -14, -38, -8,
    -- filter=50 channel=56
    -5, 8, 8, -8, 5, 4, -12, -8, -9,
    -- filter=50 channel=57
    6, 6, 8, -1, 5, -3, 1, 6, -8,
    -- filter=50 channel=58
    -3, -10, -10, 1, 5, 1, 8, 11, 15,
    -- filter=50 channel=59
    0, -10, -4, -4, 9, 6, 3, -9, -4,
    -- filter=50 channel=60
    3, -1, 6, 7, 3, -1, 1, 2, 7,
    -- filter=50 channel=61
    0, 2, 2, 2, -3, -2, -3, -4, 0,
    -- filter=50 channel=62
    0, -5, -3, 2, -6, -5, -2, 0, -6,
    -- filter=50 channel=63
    0, -3, -2, 2, -1, -5, 6, 23, 12,
    -- filter=50 channel=64
    0, 1, -4, 1, -7, 0, -9, -4, -9,
    -- filter=50 channel=65
    -2, -2, -5, 0, 0, -6, -1, 0, 3,
    -- filter=50 channel=66
    2, 11, 5, -12, -9, 4, 7, -10, -7,
    -- filter=50 channel=67
    0, -4, -6, -7, -6, -1, 1, -1, 0,
    -- filter=50 channel=68
    5, 4, 1, 0, -2, 5, -3, -6, -8,
    -- filter=50 channel=69
    -2, 4, -2, -5, -5, -3, 7, 5, -6,
    -- filter=50 channel=70
    -3, 1, -11, -5, 6, 6, -12, -12, -5,
    -- filter=50 channel=71
    3, -3, 0, 7, 2, -8, 1, 1, 9,
    -- filter=50 channel=72
    6, 1, -4, -5, 5, 12, -7, -16, -7,
    -- filter=50 channel=73
    6, 4, 2, -4, 1, 19, -6, -15, -12,
    -- filter=50 channel=74
    8, -2, 5, 3, 10, -2, -6, -16, -2,
    -- filter=50 channel=75
    -6, -21, -21, 19, 6, -10, 0, 29, 16,
    -- filter=50 channel=76
    15, 16, 5, 0, -1, 9, -21, -32, -2,
    -- filter=50 channel=77
    -3, -1, 2, 3, 0, 3, 3, -4, -2,
    -- filter=50 channel=78
    6, 1, -6, 8, 10, -4, 6, 15, 6,
    -- filter=50 channel=79
    12, 1, -13, 0, 10, 18, -18, -31, -12,
    -- filter=50 channel=80
    2, -12, -12, -6, 6, 13, -1, -3, 0,
    -- filter=50 channel=81
    5, -4, 3, 6, -3, 0, 0, 1, 0,
    -- filter=50 channel=82
    2, -7, 4, 5, 8, -1, -6, 6, 4,
    -- filter=50 channel=83
    -7, -2, -7, -7, -2, 6, 2, 0, -3,
    -- filter=50 channel=84
    1, 7, 3, -14, 10, 6, -8, -18, -11,
    -- filter=50 channel=85
    4, -6, -3, -4, -6, -5, 6, 4, 4,
    -- filter=50 channel=86
    -6, 0, -7, -4, -2, -7, -3, -4, 7,
    -- filter=50 channel=87
    10, 15, 10, -1, 12, 8, -6, -12, -3,
    -- filter=50 channel=88
    -1, 5, 5, -8, -6, 0, -4, -2, -8,
    -- filter=50 channel=89
    6, 5, -2, 2, 12, 10, -11, -20, 0,
    -- filter=50 channel=90
    10, 5, -4, 0, 9, -9, -6, -10, 0,
    -- filter=50 channel=91
    3, 8, -5, -12, 21, 17, 0, -27, -10,
    -- filter=50 channel=92
    0, 5, 0, -1, 7, 1, -4, 2, 3,
    -- filter=50 channel=93
    -15, -17, -17, -3, 8, 0, 14, 6, 4,
    -- filter=50 channel=94
    6, 0, -1, -4, -1, -3, -6, 7, 5,
    -- filter=50 channel=95
    3, -3, 1, 6, -3, 4, -5, 6, 0,
    -- filter=50 channel=96
    2, -3, 0, -1, 4, 4, 6, -8, 0,
    -- filter=50 channel=97
    1, 3, -4, 12, 9, 0, 0, 3, 10,
    -- filter=50 channel=98
    4, -12, -4, 4, 18, 4, 1, -11, 5,
    -- filter=50 channel=99
    14, 3, -1, 7, 28, 12, -11, -24, 0,
    -- filter=50 channel=100
    5, 7, 0, 6, 2, 8, 2, 0, -6,
    -- filter=50 channel=101
    -1, 9, 10, 0, 11, 1, 14, 12, -5,
    -- filter=50 channel=102
    0, 4, -7, 6, 6, 0, 2, -3, 6,
    -- filter=50 channel=103
    -9, -15, -6, 7, 10, -9, 14, 23, 13,
    -- filter=50 channel=104
    3, -7, -2, 0, 5, 0, 3, 0, -7,
    -- filter=50 channel=105
    12, 9, 5, -4, 4, 6, -13, -12, 0,
    -- filter=50 channel=106
    3, 9, 9, -9, -4, 0, -7, -14, -1,
    -- filter=50 channel=107
    0, 11, 8, 2, 4, 3, -14, -8, -5,
    -- filter=50 channel=108
    4, 5, -7, 4, 4, -2, 4, 5, 0,
    -- filter=50 channel=109
    -2, 6, 1, -10, 14, 21, -5, -26, -9,
    -- filter=50 channel=110
    10, 7, 1, 9, 13, 8, -11, -3, 9,
    -- filter=50 channel=111
    5, -1, 7, 0, -8, -6, 3, 3, -6,
    -- filter=50 channel=112
    1, -12, 0, -4, 13, 6, -3, -10, 7,
    -- filter=50 channel=113
    2, -1, -1, 5, 11, 4, -11, -3, 9,
    -- filter=50 channel=114
    7, -11, -13, -3, 9, 22, 0, -15, -13,
    -- filter=50 channel=115
    -6, -4, 7, 0, -1, -6, 4, -1, -6,
    -- filter=50 channel=116
    0, 9, -1, -5, 7, 24, 5, -22, -4,
    -- filter=50 channel=117
    4, -7, 3, -5, 0, 2, -6, -1, -11,
    -- filter=50 channel=118
    6, -3, -3, -2, 0, -3, -6, -6, -4,
    -- filter=50 channel=119
    8, 5, -4, 0, 4, -10, -11, -11, -6,
    -- filter=50 channel=120
    15, 1, 6, -1, 14, 14, -12, -31, -16,
    -- filter=50 channel=121
    8, 9, -1, -2, -5, -2, 0, -8, 2,
    -- filter=50 channel=122
    -10, -17, -19, 9, 13, -1, 14, 26, 13,
    -- filter=50 channel=123
    -1, 6, 0, -1, 8, -8, -2, 1, -5,
    -- filter=50 channel=124
    3, 10, 2, 1, 0, 9, -2, -5, -1,
    -- filter=50 channel=125
    7, 0, -6, -2, 17, 19, -2, -14, -4,
    -- filter=50 channel=126
    -3, 6, -8, -3, 7, 11, -12, -1, -9,
    -- filter=50 channel=127
    7, 7, 4, -7, -6, -2, 5, -3, 0,
    -- filter=51 channel=0
    7, 3, 0, 10, -11, 4, 1, -3, 7,
    -- filter=51 channel=1
    11, 0, 0, 9, -11, 6, -2, -8, 0,
    -- filter=51 channel=2
    4, 0, 2, -3, 0, -2, 9, 0, -8,
    -- filter=51 channel=3
    0, -8, -8, 8, -16, -5, -1, -4, 1,
    -- filter=51 channel=4
    0, -16, -4, -12, 10, -12, 16, -8, -9,
    -- filter=51 channel=5
    3, -4, 0, 6, -3, 10, 1, -10, 8,
    -- filter=51 channel=6
    2, -5, 0, -9, -1, 1, -8, 6, -2,
    -- filter=51 channel=7
    5, -1, -4, 1, -3, -1, 2, 0, -3,
    -- filter=51 channel=8
    2, 10, 5, -8, 21, -10, 4, -4, -1,
    -- filter=51 channel=9
    -4, -1, 3, -9, -4, -1, 1, 0, -6,
    -- filter=51 channel=10
    2, 0, -5, 5, -6, 15, -15, 15, 0,
    -- filter=51 channel=11
    -8, -8, 5, -4, -1, 4, 1, 0, -1,
    -- filter=51 channel=12
    11, 0, 0, 11, 7, 11, -3, 4, -12,
    -- filter=51 channel=13
    2, -7, 1, 9, -13, 4, -6, 13, -7,
    -- filter=51 channel=14
    -3, -6, 1, 0, -2, 3, 1, -4, -7,
    -- filter=51 channel=15
    3, -8, 0, -9, 6, 0, -2, 6, -2,
    -- filter=51 channel=16
    5, 3, -3, 7, -3, 10, -2, -2, -1,
    -- filter=51 channel=17
    -1, 0, 2, -4, -4, 0, 0, 4, 6,
    -- filter=51 channel=18
    12, -5, 8, -4, -14, 9, -16, 8, 1,
    -- filter=51 channel=19
    0, -7, -4, 2, -4, -4, 0, -2, -3,
    -- filter=51 channel=20
    1, -3, 10, -15, 9, -7, -13, 4, -3,
    -- filter=51 channel=21
    -1, -6, 3, 0, -4, 9, -4, 0, -9,
    -- filter=51 channel=22
    -5, 7, 3, -5, 5, -2, -1, 5, -5,
    -- filter=51 channel=23
    -10, -1, 3, -21, 18, -5, -4, 22, -22,
    -- filter=51 channel=24
    2, -1, 2, 4, 4, -4, -3, 5, 1,
    -- filter=51 channel=25
    10, -10, 12, 3, -14, 19, -7, 6, -16,
    -- filter=51 channel=26
    3, -9, 3, 4, 0, -5, 2, -9, -10,
    -- filter=51 channel=27
    6, -21, 13, -16, 13, 1, -2, 7, -19,
    -- filter=51 channel=28
    6, 3, 4, 2, 0, 3, 0, 0, -5,
    -- filter=51 channel=29
    3, 0, 3, 0, 10, 12, -7, 11, 5,
    -- filter=51 channel=30
    3, -14, 0, -8, 0, 5, -4, 1, -8,
    -- filter=51 channel=31
    0, -7, 3, -12, 1, 3, -3, 10, -15,
    -- filter=51 channel=32
    16, -7, 11, -8, -6, 11, -6, 13, -10,
    -- filter=51 channel=33
    6, -18, -2, 0, -8, 6, -9, 3, -8,
    -- filter=51 channel=34
    3, 2, -7, -7, 29, -21, 15, -2, -12,
    -- filter=51 channel=35
    -3, 1, -5, 1, 0, 0, -3, -4, -3,
    -- filter=51 channel=36
    -7, -6, -3, -9, 7, -2, 0, 13, -6,
    -- filter=51 channel=37
    15, -5, 2, 2, -7, -3, 0, -4, -4,
    -- filter=51 channel=38
    -2, -14, -1, -2, 0, 0, -12, 10, -2,
    -- filter=51 channel=39
    1, 1, 2, -3, 7, 2, 1, 3, -7,
    -- filter=51 channel=40
    -8, 2, 5, -6, -4, 7, -7, 4, 4,
    -- filter=51 channel=41
    5, 23, -6, 22, -6, 4, -3, 0, 0,
    -- filter=51 channel=42
    -6, -5, 4, -3, -9, 4, -2, -8, -4,
    -- filter=51 channel=43
    2, 2, -12, 4, -10, -1, -5, -2, -4,
    -- filter=51 channel=44
    10, -3, 13, 0, -1, -1, 7, 10, -5,
    -- filter=51 channel=45
    3, 0, 5, -8, -9, -1, 4, -7, 2,
    -- filter=51 channel=46
    3, 5, -3, 6, -3, -1, -5, 0, 7,
    -- filter=51 channel=47
    7, -9, 8, 5, -5, 13, -2, 2, -4,
    -- filter=51 channel=48
    2, -18, 10, -9, -1, 0, -1, 16, -14,
    -- filter=51 channel=49
    -10, -4, 0, -10, 1, 2, 0, 0, -3,
    -- filter=51 channel=50
    0, -7, 0, -9, 2, -10, -7, 12, -15,
    -- filter=51 channel=51
    2, -3, -7, 0, 5, 6, 0, 3, 0,
    -- filter=51 channel=52
    -4, 0, -2, -5, 23, -5, 4, 11, -15,
    -- filter=51 channel=53
    -1, 0, 1, -4, 7, -1, 0, -2, 1,
    -- filter=51 channel=54
    6, -4, -2, 0, 0, 5, 2, -6, 3,
    -- filter=51 channel=55
    9, -9, 1, -1, 2, 10, -9, 20, -2,
    -- filter=51 channel=56
    2, 11, -1, 1, 12, -10, 9, -3, 0,
    -- filter=51 channel=57
    6, -2, 0, -10, -5, -4, -5, 3, 1,
    -- filter=51 channel=58
    -1, 3, -1, 1, -7, -6, 3, 0, -1,
    -- filter=51 channel=59
    0, -16, 0, 0, -5, 20, -13, 10, 0,
    -- filter=51 channel=60
    3, -4, 3, 6, -6, -2, -7, 0, -1,
    -- filter=51 channel=61
    3, 9, -1, 3, 12, -6, 5, 7, -8,
    -- filter=51 channel=62
    6, 0, -6, -3, 3, 0, 2, -3, 4,
    -- filter=51 channel=63
    -2, 1, 3, 8, 1, 5, 4, -5, 3,
    -- filter=51 channel=64
    -3, 10, 6, 0, 6, 0, -1, -7, -1,
    -- filter=51 channel=65
    1, 1, -4, -2, 0, -5, 3, 0, 1,
    -- filter=51 channel=66
    14, 3, -7, 19, -5, 7, 4, 13, -3,
    -- filter=51 channel=67
    -2, 4, -7, 2, 6, -7, 6, 2, -6,
    -- filter=51 channel=68
    4, -12, 6, -2, -6, 4, 5, 6, -9,
    -- filter=51 channel=69
    -1, 3, -6, 0, -9, 7, -5, -3, 0,
    -- filter=51 channel=70
    1, -13, -6, -5, 3, -6, -4, 4, -15,
    -- filter=51 channel=71
    -7, 0, -7, -3, -3, -6, 0, -7, 0,
    -- filter=51 channel=72
    5, -7, 9, -5, -6, 16, -8, 14, -12,
    -- filter=51 channel=73
    7, -14, 4, -13, 13, 5, 4, 10, -6,
    -- filter=51 channel=74
    2, 2, 7, -4, 18, -26, 16, 0, -22,
    -- filter=51 channel=75
    4, 1, -4, 16, -27, 12, 1, -6, 10,
    -- filter=51 channel=76
    -7, 0, 6, -3, 4, 5, -18, 11, 7,
    -- filter=51 channel=77
    5, 0, -5, 5, -1, 3, -7, -1, 1,
    -- filter=51 channel=78
    -5, 0, 2, -5, -4, -4, 3, 0, -3,
    -- filter=51 channel=79
    7, -19, 10, -5, -18, 14, -7, 17, -3,
    -- filter=51 channel=80
    8, -9, 9, -2, -10, 21, -15, 21, -12,
    -- filter=51 channel=81
    -5, 6, 3, 2, -4, 2, -1, -4, 6,
    -- filter=51 channel=82
    5, 5, -6, -2, -2, -6, 1, 3, 6,
    -- filter=51 channel=83
    -3, 3, -4, -12, 10, -10, 4, 0, -9,
    -- filter=51 channel=84
    -3, -9, 2, -4, 10, -5, 0, 2, -4,
    -- filter=51 channel=85
    5, 1, 2, -6, -1, 4, 5, 6, -2,
    -- filter=51 channel=86
    2, -7, 5, -4, 2, -11, -3, 10, -6,
    -- filter=51 channel=87
    -4, 8, -5, -4, 18, -13, 3, 8, 0,
    -- filter=51 channel=88
    0, 5, 5, -11, 16, -9, -2, 8, -12,
    -- filter=51 channel=89
    10, -14, 4, 3, -16, 19, -13, 18, 2,
    -- filter=51 channel=90
    0, 3, -4, -4, 8, -7, 4, -1, -11,
    -- filter=51 channel=91
    1, -13, 15, -12, 13, 0, -3, 13, -5,
    -- filter=51 channel=92
    2, 0, -12, 0, 8, -4, -2, -2, 0,
    -- filter=51 channel=93
    10, 1, 0, 3, 4, -1, 3, -1, -3,
    -- filter=51 channel=94
    5, 0, 0, 1, 6, 4, 0, 0, -5,
    -- filter=51 channel=95
    -3, 1, -3, 0, 4, 0, -4, -1, 1,
    -- filter=51 channel=96
    -7, -7, -8, 3, -5, 3, -1, -2, 0,
    -- filter=51 channel=97
    -3, -7, -13, 0, -4, -4, -1, 4, 0,
    -- filter=51 channel=98
    15, -22, 13, -10, -8, 8, -13, 21, -3,
    -- filter=51 channel=99
    0, -8, 14, -15, 25, -7, 2, 29, -29,
    -- filter=51 channel=100
    2, 14, 2, -1, 5, 2, -4, -2, 3,
    -- filter=51 channel=101
    -5, -13, -9, -9, 8, -14, 13, 6, 1,
    -- filter=51 channel=102
    -6, -4, 7, -3, 1, -4, 4, 2, 0,
    -- filter=51 channel=103
    10, -2, 1, -1, -9, 9, -8, 1, 2,
    -- filter=51 channel=104
    9, -14, 11, -12, 3, 9, -8, 17, -9,
    -- filter=51 channel=105
    0, -1, 6, -6, 0, 3, -5, 9, -2,
    -- filter=51 channel=106
    -5, 7, 0, 0, 2, 0, 0, 4, 1,
    -- filter=51 channel=107
    -3, -1, 0, -3, 10, -10, -2, 12, -14,
    -- filter=51 channel=108
    5, 3, -3, 5, -9, 3, 3, 1, 9,
    -- filter=51 channel=109
    10, -17, 11, -16, 12, 6, 2, 11, -15,
    -- filter=51 channel=110
    -1, -1, 3, 2, 7, 0, -8, 3, -2,
    -- filter=51 channel=111
    -6, -1, -6, 3, -7, 3, -7, 6, 4,
    -- filter=51 channel=112
    1, -5, 9, -3, 5, -8, 3, -1, -13,
    -- filter=51 channel=113
    10, -6, -2, -3, -6, 0, -5, 6, 0,
    -- filter=51 channel=114
    15, -23, 15, -8, -6, 0, -1, 17, -15,
    -- filter=51 channel=115
    -4, 6, -2, -1, -1, -1, 5, -1, -3,
    -- filter=51 channel=116
    4, -17, 8, -17, 3, 14, -4, 11, -8,
    -- filter=51 channel=117
    5, 0, 2, 3, 1, -2, 0, 2, -1,
    -- filter=51 channel=118
    -1, 6, 3, 1, 3, -4, 5, -4, -5,
    -- filter=51 channel=119
    -4, 21, -4, -7, 31, -15, 8, -1, -7,
    -- filter=51 channel=120
    -4, -12, 10, -19, 34, -20, -1, 24, -28,
    -- filter=51 channel=121
    11, 7, 1, 4, -3, 12, -7, 0, 1,
    -- filter=51 channel=122
    13, -4, 3, 0, 3, 8, -1, 0, -9,
    -- filter=51 channel=123
    -8, 5, -10, 0, 7, -14, -1, -7, -11,
    -- filter=51 channel=124
    0, 0, 0, -6, 9, -1, -5, 7, 2,
    -- filter=51 channel=125
    0, -20, 12, -15, 7, 6, -2, 10, -10,
    -- filter=51 channel=126
    3, -1, 3, 16, -18, 7, -9, 6, 11,
    -- filter=51 channel=127
    8, 4, 1, 0, -4, 1, -1, -4, 3,
    -- filter=52 channel=0
    3, 5, 5, 1, 13, 11, 0, 12, 6,
    -- filter=52 channel=1
    -4, -3, 2, 3, 4, 12, 6, 1, 5,
    -- filter=52 channel=2
    -2, -3, 0, 6, 5, -3, 0, 0, -4,
    -- filter=52 channel=3
    1, 10, 7, 0, 7, -3, 0, 1, 4,
    -- filter=52 channel=4
    -2, 7, 5, 0, 1, 0, 5, 4, -2,
    -- filter=52 channel=5
    -7, 3, -2, 8, 9, 12, 0, 4, 11,
    -- filter=52 channel=6
    4, 0, 2, -5, -1, 7, -5, -6, 3,
    -- filter=52 channel=7
    -7, 0, 4, 0, -6, -7, 2, -7, -2,
    -- filter=52 channel=8
    3, 7, 5, 0, 0, -3, -4, 7, -4,
    -- filter=52 channel=9
    -6, -2, 0, -6, -6, -3, 5, 6, 6,
    -- filter=52 channel=10
    1, 0, 0, -2, -1, -1, 1, -4, -7,
    -- filter=52 channel=11
    -7, -7, 7, 0, 3, 5, -3, -8, 4,
    -- filter=52 channel=12
    -6, -1, 3, 4, -4, 5, 4, 2, 5,
    -- filter=52 channel=13
    1, -6, 3, -5, -3, -9, -3, -5, -3,
    -- filter=52 channel=14
    -3, 6, 2, -5, -1, 3, 0, 7, -5,
    -- filter=52 channel=15
    -2, -4, 1, 2, -7, -1, -9, 0, 2,
    -- filter=52 channel=16
    1, -3, -2, 0, -3, 1, 4, -1, 0,
    -- filter=52 channel=17
    -7, 2, 3, -4, -5, 4, 0, -4, 6,
    -- filter=52 channel=18
    0, 0, 5, -3, -3, -5, -3, 0, 3,
    -- filter=52 channel=19
    1, -1, 1, 7, -4, -2, 6, 4, 4,
    -- filter=52 channel=20
    -5, 0, 7, 0, 2, 5, -6, -7, -9,
    -- filter=52 channel=21
    4, -2, 6, -3, -1, -7, 6, -4, 3,
    -- filter=52 channel=22
    -5, 0, 1, -6, 1, 9, 7, 0, 0,
    -- filter=52 channel=23
    1, -1, 0, 2, 0, -8, -5, 1, -3,
    -- filter=52 channel=24
    -1, -3, -3, -2, -1, -2, 2, -6, 2,
    -- filter=52 channel=25
    -4, 2, 0, -1, 0, -7, 0, 0, -2,
    -- filter=52 channel=26
    4, 0, 5, 4, -1, 4, 7, 7, -2,
    -- filter=52 channel=27
    0, 0, 8, -10, -7, -2, -7, -1, -2,
    -- filter=52 channel=28
    -1, 5, -7, 4, 5, 7, -4, -3, 4,
    -- filter=52 channel=29
    -6, -5, 5, 2, -8, 6, -1, -1, -5,
    -- filter=52 channel=30
    -3, 0, -6, 0, -3, -4, -3, -2, 0,
    -- filter=52 channel=31
    -3, 3, 6, -2, -7, 0, 0, -10, -3,
    -- filter=52 channel=32
    -5, -7, 5, -8, -2, -5, 4, 1, 4,
    -- filter=52 channel=33
    -1, -3, 5, 5, -6, 7, 0, -6, -5,
    -- filter=52 channel=34
    6, 5, -6, 6, 1, 2, 6, 8, -3,
    -- filter=52 channel=35
    -1, -3, 2, -4, -3, 0, -3, -1, 2,
    -- filter=52 channel=36
    -2, -1, -6, 6, -7, -5, -7, -6, -3,
    -- filter=52 channel=37
    -6, -7, 7, 0, 11, 9, -5, 3, 8,
    -- filter=52 channel=38
    0, -3, -3, 0, -1, -4, 2, -2, -1,
    -- filter=52 channel=39
    3, -1, 0, 4, -1, 2, 0, 4, -5,
    -- filter=52 channel=40
    0, -3, 0, 5, 0, 0, 1, -2, -7,
    -- filter=52 channel=41
    -3, 1, -4, -2, -2, 0, 2, -1, 1,
    -- filter=52 channel=42
    -7, -7, -3, -8, -1, 8, 1, -5, -2,
    -- filter=52 channel=43
    -1, 5, 2, -5, -4, 8, 0, 5, 0,
    -- filter=52 channel=44
    -2, 6, 8, 5, 7, 6, 2, 5, 5,
    -- filter=52 channel=45
    0, -3, 7, -3, 0, -1, -2, -5, 0,
    -- filter=52 channel=46
    -2, -5, 2, -1, 0, 7, 0, 1, 0,
    -- filter=52 channel=47
    6, -1, 3, -1, 0, -2, -1, -6, 3,
    -- filter=52 channel=48
    -7, -3, -5, -6, -5, -2, 2, -10, -4,
    -- filter=52 channel=49
    -1, -7, 4, 3, -7, 2, -1, -7, -7,
    -- filter=52 channel=50
    0, 3, 5, -4, -9, 4, 0, -1, -7,
    -- filter=52 channel=51
    2, -2, -7, -5, 0, -2, 0, -3, -6,
    -- filter=52 channel=52
    0, -5, -1, 6, 5, -3, 7, -4, 4,
    -- filter=52 channel=53
    2, 0, -2, -8, 1, 0, 5, -7, 1,
    -- filter=52 channel=54
    5, 0, 2, 2, -1, 3, 5, 0, -6,
    -- filter=52 channel=55
    2, 4, 5, -9, 0, -2, -1, -5, -2,
    -- filter=52 channel=56
    2, -2, -6, 0, 1, 0, 1, -1, 2,
    -- filter=52 channel=57
    -6, 0, 0, 4, 5, -1, 4, 7, 0,
    -- filter=52 channel=58
    -1, 6, -3, -2, 3, 8, 0, 9, 10,
    -- filter=52 channel=59
    -7, -5, 2, -8, 2, -6, -4, -5, 3,
    -- filter=52 channel=60
    3, -5, -3, -6, -3, -2, -4, 7, 5,
    -- filter=52 channel=61
    3, 3, -7, -6, 4, -7, 3, 4, 0,
    -- filter=52 channel=62
    5, 0, -4, 0, 6, 3, -1, 0, -2,
    -- filter=52 channel=63
    -1, 4, 2, 0, 0, 0, -5, 5, 7,
    -- filter=52 channel=64
    2, 3, 3, -4, -4, -8, 6, 3, -6,
    -- filter=52 channel=65
    -6, 0, -2, 6, 0, 5, 2, 7, -1,
    -- filter=52 channel=66
    -5, 0, -6, 5, -7, -5, 0, -1, 1,
    -- filter=52 channel=67
    -3, -2, 0, 5, -2, 3, 3, 1, -1,
    -- filter=52 channel=68
    -7, -6, 3, -6, 4, -7, 2, -1, -4,
    -- filter=52 channel=69
    -5, -6, -2, 1, -5, 5, -3, 6, 6,
    -- filter=52 channel=70
    -7, 0, 1, -5, 1, -3, -8, 4, -6,
    -- filter=52 channel=71
    1, 2, 1, 7, -3, -6, -2, 4, 2,
    -- filter=52 channel=72
    2, -7, -3, -4, -9, -7, -6, -11, 2,
    -- filter=52 channel=73
    2, 3, -2, -6, 4, -6, 0, -7, 5,
    -- filter=52 channel=74
    0, 5, 0, 4, -2, 4, 4, 3, -3,
    -- filter=52 channel=75
    4, 4, 10, -5, 7, 15, 0, 13, 15,
    -- filter=52 channel=76
    -5, -1, -1, 2, -3, -6, -3, -10, 1,
    -- filter=52 channel=77
    5, -6, 5, -5, 0, 4, 7, -6, -4,
    -- filter=52 channel=78
    0, 7, -4, -6, 0, 0, -6, 4, 8,
    -- filter=52 channel=79
    -3, -3, -5, -3, -8, -5, -7, -4, -5,
    -- filter=52 channel=80
    2, 2, 0, 0, -7, -12, -8, -3, -4,
    -- filter=52 channel=81
    3, -6, -4, -3, -4, 1, 5, 4, -5,
    -- filter=52 channel=82
    -1, 7, 1, -1, 0, 2, -6, -5, 6,
    -- filter=52 channel=83
    2, 0, 5, 6, -2, 2, 0, -4, -1,
    -- filter=52 channel=84
    -8, -3, -3, 1, -3, 4, 5, -4, -7,
    -- filter=52 channel=85
    4, -5, -5, 5, 5, 6, -6, -2, -7,
    -- filter=52 channel=86
    -7, 0, -2, 3, 2, -3, -1, 8, 0,
    -- filter=52 channel=87
    -7, -1, 7, 3, 3, -6, 7, 0, -2,
    -- filter=52 channel=88
    -1, 4, 0, -6, 5, 3, -6, -8, -9,
    -- filter=52 channel=89
    4, -6, -2, -4, -9, -2, 0, 1, -10,
    -- filter=52 channel=90
    6, -3, 2, -4, 3, -3, 6, -3, 4,
    -- filter=52 channel=91
    -4, -8, -1, 3, 1, 0, -10, -4, 0,
    -- filter=52 channel=92
    1, -5, 1, -1, -1, -6, -5, 7, 6,
    -- filter=52 channel=93
    4, -6, 0, 0, 8, 0, 0, 9, 1,
    -- filter=52 channel=94
    -2, 1, -6, 6, 2, -4, -5, 6, 5,
    -- filter=52 channel=95
    -7, 6, -4, 2, -7, -2, 0, -6, -3,
    -- filter=52 channel=96
    -1, -5, 1, -4, -7, 0, -4, -3, -6,
    -- filter=52 channel=97
    5, -3, 5, -7, 1, 7, 6, 3, -6,
    -- filter=52 channel=98
    -6, 2, 5, -7, 1, 2, -3, -7, 3,
    -- filter=52 channel=99
    -5, 4, -4, 0, -7, -7, -1, 0, -7,
    -- filter=52 channel=100
    -4, -2, 4, 2, 7, 6, 6, -4, -4,
    -- filter=52 channel=101
    3, 0, 1, -6, -4, 5, -6, 0, 0,
    -- filter=52 channel=102
    6, 0, 0, 2, 0, 2, 0, 2, 4,
    -- filter=52 channel=103
    -3, -5, 3, -1, 3, 2, 0, -3, -3,
    -- filter=52 channel=104
    5, -1, -1, -4, -5, 1, -4, -1, -8,
    -- filter=52 channel=105
    -3, -1, -4, -6, 0, -6, -2, -5, 0,
    -- filter=52 channel=106
    -4, 3, 5, 1, -5, -7, -2, -9, -1,
    -- filter=52 channel=107
    0, 0, 2, -4, 0, -5, 2, 5, 5,
    -- filter=52 channel=108
    0, -1, 4, 1, 6, 6, 0, -3, 5,
    -- filter=52 channel=109
    -1, -4, 0, 0, 1, -8, -5, 3, -5,
    -- filter=52 channel=110
    -6, -5, -5, -5, -4, 6, -2, -3, 1,
    -- filter=52 channel=111
    -5, -3, -3, -4, -2, 6, -4, -5, -2,
    -- filter=52 channel=112
    -5, 6, -6, 3, 3, 1, 4, 4, 1,
    -- filter=52 channel=113
    3, 0, 5, 1, 4, -3, 5, -1, 0,
    -- filter=52 channel=114
    -4, -8, 6, -5, 4, 7, 0, 6, 8,
    -- filter=52 channel=115
    -6, 0, -2, 1, 1, 5, 0, 1, -4,
    -- filter=52 channel=116
    -1, 1, -3, -7, -5, -6, 0, -1, -3,
    -- filter=52 channel=117
    5, -3, 5, 5, -7, -5, 6, -4, 0,
    -- filter=52 channel=118
    5, 5, 1, 5, 1, -3, 2, 3, 2,
    -- filter=52 channel=119
    0, -3, 4, 1, 1, 5, -5, 4, -5,
    -- filter=52 channel=120
    -2, 1, -3, 1, -7, -5, -9, 2, 3,
    -- filter=52 channel=121
    -1, -2, -2, -2, 0, -6, -7, -8, -7,
    -- filter=52 channel=122
    0, 2, -4, 5, -6, 0, 5, -8, -3,
    -- filter=52 channel=123
    3, -4, 1, -3, 2, -1, -2, -4, -1,
    -- filter=52 channel=124
    0, -3, 1, 1, -3, -3, -6, 0, 5,
    -- filter=52 channel=125
    6, 5, 7, 0, -2, 2, -5, -10, -4,
    -- filter=52 channel=126
    5, 5, 2, -2, 4, -4, -3, -7, 0,
    -- filter=52 channel=127
    4, 5, 3, 0, -2, -4, 4, -5, -5,
    -- filter=53 channel=0
    9, 0, -5, 0, 4, -4, 0, 0, -14,
    -- filter=53 channel=1
    -2, -4, -9, 9, 10, 4, 6, 8, -8,
    -- filter=53 channel=2
    -2, -7, -2, 2, 6, 1, -1, 2, 5,
    -- filter=53 channel=3
    3, 1, -2, -2, 3, 0, 3, 9, -4,
    -- filter=53 channel=4
    -11, 4, -5, -10, 6, 5, 1, -3, 0,
    -- filter=53 channel=5
    11, 3, -8, 13, 9, -3, 6, 5, -8,
    -- filter=53 channel=6
    -6, -2, -7, -11, -4, 3, -8, -10, 0,
    -- filter=53 channel=7
    0, -2, 6, 3, 1, 1, 3, 3, 3,
    -- filter=53 channel=8
    6, -3, -2, 8, 3, -2, 5, 3, 6,
    -- filter=53 channel=9
    -4, -3, 0, -1, 1, 3, -2, 8, 0,
    -- filter=53 channel=10
    -1, -3, 0, -4, 1, 5, -5, 8, -3,
    -- filter=53 channel=11
    2, -5, 0, -16, -11, -1, -11, 1, 1,
    -- filter=53 channel=12
    1, -2, 3, 0, -7, 5, -2, -5, 7,
    -- filter=53 channel=13
    -11, -7, 1, -21, -5, 2, -8, 4, 11,
    -- filter=53 channel=14
    2, -4, 3, -3, -6, -1, -6, 3, 5,
    -- filter=53 channel=15
    5, 7, -2, -10, -10, -5, -1, -2, 2,
    -- filter=53 channel=16
    -3, -11, -7, -1, -1, 3, 7, 7, 1,
    -- filter=53 channel=17
    1, -6, -1, -1, 2, 2, -6, 0, 0,
    -- filter=53 channel=18
    -7, 7, 3, -17, -2, 2, -14, -2, 0,
    -- filter=53 channel=19
    -1, -3, 3, 7, 3, -3, -6, 3, -4,
    -- filter=53 channel=20
    -5, -11, -2, -17, -17, -1, -19, -10, -1,
    -- filter=53 channel=21
    -5, -1, -6, -2, 11, 0, -2, -1, -12,
    -- filter=53 channel=22
    -3, -2, -7, -5, -9, -1, 2, -1, 0,
    -- filter=53 channel=23
    -3, 7, -2, -8, -10, -9, -9, 0, -5,
    -- filter=53 channel=24
    2, -5, -7, -5, -3, -6, 5, 1, 0,
    -- filter=53 channel=25
    0, 9, 6, -1, 11, 7, 6, 4, 1,
    -- filter=53 channel=26
    -1, -8, -5, 12, 7, -9, 4, -4, -9,
    -- filter=53 channel=27
    3, 11, 8, -8, 9, -4, -2, 12, -4,
    -- filter=53 channel=28
    -7, 1, 4, 6, -4, -4, -4, 6, 0,
    -- filter=53 channel=29
    -9, 4, 5, -7, -6, -2, -13, -12, 1,
    -- filter=53 channel=30
    3, -7, -6, 0, 5, 2, 4, 3, 0,
    -- filter=53 channel=31
    4, -5, 7, -7, 4, -2, 1, 6, -15,
    -- filter=53 channel=32
    4, 10, 5, -18, -2, 2, -3, 3, -4,
    -- filter=53 channel=33
    4, 10, 0, -5, 9, 8, 4, 12, 3,
    -- filter=53 channel=34
    0, 3, -3, 2, -5, -2, -1, 0, -7,
    -- filter=53 channel=35
    -3, 4, -5, -4, 0, -4, -6, 6, 5,
    -- filter=53 channel=36
    -2, -13, -1, -7, -11, -1, 2, -9, -10,
    -- filter=53 channel=37
    1, -7, -11, 13, 13, -9, 3, 10, -15,
    -- filter=53 channel=38
    3, 3, -2, 2, 9, 3, -3, 5, -6,
    -- filter=53 channel=39
    -1, 0, -3, -4, -7, -8, 0, -10, -3,
    -- filter=53 channel=40
    -1, -3, 2, -11, -13, -2, -11, -10, 3,
    -- filter=53 channel=41
    -9, -10, -5, -16, -10, 1, -16, -7, 7,
    -- filter=53 channel=42
    0, -1, -1, -4, 9, -2, -1, 7, -8,
    -- filter=53 channel=43
    0, 0, 0, -12, -6, 3, -5, -1, -6,
    -- filter=53 channel=44
    7, 4, 0, 4, 14, 3, 14, 11, -10,
    -- filter=53 channel=45
    5, 0, -1, 1, -2, -7, 0, 0, -8,
    -- filter=53 channel=46
    0, -8, 2, -7, -1, 0, -1, 4, 1,
    -- filter=53 channel=47
    5, 0, -1, 1, 19, 0, 14, 5, -5,
    -- filter=53 channel=48
    -8, 1, -6, -1, 5, 7, 12, 6, 3,
    -- filter=53 channel=49
    -9, 7, 0, -11, 4, -3, -5, 4, 6,
    -- filter=53 channel=50
    5, 2, 2, -8, 6, -5, 7, 5, -10,
    -- filter=53 channel=51
    -3, 0, 3, 4, -5, 0, 1, 6, -7,
    -- filter=53 channel=52
    0, 5, 5, -3, 0, -3, -2, -7, -7,
    -- filter=53 channel=53
    -8, -4, 7, -5, -10, -7, -8, -1, -7,
    -- filter=53 channel=54
    -5, -6, -4, 3, 3, 2, 2, 3, 3,
    -- filter=53 channel=55
    -10, 3, 11, -12, -7, -5, -17, -7, 6,
    -- filter=53 channel=56
    -5, 2, -8, -4, -7, -2, -5, 2, 3,
    -- filter=53 channel=57
    -2, 5, -6, -6, -3, 1, 4, -4, 0,
    -- filter=53 channel=58
    6, 3, -9, 11, -3, 0, 4, -1, -12,
    -- filter=53 channel=59
    -3, 2, 0, -5, 12, -1, -5, 2, -6,
    -- filter=53 channel=60
    -4, 1, 5, 0, 7, -4, 2, 1, -4,
    -- filter=53 channel=61
    -6, -4, 2, -7, 0, -4, 3, -6, 5,
    -- filter=53 channel=62
    -1, 1, 3, 4, -8, -5, -2, -6, -6,
    -- filter=53 channel=63
    0, -1, -3, 2, -3, -5, 9, 1, -5,
    -- filter=53 channel=64
    -3, -1, -2, -3, -11, 3, -1, -8, 6,
    -- filter=53 channel=65
    4, -4, 0, -2, -1, -5, -2, 0, -3,
    -- filter=53 channel=66
    -2, -8, -5, -13, 1, -6, -11, -6, -4,
    -- filter=53 channel=67
    0, -5, 5, 6, -6, 0, -1, -4, -7,
    -- filter=53 channel=68
    2, 3, 0, -4, 1, -1, 3, 5, -6,
    -- filter=53 channel=69
    -9, -7, -2, -8, -3, -6, 0, 3, -5,
    -- filter=53 channel=70
    -4, 12, 8, -5, -5, 5, 0, 0, 0,
    -- filter=53 channel=71
    -4, 6, 0, -8, -6, 2, -3, -1, -6,
    -- filter=53 channel=72
    -12, -3, 0, -3, 2, 5, 1, 6, -2,
    -- filter=53 channel=73
    0, -3, 0, -2, -1, 9, 5, -4, 8,
    -- filter=53 channel=74
    0, 5, -7, 4, 5, -12, 0, -3, 1,
    -- filter=53 channel=75
    0, 2, -8, 1, 8, -7, 5, -1, -10,
    -- filter=53 channel=76
    -11, -2, 0, -8, -9, -1, -12, -6, 3,
    -- filter=53 channel=77
    -5, -7, 0, -3, -7, 7, 0, 0, 3,
    -- filter=53 channel=78
    7, -3, -8, 11, 8, -2, 2, 8, 3,
    -- filter=53 channel=79
    -5, 5, 0, -21, -8, -1, -6, 6, 12,
    -- filter=53 channel=80
    0, 5, -4, -3, 12, 11, 10, 4, -4,
    -- filter=53 channel=81
    7, 0, 6, 3, 3, 6, -2, 6, 0,
    -- filter=53 channel=82
    -1, -5, 3, 0, 6, 4, 3, -7, -8,
    -- filter=53 channel=83
    2, 5, 4, 2, -4, 2, 5, 6, -2,
    -- filter=53 channel=84
    -6, -5, 4, -2, 3, 4, -6, 0, 4,
    -- filter=53 channel=85
    -1, -3, -7, 5, -3, 1, -3, -3, -6,
    -- filter=53 channel=86
    7, 0, 4, 4, 0, 2, -2, -1, -1,
    -- filter=53 channel=87
    4, -2, -1, -3, -4, -11, -7, -7, 0,
    -- filter=53 channel=88
    -5, -13, -1, 1, -2, -5, -3, -14, 2,
    -- filter=53 channel=89
    -4, -6, 12, -22, 4, 3, -13, -2, 0,
    -- filter=53 channel=90
    -7, -1, -6, 2, -6, -10, -5, -5, -2,
    -- filter=53 channel=91
    4, 2, 4, -9, 1, -6, 1, 2, 5,
    -- filter=53 channel=92
    -4, -7, 3, -6, -1, 0, 0, -9, 3,
    -- filter=53 channel=93
    -2, -2, -12, 12, 11, 3, 16, 3, 0,
    -- filter=53 channel=94
    5, -6, 2, -1, 0, -5, 7, -6, 4,
    -- filter=53 channel=95
    0, -4, -4, -2, -5, 2, 7, 1, 6,
    -- filter=53 channel=96
    3, 4, 4, -6, 2, -4, -7, 7, 4,
    -- filter=53 channel=97
    -3, -4, -8, 6, 5, 0, -4, 6, -8,
    -- filter=53 channel=98
    3, 0, 4, -8, 10, 8, 9, 10, 9,
    -- filter=53 channel=99
    -1, -2, 6, -10, 1, -7, -7, -8, 1,
    -- filter=53 channel=100
    6, -6, 5, -4, -4, -1, 3, 3, -2,
    -- filter=53 channel=101
    -9, 4, 3, -8, 6, -5, 5, 5, 7,
    -- filter=53 channel=102
    0, 4, 1, 0, -2, -5, 7, -5, 4,
    -- filter=53 channel=103
    4, -3, -2, 11, 17, -5, 5, 4, -5,
    -- filter=53 channel=104
    -10, 3, 5, -6, 0, -6, 3, 6, -4,
    -- filter=53 channel=105
    3, -6, 0, -7, -5, -9, -6, 0, 7,
    -- filter=53 channel=106
    -8, 0, 1, -9, -5, -6, -4, 0, -1,
    -- filter=53 channel=107
    -7, -5, 2, 0, -13, -6, -7, -14, -4,
    -- filter=53 channel=108
    -6, -1, 1, 1, -5, -4, 2, 4, 3,
    -- filter=53 channel=109
    -6, 2, 3, -1, 8, 10, 12, 9, -1,
    -- filter=53 channel=110
    0, -6, 4, -10, 0, 2, 2, -2, 6,
    -- filter=53 channel=111
    3, -2, -2, -3, -6, 0, -7, -9, -1,
    -- filter=53 channel=112
    0, 6, 1, 12, 7, 3, 12, 0, -2,
    -- filter=53 channel=113
    4, -4, -1, 2, 3, -3, -5, -2, 6,
    -- filter=53 channel=114
    2, 6, -3, -9, -1, 2, 4, 4, -7,
    -- filter=53 channel=115
    0, 1, -3, 3, -6, 0, 2, -1, 4,
    -- filter=53 channel=116
    -8, 4, 3, -11, -1, 7, 4, 0, 5,
    -- filter=53 channel=117
    -3, 5, 3, -11, -7, 8, 5, 2, -6,
    -- filter=53 channel=118
    3, -7, 0, 7, -7, 5, -1, 6, 7,
    -- filter=53 channel=119
    4, 0, 2, 6, -10, -1, -3, 0, 0,
    -- filter=53 channel=120
    -6, 3, 0, -6, 2, -1, 0, 4, -4,
    -- filter=53 channel=121
    -5, -5, -5, -5, -4, -3, -2, 1, 1,
    -- filter=53 channel=122
    -6, -7, -12, 9, 18, -6, 12, 0, -15,
    -- filter=53 channel=123
    7, 5, 0, 7, -1, -5, -5, -9, 0,
    -- filter=53 channel=124
    -5, 2, 2, -7, 0, 4, 0, 1, -4,
    -- filter=53 channel=125
    1, 1, 6, -7, 9, -5, 1, -3, -6,
    -- filter=53 channel=126
    0, 1, 0, -1, 0, 2, -12, 2, 7,
    -- filter=53 channel=127
    -9, 0, -2, -2, -4, -3, 2, 0, -2,
    -- filter=54 channel=0
    0, 5, 0, 9, 14, 0, 4, 1, -1,
    -- filter=54 channel=1
    0, -4, -11, 14, 12, 0, 9, 0, -6,
    -- filter=54 channel=2
    0, 2, -7, 2, 6, 0, 2, 5, -2,
    -- filter=54 channel=3
    6, 3, -7, -5, 0, -2, -3, 6, 4,
    -- filter=54 channel=4
    0, -4, -2, 0, 0, 3, -2, 4, 3,
    -- filter=54 channel=5
    1, -6, -7, 12, 7, -11, 9, -1, -12,
    -- filter=54 channel=6
    1, 3, -1, 1, 5, -1, -2, -5, -5,
    -- filter=54 channel=7
    -6, -5, -3, 5, -3, -6, 1, -1, 5,
    -- filter=54 channel=8
    2, -6, -5, -7, -5, 4, 7, -1, 5,
    -- filter=54 channel=9
    6, -2, 4, -3, 0, -3, 0, 3, 1,
    -- filter=54 channel=10
    -8, 0, -3, -6, -8, -6, 6, 6, 0,
    -- filter=54 channel=11
    -11, 2, 8, -12, -4, 0, -13, 3, 2,
    -- filter=54 channel=12
    -6, -5, 4, 0, 0, -7, -2, 0, 0,
    -- filter=54 channel=13
    5, 8, -1, -9, 1, 0, -5, -1, -4,
    -- filter=54 channel=14
    -7, -2, -1, 0, 6, -5, 4, -4, -2,
    -- filter=54 channel=15
    4, 8, 1, -11, 5, 4, -9, -4, -4,
    -- filter=54 channel=16
    3, 0, -11, 0, 0, -6, 4, -2, 0,
    -- filter=54 channel=17
    0, 7, 2, -4, 7, 3, -7, -3, 5,
    -- filter=54 channel=18
    2, 11, 11, -13, 4, 9, -13, -3, 12,
    -- filter=54 channel=19
    -3, 1, -4, 5, 5, -5, 4, 3, 6,
    -- filter=54 channel=20
    -3, 2, 6, -19, -14, 0, -12, -11, -6,
    -- filter=54 channel=21
    -1, -1, 2, 2, -4, 1, 7, -9, -4,
    -- filter=54 channel=22
    1, 8, 3, 0, 8, 5, -4, 2, 5,
    -- filter=54 channel=23
    -2, 11, 11, -12, -8, 2, -4, 6, -1,
    -- filter=54 channel=24
    1, -4, 0, -4, 0, -5, -5, -6, -5,
    -- filter=54 channel=25
    2, 4, 0, 5, 7, -6, 0, 4, -2,
    -- filter=54 channel=26
    -4, -10, 1, 6, -5, 0, 0, -1, -7,
    -- filter=54 channel=27
    8, 7, 8, 4, 0, 0, 1, 13, -4,
    -- filter=54 channel=28
    -4, 1, -6, 1, -3, -6, -1, 0, -1,
    -- filter=54 channel=29
    -7, -3, 3, -18, -5, 3, -13, -4, 7,
    -- filter=54 channel=30
    -2, -2, -2, -3, -1, -6, 8, 5, -4,
    -- filter=54 channel=31
    -7, -9, 12, -6, -8, 2, 1, -3, 1,
    -- filter=54 channel=32
    2, 5, 1, 0, -1, 5, -3, 1, -1,
    -- filter=54 channel=33
    2, -2, 4, 5, 2, -6, 1, 0, -3,
    -- filter=54 channel=34
    3, 0, 2, 2, 0, -3, 0, -6, -11,
    -- filter=54 channel=35
    -2, -2, -3, 0, 0, 2, -5, 4, 6,
    -- filter=54 channel=36
    -5, -9, 6, -11, -2, 4, 0, 1, 2,
    -- filter=54 channel=37
    -2, 2, -3, 16, 12, -3, 5, 7, 0,
    -- filter=54 channel=38
    3, 7, 7, -1, 4, -4, 6, 0, -6,
    -- filter=54 channel=39
    -7, -2, -5, -9, -9, 1, 0, -2, -5,
    -- filter=54 channel=40
    5, -6, 5, -3, -3, -2, -8, 0, -6,
    -- filter=54 channel=41
    -5, 3, -1, -11, -4, -4, -13, 0, -5,
    -- filter=54 channel=42
    0, -3, 2, 7, 7, -1, 1, -5, -5,
    -- filter=54 channel=43
    0, -1, 0, 0, -6, -3, -6, -3, 0,
    -- filter=54 channel=44
    -1, -1, -9, 10, 6, -10, 4, 7, 1,
    -- filter=54 channel=45
    -3, 2, 3, 0, -5, -7, 2, -2, -4,
    -- filter=54 channel=46
    -2, -6, -4, 0, -5, 3, -2, -6, 0,
    -- filter=54 channel=47
    0, -6, -9, 8, -1, -6, 11, -1, 2,
    -- filter=54 channel=48
    7, -4, -3, 0, 6, -4, 15, -5, 3,
    -- filter=54 channel=49
    -2, -3, -1, -9, 6, 2, -4, 8, 11,
    -- filter=54 channel=50
    -2, -5, 10, 6, -1, 2, 1, -2, 5,
    -- filter=54 channel=51
    5, -1, -4, -3, 2, -6, -1, 5, 7,
    -- filter=54 channel=52
    0, 4, 6, 2, 5, -6, -6, -4, 0,
    -- filter=54 channel=53
    -5, 4, 0, -9, 1, 5, -4, 5, -3,
    -- filter=54 channel=54
    4, 5, 2, -4, 1, -6, 4, 6, -3,
    -- filter=54 channel=55
    2, -3, 8, -13, -3, 1, -4, 4, 0,
    -- filter=54 channel=56
    7, 0, 0, 2, 6, 0, -3, 5, -10,
    -- filter=54 channel=57
    -7, 0, 6, 6, 0, 2, -2, -4, 2,
    -- filter=54 channel=58
    -5, -11, -1, 1, 0, -2, 2, -6, -5,
    -- filter=54 channel=59
    -1, 2, 5, 3, 3, 5, 10, 0, 8,
    -- filter=54 channel=60
    -7, 2, 1, 0, -5, 4, 6, -1, 2,
    -- filter=54 channel=61
    -4, 6, -5, -5, -4, -7, 2, 3, 1,
    -- filter=54 channel=62
    2, -4, 6, -6, 3, 1, -5, -3, -6,
    -- filter=54 channel=63
    -7, -11, 0, 3, -10, 1, -3, -9, -4,
    -- filter=54 channel=64
    4, -6, -1, -6, -4, 0, -8, -2, 0,
    -- filter=54 channel=65
    1, 5, 3, -1, 2, -7, -2, 0, 7,
    -- filter=54 channel=66
    -2, -1, -6, -7, 3, -7, -10, 7, -2,
    -- filter=54 channel=67
    0, -6, -5, -6, -3, 2, -2, -5, -6,
    -- filter=54 channel=68
    -5, -4, 0, -8, -7, -5, -3, 2, 7,
    -- filter=54 channel=69
    5, -2, 2, -5, 1, 2, 0, 6, -6,
    -- filter=54 channel=70
    -2, 6, 4, 3, 5, -4, 5, 3, -4,
    -- filter=54 channel=71
    4, -5, 5, 4, 2, 7, 7, 3, -3,
    -- filter=54 channel=72
    -10, -8, -2, -7, -7, -5, 4, -6, 3,
    -- filter=54 channel=73
    -2, -3, 3, -7, -3, 0, -6, 9, 4,
    -- filter=54 channel=74
    6, 5, 2, -6, 9, -12, 6, 0, -9,
    -- filter=54 channel=75
    10, -6, -8, 17, 11, 7, 1, -3, 0,
    -- filter=54 channel=76
    -10, -5, -2, -17, -13, 6, -14, 0, 6,
    -- filter=54 channel=77
    -5, 3, -6, -5, 4, -5, -2, 5, -7,
    -- filter=54 channel=78
    -4, -4, -7, -3, -2, -8, -2, -6, -8,
    -- filter=54 channel=79
    -2, 12, 12, -9, 7, 11, -4, 3, 8,
    -- filter=54 channel=80
    2, -10, -1, -4, -9, -10, 8, 3, -1,
    -- filter=54 channel=81
    6, 7, 2, -1, 4, 3, -6, 1, 4,
    -- filter=54 channel=82
    7, -2, 2, -3, 5, 3, -1, 3, 1,
    -- filter=54 channel=83
    -5, -7, -4, 2, 0, -6, 4, -3, 4,
    -- filter=54 channel=84
    1, 1, -4, -6, 6, 3, -1, 8, 1,
    -- filter=54 channel=85
    1, 0, 6, 0, 1, 0, 3, 6, 4,
    -- filter=54 channel=86
    7, -6, 3, -3, 0, 0, 0, -3, -6,
    -- filter=54 channel=87
    -2, 5, 3, -3, -2, 1, 0, -6, -5,
    -- filter=54 channel=88
    -8, -4, -2, -9, -8, -4, -2, -3, 1,
    -- filter=54 channel=89
    -1, 3, 6, -3, -1, 4, -9, 0, 1,
    -- filter=54 channel=90
    5, 4, -2, -6, -12, 4, 1, -10, 0,
    -- filter=54 channel=91
    6, 3, 1, 1, 1, 5, -2, 4, 0,
    -- filter=54 channel=92
    -2, -5, 1, 0, 1, -7, 2, 5, -3,
    -- filter=54 channel=93
    -1, -2, 1, 13, 10, -7, 5, -1, -3,
    -- filter=54 channel=94
    2, 5, -4, -2, -2, 3, -4, -5, 0,
    -- filter=54 channel=95
    5, -3, 5, 4, -4, 2, 3, 2, -8,
    -- filter=54 channel=96
    1, 6, -6, -4, -5, 4, -2, 0, -3,
    -- filter=54 channel=97
    5, 8, 4, 1, 6, 0, -1, 3, -2,
    -- filter=54 channel=98
    -4, -3, 4, -4, 4, -7, 5, 6, 0,
    -- filter=54 channel=99
    0, -5, 1, -10, -9, -9, -6, 4, 6,
    -- filter=54 channel=100
    -5, 6, 0, 0, 3, -6, -1, 3, -8,
    -- filter=54 channel=101
    3, 2, 4, 5, -1, -2, 4, 0, 6,
    -- filter=54 channel=102
    -4, -6, 3, 2, 7, -5, -7, 2, -3,
    -- filter=54 channel=103
    7, -9, -5, 6, -2, -1, 10, 7, -4,
    -- filter=54 channel=104
    -8, -11, -1, -2, 0, -10, 12, 5, 4,
    -- filter=54 channel=105
    -6, -2, -5, -6, 1, 0, -3, 0, 0,
    -- filter=54 channel=106
    0, 6, -1, -9, -4, 1, -9, -2, 7,
    -- filter=54 channel=107
    2, 1, 4, -10, -2, 7, -14, -9, -3,
    -- filter=54 channel=108
    -5, -7, -2, -1, 0, 5, -2, 1, 5,
    -- filter=54 channel=109
    2, 0, 3, 0, 6, -7, 9, -1, -2,
    -- filter=54 channel=110
    5, -1, -2, -11, -5, -1, 1, 0, -2,
    -- filter=54 channel=111
    -2, -2, 1, 6, -1, 3, 0, 5, 3,
    -- filter=54 channel=112
    -4, -3, 4, -1, -1, -9, -2, -2, -7,
    -- filter=54 channel=113
    -5, 8, -6, 2, 1, 4, 0, 5, -1,
    -- filter=54 channel=114
    0, 2, 2, 0, 15, 3, -7, 8, -2,
    -- filter=54 channel=115
    -2, -1, -6, -3, 2, 0, 0, -2, -2,
    -- filter=54 channel=116
    1, 6, 11, -3, -8, -2, 0, 9, 10,
    -- filter=54 channel=117
    4, -5, -3, -4, 3, -4, -1, 5, 7,
    -- filter=54 channel=118
    0, -3, 0, -1, -6, -2, -7, -1, 6,
    -- filter=54 channel=119
    1, -4, 0, 3, 5, -5, 0, 0, -9,
    -- filter=54 channel=120
    -7, 6, 2, -12, -1, -9, -1, 6, 8,
    -- filter=54 channel=121
    -7, 0, 3, 0, 1, -7, 3, 0, -2,
    -- filter=54 channel=122
    2, -7, -8, 8, -9, -12, 12, -7, -8,
    -- filter=54 channel=123
    2, 3, -6, 2, 3, -8, -3, -6, -7,
    -- filter=54 channel=124
    -6, 2, -3, -9, 0, 3, 4, -5, 1,
    -- filter=54 channel=125
    -5, -9, -3, 3, -10, 0, 5, 4, 8,
    -- filter=54 channel=126
    0, 8, 5, -10, 5, 10, -8, 2, -5,
    -- filter=54 channel=127
    -6, -6, 2, 1, 5, -3, -1, -4, 5,
    -- filter=55 channel=0
    2, 4, 3, 2, -4, 7, 1, -2, -8,
    -- filter=55 channel=1
    3, 3, 8, -3, -1, -4, -2, -1, 3,
    -- filter=55 channel=2
    -2, -3, -2, 2, 2, -5, 2, -1, -4,
    -- filter=55 channel=3
    0, 0, -3, 1, 6, 4, -6, -8, 0,
    -- filter=55 channel=4
    -5, 2, 0, -5, -1, 4, -1, 7, -1,
    -- filter=55 channel=5
    -1, 7, 7, 7, 2, 10, -8, -7, -4,
    -- filter=55 channel=6
    -1, 1, 2, 6, 0, -3, 0, 5, 6,
    -- filter=55 channel=7
    -2, -1, 3, 3, -1, -5, 7, 0, 4,
    -- filter=55 channel=8
    2, 2, 3, -5, -6, 1, -5, -4, 0,
    -- filter=55 channel=9
    -5, 4, 3, -1, -5, 2, 3, -5, 4,
    -- filter=55 channel=10
    1, -6, 0, -5, 5, 5, -4, -2, -5,
    -- filter=55 channel=11
    0, 0, 1, 5, 7, 0, 6, -7, 6,
    -- filter=55 channel=12
    6, 7, -3, 7, 0, 3, -4, -7, 2,
    -- filter=55 channel=13
    -6, -3, 3, -1, 0, -3, -1, -6, -3,
    -- filter=55 channel=14
    0, -1, -3, 0, 4, -4, 4, -5, 2,
    -- filter=55 channel=15
    -1, 0, -6, 4, 3, -5, 0, -3, -4,
    -- filter=55 channel=16
    -3, 5, 0, -2, 2, 3, 8, 3, 3,
    -- filter=55 channel=17
    -6, 4, 7, 6, 3, 6, 0, 2, -2,
    -- filter=55 channel=18
    -5, 4, -3, -4, -8, -5, 3, 4, -6,
    -- filter=55 channel=19
    2, 6, -6, 3, 0, -4, 0, -4, -2,
    -- filter=55 channel=20
    0, 1, 4, -1, -3, -2, -1, 5, -5,
    -- filter=55 channel=21
    -4, -2, 1, 4, -7, -3, 4, -4, 1,
    -- filter=55 channel=22
    6, 3, 3, -5, 5, 6, -8, 6, 6,
    -- filter=55 channel=23
    0, -5, 0, 3, -2, -2, -4, -8, -7,
    -- filter=55 channel=24
    -1, -3, -5, -4, -2, 0, 4, 2, 7,
    -- filter=55 channel=25
    4, -3, -5, 5, -9, 5, -4, 0, -7,
    -- filter=55 channel=26
    5, 7, -4, 6, 5, 1, 1, 8, -3,
    -- filter=55 channel=27
    -4, 4, 2, -6, -1, 0, -6, 3, -8,
    -- filter=55 channel=28
    3, -6, -5, -1, 0, 2, 6, -1, -5,
    -- filter=55 channel=29
    -6, 4, 5, -5, 0, 5, 1, 1, 3,
    -- filter=55 channel=30
    0, -1, -1, 5, -5, 5, -1, -7, 0,
    -- filter=55 channel=31
    4, 0, 0, -10, 0, 5, -1, -6, 7,
    -- filter=55 channel=32
    5, 5, 7, 0, 1, -6, -6, -6, 0,
    -- filter=55 channel=33
    -5, -3, 5, 3, 1, 5, -5, 0, -3,
    -- filter=55 channel=34
    7, 0, 2, 0, 1, 9, 0, -4, -3,
    -- filter=55 channel=35
    -1, 0, 6, 4, -2, -5, -2, 4, 5,
    -- filter=55 channel=36
    -6, -8, -3, 1, 2, -7, 6, -2, 0,
    -- filter=55 channel=37
    2, -3, 5, 6, -4, -2, -8, 0, 3,
    -- filter=55 channel=38
    -1, 6, 5, -6, 3, -6, 0, -6, 1,
    -- filter=55 channel=39
    5, -5, 1, 7, -2, -2, -1, 3, -6,
    -- filter=55 channel=40
    3, 5, -7, -5, -5, -1, 0, -1, -2,
    -- filter=55 channel=41
    4, -1, 0, -2, 5, -3, 8, -5, 2,
    -- filter=55 channel=42
    -2, 3, 7, -6, 1, -4, 0, -8, -7,
    -- filter=55 channel=43
    -4, 4, -2, 5, 2, 1, 3, -3, 4,
    -- filter=55 channel=44
    2, 3, -5, -6, -4, 0, -3, 0, -7,
    -- filter=55 channel=45
    -3, -1, -6, 1, -3, 0, -7, -4, -6,
    -- filter=55 channel=46
    -6, -5, -1, 0, 3, -2, -5, -4, -7,
    -- filter=55 channel=47
    3, 7, 0, 6, -5, 6, 7, -5, -2,
    -- filter=55 channel=48
    6, -7, 1, -1, 0, 3, 5, 3, 0,
    -- filter=55 channel=49
    -7, 0, -2, 6, 5, -5, 5, 2, 0,
    -- filter=55 channel=50
    0, 5, 0, -3, -7, 6, -3, 5, 2,
    -- filter=55 channel=51
    0, -3, -7, 7, 0, 0, -1, 5, 2,
    -- filter=55 channel=52
    2, 0, 0, -1, 2, 2, 4, -5, 0,
    -- filter=55 channel=53
    -4, 1, 0, -1, -7, 4, -6, 1, 6,
    -- filter=55 channel=54
    0, 6, 6, 0, 7, -4, -3, 3, 6,
    -- filter=55 channel=55
    -3, 2, -7, -6, -6, -2, 5, 0, -3,
    -- filter=55 channel=56
    1, -3, 4, 2, 7, 0, 0, -6, 5,
    -- filter=55 channel=57
    -7, -7, 4, 5, 3, 5, 4, 2, 1,
    -- filter=55 channel=58
    4, 0, 4, -4, 4, 0, -6, 3, -5,
    -- filter=55 channel=59
    -2, -2, -3, 0, -6, 4, 5, 2, -5,
    -- filter=55 channel=60
    -1, 2, 5, 7, 5, 3, 1, 5, -4,
    -- filter=55 channel=61
    6, 1, 1, 4, -3, 8, 0, 1, 0,
    -- filter=55 channel=62
    2, 3, 4, 1, 3, 4, -3, 3, -4,
    -- filter=55 channel=63
    7, 2, 3, 6, 3, -4, 6, 6, 4,
    -- filter=55 channel=64
    -1, 2, 0, -2, -1, -2, -4, 7, 6,
    -- filter=55 channel=65
    7, 0, 3, -4, -3, 2, 5, 0, -7,
    -- filter=55 channel=66
    3, -4, 1, 3, -2, -7, 1, -2, -5,
    -- filter=55 channel=67
    -2, 2, 1, 3, 6, -5, 2, 1, -4,
    -- filter=55 channel=68
    -7, 0, -5, -6, 1, -7, 6, 6, 1,
    -- filter=55 channel=69
    -4, -3, 1, 0, 6, 3, 1, -2, -6,
    -- filter=55 channel=70
    4, 0, 2, 0, -4, 4, -4, -5, -5,
    -- filter=55 channel=71
    -2, 6, -5, 2, -5, -4, -5, -1, -2,
    -- filter=55 channel=72
    -8, -2, -2, -8, -3, -5, 3, -5, 4,
    -- filter=55 channel=73
    4, 6, 0, -5, -6, 1, 0, -7, -7,
    -- filter=55 channel=74
    -3, 1, -4, -4, -5, 2, 3, 5, 3,
    -- filter=55 channel=75
    -2, 5, 12, -5, 5, 0, -3, -7, 4,
    -- filter=55 channel=76
    -1, -7, 0, -6, 0, 3, -4, 0, 7,
    -- filter=55 channel=77
    0, 6, -4, -4, 1, -2, 0, 0, -1,
    -- filter=55 channel=78
    0, -2, 4, 0, -5, 5, 4, 6, 6,
    -- filter=55 channel=79
    -6, -8, 5, -7, -4, -3, -9, -3, -8,
    -- filter=55 channel=80
    -9, 5, 5, -1, -7, -1, 7, 1, -1,
    -- filter=55 channel=81
    -6, -7, 5, -5, -5, 0, -7, -3, 4,
    -- filter=55 channel=82
    -6, -2, -2, -6, 1, 7, -2, 5, 0,
    -- filter=55 channel=83
    0, 1, -2, 1, 2, -6, 2, -3, -6,
    -- filter=55 channel=84
    -5, -3, 1, 0, -2, 4, -3, -5, 0,
    -- filter=55 channel=85
    7, 6, -2, 1, 2, -3, -3, 7, 1,
    -- filter=55 channel=86
    5, 4, 6, 2, 1, 2, -2, -4, -6,
    -- filter=55 channel=87
    7, 4, -7, -5, 2, 2, 6, -3, 0,
    -- filter=55 channel=88
    -5, 1, -6, -4, 5, 4, 2, -3, -3,
    -- filter=55 channel=89
    -7, 3, -7, -1, -2, -4, -1, -1, 0,
    -- filter=55 channel=90
    0, 6, -1, -6, 7, 0, 0, 0, 6,
    -- filter=55 channel=91
    4, -4, 1, 0, 1, 4, -6, 1, -7,
    -- filter=55 channel=92
    0, 0, 4, -2, -5, 5, -1, 2, -6,
    -- filter=55 channel=93
    5, 6, 4, -6, 4, -4, 0, 1, -7,
    -- filter=55 channel=94
    -6, -2, -4, -3, -5, -4, -6, -7, -2,
    -- filter=55 channel=95
    -5, 7, -5, 3, 7, -1, 4, 2, 0,
    -- filter=55 channel=96
    -7, 5, 2, 4, -3, 2, 1, 2, -3,
    -- filter=55 channel=97
    -1, -4, 2, -4, 6, 3, -2, 0, 5,
    -- filter=55 channel=98
    -5, -1, 0, 3, 4, -5, -5, 0, -2,
    -- filter=55 channel=99
    0, 4, 0, 0, 2, 3, 8, 0, -3,
    -- filter=55 channel=100
    -6, -5, -4, 3, 4, -6, 7, -6, 1,
    -- filter=55 channel=101
    1, 2, -6, 2, 2, 0, 8, 0, 1,
    -- filter=55 channel=102
    -5, 0, 2, 2, -5, -1, 3, -3, 4,
    -- filter=55 channel=103
    -3, -3, 8, 5, -6, 7, 6, 0, 3,
    -- filter=55 channel=104
    -3, -4, 6, -1, -8, 5, 6, 8, 0,
    -- filter=55 channel=105
    -3, -2, -6, 6, -6, -1, -5, 5, 0,
    -- filter=55 channel=106
    -4, 3, 4, 0, 5, 5, -5, 1, 0,
    -- filter=55 channel=107
    5, -5, 0, 3, -3, 2, 3, -7, -3,
    -- filter=55 channel=108
    0, -6, -2, 6, 5, 5, 3, 6, -1,
    -- filter=55 channel=109
    -5, 6, -3, 5, -2, 5, 1, -6, 3,
    -- filter=55 channel=110
    2, 5, 6, -3, -5, -2, 6, -4, 6,
    -- filter=55 channel=111
    4, 6, 2, -1, 1, 6, 3, 2, -2,
    -- filter=55 channel=112
    -5, -5, 0, 5, 1, 5, -4, -3, 4,
    -- filter=55 channel=113
    2, 1, 7, 0, -3, 3, 4, -9, 3,
    -- filter=55 channel=114
    -2, 1, -6, -2, -4, -6, -9, 0, 2,
    -- filter=55 channel=115
    2, -6, 0, -3, 1, -1, -6, 4, -6,
    -- filter=55 channel=116
    3, 0, -1, 2, -3, 0, 2, -1, 5,
    -- filter=55 channel=117
    -3, 3, 3, -5, 0, 2, 6, -2, -2,
    -- filter=55 channel=118
    6, -5, 1, -2, -4, 3, -3, 5, -5,
    -- filter=55 channel=119
    4, 0, 3, 0, -5, 9, 0, 0, 0,
    -- filter=55 channel=120
    3, -4, 0, -2, -6, -1, -5, 1, 0,
    -- filter=55 channel=121
    5, 1, 1, -4, 1, -3, 4, -3, 3,
    -- filter=55 channel=122
    -2, 0, 8, -4, -2, -1, 2, 6, -4,
    -- filter=55 channel=123
    -6, 2, 0, -4, 3, -4, 5, 6, -3,
    -- filter=55 channel=124
    4, 3, -7, 3, 5, -4, -5, -2, 4,
    -- filter=55 channel=125
    -3, -8, -8, -7, 1, 2, 7, 3, -1,
    -- filter=55 channel=126
    3, 7, -3, -5, -1, -3, -4, 0, -7,
    -- filter=55 channel=127
    0, 1, 0, 2, 6, 0, -3, 7, -7,
    -- filter=56 channel=0
    6, -5, -4, -3, 4, 1, 8, -1, 1,
    -- filter=56 channel=1
    1, 7, -4, 3, -2, -7, 10, 9, -7,
    -- filter=56 channel=2
    0, 6, -5, -1, 5, -3, -1, 0, 1,
    -- filter=56 channel=3
    5, -3, 1, 3, -3, -5, 5, 5, 5,
    -- filter=56 channel=4
    7, 6, 6, 0, 7, -4, 0, 1, 6,
    -- filter=56 channel=5
    -4, 5, -8, 8, 4, -8, 0, -3, -6,
    -- filter=56 channel=6
    4, 6, 4, 0, -1, 2, 5, -7, 1,
    -- filter=56 channel=7
    -5, 0, -1, -5, 1, 4, 4, -4, -2,
    -- filter=56 channel=8
    3, -6, 1, -5, 3, 1, -1, -5, -1,
    -- filter=56 channel=9
    -2, 6, -4, 4, -6, 0, -5, 0, -4,
    -- filter=56 channel=10
    -2, -5, 6, -7, -4, 6, 4, 0, -2,
    -- filter=56 channel=11
    -5, 0, 1, 7, 1, -7, -2, -2, -3,
    -- filter=56 channel=12
    6, 0, 0, 0, 0, 4, -5, -3, -3,
    -- filter=56 channel=13
    -7, 3, -1, -2, -1, 5, 5, -2, 2,
    -- filter=56 channel=14
    2, 4, 6, -6, -7, 1, 6, -3, -6,
    -- filter=56 channel=15
    -3, 3, 0, -3, 6, 5, 1, -7, 6,
    -- filter=56 channel=16
    -2, -6, -2, 3, -4, -4, 0, -5, -4,
    -- filter=56 channel=17
    4, -2, 3, -2, -3, -6, 6, -3, -3,
    -- filter=56 channel=18
    -4, -7, 2, 2, 0, -3, 3, -4, -6,
    -- filter=56 channel=19
    0, 0, -1, 4, 4, -4, -5, -3, 6,
    -- filter=56 channel=20
    -1, -5, -4, -6, -1, -3, -6, 2, 7,
    -- filter=56 channel=21
    -3, 4, 0, 3, 2, 0, -2, 0, -3,
    -- filter=56 channel=22
    -2, 0, -5, 5, -1, 1, -3, 7, 2,
    -- filter=56 channel=23
    -5, 5, 6, -4, -5, -3, -5, 7, 3,
    -- filter=56 channel=24
    5, -5, -1, 0, 2, -6, 4, 0, 7,
    -- filter=56 channel=25
    3, -5, 7, -7, 5, -6, -3, -2, -1,
    -- filter=56 channel=26
    2, 3, 5, 1, 6, -3, 4, 4, 5,
    -- filter=56 channel=27
    1, -8, 5, 0, -2, 7, 0, -5, -10,
    -- filter=56 channel=28
    -4, -7, -1, 0, -5, 1, -6, 5, 0,
    -- filter=56 channel=29
    6, 5, 4, 0, 1, 2, -5, 1, -1,
    -- filter=56 channel=30
    0, 4, 0, 0, 1, 0, 3, -3, 5,
    -- filter=56 channel=31
    -1, -4, 2, 3, 0, 2, 4, -5, -7,
    -- filter=56 channel=32
    -4, 3, 3, -2, -2, -6, 0, -6, -8,
    -- filter=56 channel=33
    4, 0, 1, 4, 0, 6, -4, 0, 3,
    -- filter=56 channel=34
    4, 3, 8, -2, 6, 4, -5, 1, 5,
    -- filter=56 channel=35
    -3, -1, -3, 0, 0, 7, 0, 1, 2,
    -- filter=56 channel=36
    2, 0, 5, 4, -3, -4, -4, 5, 2,
    -- filter=56 channel=37
    7, 3, 4, 3, 2, 5, 2, 6, -7,
    -- filter=56 channel=38
    5, -3, 4, -1, -8, -1, -1, 0, -1,
    -- filter=56 channel=39
    6, 0, 1, -5, -1, -4, -6, -5, -1,
    -- filter=56 channel=40
    -1, -2, 5, -4, -3, 6, -4, 2, 3,
    -- filter=56 channel=41
    0, 7, -8, -2, 7, -6, 5, 5, 7,
    -- filter=56 channel=42
    5, -4, -6, 6, -7, 1, 8, -4, -1,
    -- filter=56 channel=43
    2, 4, 0, 3, -3, -4, 0, 3, -5,
    -- filter=56 channel=44
    -6, 1, -2, -1, 5, 6, 8, 4, -5,
    -- filter=56 channel=45
    0, -5, -6, 6, -2, 0, -3, -1, -6,
    -- filter=56 channel=46
    6, 3, 5, 5, 1, 1, -2, 1, 7,
    -- filter=56 channel=47
    -3, 2, 2, 3, -5, 0, -4, -6, 2,
    -- filter=56 channel=48
    -4, 1, -2, 3, 5, -4, -7, 0, 3,
    -- filter=56 channel=49
    4, -8, -6, -5, -2, -3, -6, -3, 0,
    -- filter=56 channel=50
    1, -3, -5, 6, 4, -4, 0, -6, -4,
    -- filter=56 channel=51
    5, 5, -5, 2, -5, -5, 0, -1, 0,
    -- filter=56 channel=52
    5, -3, -4, 3, 1, 1, 1, -5, -5,
    -- filter=56 channel=53
    3, -2, 6, -2, -4, -3, 2, -6, -6,
    -- filter=56 channel=54
    5, -4, 4, 2, 1, 5, -2, 0, -3,
    -- filter=56 channel=55
    -5, 4, -5, 5, 4, -1, -8, -3, 2,
    -- filter=56 channel=56
    7, -4, 0, 1, 0, 1, 5, -4, 6,
    -- filter=56 channel=57
    4, -5, -7, -6, -1, 4, -2, -7, 6,
    -- filter=56 channel=58
    5, -1, -4, 8, 3, -1, 1, -5, 0,
    -- filter=56 channel=59
    -1, -4, -3, 5, 2, -7, -4, -4, -4,
    -- filter=56 channel=60
    6, 4, 0, -4, -2, -1, -2, 2, -2,
    -- filter=56 channel=61
    3, -3, -1, -5, 4, 5, -7, -6, 3,
    -- filter=56 channel=62
    0, 4, -2, -6, 5, -2, -7, -4, 5,
    -- filter=56 channel=63
    -2, -7, -4, 0, 3, -3, 0, 6, 0,
    -- filter=56 channel=64
    -5, -2, 3, -7, -4, 4, -5, -6, 3,
    -- filter=56 channel=65
    -7, -6, 1, 0, 3, -7, 0, 4, 1,
    -- filter=56 channel=66
    -5, 1, -6, -3, -1, -2, 6, 2, 1,
    -- filter=56 channel=67
    0, -6, 4, -2, 6, -4, -6, 1, 3,
    -- filter=56 channel=68
    -5, -7, 0, 0, 0, 3, -2, 3, 7,
    -- filter=56 channel=69
    -4, 0, -6, 0, -1, -2, 1, 6, 1,
    -- filter=56 channel=70
    1, 7, 10, -2, -7, 1, 3, -6, -1,
    -- filter=56 channel=71
    -7, 1, 8, 2, 4, 1, 0, 2, -3,
    -- filter=56 channel=72
    -1, 2, 3, 1, 5, 3, 3, 6, -8,
    -- filter=56 channel=73
    0, 2, 4, 0, 6, 0, -7, 6, -2,
    -- filter=56 channel=74
    0, 7, 0, 4, 0, -3, 1, -2, -6,
    -- filter=56 channel=75
    6, -3, 1, 8, -3, -6, 9, -1, 2,
    -- filter=56 channel=76
    1, 8, 5, 0, -2, -6, 2, 2, -6,
    -- filter=56 channel=77
    2, -2, -4, 1, 0, -5, -5, 4, 0,
    -- filter=56 channel=78
    0, 7, 4, -5, 1, 2, 7, 4, 3,
    -- filter=56 channel=79
    2, 0, -5, 4, -1, -4, -1, 1, -3,
    -- filter=56 channel=80
    -4, -5, 0, -2, 5, -3, -3, -6, 1,
    -- filter=56 channel=81
    -1, -6, -4, -5, -4, -7, -2, -5, -5,
    -- filter=56 channel=82
    6, 3, 2, -5, 2, 7, 5, -7, 6,
    -- filter=56 channel=83
    0, 4, 3, 6, -4, 1, 6, -2, -7,
    -- filter=56 channel=84
    -4, 4, -5, -5, 5, 1, 1, 6, 2,
    -- filter=56 channel=85
    -1, -3, 0, -4, 0, -6, -7, -2, -7,
    -- filter=56 channel=86
    7, 0, 6, -2, 4, -4, -4, -3, -4,
    -- filter=56 channel=87
    -2, 3, 3, 0, -6, 4, 1, -1, 4,
    -- filter=56 channel=88
    -3, 0, 7, -5, 2, 0, -2, 1, -2,
    -- filter=56 channel=89
    3, -6, -4, 2, 1, 6, -4, -2, -6,
    -- filter=56 channel=90
    -4, 3, 10, -6, 3, 2, -6, 3, 6,
    -- filter=56 channel=91
    0, -8, 8, 8, 0, 0, -6, 0, 2,
    -- filter=56 channel=92
    0, -3, -3, -6, -5, 8, -6, -3, 0,
    -- filter=56 channel=93
    0, -1, 0, 0, 5, -1, -2, -7, -8,
    -- filter=56 channel=94
    -1, -3, 5, -6, 5, -4, -3, -1, -3,
    -- filter=56 channel=95
    7, -3, 0, -1, -2, -7, 4, 0, 0,
    -- filter=56 channel=96
    -2, 4, -7, 6, -1, -3, 6, 2, 5,
    -- filter=56 channel=97
    2, 6, 3, 2, -3, -1, -4, 7, 7,
    -- filter=56 channel=98
    0, -7, -2, -5, -7, -8, -7, 2, -10,
    -- filter=56 channel=99
    -8, 8, 6, 4, 2, 8, -8, 3, 0,
    -- filter=56 channel=100
    0, -6, 6, 0, 1, 5, -6, 6, 1,
    -- filter=56 channel=101
    -6, 0, 0, 8, 2, -3, -1, 6, 7,
    -- filter=56 channel=102
    4, 4, -3, 4, -3, -2, -4, 1, 1,
    -- filter=56 channel=103
    0, 0, 3, -7, -3, -7, 1, 1, -5,
    -- filter=56 channel=104
    -5, -9, 7, -5, 1, 1, -2, -1, -3,
    -- filter=56 channel=105
    -3, 4, 3, 4, -8, 3, -3, 3, -1,
    -- filter=56 channel=106
    -6, 7, -4, 0, 3, 0, -1, 5, 0,
    -- filter=56 channel=107
    5, 5, -1, 5, 4, -2, 5, 8, 0,
    -- filter=56 channel=108
    -3, -6, -1, -1, 0, -6, 1, 1, -2,
    -- filter=56 channel=109
    -9, -7, 7, -1, -1, 6, -1, -2, -4,
    -- filter=56 channel=110
    3, -2, 5, -1, -5, -4, -3, 5, -5,
    -- filter=56 channel=111
    -3, 0, 0, 6, -6, -1, -6, 3, 1,
    -- filter=56 channel=112
    2, 1, 0, -6, 3, 4, 6, -7, -3,
    -- filter=56 channel=113
    -8, 0, 0, -7, -6, -3, 5, -3, -2,
    -- filter=56 channel=114
    3, 0, 0, 2, 1, 4, 5, -2, -5,
    -- filter=56 channel=115
    -7, 7, -5, 6, -1, -3, -5, -6, 1,
    -- filter=56 channel=116
    -3, -5, 1, -3, -4, -4, 0, 2, -2,
    -- filter=56 channel=117
    4, 6, -1, 0, 4, 2, 0, -5, -2,
    -- filter=56 channel=118
    -1, 5, 6, -3, -6, 5, -4, 4, 0,
    -- filter=56 channel=119
    4, 7, -3, 5, 5, 7, -7, -6, 1,
    -- filter=56 channel=120
    -4, 0, -2, -4, 4, -1, -8, -2, 3,
    -- filter=56 channel=121
    -2, -3, -3, -6, 3, -7, 5, 4, -3,
    -- filter=56 channel=122
    6, -2, 8, -2, 1, 7, 0, -2, -6,
    -- filter=56 channel=123
    -5, 1, 0, 5, 0, 7, -1, 0, 3,
    -- filter=56 channel=124
    0, 3, -5, -5, 0, 0, -3, 0, -3,
    -- filter=56 channel=125
    -1, -9, 3, 3, -3, 1, 3, -5, 1,
    -- filter=56 channel=126
    -6, 0, -1, 3, 2, -5, 0, 0, 3,
    -- filter=56 channel=127
    -1, -6, -4, -6, 5, 7, 0, 0, 0,
    -- filter=57 channel=0
    4, -11, -8, 9, 10, -3, 0, -8, -5,
    -- filter=57 channel=1
    -3, -2, -12, -10, -3, 7, 4, -7, 3,
    -- filter=57 channel=2
    -1, 0, 5, -6, -7, 6, 2, 9, -5,
    -- filter=57 channel=3
    2, -1, -12, 14, 14, -8, -5, 12, 4,
    -- filter=57 channel=4
    -3, 2, -11, 3, 0, 8, 18, 18, -3,
    -- filter=57 channel=5
    -2, -8, -1, 2, 8, -1, -3, 6, 7,
    -- filter=57 channel=6
    -9, 5, -3, 0, -7, -8, 1, 0, 2,
    -- filter=57 channel=7
    -7, 1, 7, 4, 3, -5, -5, -2, -5,
    -- filter=57 channel=8
    0, 0, -6, -1, -7, 2, 0, 5, 0,
    -- filter=57 channel=9
    5, 3, 0, 0, 11, -1, -8, -3, -3,
    -- filter=57 channel=10
    4, -1, -1, -2, 15, 7, -11, -13, -1,
    -- filter=57 channel=11
    0, -4, 5, -2, 1, 4, 1, 0, 0,
    -- filter=57 channel=12
    -7, 4, -7, -11, -5, -4, -7, -9, -1,
    -- filter=57 channel=13
    9, 3, -9, -1, 11, 0, -11, -18, -10,
    -- filter=57 channel=14
    3, -2, -6, -1, 7, 3, -1, 5, -3,
    -- filter=57 channel=15
    10, -5, 0, 2, 1, 7, -4, -5, -3,
    -- filter=57 channel=16
    4, 5, -9, 2, 2, -2, -8, -2, 0,
    -- filter=57 channel=17
    -7, -4, 0, 4, 0, -3, 1, -4, 5,
    -- filter=57 channel=18
    1, -1, -4, -1, 4, 10, -5, -14, -4,
    -- filter=57 channel=19
    -5, 1, -3, -7, 4, 3, 1, 2, -1,
    -- filter=57 channel=20
    0, 1, -6, 0, -3, -8, -6, -7, -5,
    -- filter=57 channel=21
    8, 4, -3, 2, 4, 3, -11, -1, -9,
    -- filter=57 channel=22
    -2, 1, -1, 7, 10, 0, -10, -7, 4,
    -- filter=57 channel=23
    3, -8, -6, 19, 23, 6, -22, -14, 0,
    -- filter=57 channel=24
    -7, -5, 4, -4, 3, 0, -3, 3, 5,
    -- filter=57 channel=25
    4, 10, 1, -7, 17, 11, -10, -20, -10,
    -- filter=57 channel=26
    1, -3, -1, -3, 0, 2, 8, -6, 5,
    -- filter=57 channel=27
    14, -1, -7, -3, 20, 10, -13, -21, 5,
    -- filter=57 channel=28
    -1, 5, -5, 4, -4, -6, -3, 5, -4,
    -- filter=57 channel=29
    -2, -7, -8, -10, -5, -4, 3, -5, -7,
    -- filter=57 channel=30
    9, -7, 0, -4, 4, 9, -9, -16, -6,
    -- filter=57 channel=31
    10, 7, 1, 5, 24, 13, -23, -10, -3,
    -- filter=57 channel=32
    0, 1, -5, -5, 17, 10, -8, -15, 1,
    -- filter=57 channel=33
    0, 4, 0, 9, 24, -5, -21, -16, 6,
    -- filter=57 channel=34
    1, -15, -3, 3, 4, 2, -15, 0, 6,
    -- filter=57 channel=35
    -2, 6, -5, 3, 0, -2, -1, -4, 0,
    -- filter=57 channel=36
    0, 2, 0, -2, -4, 0, -2, -1, 2,
    -- filter=57 channel=37
    6, -2, -2, 3, -2, 3, 0, -1, 0,
    -- filter=57 channel=38
    1, -5, -3, 0, 15, -1, -3, -6, -2,
    -- filter=57 channel=39
    2, -7, -1, -7, -4, 1, 6, -1, -2,
    -- filter=57 channel=40
    0, -2, 3, -5, 0, 2, 1, -4, 0,
    -- filter=57 channel=41
    -8, 1, 3, -23, -14, 8, 7, -7, -7,
    -- filter=57 channel=42
    5, 0, 2, 0, 4, 0, -7, -1, -1,
    -- filter=57 channel=43
    4, 0, -1, 6, -2, -5, -13, -3, -1,
    -- filter=57 channel=44
    -3, 3, 1, 3, 8, 8, 1, -3, 4,
    -- filter=57 channel=45
    2, -5, 0, 7, 4, -7, -5, -4, -4,
    -- filter=57 channel=46
    1, 2, -2, -5, -8, 7, -5, 0, -3,
    -- filter=57 channel=47
    6, 2, -9, 12, 8, 4, -14, -3, -2,
    -- filter=57 channel=48
    4, -1, -1, -8, 2, 5, -2, -19, -10,
    -- filter=57 channel=49
    1, 3, -10, -12, 7, 5, 8, 6, -4,
    -- filter=57 channel=50
    5, 6, -5, 10, 20, 0, -8, -10, 6,
    -- filter=57 channel=51
    6, 3, 4, 4, 3, 2, 3, -7, -6,
    -- filter=57 channel=52
    1, -6, 0, 0, -5, 0, -2, 3, 7,
    -- filter=57 channel=53
    0, -1, 0, 0, 6, 2, -2, 3, 0,
    -- filter=57 channel=54
    3, -3, 0, 2, 0, -3, -4, 5, 3,
    -- filter=57 channel=55
    11, -3, 0, 0, 10, -1, -16, -10, -8,
    -- filter=57 channel=56
    6, -9, -3, 3, -2, 0, 0, -3, -8,
    -- filter=57 channel=57
    4, 3, 5, -2, -5, 8, 0, 6, -7,
    -- filter=57 channel=58
    -4, 4, -2, -2, 2, 5, -1, 0, -6,
    -- filter=57 channel=59
    7, 15, 4, 1, 14, 13, -11, -13, -7,
    -- filter=57 channel=60
    -5, 6, -4, -5, -1, 0, -3, -6, -4,
    -- filter=57 channel=61
    0, -8, -5, -9, -6, -7, 6, -3, -5,
    -- filter=57 channel=62
    -6, 6, 1, -1, 4, 6, -3, 5, -5,
    -- filter=57 channel=63
    3, -3, 5, -5, -6, -4, -2, -7, -9,
    -- filter=57 channel=64
    4, -6, 2, -1, 0, 7, 6, -4, -7,
    -- filter=57 channel=65
    4, 1, -5, 7, -6, 0, -2, -4, 5,
    -- filter=57 channel=66
    -1, 0, 0, -9, 1, -5, -6, -11, -3,
    -- filter=57 channel=67
    5, -3, -2, -2, -6, 5, -6, 0, -1,
    -- filter=57 channel=68
    6, 1, 2, -2, 1, 5, 11, -2, -7,
    -- filter=57 channel=69
    6, -5, -4, -4, 2, 2, -5, 0, 2,
    -- filter=57 channel=70
    2, 3, -5, 4, 14, 4, -8, -9, 1,
    -- filter=57 channel=71
    0, -7, 0, 8, 2, 4, -11, 6, -1,
    -- filter=57 channel=72
    8, 2, 1, -2, 17, 0, -9, -17, 1,
    -- filter=57 channel=73
    2, -3, -5, -13, 0, 3, 2, -1, 4,
    -- filter=57 channel=74
    1, -3, -7, 8, 9, 3, -12, -1, 5,
    -- filter=57 channel=75
    0, -5, -13, 10, 19, 0, -16, -15, -7,
    -- filter=57 channel=76
    -2, -3, 5, -8, -2, 1, 0, -7, -11,
    -- filter=57 channel=77
    0, 2, 5, -3, -5, 2, 2, 0, 0,
    -- filter=57 channel=78
    0, 4, -4, -1, -4, 0, -4, -3, 6,
    -- filter=57 channel=79
    2, -3, -2, -6, 20, 12, -18, -18, -6,
    -- filter=57 channel=80
    12, 10, -7, 0, 14, 9, -6, -27, -2,
    -- filter=57 channel=81
    -3, 4, -2, -4, 1, -6, 4, 0, -5,
    -- filter=57 channel=82
    -4, -8, 1, 5, -3, -3, 3, 4, 0,
    -- filter=57 channel=83
    9, 11, -1, -6, 1, 0, 6, -7, 2,
    -- filter=57 channel=84
    -3, -3, -8, -5, -1, -3, -3, -5, -7,
    -- filter=57 channel=85
    6, 3, 2, 2, 2, -3, 6, -2, 1,
    -- filter=57 channel=86
    0, -6, -7, -1, 2, 1, -1, -8, -3,
    -- filter=57 channel=87
    -6, -4, -6, 4, -2, 2, 3, -2, -2,
    -- filter=57 channel=88
    -5, 0, 6, -5, -8, 6, 0, 0, -6,
    -- filter=57 channel=89
    0, 6, -6, 3, 18, 0, -14, -9, 1,
    -- filter=57 channel=90
    0, -6, 9, 0, 0, 3, -10, -5, 9,
    -- filter=57 channel=91
    11, 6, -4, -15, 6, 14, -3, -6, -1,
    -- filter=57 channel=92
    0, -3, -3, 4, 6, 1, -7, -1, 8,
    -- filter=57 channel=93
    8, 2, -3, 0, 0, -3, 0, -9, -6,
    -- filter=57 channel=94
    -1, 0, -6, -6, -5, 0, 3, -6, -4,
    -- filter=57 channel=95
    2, -6, 1, 6, 5, 1, -5, -5, -1,
    -- filter=57 channel=96
    1, 5, 3, -1, -3, 0, -5, 4, -5,
    -- filter=57 channel=97
    0, -5, -8, 13, 14, -6, -13, 0, 12,
    -- filter=57 channel=98
    2, -1, -3, 3, 24, 10, -9, -7, -6,
    -- filter=57 channel=99
    12, 3, -3, 2, 12, 1, -20, -17, -1,
    -- filter=57 channel=100
    0, 0, 3, 5, -9, -3, -8, -6, 5,
    -- filter=57 channel=101
    0, 1, -5, 1, 1, 2, 15, 3, 6,
    -- filter=57 channel=102
    -4, 4, 2, 5, -1, -3, -6, 7, 6,
    -- filter=57 channel=103
    9, 1, -11, 17, 9, 3, -16, -3, -5,
    -- filter=57 channel=104
    1, 5, -3, -1, 3, 1, -8, -14, 4,
    -- filter=57 channel=105
    4, 0, 6, -8, -8, -7, -7, -8, 0,
    -- filter=57 channel=106
    -8, 0, 2, 3, -6, 7, 7, 0, 0,
    -- filter=57 channel=107
    -1, -1, 1, 3, 3, -1, -9, 0, -5,
    -- filter=57 channel=108
    -5, 0, 4, -5, -1, 2, 3, -2, -9,
    -- filter=57 channel=109
    12, 7, 3, -9, 14, 10, -13, -10, -1,
    -- filter=57 channel=110
    0, 0, -1, 0, 1, -1, -7, -1, -1,
    -- filter=57 channel=111
    1, 1, -1, 1, -3, -4, 3, 1, 5,
    -- filter=57 channel=112
    6, -8, 0, 5, 10, 3, -1, -2, 1,
    -- filter=57 channel=113
    1, 0, -9, 17, 20, 2, -15, -4, 7,
    -- filter=57 channel=114
    0, 2, -12, -8, 10, 10, 1, -16, -5,
    -- filter=57 channel=115
    1, 6, -2, 0, -3, -3, -4, 0, -5,
    -- filter=57 channel=116
    0, 12, -6, -16, 8, 14, 3, -9, 0,
    -- filter=57 channel=117
    6, 0, 2, 2, -4, 4, 2, -6, 0,
    -- filter=57 channel=118
    0, 2, 6, -7, 1, -2, -6, -5, -1,
    -- filter=57 channel=119
    3, -7, -3, 4, -9, -8, -3, -2, 0,
    -- filter=57 channel=120
    0, 2, -5, -3, 4, 8, -1, -3, 0,
    -- filter=57 channel=121
    2, 0, -5, 6, -3, 3, -6, -2, -4,
    -- filter=57 channel=122
    0, 0, 3, -2, 7, 1, -14, -17, -6,
    -- filter=57 channel=123
    0, 2, 2, 11, 6, 1, -10, 11, 3,
    -- filter=57 channel=124
    -3, -9, -1, -2, -2, -6, 0, -1, 2,
    -- filter=57 channel=125
    2, 4, 3, -10, 0, 9, -1, -10, -2,
    -- filter=57 channel=126
    2, -2, 4, -3, 9, 7, -16, -14, -2,
    -- filter=57 channel=127
    -5, 1, 0, -1, -1, 5, -7, -6, -6,
    -- filter=58 channel=0
    -21, -18, -3, 9, 2, 6, 13, 5, 14,
    -- filter=58 channel=1
    -13, -12, -8, 6, 3, 1, 19, 12, 9,
    -- filter=58 channel=2
    10, 12, -3, 4, -2, -4, 4, 5, 2,
    -- filter=58 channel=3
    17, 16, 7, 20, 31, -5, 3, 4, 8,
    -- filter=58 channel=4
    21, 14, -3, 9, -4, 8, 9, 22, 1,
    -- filter=58 channel=5
    -21, -7, -1, 8, 19, 3, 5, 14, 11,
    -- filter=58 channel=6
    10, 6, -1, 2, -5, -4, -1, -8, -7,
    -- filter=58 channel=7
    -3, 0, -2, -1, -5, 4, 1, -1, 3,
    -- filter=58 channel=8
    5, 8, -5, -5, -2, 0, 5, 10, 10,
    -- filter=58 channel=9
    0, -5, 3, 3, 6, 6, -7, 6, -1,
    -- filter=58 channel=10
    14, 15, 0, 9, 15, 0, -4, -20, -6,
    -- filter=58 channel=11
    20, 17, 8, 1, 4, 3, -21, -7, 2,
    -- filter=58 channel=12
    -9, -1, -1, 2, -12, -11, 0, -13, 5,
    -- filter=58 channel=13
    9, 20, 0, -8, 0, -6, -6, -28, -4,
    -- filter=58 channel=14
    0, 7, 3, -3, 7, 2, 6, 6, 0,
    -- filter=58 channel=15
    14, 12, -7, 0, 4, 7, -19, -32, -5,
    -- filter=58 channel=16
    -14, -11, 0, 10, 14, 2, 0, 1, 7,
    -- filter=58 channel=17
    -5, 6, 3, -2, 1, 3, 3, 3, 0,
    -- filter=58 channel=18
    18, 26, 5, 0, -2, 4, -16, -37, -9,
    -- filter=58 channel=19
    7, -1, 2, -6, -5, 2, -4, 7, -2,
    -- filter=58 channel=20
    27, 24, 0, 6, 3, -1, -23, -19, -3,
    -- filter=58 channel=21
    -4, -2, -10, -2, 6, -1, 7, 8, 3,
    -- filter=58 channel=22
    7, -7, 0, 7, -1, 0, -5, -3, 2,
    -- filter=58 channel=23
    24, 4, -5, 17, 15, -3, -30, -33, -7,
    -- filter=58 channel=24
    2, -2, -6, -2, 3, -3, -3, 5, -1,
    -- filter=58 channel=25
    0, 7, 0, 2, 4, -9, -10, -9, -5,
    -- filter=58 channel=26
    -3, -5, -1, 0, -1, -3, 0, 9, 7,
    -- filter=58 channel=27
    15, 18, -6, 1, -8, 2, -20, -24, -2,
    -- filter=58 channel=28
    0, 1, -2, 0, 2, -5, 0, 0, -2,
    -- filter=58 channel=29
    29, 21, 12, -7, -10, 0, -17, -13, 1,
    -- filter=58 channel=30
    -6, 3, 0, -6, -10, -1, -3, 7, 0,
    -- filter=58 channel=31
    11, 7, -6, 15, 1, 5, -18, -13, -4,
    -- filter=58 channel=32
    11, 19, -4, 7, -4, -3, -8, -25, -6,
    -- filter=58 channel=33
    0, 6, 1, 10, 17, 3, 1, -22, -4,
    -- filter=58 channel=34
    -13, -8, -4, 0, -6, 0, -1, -1, 0,
    -- filter=58 channel=35
    0, 0, 4, -3, 0, -1, 0, 3, -4,
    -- filter=58 channel=36
    0, 11, 7, -8, -13, -1, -5, -5, 9,
    -- filter=58 channel=37
    -19, -23, -6, -9, -2, -3, 9, 20, 6,
    -- filter=58 channel=38
    0, 6, 1, 9, 9, 4, -4, -14, 2,
    -- filter=58 channel=39
    10, 14, 6, -2, 0, 7, -2, -13, 1,
    -- filter=58 channel=40
    -3, -2, 1, 5, 5, 5, -9, -13, -10,
    -- filter=58 channel=41
    -3, 0, 1, -26, -13, -11, 10, -12, -16,
    -- filter=58 channel=42
    3, -5, -6, 0, 5, 5, 0, 5, -2,
    -- filter=58 channel=43
    -3, 0, -6, 14, 16, -1, 1, -12, -6,
    -- filter=58 channel=44
    -18, -7, -12, 5, 2, -3, 6, 12, 7,
    -- filter=58 channel=45
    -8, -8, -9, 5, -7, -7, -1, 6, 4,
    -- filter=58 channel=46
    -4, 6, -5, -2, -5, 0, 9, -5, 2,
    -- filter=58 channel=47
    -23, -9, -14, 12, 16, 3, 0, 6, 3,
    -- filter=58 channel=48
    -6, 0, -8, -10, -11, -13, -15, -5, 4,
    -- filter=58 channel=49
    17, 10, -1, -5, -13, -1, -9, -7, 8,
    -- filter=58 channel=50
    0, 8, -1, -4, -1, -3, -10, 0, -8,
    -- filter=58 channel=51
    1, 2, 7, 0, -4, 0, -5, 0, 0,
    -- filter=58 channel=52
    11, 6, -4, 4, -10, 0, -9, 1, -3,
    -- filter=58 channel=53
    12, 16, -5, 1, 7, 5, -10, -10, 3,
    -- filter=58 channel=54
    4, 1, 2, -4, -1, -4, 1, 6, 0,
    -- filter=58 channel=55
    22, 28, 4, 5, 12, 0, -36, -43, -7,
    -- filter=58 channel=56
    5, -1, 0, 2, -4, -1, -5, 4, -3,
    -- filter=58 channel=57
    -9, 5, 5, -8, -11, 4, 4, -5, -6,
    -- filter=58 channel=58
    0, -5, -7, -1, 13, 9, 5, 12, 11,
    -- filter=58 channel=59
    4, 9, 6, -2, 6, -2, -3, -8, -12,
    -- filter=58 channel=60
    -4, 4, 6, 6, 4, -4, -3, 4, 2,
    -- filter=58 channel=61
    5, 8, 1, -8, -5, 6, -5, 0, 5,
    -- filter=58 channel=62
    3, 8, 2, 9, 8, 3, -4, -8, -6,
    -- filter=58 channel=63
    -13, -7, -8, -2, 10, 9, 2, 7, 3,
    -- filter=58 channel=64
    6, 3, 0, -5, 2, -1, -4, -6, 2,
    -- filter=58 channel=65
    0, 3, 0, 3, 1, 0, -4, 2, 2,
    -- filter=58 channel=66
    -7, 5, 7, -2, -1, -3, 6, -10, 1,
    -- filter=58 channel=67
    2, 3, -9, 3, -5, 6, 2, -6, 2,
    -- filter=58 channel=68
    -6, 5, -9, -7, -2, -5, 2, 4, 5,
    -- filter=58 channel=69
    -10, 1, -7, -2, -1, -2, 8, 2, 7,
    -- filter=58 channel=70
    12, -1, 0, 5, -3, -9, -14, -9, -6,
    -- filter=58 channel=71
    0, 1, -3, 2, 13, 5, 5, -7, -7,
    -- filter=58 channel=72
    6, 18, -1, 5, 4, 7, -13, -17, -4,
    -- filter=58 channel=73
    14, 24, -3, -3, -15, -4, -18, -17, 3,
    -- filter=58 channel=74
    3, -9, -11, 4, -16, -5, -2, -4, 3,
    -- filter=58 channel=75
    -18, 0, -4, 9, 24, -6, 12, -3, -4,
    -- filter=58 channel=76
    11, 14, 6, 5, -4, 1, -14, -27, -12,
    -- filter=58 channel=77
    -7, 0, 3, 5, 1, 6, 0, 0, -7,
    -- filter=58 channel=78
    -4, -2, -3, 10, 6, 10, 0, 1, 11,
    -- filter=58 channel=79
    18, 23, 4, 14, 5, -8, -20, -43, 0,
    -- filter=58 channel=80
    -7, 9, 1, 0, 14, -5, -17, -9, 4,
    -- filter=58 channel=81
    5, 0, -3, 4, 5, -3, 6, -2, 5,
    -- filter=58 channel=82
    -3, -7, -4, 3, 9, 5, -3, 4, 0,
    -- filter=58 channel=83
    -1, 9, -9, -14, -3, -7, -2, 0, 0,
    -- filter=58 channel=84
    15, 14, 4, -9, -13, 3, -3, -9, 9,
    -- filter=58 channel=85
    0, 0, 3, 6, 0, 3, -1, -1, -3,
    -- filter=58 channel=86
    -1, -12, 0, 0, -1, 0, 1, -4, 9,
    -- filter=58 channel=87
    16, 13, 0, -4, 4, -2, -13, -1, -6,
    -- filter=58 channel=88
    2, 4, -3, -2, -15, -6, 4, 3, -1,
    -- filter=58 channel=89
    18, 29, 6, 15, 4, 2, -23, -41, -8,
    -- filter=58 channel=90
    4, 0, -7, 3, 2, 1, -7, -5, 4,
    -- filter=58 channel=91
    19, 19, -11, -5, -16, 7, -21, -20, -2,
    -- filter=58 channel=92
    -4, 2, -8, 3, 1, -5, -7, -1, 3,
    -- filter=58 channel=93
    -21, -7, -18, 0, -8, 0, -2, 8, 10,
    -- filter=58 channel=94
    4, 6, -4, 1, 3, 0, 2, 4, 0,
    -- filter=58 channel=95
    6, 5, 3, -1, -1, -8, 1, -7, 2,
    -- filter=58 channel=96
    -4, -3, -7, -4, 1, -5, -4, -3, 3,
    -- filter=58 channel=97
    4, 2, 3, 8, 21, -1, 5, 1, -4,
    -- filter=58 channel=98
    0, 16, -4, 8, 14, 3, -12, -19, 3,
    -- filter=58 channel=99
    16, 25, 1, 8, 0, 6, -19, -16, 4,
    -- filter=58 channel=100
    -4, -5, -4, 0, -7, 0, -1, 4, 2,
    -- filter=58 channel=101
    7, 18, -4, 7, 7, -2, 1, 6, 1,
    -- filter=58 channel=102
    5, 6, 5, -4, -2, 1, -5, -4, -4,
    -- filter=58 channel=103
    -8, -13, 0, 17, 19, 2, -1, 5, -1,
    -- filter=58 channel=104
    0, 9, 3, 2, -5, -3, -3, -10, 5,
    -- filter=58 channel=105
    10, 11, 3, 0, 0, 4, -5, -20, 3,
    -- filter=58 channel=106
    0, 4, -4, -3, 0, -3, -3, -5, 3,
    -- filter=58 channel=107
    12, 8, -9, 9, 0, 4, -8, -21, -1,
    -- filter=58 channel=108
    0, 4, -3, -2, 1, 3, 2, -4, 4,
    -- filter=58 channel=109
    16, 30, 4, 5, -13, 1, -22, -16, 7,
    -- filter=58 channel=110
    6, 2, -1, 7, 13, 0, -4, -10, 3,
    -- filter=58 channel=111
    6, 0, 0, -5, 4, -1, -1, -3, -1,
    -- filter=58 channel=112
    4, -5, -11, 6, 1, -5, -3, 0, -3,
    -- filter=58 channel=113
    -5, 1, -6, 12, 21, -6, -8, -19, 1,
    -- filter=58 channel=114
    10, 21, -1, 0, -2, -8, -15, -14, 5,
    -- filter=58 channel=115
    0, -6, -6, -1, 4, 4, -4, 0, 1,
    -- filter=58 channel=116
    10, 30, -2, -7, -11, -5, -16, -20, -5,
    -- filter=58 channel=117
    5, 0, -3, -7, -3, -1, 0, -6, 1,
    -- filter=58 channel=118
    3, -4, 0, 3, -2, 5, 0, -4, 3,
    -- filter=58 channel=119
    4, -2, -6, -7, -15, -3, -4, 3, -4,
    -- filter=58 channel=120
    22, 26, -7, 0, -22, 4, -23, -20, 0,
    -- filter=58 channel=121
    8, 0, 9, 7, 14, 3, -1, -7, -1,
    -- filter=58 channel=122
    -22, -21, -20, 7, 13, 4, 5, 23, 12,
    -- filter=58 channel=123
    1, -8, 2, 2, 8, -6, -1, 4, -2,
    -- filter=58 channel=124
    3, 0, 0, -2, 1, 0, 0, -13, -1,
    -- filter=58 channel=125
    12, 17, 2, 5, -3, -4, -8, -18, 7,
    -- filter=58 channel=126
    3, 2, -4, 18, 19, 8, -6, -12, -10,
    -- filter=58 channel=127
    -1, 6, 0, -4, 2, 0, 1, -5, -3,
    -- filter=59 channel=0
    -2, -4, -6, 2, 0, 0, 13, 0, 1,
    -- filter=59 channel=1
    7, -6, 5, 0, -8, -3, 2, -6, 9,
    -- filter=59 channel=2
    -5, -2, 5, -5, 0, -3, -9, 0, -3,
    -- filter=59 channel=3
    0, -8, -4, 3, 0, 0, 8, -7, -9,
    -- filter=59 channel=4
    3, -14, -7, -1, -7, -8, -7, -15, -9,
    -- filter=59 channel=5
    -2, -6, 13, -7, -11, 10, -14, 0, 18,
    -- filter=59 channel=6
    -1, 0, -5, 7, -6, -6, -5, 3, -15,
    -- filter=59 channel=7
    -6, -5, -6, -6, -3, -2, 2, -1, 7,
    -- filter=59 channel=8
    -6, 0, -4, 2, 2, -7, 4, -5, -1,
    -- filter=59 channel=9
    -1, -1, 3, 0, -3, 2, -3, 0, 5,
    -- filter=59 channel=10
    -4, 2, 0, -1, -8, 0, -1, -15, 4,
    -- filter=59 channel=11
    0, -1, -4, 4, 0, -12, -2, -2, -7,
    -- filter=59 channel=12
    -2, -1, 0, 3, -3, -9, 13, -2, -7,
    -- filter=59 channel=13
    14, -7, -8, 9, 5, -6, 2, 0, -10,
    -- filter=59 channel=14
    7, 6, 3, -3, -6, 0, 6, 0, 1,
    -- filter=59 channel=15
    3, -4, -14, 15, 7, -11, 6, 8, -12,
    -- filter=59 channel=16
    1, -3, 7, -1, -1, 6, -7, -14, 5,
    -- filter=59 channel=17
    2, 2, 2, -6, 6, -1, -5, 3, -3,
    -- filter=59 channel=18
    11, 7, -17, 16, 1, -13, 9, 7, -21,
    -- filter=59 channel=19
    -7, 0, 3, 2, 0, 7, 0, 5, 6,
    -- filter=59 channel=20
    -10, -8, -21, 3, 3, -14, -6, 2, -13,
    -- filter=59 channel=21
    -9, -9, 18, -1, -5, 26, -6, -16, 19,
    -- filter=59 channel=22
    -1, -6, 0, 6, 4, -10, 5, -1, -1,
    -- filter=59 channel=23
    -2, -9, 0, 13, 4, 0, 1, -10, -5,
    -- filter=59 channel=24
    -1, -2, 6, 0, 2, 1, 3, 2, 6,
    -- filter=59 channel=25
    -1, -10, 6, 10, 0, 7, -2, -3, 12,
    -- filter=59 channel=26
    -8, -1, 5, -9, -6, 4, -5, -6, 5,
    -- filter=59 channel=27
    1, 0, 9, 7, 6, 9, 6, -9, 12,
    -- filter=59 channel=28
    -5, 4, -5, 1, 6, -1, 2, 2, -5,
    -- filter=59 channel=29
    -9, 0, -19, 5, 13, -8, 1, -1, -20,
    -- filter=59 channel=30
    0, 3, -3, 1, -1, 1, 1, 0, 12,
    -- filter=59 channel=31
    -1, 1, 29, -3, -2, 34, -20, -20, 16,
    -- filter=59 channel=32
    1, -2, -2, 11, 0, -4, 3, -7, -17,
    -- filter=59 channel=33
    3, -4, 5, 4, 5, 4, 3, 1, 5,
    -- filter=59 channel=34
    3, -7, 0, -5, -6, 0, 4, -6, 4,
    -- filter=59 channel=35
    0, -6, 1, 6, 4, -2, -1, 7, -4,
    -- filter=59 channel=36
    -8, 0, 6, -11, 0, 9, -3, -6, -6,
    -- filter=59 channel=37
    0, -10, 3, 0, -18, 4, -9, -6, 6,
    -- filter=59 channel=38
    0, -3, -4, 9, 3, 1, -3, -5, 9,
    -- filter=59 channel=39
    -2, 3, -1, -1, 3, 0, 0, 0, -13,
    -- filter=59 channel=40
    -1, 3, 0, -4, -4, 1, 0, -3, -2,
    -- filter=59 channel=41
    7, -11, -17, 8, -3, -5, 7, -7, -13,
    -- filter=59 channel=42
    2, -1, 0, -2, 1, 7, -2, 5, 0,
    -- filter=59 channel=43
    0, -5, -9, 13, -2, -5, 0, 0, -12,
    -- filter=59 channel=44
    5, 2, 17, -8, -6, 21, -11, -11, 14,
    -- filter=59 channel=45
    6, -5, -4, 4, 2, 0, 1, 3, -7,
    -- filter=59 channel=46
    -2, 3, -2, -2, 6, -3, 0, 7, 1,
    -- filter=59 channel=47
    -12, 2, 21, -2, -3, 19, -9, -16, 18,
    -- filter=59 channel=48
    -7, 5, 15, -4, 0, 23, -6, -15, 7,
    -- filter=59 channel=49
    5, 1, -11, 10, -3, -15, 9, -4, -16,
    -- filter=59 channel=50
    -6, 5, 3, 2, 3, 9, -6, 5, 10,
    -- filter=59 channel=51
    1, -3, 6, 0, 3, 4, -6, 4, -7,
    -- filter=59 channel=52
    7, -8, -4, -1, -5, -7, -4, -3, 0,
    -- filter=59 channel=53
    -5, -6, -7, 0, -6, -4, -4, 2, 0,
    -- filter=59 channel=54
    1, 7, -3, -6, 0, 0, -6, 1, 3,
    -- filter=59 channel=55
    7, -2, -11, 6, 4, -10, 3, -7, -15,
    -- filter=59 channel=56
    -7, 0, 3, -3, 2, 7, 2, -7, 3,
    -- filter=59 channel=57
    5, -8, -6, 1, 0, -3, -1, 0, -3,
    -- filter=59 channel=58
    -8, -1, 9, -7, -5, 2, -13, 4, 8,
    -- filter=59 channel=59
    -2, -8, 14, 7, -9, 9, 5, -16, 8,
    -- filter=59 channel=60
    -4, -7, -1, -5, -7, -4, 3, -1, 1,
    -- filter=59 channel=61
    5, -1, 0, -8, -1, 0, -2, -5, 6,
    -- filter=59 channel=62
    -4, 2, 0, 5, -7, 0, -4, -2, -5,
    -- filter=59 channel=63
    -14, -10, 2, -8, 0, 6, -7, -9, 3,
    -- filter=59 channel=64
    -9, 0, -2, -1, 1, 1, -6, -4, 2,
    -- filter=59 channel=65
    -6, 7, 6, -3, 0, 0, -4, 6, -7,
    -- filter=59 channel=66
    0, -3, 4, 7, -3, -1, 15, 0, -4,
    -- filter=59 channel=67
    -7, 1, 1, 0, 0, -5, 6, 9, 2,
    -- filter=59 channel=68
    -2, 3, 3, -4, 1, -10, 0, -4, -3,
    -- filter=59 channel=69
    5, 4, 5, 5, -5, 0, -1, -8, -7,
    -- filter=59 channel=70
    10, -3, 8, 9, -4, -3, 5, 0, -1,
    -- filter=59 channel=71
    -2, 2, 4, 0, -2, 0, 5, -2, 3,
    -- filter=59 channel=72
    -9, 1, 16, 0, 0, 18, -4, -13, 1,
    -- filter=59 channel=73
    -1, -3, -3, 3, 0, -12, -1, -6, -3,
    -- filter=59 channel=74
    1, 2, 10, -7, 2, 11, -5, -3, 14,
    -- filter=59 channel=75
    -5, 0, 9, 7, -11, -6, 9, -8, 10,
    -- filter=59 channel=76
    -8, -9, -18, 4, 0, -17, 7, 0, -17,
    -- filter=59 channel=77
    1, -1, 0, 5, 0, 3, 6, 3, -3,
    -- filter=59 channel=78
    -6, 1, 0, -11, -6, 0, -1, -4, 8,
    -- filter=59 channel=79
    13, 0, -16, 22, 1, -14, 11, -4, -12,
    -- filter=59 channel=80
    -4, 4, 19, -8, -9, 24, -2, -25, 19,
    -- filter=59 channel=81
    -5, 2, -6, 1, -6, -4, -2, -7, 0,
    -- filter=59 channel=82
    -1, -3, 7, -4, 0, 2, -3, 0, 6,
    -- filter=59 channel=83
    2, 5, 9, -5, 5, 4, -5, -8, 4,
    -- filter=59 channel=84
    4, -5, -10, 11, -3, -2, -5, -8, -16,
    -- filter=59 channel=85
    6, -1, 5, 5, -1, -5, -4, -3, -1,
    -- filter=59 channel=86
    1, -8, 0, -4, -4, 1, -1, -3, 5,
    -- filter=59 channel=87
    -6, -6, -16, 4, -5, -6, -3, -6, -13,
    -- filter=59 channel=88
    -9, -6, 4, -4, 0, 9, -14, -9, 4,
    -- filter=59 channel=89
    7, -10, 0, 12, 3, -3, 12, -2, 0,
    -- filter=59 channel=90
    -10, 2, 0, -2, -11, 11, -13, -6, -1,
    -- filter=59 channel=91
    -2, -5, 1, 0, -3, -4, 3, 0, 0,
    -- filter=59 channel=92
    -2, 4, 9, 6, -2, 6, -8, 1, 0,
    -- filter=59 channel=93
    -2, -10, 10, -10, -16, 16, -15, -14, 12,
    -- filter=59 channel=94
    -6, 0, 6, 0, 2, 2, 2, 3, 7,
    -- filter=59 channel=95
    2, 4, -4, 0, -3, -3, -6, 0, -8,
    -- filter=59 channel=96
    -2, -4, -8, 4, 1, 3, -4, 4, 2,
    -- filter=59 channel=97
    0, 5, -3, 0, -3, 8, 2, -2, 9,
    -- filter=59 channel=98
    5, -5, 11, 0, -2, 13, -7, -17, 8,
    -- filter=59 channel=99
    -6, -5, 7, -13, -11, 6, -8, -10, 3,
    -- filter=59 channel=100
    0, 3, 3, -8, 2, 2, -8, -4, -1,
    -- filter=59 channel=101
    -5, -2, -5, 6, -9, -10, -6, -11, -4,
    -- filter=59 channel=102
    -3, 6, -7, 4, -2, 5, 4, 6, -5,
    -- filter=59 channel=103
    1, 5, 30, -8, 0, 25, -14, -9, 22,
    -- filter=59 channel=104
    -10, 0, 23, -8, -2, 25, -16, -20, 10,
    -- filter=59 channel=105
    -11, -8, -3, 6, 5, -2, 4, -1, -5,
    -- filter=59 channel=106
    -1, -6, -12, 0, 6, -11, -7, 5, -10,
    -- filter=59 channel=107
    5, 0, -17, 3, -2, -20, 12, 7, -10,
    -- filter=59 channel=108
    3, -9, -12, -9, -2, -9, -2, 0, -6,
    -- filter=59 channel=109
    0, -8, 5, 3, 0, -1, -8, -10, -6,
    -- filter=59 channel=110
    2, 4, -1, -4, 1, 6, -11, -15, -5,
    -- filter=59 channel=111
    2, -4, 0, 0, 5, -1, 0, -2, -4,
    -- filter=59 channel=112
    0, 5, 8, -2, -1, 10, -6, -7, 12,
    -- filter=59 channel=113
    -6, -7, 7, 0, 1, 9, -7, -4, 5,
    -- filter=59 channel=114
    1, 2, -13, 13, 8, -13, 17, -1, -13,
    -- filter=59 channel=115
    3, -5, 4, -2, 3, 2, 5, -2, -1,
    -- filter=59 channel=116
    -7, -4, 3, 9, -3, -3, -9, -3, -11,
    -- filter=59 channel=117
    1, -3, -7, 0, 1, -3, 0, -6, 3,
    -- filter=59 channel=118
    1, 5, -7, -7, -3, -5, 2, 6, 1,
    -- filter=59 channel=119
    3, 0, 2, -7, -5, 13, -9, -1, 3,
    -- filter=59 channel=120
    6, -11, 0, 10, -7, 5, 5, -7, -3,
    -- filter=59 channel=121
    0, -3, -5, 8, 0, 1, 6, -8, -3,
    -- filter=59 channel=122
    -10, 2, 29, -19, -17, 45, -27, -20, 34,
    -- filter=59 channel=123
    -7, 4, 8, -4, 6, 7, -4, 0, 9,
    -- filter=59 channel=124
    4, 0, -9, 6, 5, -11, 6, 3, -11,
    -- filter=59 channel=125
    -1, 1, 8, 1, -6, 7, -12, -15, 1,
    -- filter=59 channel=126
    0, 6, -10, 8, -6, -5, 11, -2, -9,
    -- filter=59 channel=127
    7, -2, 4, -3, 0, -8, -4, 0, -7,
    -- filter=60 channel=0
    -6, -2, 3, -3, 0, 2, -4, 0, 0,
    -- filter=60 channel=1
    0, 0, -1, 6, -9, -7, -2, -13, -2,
    -- filter=60 channel=2
    2, 1, 0, -6, -1, 0, 2, 1, -8,
    -- filter=60 channel=3
    -2, -2, 2, 0, -5, 4, -7, 0, -1,
    -- filter=60 channel=4
    0, -6, 8, 0, -12, -3, -2, -6, -1,
    -- filter=60 channel=5
    -1, 2, -4, 10, 5, 3, -1, 9, -1,
    -- filter=60 channel=6
    -7, -1, 6, -5, 5, 11, -3, 2, -2,
    -- filter=60 channel=7
    7, 3, 5, -1, 4, -6, 0, 1, -7,
    -- filter=60 channel=8
    -4, -4, 7, -12, -5, 8, -1, -4, -6,
    -- filter=60 channel=9
    8, 4, 3, -2, 4, -2, 2, -2, 2,
    -- filter=60 channel=10
    -3, 8, 8, -3, -4, -4, -4, -2, -2,
    -- filter=60 channel=11
    -10, -6, 1, -5, 7, 4, -5, -5, 3,
    -- filter=60 channel=12
    0, 0, 2, -8, 5, -6, -11, -8, 6,
    -- filter=60 channel=13
    -14, -6, 4, 3, 3, 5, -2, -9, -9,
    -- filter=60 channel=14
    -3, 5, 3, 1, 3, 2, 1, -6, 5,
    -- filter=60 channel=15
    -11, 4, 10, -2, 8, 17, -16, -7, -2,
    -- filter=60 channel=16
    1, -1, -1, 7, 3, -5, 2, 11, 0,
    -- filter=60 channel=17
    -3, -6, -6, -6, 0, -6, 4, 6, -3,
    -- filter=60 channel=18
    -6, 13, 17, -7, 8, 28, -13, -8, 3,
    -- filter=60 channel=19
    -5, -2, 5, -2, -2, -1, 0, 0, 0,
    -- filter=60 channel=20
    -16, -4, 5, -17, 8, 5, -9, 1, 1,
    -- filter=60 channel=21
    9, -10, -12, 1, -9, -6, 17, 2, -7,
    -- filter=60 channel=22
    1, 8, 0, -5, 9, 14, -8, -1, -4,
    -- filter=60 channel=23
    -16, 5, 13, -4, 2, 21, -6, -5, 2,
    -- filter=60 channel=24
    6, -4, 0, 2, -3, -1, -3, 7, 0,
    -- filter=60 channel=25
    -11, -5, -2, 0, 3, 7, -6, -3, -10,
    -- filter=60 channel=26
    -2, 3, 1, 7, 0, -7, 4, 4, 6,
    -- filter=60 channel=27
    1, 0, 9, 1, 3, 20, -13, -3, -8,
    -- filter=60 channel=28
    -3, 6, 2, 1, 0, -2, 4, 6, 4,
    -- filter=60 channel=29
    0, 1, 3, -7, 12, 9, -8, -5, 4,
    -- filter=60 channel=30
    0, 6, -1, -3, 1, 10, 5, 1, -11,
    -- filter=60 channel=31
    -4, -6, -5, 1, -1, 4, 13, 11, -6,
    -- filter=60 channel=32
    -5, 7, 8, -10, 5, 12, -13, -15, 2,
    -- filter=60 channel=33
    0, 7, 1, 10, 8, 10, -11, -7, -6,
    -- filter=60 channel=34
    -5, -1, 11, -5, 3, 3, -10, 6, 13,
    -- filter=60 channel=35
    6, 2, -6, 0, -4, 2, 6, 3, -4,
    -- filter=60 channel=36
    2, -11, -6, 1, -7, -9, -1, -7, 0,
    -- filter=60 channel=37
    11, 0, 5, 0, -2, -3, 5, -5, 5,
    -- filter=60 channel=38
    2, -2, -2, 10, -3, 8, -5, 7, 4,
    -- filter=60 channel=39
    0, -3, 5, -8, 3, 6, -8, -8, -4,
    -- filter=60 channel=40
    -11, 3, 0, -8, -4, 9, -4, -8, -4,
    -- filter=60 channel=41
    -20, 6, 5, -15, 0, -1, -19, -7, 8,
    -- filter=60 channel=42
    3, 5, 0, -1, 0, 6, 3, -3, 3,
    -- filter=60 channel=43
    -15, 8, 8, -7, 6, 12, -7, 2, -3,
    -- filter=60 channel=44
    3, -6, 0, 0, -6, 2, 2, 1, 6,
    -- filter=60 channel=45
    0, -2, 4, -1, 0, 0, -3, 3, 0,
    -- filter=60 channel=46
    4, -4, 0, 1, 0, -1, -5, -7, 1,
    -- filter=60 channel=47
    11, 2, -9, 4, -8, 1, 4, 14, -3,
    -- filter=60 channel=48
    6, -3, 6, 8, -7, 3, -6, -7, -10,
    -- filter=60 channel=49
    0, 2, 5, -5, 0, 3, -3, -5, -1,
    -- filter=60 channel=50
    7, -4, -3, 1, -5, 3, 0, -6, -4,
    -- filter=60 channel=51
    2, 0, -1, -6, 2, -4, 6, -1, 2,
    -- filter=60 channel=52
    -8, -7, 8, 0, -2, 4, -10, 2, 5,
    -- filter=60 channel=53
    2, -3, -3, -4, 8, 6, -7, 1, 2,
    -- filter=60 channel=54
    7, -4, -5, 0, -2, 4, 3, 1, 0,
    -- filter=60 channel=55
    -14, 9, 8, -4, 14, 11, -5, -5, 0,
    -- filter=60 channel=56
    0, -3, 7, -12, -1, 2, -5, 2, 9,
    -- filter=60 channel=57
    -4, -2, 2, 5, 4, -1, -9, 3, -3,
    -- filter=60 channel=58
    4, 0, 3, -4, -6, -7, -4, 0, 6,
    -- filter=60 channel=59
    5, -4, 0, 7, -6, 5, 2, 1, 0,
    -- filter=60 channel=60
    1, 0, 5, 1, 6, -4, 3, 1, 3,
    -- filter=60 channel=61
    -2, 0, 0, -5, -2, 2, -6, -3, -1,
    -- filter=60 channel=62
    4, 0, -1, -4, -1, -3, -1, 0, 6,
    -- filter=60 channel=63
    5, 4, -2, 1, -2, -2, -1, 0, 1,
    -- filter=60 channel=64
    4, -1, -6, -4, -2, -1, 2, 3, -6,
    -- filter=60 channel=65
    5, 5, -7, 5, -2, -6, 6, 4, -6,
    -- filter=60 channel=66
    -7, -3, 4, -3, -4, 3, -10, -5, -2,
    -- filter=60 channel=67
    2, -2, -4, 5, 3, -7, 0, -8, 0,
    -- filter=60 channel=68
    -3, -4, 2, -9, -3, -4, -7, 4, -8,
    -- filter=60 channel=69
    -3, -5, 4, -8, -1, -2, -6, -1, 4,
    -- filter=60 channel=70
    0, -3, 4, 1, 5, 13, -2, -12, 8,
    -- filter=60 channel=71
    5, -4, -6, 3, 0, 3, 2, -5, 0,
    -- filter=60 channel=72
    -1, 0, -2, -5, -6, -2, 6, -4, -6,
    -- filter=60 channel=73
    2, 0, 6, -11, 7, 11, -13, -3, -7,
    -- filter=60 channel=74
    -6, 4, 0, -9, -3, 14, -8, -7, 9,
    -- filter=60 channel=75
    0, -2, 0, 6, -5, 4, 0, -5, 11,
    -- filter=60 channel=76
    -15, 3, 1, 1, 11, 4, 0, -8, -4,
    -- filter=60 channel=77
    -4, -1, 4, -5, -1, -8, 6, 0, 4,
    -- filter=60 channel=78
    0, -6, -2, 4, 8, -1, -2, 4, 5,
    -- filter=60 channel=79
    -17, 3, 13, 0, 12, 22, -20, -16, -5,
    -- filter=60 channel=80
    0, 2, 0, 12, -11, -11, 8, 2, -4,
    -- filter=60 channel=81
    7, -7, 3, -6, 7, -4, -5, 5, -5,
    -- filter=60 channel=82
    7, 2, 0, -6, 7, 8, 2, -4, -3,
    -- filter=60 channel=83
    0, 1, 0, 7, -5, -2, 5, -5, 0,
    -- filter=60 channel=84
    -7, 5, 12, -12, 4, 15, -3, -5, 2,
    -- filter=60 channel=85
    0, 3, -4, -2, 1, -4, 0, 4, -7,
    -- filter=60 channel=86
    1, -1, 2, 4, -5, -2, -8, -3, 0,
    -- filter=60 channel=87
    -5, 2, -6, -15, -6, 11, -7, -11, -5,
    -- filter=60 channel=88
    -4, 1, -1, 2, 1, -10, 9, 3, -10,
    -- filter=60 channel=89
    -14, 3, 5, 3, -2, 12, 1, -10, -9,
    -- filter=60 channel=90
    -8, 5, -8, 1, -7, -2, 2, 8, 5,
    -- filter=60 channel=91
    -7, 0, 11, 1, 9, 7, -10, -10, 1,
    -- filter=60 channel=92
    -3, 1, 0, -4, 2, 12, -2, -6, 4,
    -- filter=60 channel=93
    6, 0, -5, -1, -3, -8, 2, -6, -8,
    -- filter=60 channel=94
    -4, 0, -7, -5, -2, 3, -5, 6, -1,
    -- filter=60 channel=95
    6, 6, 3, 6, -6, -3, -6, -5, -5,
    -- filter=60 channel=96
    0, 6, -6, -7, -6, -1, 6, -6, -4,
    -- filter=60 channel=97
    -1, 1, 1, 3, 5, -6, -1, 0, 8,
    -- filter=60 channel=98
    4, 4, 0, -1, -5, 10, -8, 0, -8,
    -- filter=60 channel=99
    -1, 6, 7, -3, 1, 11, -1, 5, -5,
    -- filter=60 channel=100
    -4, -1, -2, -11, 7, 5, 2, -4, 0,
    -- filter=60 channel=101
    -4, 0, 8, -3, -10, -6, -9, -2, 1,
    -- filter=60 channel=102
    0, 0, 0, 4, 6, -4, 0, 0, -5,
    -- filter=60 channel=103
    8, -1, -7, 15, -3, -12, 12, 15, 9,
    -- filter=60 channel=104
    6, 4, -6, 5, -9, 1, 7, 4, 0,
    -- filter=60 channel=105
    -11, -2, -4, -9, 6, 5, -3, 0, 7,
    -- filter=60 channel=106
    3, -6, -7, -9, 2, -7, 2, -6, -4,
    -- filter=60 channel=107
    -12, 8, 8, -14, -1, 9, -14, 0, 2,
    -- filter=60 channel=108
    -4, -2, 0, -5, -2, -2, 1, -7, -4,
    -- filter=60 channel=109
    0, 9, 5, -8, 3, 23, -15, -13, 1,
    -- filter=60 channel=110
    -1, -7, -5, -3, 3, 0, 2, 4, -3,
    -- filter=60 channel=111
    4, 4, 0, -3, 0, 0, 0, -5, -1,
    -- filter=60 channel=112
    -1, -4, -1, 8, 8, 3, -5, -8, -4,
    -- filter=60 channel=113
    4, -2, -3, -1, 8, 7, 1, 3, 4,
    -- filter=60 channel=114
    -14, -1, 14, -1, 13, 19, -12, -16, -2,
    -- filter=60 channel=115
    -6, -5, -1, 3, 4, -4, -2, -5, 0,
    -- filter=60 channel=116
    -9, 5, 2, 1, 0, 5, -3, -7, -15,
    -- filter=60 channel=117
    0, -4, -9, 0, 4, -3, -6, 1, 1,
    -- filter=60 channel=118
    -7, 0, -4, -5, -1, -1, 1, -6, -1,
    -- filter=60 channel=119
    -11, 1, 0, -10, -2, 11, -14, -5, 14,
    -- filter=60 channel=120
    -7, -3, 7, 0, 12, 21, -10, -7, 0,
    -- filter=60 channel=121
    -4, 5, -5, 4, -9, 2, -10, -3, 7,
    -- filter=60 channel=122
    6, -9, -10, 11, -3, -15, 15, 6, 0,
    -- filter=60 channel=123
    -7, 0, 8, -2, 5, -2, -3, -5, 3,
    -- filter=60 channel=124
    -8, 5, 6, 0, 8, 0, -10, 3, -2,
    -- filter=60 channel=125
    0, -5, 2, 6, -5, 8, 1, -5, -11,
    -- filter=60 channel=126
    -5, 0, 6, 1, -4, -4, 0, -1, -6,
    -- filter=60 channel=127
    -3, -2, 5, -7, -5, 0, -6, 3, -3,
    -- filter=61 channel=0
    -9, -5, 0, -1, -5, -6, 8, 2, 10,
    -- filter=61 channel=1
    3, 0, 8, -10, -9, 6, 10, -4, 5,
    -- filter=61 channel=2
    4, 0, -5, 7, 2, -6, -9, 0, -1,
    -- filter=61 channel=3
    -7, -8, -3, -6, -2, -7, -5, 1, 3,
    -- filter=61 channel=4
    1, 1, -6, 4, -10, -13, -11, -12, 0,
    -- filter=61 channel=5
    -10, -11, 0, -7, -5, -5, -2, -6, 2,
    -- filter=61 channel=6
    -3, 2, 1, 7, 4, 0, 2, -1, 0,
    -- filter=61 channel=7
    -6, 3, 4, -5, -1, 3, -2, -4, 2,
    -- filter=61 channel=8
    2, -3, 0, 6, 0, 6, -2, -4, 6,
    -- filter=61 channel=9
    -5, -7, 7, -1, 5, -6, 2, -1, -7,
    -- filter=61 channel=10
    4, -7, -4, 0, 14, 7, -5, -3, -4,
    -- filter=61 channel=11
    0, -1, 0, 3, 13, -5, -6, 2, -3,
    -- filter=61 channel=12
    6, -1, 1, -3, 9, -4, 2, -7, 6,
    -- filter=61 channel=13
    -2, 6, 2, -4, 11, 6, -2, 0, -5,
    -- filter=61 channel=14
    -7, 6, 1, 6, -4, -5, -1, -6, -5,
    -- filter=61 channel=15
    -13, -8, -5, 5, 14, 0, -5, 2, -10,
    -- filter=61 channel=16
    4, -3, -3, 0, 2, 3, 3, 0, 6,
    -- filter=61 channel=17
    -2, 1, -4, 5, 3, -7, 5, -6, 7,
    -- filter=61 channel=18
    -15, 5, -3, -11, 18, 3, 4, 5, -8,
    -- filter=61 channel=19
    6, -2, -6, 4, 5, 7, 4, -6, 0,
    -- filter=61 channel=20
    -13, -2, -14, 4, 16, -10, 0, -6, -13,
    -- filter=61 channel=21
    1, -6, 0, -1, -2, 7, -6, 1, -2,
    -- filter=61 channel=22
    0, -5, -1, 0, 0, 0, 1, -2, -4,
    -- filter=61 channel=23
    -12, 5, 0, 8, 11, 0, 3, -9, -13,
    -- filter=61 channel=24
    4, 5, -2, 1, 0, 5, -6, -3, -1,
    -- filter=61 channel=25
    -7, 0, 11, 0, 3, -1, 5, 0, -1,
    -- filter=61 channel=26
    1, 4, 6, -6, -2, -1, -5, -1, -5,
    -- filter=61 channel=27
    -11, 4, 9, 2, 16, 7, 2, -10, -13,
    -- filter=61 channel=28
    -4, -1, -6, 6, 7, -2, 4, 7, 1,
    -- filter=61 channel=29
    -8, 1, -2, 3, 17, 3, -7, -8, -2,
    -- filter=61 channel=30
    -10, -4, 4, -5, -2, 1, 8, -4, -10,
    -- filter=61 channel=31
    4, 3, 15, 3, 0, 1, 6, -3, -19,
    -- filter=61 channel=32
    -10, 7, 0, -13, 3, -2, -5, 2, 0,
    -- filter=61 channel=33
    -7, -7, 9, -2, 9, 5, 0, 8, 2,
    -- filter=61 channel=34
    0, 0, 9, 0, -8, 2, 1, -11, 3,
    -- filter=61 channel=35
    -5, 0, 4, -6, -4, 3, 0, 2, 2,
    -- filter=61 channel=36
    3, 0, -1, 4, 4, 2, -2, -5, -14,
    -- filter=61 channel=37
    0, -7, 11, 3, -4, -5, 5, -7, 2,
    -- filter=61 channel=38
    -4, 2, -3, -1, 7, -2, 6, -6, -8,
    -- filter=61 channel=39
    -4, -3, 1, 6, 10, -5, 0, 4, -8,
    -- filter=61 channel=40
    -7, 2, -9, 2, 3, 2, 1, -5, 4,
    -- filter=61 channel=41
    1, 3, -1, -2, 0, 7, -9, -8, 14,
    -- filter=61 channel=42
    -4, -5, -1, -4, -7, -2, 0, 6, -9,
    -- filter=61 channel=43
    -2, 1, -5, -2, 5, -6, -5, -4, -5,
    -- filter=61 channel=44
    0, 0, 2, -7, -10, -4, 0, -4, 0,
    -- filter=61 channel=45
    -8, -3, -6, -6, 3, -1, -7, 1, 1,
    -- filter=61 channel=46
    5, 3, 0, 4, -6, -7, 5, 5, 5,
    -- filter=61 channel=47
    -7, 1, 3, 0, -10, -1, 5, 1, -3,
    -- filter=61 channel=48
    -7, 2, 10, 1, 0, 3, 9, -6, -15,
    -- filter=61 channel=49
    -9, 1, 2, 3, -3, -8, 1, -6, 0,
    -- filter=61 channel=50
    -7, -4, 3, -5, -1, 2, 1, 4, -3,
    -- filter=61 channel=51
    -1, -6, -4, -4, 2, 4, 5, 4, -2,
    -- filter=61 channel=52
    4, -3, 0, -3, -5, -5, -6, 2, -5,
    -- filter=61 channel=53
    -8, 0, 4, 5, 9, -3, -6, -2, 0,
    -- filter=61 channel=54
    -4, -3, 2, -7, -1, 1, -3, -6, 1,
    -- filter=61 channel=55
    -2, -5, -6, 1, 21, 1, -5, 6, -13,
    -- filter=61 channel=56
    -1, 2, 0, 1, 2, 0, 3, 1, 5,
    -- filter=61 channel=57
    -5, -2, -6, -2, 2, -3, 5, -5, 0,
    -- filter=61 channel=58
    0, -8, -6, -4, -8, 1, -3, -1, -6,
    -- filter=61 channel=59
    0, 6, 7, -2, 15, 7, 4, 0, -2,
    -- filter=61 channel=60
    -2, 3, 6, 3, 0, 5, -5, -5, 1,
    -- filter=61 channel=61
    7, 3, 0, -6, -4, -1, -2, -9, -7,
    -- filter=61 channel=62
    0, -3, 0, 0, 4, 0, -6, -3, -3,
    -- filter=61 channel=63
    -4, -6, 5, -8, -10, 4, -5, -2, 3,
    -- filter=61 channel=64
    4, 0, -4, 8, 3, -7, -4, 1, -1,
    -- filter=61 channel=65
    -6, 6, 0, 4, -5, -4, -1, -6, -3,
    -- filter=61 channel=66
    -4, 5, 1, 0, 6, 1, 1, -5, 1,
    -- filter=61 channel=67
    6, -1, 5, 7, 5, -3, 6, 4, 4,
    -- filter=61 channel=68
    0, -3, -7, 5, 1, 4, -1, 2, -2,
    -- filter=61 channel=69
    -6, -6, -3, -4, 0, 5, -3, 2, -5,
    -- filter=61 channel=70
    1, -3, 5, 7, -1, -7, 2, 3, -8,
    -- filter=61 channel=71
    -1, 4, 5, 0, 5, 1, -1, -3, 6,
    -- filter=61 channel=72
    4, -1, 4, 1, 9, 2, 0, 2, -15,
    -- filter=61 channel=73
    -10, 3, -3, 3, 9, -7, -5, -1, -8,
    -- filter=61 channel=74
    7, 3, 1, 6, 6, 3, -2, -11, -6,
    -- filter=61 channel=75
    -5, -18, 6, -9, 0, 7, 3, 1, 3,
    -- filter=61 channel=76
    -9, 0, -15, 0, 15, 0, 1, 3, -1,
    -- filter=61 channel=77
    -2, -3, 5, -6, 6, 3, 5, 5, 1,
    -- filter=61 channel=78
    -5, -7, 3, 6, 3, 4, 6, -8, 5,
    -- filter=61 channel=79
    -6, 3, -1, -1, 7, 7, 0, 0, -10,
    -- filter=61 channel=80
    -5, 0, 13, -6, 10, -2, 0, -1, -10,
    -- filter=61 channel=81
    4, 0, 2, 0, -6, 0, 0, -2, -5,
    -- filter=61 channel=82
    0, -6, 5, 1, -1, -6, 5, -2, -4,
    -- filter=61 channel=83
    4, 5, 5, -3, 7, -1, 5, -10, 0,
    -- filter=61 channel=84
    2, 10, -8, 0, 12, 4, -10, -4, 0,
    -- filter=61 channel=85
    3, 0, 5, -6, 6, -1, -6, 5, -1,
    -- filter=61 channel=86
    -2, -8, 0, 4, -9, 2, 0, 0, -5,
    -- filter=61 channel=87
    0, 0, 5, -3, -2, -1, 0, -10, -9,
    -- filter=61 channel=88
    4, 0, 2, 9, -2, -8, -3, -2, -4,
    -- filter=61 channel=89
    -8, 6, -6, 6, 22, -1, 1, -1, -4,
    -- filter=61 channel=90
    9, -8, 7, 1, 5, 0, -5, -11, -1,
    -- filter=61 channel=91
    -12, 1, 4, 3, 10, -7, 4, 0, -7,
    -- filter=61 channel=92
    -4, 0, 4, 2, -9, 5, -1, 2, -6,
    -- filter=61 channel=93
    -9, 1, 8, -5, -14, 0, -1, -4, -6,
    -- filter=61 channel=94
    0, 4, 4, 0, -5, -4, -2, -3, -4,
    -- filter=61 channel=95
    -5, -3, 1, -6, -1, -2, -1, -5, 0,
    -- filter=61 channel=96
    -1, 1, 2, 2, -3, -2, 0, -4, 3,
    -- filter=61 channel=97
    4, -5, 7, -9, -7, 1, -3, 2, 0,
    -- filter=61 channel=98
    -7, 0, 6, 0, 8, 6, 6, -8, -14,
    -- filter=61 channel=99
    0, 9, 11, 12, 10, -5, 2, -13, -22,
    -- filter=61 channel=100
    -1, -2, -7, -4, -6, 3, 5, -4, -1,
    -- filter=61 channel=101
    4, -7, -2, -8, -10, -8, -8, -6, 0,
    -- filter=61 channel=102
    -5, -1, 5, 1, -2, -1, 5, -4, -3,
    -- filter=61 channel=103
    -3, -14, 7, -6, 2, 4, -3, 3, -3,
    -- filter=61 channel=104
    -1, 7, 10, 7, 2, -7, -1, 0, -6,
    -- filter=61 channel=105
    -12, 1, 0, -4, 2, -4, -1, 2, 1,
    -- filter=61 channel=106
    4, 6, 1, 5, -3, -5, -7, -6, -4,
    -- filter=61 channel=107
    -10, -3, -9, 5, 11, 0, -8, -4, -3,
    -- filter=61 channel=108
    -5, 0, -4, 3, 2, -6, -4, 2, 3,
    -- filter=61 channel=109
    -14, 8, 9, 8, 18, 8, 3, -13, -15,
    -- filter=61 channel=110
    8, -7, 5, -1, 1, -2, -3, 4, -13,
    -- filter=61 channel=111
    0, -2, 1, -5, 0, 7, -1, -1, 0,
    -- filter=61 channel=112
    3, -1, 1, 0, 3, 1, 0, -5, -8,
    -- filter=61 channel=113
    1, -9, 10, -4, 0, 3, -1, -1, 0,
    -- filter=61 channel=114
    -9, -2, 1, -8, 9, -2, 5, -9, -11,
    -- filter=61 channel=115
    0, -1, 4, 6, 4, 6, 5, -2, 2,
    -- filter=61 channel=116
    -2, 8, -1, -4, 6, -3, -6, -6, -13,
    -- filter=61 channel=117
    -6, 2, 6, 3, -3, -3, 7, -4, -8,
    -- filter=61 channel=118
    2, 1, 6, -7, 2, 3, -3, -2, 4,
    -- filter=61 channel=119
    5, 0, 3, 4, 2, 5, 1, -3, -3,
    -- filter=61 channel=120
    -12, 7, 6, 13, 15, -4, 0, -10, -19,
    -- filter=61 channel=121
    5, 2, 6, -8, 4, 3, 0, 7, 3,
    -- filter=61 channel=122
    -4, -4, 15, -12, 0, 7, 1, 0, -8,
    -- filter=61 channel=123
    2, -4, 7, -4, -2, -7, 0, -8, -6,
    -- filter=61 channel=124
    -2, 3, -7, 0, 9, 0, -7, 3, -5,
    -- filter=61 channel=125
    -4, 4, 10, 7, 8, -7, -3, -4, -9,
    -- filter=61 channel=126
    -4, -9, 0, -7, 3, 2, -2, -1, 7,
    -- filter=61 channel=127
    2, 5, -7, 2, -2, -5, -6, 0, 3,
    -- filter=62 channel=0
    4, 7, 0, -1, -27, -20, -6, -25, -27,
    -- filter=62 channel=1
    4, -1, 3, -4, -16, -18, -4, -16, -15,
    -- filter=62 channel=2
    3, -2, 1, 7, -6, -6, 4, 0, 9,
    -- filter=62 channel=3
    4, -11, 5, -9, -10, -11, 3, -2, 10,
    -- filter=62 channel=4
    -4, -6, -10, 3, -2, 5, 8, -6, -3,
    -- filter=62 channel=5
    0, 3, -1, 0, -22, -15, -9, -17, -11,
    -- filter=62 channel=6
    1, -1, 2, 0, -5, -2, -7, 0, 4,
    -- filter=62 channel=7
    -6, -6, -5, -3, -4, 1, 1, 2, 0,
    -- filter=62 channel=8
    -7, 1, 3, -5, -4, -1, -3, -2, 0,
    -- filter=62 channel=9
    0, 5, -9, 4, -9, -4, 0, -4, 5,
    -- filter=62 channel=10
    -8, -6, 7, -7, 7, 6, 6, 5, 8,
    -- filter=62 channel=11
    -6, -4, -8, -2, 5, 4, -5, 8, 11,
    -- filter=62 channel=12
    5, 5, 5, 6, 0, -5, 3, 10, 8,
    -- filter=62 channel=13
    6, -1, -1, -5, 8, 3, 5, 2, 6,
    -- filter=62 channel=14
    2, -6, -2, 1, 1, -5, 1, -5, 3,
    -- filter=62 channel=15
    4, -9, -1, -4, 0, 0, -9, 0, 2,
    -- filter=62 channel=16
    2, -4, 7, -7, -6, -3, 0, 2, 0,
    -- filter=62 channel=17
    2, -6, 1, 5, 4, 3, 1, -2, 6,
    -- filter=62 channel=18
    3, -10, 2, -14, 5, -2, -3, -4, -3,
    -- filter=62 channel=19
    -5, 5, 3, 3, -5, -3, 7, 2, -7,
    -- filter=62 channel=20
    -14, -1, -13, 1, 22, 21, -7, 5, 18,
    -- filter=62 channel=21
    3, 8, 3, 13, 5, -3, 15, 11, 5,
    -- filter=62 channel=22
    -7, 0, -8, -6, -10, -8, 0, -5, -6,
    -- filter=62 channel=23
    -1, 2, -4, 3, 14, -1, 1, 12, 17,
    -- filter=62 channel=24
    2, 6, 5, -3, 6, 5, 7, -6, -6,
    -- filter=62 channel=25
    -7, 4, 0, -5, 2, -6, 2, -3, -10,
    -- filter=62 channel=26
    0, 6, 6, 7, -11, 4, -6, 0, -5,
    -- filter=62 channel=27
    -6, 11, -11, -3, 4, 1, 0, 2, -6,
    -- filter=62 channel=28
    0, 3, 6, 6, -3, -4, 4, -4, -2,
    -- filter=62 channel=29
    -17, -13, -13, 5, 12, 9, -2, 0, -2,
    -- filter=62 channel=30
    8, -1, -1, -2, -1, -11, 7, -1, -4,
    -- filter=62 channel=31
    6, 0, -7, 13, 17, -8, 18, 18, -5,
    -- filter=62 channel=32
    -8, 0, 0, -13, 4, 1, -6, -1, 3,
    -- filter=62 channel=33
    6, -3, 9, -11, 5, 0, 5, -5, -3,
    -- filter=62 channel=34
    -11, 1, 4, -11, -1, -3, -18, 0, 6,
    -- filter=62 channel=35
    1, -3, -2, -3, 2, 5, -2, -5, 3,
    -- filter=62 channel=36
    1, 0, -2, 4, 16, 2, 0, 9, 13,
    -- filter=62 channel=37
    10, 7, 8, -4, -22, -14, -3, -12, -3,
    -- filter=62 channel=38
    -2, -1, -4, -1, 8, -1, 3, 0, 6,
    -- filter=62 channel=39
    0, 3, -6, -3, 12, 11, 3, 11, -3,
    -- filter=62 channel=40
    0, 4, 4, 8, 12, 8, -3, 9, 1,
    -- filter=62 channel=41
    -17, -2, 11, -12, 7, -1, -8, 0, -4,
    -- filter=62 channel=42
    -3, -2, 6, -3, -9, -12, 6, -6, 2,
    -- filter=62 channel=43
    -3, -6, -5, 0, 4, -8, -8, 2, 0,
    -- filter=62 channel=44
    1, 9, -3, -8, -13, -15, 8, -13, -6,
    -- filter=62 channel=45
    2, 4, -1, 11, 6, 3, -2, 0, 6,
    -- filter=62 channel=46
    5, 5, 7, -9, -5, -8, -6, 2, 5,
    -- filter=62 channel=47
    3, 7, 10, -11, -10, -9, 2, -5, 2,
    -- filter=62 channel=48
    0, 1, -1, 3, -4, -9, 4, -5, -5,
    -- filter=62 channel=49
    -2, 0, -11, -5, -1, 3, -7, 0, 1,
    -- filter=62 channel=50
    1, 9, -7, 6, 7, -8, 4, 2, 0,
    -- filter=62 channel=51
    -1, -5, 5, -1, 0, -6, 0, 5, -4,
    -- filter=62 channel=52
    -1, 5, -2, -1, 5, 0, -1, 9, 7,
    -- filter=62 channel=53
    -7, 0, -1, 7, 6, 9, -2, -1, -3,
    -- filter=62 channel=54
    2, 0, -4, -3, 2, 1, -7, 2, -3,
    -- filter=62 channel=55
    -13, -1, -3, 3, 15, 13, -6, 17, 16,
    -- filter=62 channel=56
    4, 4, -3, 2, 0, -3, -6, 0, 0,
    -- filter=62 channel=57
    -8, -3, -6, 3, 0, -1, -2, 3, 0,
    -- filter=62 channel=58
    -1, 1, 0, -9, -9, -7, -5, -11, -7,
    -- filter=62 channel=59
    1, 2, 2, 1, -5, -1, -1, 1, 4,
    -- filter=62 channel=60
    7, 6, -1, 5, -3, -5, 6, 3, 2,
    -- filter=62 channel=61
    3, 4, 4, 0, -1, 11, -1, 2, 0,
    -- filter=62 channel=62
    -1, -3, 2, -2, 2, 0, 7, -4, 3,
    -- filter=62 channel=63
    1, 0, 5, 6, -9, -3, 4, 2, -9,
    -- filter=62 channel=64
    0, 4, -3, 8, 9, 0, -3, 2, 0,
    -- filter=62 channel=65
    1, 5, -2, 0, -3, -3, 4, -4, -1,
    -- filter=62 channel=66
    -2, 7, 5, -2, 4, 8, 0, 5, 1,
    -- filter=62 channel=67
    5, -4, -7, 6, -4, -3, -6, -3, -5,
    -- filter=62 channel=68
    0, 7, -3, -1, 4, -1, 2, 2, 0,
    -- filter=62 channel=69
    1, -5, 6, 3, -3, 0, 0, -2, 6,
    -- filter=62 channel=70
    3, 1, 7, -2, 2, -3, 2, -8, 0,
    -- filter=62 channel=71
    0, -7, 6, 8, 7, 4, 0, -1, 0,
    -- filter=62 channel=72
    0, 7, -5, 9, 9, 5, 17, 18, 8,
    -- filter=62 channel=73
    -9, 1, -8, 2, 10, 3, -9, 2, 7,
    -- filter=62 channel=74
    -4, 9, 0, 1, 5, 2, -2, -1, -5,
    -- filter=62 channel=75
    6, -3, 8, -11, -22, -16, -1, -10, -20,
    -- filter=62 channel=76
    -9, 2, 4, 3, 20, 20, 1, 5, 17,
    -- filter=62 channel=77
    2, -5, 6, 0, 6, 3, -6, 3, -4,
    -- filter=62 channel=78
    2, 2, -1, -7, 2, -11, 6, -4, 0,
    -- filter=62 channel=79
    -1, 1, -1, -12, 5, -4, -4, 0, 4,
    -- filter=62 channel=80
    -2, 7, 2, 0, 2, -14, 6, 19, -5,
    -- filter=62 channel=81
    -6, 6, -6, 6, -6, 2, -4, 0, 0,
    -- filter=62 channel=82
    7, 0, 3, 1, -3, 0, -6, 0, 2,
    -- filter=62 channel=83
    -5, -4, -1, 6, -6, 0, -4, -1, 5,
    -- filter=62 channel=84
    -4, 5, 0, 1, 3, 5, -9, -4, 4,
    -- filter=62 channel=85
    -1, -7, 6, -2, -1, 5, -5, -6, -6,
    -- filter=62 channel=86
    1, 6, 10, -9, -8, -1, 0, -2, 6,
    -- filter=62 channel=87
    -6, -5, -1, 5, 13, 11, -2, -1, 9,
    -- filter=62 channel=88
    -8, 6, 5, 5, 17, 9, 8, 10, 6,
    -- filter=62 channel=89
    -1, 1, -8, 5, 15, 7, 10, 15, 10,
    -- filter=62 channel=90
    -4, -2, -4, 4, 18, -2, 9, 15, 5,
    -- filter=62 channel=91
    -1, -2, -7, 7, 1, -1, 1, 3, 7,
    -- filter=62 channel=92
    5, -3, 5, -7, 3, -6, 0, -8, 2,
    -- filter=62 channel=93
    -8, 0, 1, -8, -17, -21, 6, -10, -2,
    -- filter=62 channel=94
    -4, 6, -1, -5, -3, 3, -3, -4, -4,
    -- filter=62 channel=95
    -3, -3, 1, -3, 5, 0, -3, -2, -4,
    -- filter=62 channel=96
    7, -4, -7, -2, 0, 2, -3, -2, 2,
    -- filter=62 channel=97
    9, -8, -5, -3, -7, -5, 4, -7, 1,
    -- filter=62 channel=98
    -1, -4, 1, -2, -3, -4, -1, 7, -14,
    -- filter=62 channel=99
    -15, 3, -11, 0, 25, 0, 4, 15, 6,
    -- filter=62 channel=100
    0, 1, 0, -1, 4, 0, -3, 7, -3,
    -- filter=62 channel=101
    1, 2, -10, -2, -5, 6, 1, 5, 1,
    -- filter=62 channel=102
    7, -3, 3, 1, 0, -4, 2, 4, 7,
    -- filter=62 channel=103
    -2, -5, 8, 3, -17, -10, 8, -10, -13,
    -- filter=62 channel=104
    -5, 1, -10, 2, 1, 0, 4, 17, -4,
    -- filter=62 channel=105
    0, -2, 0, -8, 7, 2, -9, 0, 13,
    -- filter=62 channel=106
    -5, 2, -4, 6, 9, 7, 7, 7, 4,
    -- filter=62 channel=107
    -13, 0, 0, -7, 2, 2, -8, -7, 4,
    -- filter=62 channel=108
    -8, 2, 1, 0, 4, -7, 4, -7, 0,
    -- filter=62 channel=109
    -6, 2, -4, -15, 0, 0, -2, 4, -6,
    -- filter=62 channel=110
    4, -1, 1, -3, 3, 5, -1, 15, -1,
    -- filter=62 channel=111
    -8, -2, 9, 0, -1, -1, -3, -4, 9,
    -- filter=62 channel=112
    -1, 5, 8, 0, -4, 3, -3, -10, -1,
    -- filter=62 channel=113
    6, -5, -2, -7, 5, 5, -4, 0, 1,
    -- filter=62 channel=114
    -8, 0, -7, -18, -23, -16, -6, -13, -13,
    -- filter=62 channel=115
    3, -1, 3, -6, 4, -3, 3, 0, 3,
    -- filter=62 channel=116
    0, -7, -12, -6, 11, 0, 8, 7, -1,
    -- filter=62 channel=117
    -5, -4, 2, 3, 1, 0, 5, 8, -1,
    -- filter=62 channel=118
    5, -2, -4, 3, -5, 3, 1, -4, -4,
    -- filter=62 channel=119
    -9, 7, 8, -4, 5, -4, -7, 1, 0,
    -- filter=62 channel=120
    -4, 3, -5, 6, 6, 4, -8, 3, 8,
    -- filter=62 channel=121
    -1, 7, 5, -1, 4, 8, 2, 8, 7,
    -- filter=62 channel=122
    7, 10, 13, -4, -1, -9, 18, 10, -2,
    -- filter=62 channel=123
    -4, 8, 2, 2, 0, -3, -4, -3, 2,
    -- filter=62 channel=124
    -11, 0, -6, -4, 5, 3, -4, -7, 3,
    -- filter=62 channel=125
    -10, 0, -8, -6, 18, 1, 0, 15, -3,
    -- filter=62 channel=126
    0, 2, 0, 1, 9, 1, 2, 4, -6,
    -- filter=62 channel=127
    0, 5, 5, -5, 0, 3, 6, 6, -1,
    -- filter=63 channel=0
    8, -4, 7, -3, -7, 7, 6, 0, 7,
    -- filter=63 channel=1
    7, 2, 9, -6, -18, 6, 8, -14, 4,
    -- filter=63 channel=2
    -3, -7, 0, -5, -4, -2, 4, 1, 0,
    -- filter=63 channel=3
    0, 0, -11, 5, -4, -4, 0, -7, -7,
    -- filter=63 channel=4
    -8, -12, -3, 1, -10, -18, 1, -9, -15,
    -- filter=63 channel=5
    -4, -4, 9, -12, -15, 10, 6, -8, 2,
    -- filter=63 channel=6
    2, -1, 3, 1, 0, 0, 4, 2, 2,
    -- filter=63 channel=7
    6, -1, 0, 0, 0, 6, 3, 6, 1,
    -- filter=63 channel=8
    -6, 0, 0, -3, 4, -2, 2, -1, 2,
    -- filter=63 channel=9
    -1, -8, 0, -5, -4, 0, -1, 0, 11,
    -- filter=63 channel=10
    10, 0, -10, 3, 0, 15, -8, -1, 13,
    -- filter=63 channel=11
    0, -6, -3, -3, 2, -1, -4, 3, 0,
    -- filter=63 channel=12
    -5, 0, 6, 1, 0, 5, 2, -3, 6,
    -- filter=63 channel=13
    0, -3, -5, 4, -2, 5, 2, -3, 6,
    -- filter=63 channel=14
    5, -2, 7, 0, 4, -4, -5, 5, -2,
    -- filter=63 channel=15
    9, 5, 4, 2, -6, -6, -9, -6, 5,
    -- filter=63 channel=16
    -4, 2, -1, -3, -10, 16, -4, -5, 15,
    -- filter=63 channel=17
    1, -6, 2, -2, -1, -2, 1, -2, -2,
    -- filter=63 channel=18
    6, -8, -3, -6, -2, 14, -9, 0, 7,
    -- filter=63 channel=19
    -2, 4, -3, 4, -2, 0, -7, -6, 4,
    -- filter=63 channel=20
    4, -1, 8, -3, 12, -4, -4, 6, -2,
    -- filter=63 channel=21
    -6, -6, -7, -9, -12, 4, -2, -6, 6,
    -- filter=63 channel=22
    5, 6, -4, -2, 0, -6, -5, -5, -4,
    -- filter=63 channel=23
    4, -15, -10, -13, -5, 4, -11, 6, -9,
    -- filter=63 channel=24
    -3, -2, -2, 0, 4, -5, -1, -2, -4,
    -- filter=63 channel=25
    5, -7, 10, 0, -18, 28, 2, -3, 18,
    -- filter=63 channel=26
    1, -2, -1, -7, -8, 1, -5, 1, 6,
    -- filter=63 channel=27
    -1, -17, 13, -9, -9, 21, -6, -2, 10,
    -- filter=63 channel=28
    0, 7, -1, -1, 4, 0, 1, 0, 5,
    -- filter=63 channel=29
    6, 0, 2, 9, -1, 9, -6, 1, 0,
    -- filter=63 channel=30
    -3, -4, 0, 1, -6, 6, 1, -4, 10,
    -- filter=63 channel=31
    -8, -19, -7, -25, 0, 13, -10, 15, 15,
    -- filter=63 channel=32
    9, -4, 5, 3, -15, 8, -9, 2, 9,
    -- filter=63 channel=33
    7, -6, 0, -8, -10, 7, -3, 0, 10,
    -- filter=63 channel=34
    -17, 7, 13, -12, 8, -4, 1, 17, 0,
    -- filter=63 channel=35
    -1, -6, 0, 5, -6, 5, 1, -5, -3,
    -- filter=63 channel=36
    -5, -6, -3, -9, 2, -1, -4, 7, 4,
    -- filter=63 channel=37
    -6, -13, 11, -12, -13, 3, 3, -6, -3,
    -- filter=63 channel=38
    9, 0, 0, -6, 0, 9, -4, 3, 13,
    -- filter=63 channel=39
    -6, 4, 2, 2, 5, 2, -2, 0, 2,
    -- filter=63 channel=40
    0, -1, -2, -7, -2, 0, -3, 2, -1,
    -- filter=63 channel=41
    -10, 10, 4, -8, 4, 19, 4, 5, 6,
    -- filter=63 channel=42
    9, -9, -7, 6, -1, 2, -3, -2, 6,
    -- filter=63 channel=43
    2, -3, -4, -3, 1, -9, -6, 3, 4,
    -- filter=63 channel=44
    -7, -8, 0, -15, 0, 8, -5, 4, 13,
    -- filter=63 channel=45
    -2, -2, -3, -3, -6, 4, 0, 0, 5,
    -- filter=63 channel=46
    -4, 3, 0, -5, 7, -2, -7, -2, -5,
    -- filter=63 channel=47
    5, -5, 0, -7, -18, 16, 6, 3, 20,
    -- filter=63 channel=48
    -1, -10, 10, -11, -10, 14, -7, -6, 8,
    -- filter=63 channel=49
    -3, -2, 3, -10, 7, 0, 0, 6, 5,
    -- filter=63 channel=50
    2, -1, 8, -1, 4, 1, -14, -3, 7,
    -- filter=63 channel=51
    2, 4, 3, -7, -1, -4, 4, 0, 7,
    -- filter=63 channel=52
    -5, 1, 6, -7, 4, 2, -3, -1, -8,
    -- filter=63 channel=53
    -4, 4, 0, 5, 0, 1, -6, 4, -7,
    -- filter=63 channel=54
    4, 1, 0, -6, 3, 6, -2, -2, -7,
    -- filter=63 channel=55
    10, -6, -6, -5, -9, 7, 0, -6, 6,
    -- filter=63 channel=56
    -7, 8, 6, 4, 15, 6, 1, 4, -1,
    -- filter=63 channel=57
    -5, -1, 2, -6, -8, -1, -4, -2, 1,
    -- filter=63 channel=58
    -5, 1, -3, -5, -8, -3, -3, -6, 2,
    -- filter=63 channel=59
    -3, -2, 2, -1, -10, 19, 0, -3, 20,
    -- filter=63 channel=60
    6, -1, 4, -3, 0, 7, -6, 5, 0,
    -- filter=63 channel=61
    4, 1, 0, 5, 10, 3, 7, 10, 4,
    -- filter=63 channel=62
    2, -5, -2, 7, 2, -7, -4, -7, -3,
    -- filter=63 channel=63
    7, 3, -1, -8, -7, 9, -1, 1, 6,
    -- filter=63 channel=64
    1, -5, 3, 0, 7, 0, -1, -5, -5,
    -- filter=63 channel=65
    -3, -4, -6, 0, -4, 5, 0, -5, -3,
    -- filter=63 channel=66
    3, 7, 6, -3, 8, 15, 7, 4, 10,
    -- filter=63 channel=67
    2, 0, -4, -2, -4, -1, -3, 3, -4,
    -- filter=63 channel=68
    1, -8, -7, -6, -9, -1, 5, 1, -7,
    -- filter=63 channel=69
    2, 5, 7, -3, 6, 8, 0, 6, 1,
    -- filter=63 channel=70
    -8, -14, -3, -15, 3, 1, 0, 4, -4,
    -- filter=63 channel=71
    0, -8, -6, 4, -4, 0, 5, -9, 0,
    -- filter=63 channel=72
    6, -6, -5, -7, -8, 12, -11, -8, 9,
    -- filter=63 channel=73
    1, -9, 5, -2, -5, 12, 0, 7, -1,
    -- filter=63 channel=74
    -15, -5, 7, -6, 4, 6, -9, 6, 0,
    -- filter=63 channel=75
    14, -2, -2, -3, -12, 11, 7, -10, 11,
    -- filter=63 channel=76
    -2, -3, -5, -4, -2, 1, 0, -6, -3,
    -- filter=63 channel=77
    -4, 0, 1, 3, 5, -1, 0, 0, 0,
    -- filter=63 channel=78
    0, 1, 9, -9, 3, 5, 2, 6, 9,
    -- filter=63 channel=79
    0, 0, 5, -3, -19, 11, -1, -6, 16,
    -- filter=63 channel=80
    7, -15, 3, -7, -18, 26, -9, 8, 30,
    -- filter=63 channel=81
    0, 2, 5, -5, 6, -1, 4, 2, 3,
    -- filter=63 channel=82
    -5, 5, 3, 2, 0, -1, 3, 5, -6,
    -- filter=63 channel=83
    3, -1, 4, -7, 2, -3, -4, 2, 5,
    -- filter=63 channel=84
    -10, 2, 1, 0, 3, 10, 1, 5, -1,
    -- filter=63 channel=85
    -2, -4, 7, 6, 4, 2, 0, -3, 3,
    -- filter=63 channel=86
    1, -2, 12, -6, -1, 1, 3, -3, 2,
    -- filter=63 channel=87
    0, 7, 2, 3, 11, 5, 3, -1, -2,
    -- filter=63 channel=88
    -8, 0, 0, -10, 9, 6, -4, 0, -4,
    -- filter=63 channel=89
    6, -1, -9, -2, -21, 17, -4, -2, 12,
    -- filter=63 channel=90
    -1, -6, 4, -15, 9, -2, -6, 11, -1,
    -- filter=63 channel=91
    0, -18, 3, -14, 0, 10, -2, 0, 5,
    -- filter=63 channel=92
    -3, -7, -5, -2, 5, -8, 3, 1, -1,
    -- filter=63 channel=93
    2, -9, 0, -14, -15, 15, 6, 0, 8,
    -- filter=63 channel=94
    2, -4, -6, -5, -5, -2, -5, 0, -4,
    -- filter=63 channel=95
    8, -3, -7, 4, -1, 1, 1, -3, 0,
    -- filter=63 channel=96
    0, 5, 4, 5, -9, 4, 1, -6, 6,
    -- filter=63 channel=97
    -4, 3, -7, 2, -10, -11, 1, -4, 3,
    -- filter=63 channel=98
    0, -4, 1, -13, -15, 27, -7, 1, 25,
    -- filter=63 channel=99
    -9, -11, 0, -16, 0, 14, -5, 18, 2,
    -- filter=63 channel=100
    -3, -3, 0, -3, 3, 4, -5, 3, -6,
    -- filter=63 channel=101
    -5, -1, -6, -1, 3, -1, -5, -2, -10,
    -- filter=63 channel=102
    -2, -7, 3, -4, 3, 4, 4, 2, -6,
    -- filter=63 channel=103
    4, -8, 2, -11, -19, 24, 6, -2, 14,
    -- filter=63 channel=104
    0, -13, 9, -8, 1, 13, -7, 0, 15,
    -- filter=63 channel=105
    5, 1, 4, 9, -2, 3, -5, -2, -8,
    -- filter=63 channel=106
    -2, 4, -5, -5, 5, -7, 1, 3, -6,
    -- filter=63 channel=107
    2, 3, 0, -2, 0, 2, -6, 4, -11,
    -- filter=63 channel=108
    5, 9, 4, 3, -5, 8, -2, -7, 3,
    -- filter=63 channel=109
    -6, -12, 3, -8, -1, 25, -11, -3, 11,
    -- filter=63 channel=110
    -1, -1, 1, -9, -5, 8, -8, -2, 6,
    -- filter=63 channel=111
    4, -3, 6, -5, 2, -4, 0, 2, 7,
    -- filter=63 channel=112
    -8, 0, 0, -5, -5, 9, -7, -1, -2,
    -- filter=63 channel=113
    8, -12, -6, -7, -7, -2, -2, 0, 1,
    -- filter=63 channel=114
    6, -8, 14, -9, -8, 13, -9, 0, 13,
    -- filter=63 channel=115
    6, -1, 6, 2, -3, 1, 1, 0, 6,
    -- filter=63 channel=116
    -8, -16, -3, -5, -3, 20, -12, -8, 11,
    -- filter=63 channel=117
    3, 4, -6, -5, -5, -1, -6, -2, 6,
    -- filter=63 channel=118
    -5, 0, 3, -7, -1, -2, 1, 5, -5,
    -- filter=63 channel=119
    -18, 7, 13, -8, 19, 5, -6, 10, 6,
    -- filter=63 channel=120
    -8, -16, 17, -13, 10, 6, -22, 13, 3,
    -- filter=63 channel=121
    6, -5, 1, 5, -4, 9, 6, 1, 0,
    -- filter=63 channel=122
    3, -12, 7, -8, -12, 26, 1, -3, 24,
    -- filter=63 channel=123
    -5, 1, 6, -4, 5, 1, -3, -3, -5,
    -- filter=63 channel=124
    4, -1, -4, 0, 7, 3, -3, -4, -4,
    -- filter=63 channel=125
    -8, -8, 7, -3, -9, 14, -10, -5, 12,
    -- filter=63 channel=126
    1, 1, -2, -3, -14, 8, -4, 0, 8,
    -- filter=63 channel=127
    -5, -2, 8, 5, 7, 0, 5, 0, 6,
    -- filter=64 channel=0
    -3, -13, -1, 2, 14, 9, 8, 20, 11,
    -- filter=64 channel=1
    -9, -1, -9, -3, 7, 5, 14, 8, 14,
    -- filter=64 channel=2
    0, 8, 6, -4, 5, -6, 2, 0, -8,
    -- filter=64 channel=3
    4, 3, 4, -1, 7, -3, -2, -2, -3,
    -- filter=64 channel=4
    7, 2, 2, 0, -6, -4, -3, 0, 6,
    -- filter=64 channel=5
    -1, -11, -9, 7, 10, -3, 14, 10, 15,
    -- filter=64 channel=6
    -1, 2, -5, 4, 3, 6, 0, 5, -1,
    -- filter=64 channel=7
    2, 2, -5, 0, 5, 0, 1, 0, 2,
    -- filter=64 channel=8
    -6, 3, 1, -5, -4, -2, -6, 2, -1,
    -- filter=64 channel=9
    -2, 5, 1, -2, -1, 8, 5, -9, 2,
    -- filter=64 channel=10
    1, 6, -6, 1, 2, 1, 1, -7, 3,
    -- filter=64 channel=11
    -1, 1, -5, -1, 7, 2, -4, -5, -12,
    -- filter=64 channel=12
    -1, 4, 2, 2, 4, -2, 4, 0, 4,
    -- filter=64 channel=13
    0, 0, -8, 0, -4, 6, 4, -10, -3,
    -- filter=64 channel=14
    3, 3, -1, 1, -5, -3, 4, -6, 1,
    -- filter=64 channel=15
    12, 7, -4, -6, 5, 3, -4, -14, -7,
    -- filter=64 channel=16
    -11, -6, -3, -5, -2, -7, 2, -12, 4,
    -- filter=64 channel=17
    3, 6, -4, 2, 4, -4, 0, 0, -2,
    -- filter=64 channel=18
    11, 8, -3, 10, 6, 15, -3, -11, 1,
    -- filter=64 channel=19
    0, 4, -5, 3, -1, -6, 5, 5, -7,
    -- filter=64 channel=20
    11, -4, 0, 11, 6, -10, 0, -12, -14,
    -- filter=64 channel=21
    -10, -13, -16, -8, -13, -1, -11, -10, -1,
    -- filter=64 channel=22
    3, -1, -7, 2, 3, 3, -5, 1, 1,
    -- filter=64 channel=23
    9, 6, 6, -12, 13, 7, -16, -6, 6,
    -- filter=64 channel=24
    3, 3, 5, 0, 6, -3, -1, 3, -3,
    -- filter=64 channel=25
    3, 0, -4, -5, 1, 5, 1, -6, 0,
    -- filter=64 channel=26
    0, -8, 0, -1, -11, -4, 1, -3, -3,
    -- filter=64 channel=27
    8, -7, 1, -14, 7, 19, 3, -16, 15,
    -- filter=64 channel=28
    6, -2, -7, 6, 5, 5, 4, 6, 4,
    -- filter=64 channel=29
    11, 4, 6, 11, 4, 3, 0, -3, -15,
    -- filter=64 channel=30
    -2, -2, -5, -4, 0, 5, 8, 7, 9,
    -- filter=64 channel=31
    6, -3, -14, -15, 0, -2, -10, -14, 6,
    -- filter=64 channel=32
    11, 4, 0, 2, -1, 12, 2, -14, 9,
    -- filter=64 channel=33
    5, 5, 5, 1, 9, 1, 0, -11, 10,
    -- filter=64 channel=34
    9, -4, 1, 0, 9, 2, -6, 17, 7,
    -- filter=64 channel=35
    5, -3, 0, -5, 5, -7, 1, 2, 6,
    -- filter=64 channel=36
    4, -3, -6, -6, -8, -1, 2, -11, -4,
    -- filter=64 channel=37
    -6, -9, -12, -4, 6, 1, 0, 15, 16,
    -- filter=64 channel=38
    -1, 0, 4, -8, 2, 3, -5, -10, 9,
    -- filter=64 channel=39
    7, -2, 1, 7, -5, -4, -8, -1, -2,
    -- filter=64 channel=40
    5, 0, -11, 0, 1, -8, 2, -2, -3,
    -- filter=64 channel=41
    7, 11, -3, 0, -1, -2, -3, 6, 2,
    -- filter=64 channel=42
    0, 3, -5, 0, -9, -1, 4, -1, 1,
    -- filter=64 channel=43
    2, -2, 0, 3, 15, 2, 6, -4, -8,
    -- filter=64 channel=44
    -13, -10, -12, -3, -9, -5, 1, -4, 11,
    -- filter=64 channel=45
    -9, -10, -1, 4, 5, 4, 5, 6, 6,
    -- filter=64 channel=46
    1, 3, 3, -4, -1, -5, 0, 9, -3,
    -- filter=64 channel=47
    -15, -19, -16, -7, -11, 1, 1, -7, -4,
    -- filter=64 channel=48
    -9, -2, -3, -7, -12, 8, -1, -6, 7,
    -- filter=64 channel=49
    -3, 0, -1, -4, -6, 5, 2, 0, 4,
    -- filter=64 channel=50
    2, 1, -9, -10, 5, 9, -8, -6, 1,
    -- filter=64 channel=51
    5, 5, 5, -3, 1, 5, 2, 6, 7,
    -- filter=64 channel=52
    0, 0, 2, 1, -1, 5, 3, -5, -3,
    -- filter=64 channel=53
    10, 6, 0, 9, 7, 0, 1, -10, 4,
    -- filter=64 channel=54
    -3, -3, 4, 1, 5, 0, 6, 1, 0,
    -- filter=64 channel=55
    5, 0, 4, 2, 1, 6, -4, -16, -11,
    -- filter=64 channel=56
    3, 0, 3, 2, 5, 8, -3, 2, -1,
    -- filter=64 channel=57
    5, 8, 8, 7, 4, 3, 2, 4, 7,
    -- filter=64 channel=58
    6, -3, 1, 8, 5, 2, 10, 5, 3,
    -- filter=64 channel=59
    -8, -3, -3, -5, -12, 6, -2, -11, 2,
    -- filter=64 channel=60
    1, 3, 6, 0, -1, -4, -5, 5, 7,
    -- filter=64 channel=61
    -7, -7, -5, -5, 2, 0, -5, -6, -4,
    -- filter=64 channel=62
    7, 0, -5, -6, 5, -1, -4, 0, -4,
    -- filter=64 channel=63
    5, -5, -7, 9, 1, 8, 0, 2, 8,
    -- filter=64 channel=64
    7, 0, 0, -3, -3, 1, 1, -1, -4,
    -- filter=64 channel=65
    1, 5, -1, 3, 0, -3, 1, -6, -1,
    -- filter=64 channel=66
    5, -6, -3, -3, 3, 8, 0, -5, -1,
    -- filter=64 channel=67
    3, 0, 0, -6, 6, -6, -3, 0, -3,
    -- filter=64 channel=68
    -2, 0, -1, -3, 2, -3, 0, -10, -7,
    -- filter=64 channel=69
    6, -4, 6, 6, 6, -3, 0, -1, 3,
    -- filter=64 channel=70
    -1, 2, -4, -13, 9, 3, -5, -2, 9,
    -- filter=64 channel=71
    -6, -3, 0, -3, 5, -9, -5, -6, -1,
    -- filter=64 channel=72
    4, 7, -3, -4, -4, -1, 0, -14, 4,
    -- filter=64 channel=73
    4, 1, 3, 3, 0, 0, 1, -3, -3,
    -- filter=64 channel=74
    -2, 0, -6, -15, 6, -4, -7, -7, 14,
    -- filter=64 channel=75
    -5, -6, -11, 6, 10, 7, 4, 18, 2,
    -- filter=64 channel=76
    11, -3, -6, 6, -2, -5, -1, -6, -19,
    -- filter=64 channel=77
    0, 0, -1, -2, 6, 6, -1, 5, -4,
    -- filter=64 channel=78
    -2, -3, -2, 1, 1, -4, -5, -3, 1,
    -- filter=64 channel=79
    7, -3, 0, 6, -1, 8, 2, -4, 0,
    -- filter=64 channel=80
    1, -3, -6, -8, -18, -3, -10, -20, -2,
    -- filter=64 channel=81
    -7, 2, -3, 1, 1, 1, -1, 4, -7,
    -- filter=64 channel=82
    -5, -3, 2, 1, 3, -5, 1, 5, 5,
    -- filter=64 channel=83
    -8, -2, 7, -9, 2, -7, -3, -3, 5,
    -- filter=64 channel=84
    0, 2, 8, -2, 3, 3, 7, -5, -1,
    -- filter=64 channel=85
    -1, 1, 1, 0, 0, 0, -1, 5, -3,
    -- filter=64 channel=86
    -2, -3, 4, -4, 8, 1, 8, -1, 7,
    -- filter=64 channel=87
    2, 5, 0, -5, 2, 6, 0, 4, -3,
    -- filter=64 channel=88
    -10, -8, 1, 1, 2, -6, -10, -5, -11,
    -- filter=64 channel=89
    12, 13, 2, -2, -6, 2, 0, -17, -5,
    -- filter=64 channel=90
    -7, 2, -5, -5, 2, 0, -1, -8, -1,
    -- filter=64 channel=91
    -4, -4, -3, -9, -2, 7, -2, -11, -3,
    -- filter=64 channel=92
    5, 6, 3, -1, 10, 4, 0, 7, 8,
    -- filter=64 channel=93
    -8, -10, 0, -5, 4, 6, -4, -2, 11,
    -- filter=64 channel=94
    2, 3, -2, 6, 3, 0, -1, -5, -5,
    -- filter=64 channel=95
    -2, -2, -6, -2, 0, 3, 0, -5, -6,
    -- filter=64 channel=96
    -1, 4, 5, -6, -3, -4, -6, -9, 5,
    -- filter=64 channel=97
    -5, -9, 1, 1, 6, -4, 5, -2, 3,
    -- filter=64 channel=98
    0, -2, 5, -2, -8, 1, -6, -14, -1,
    -- filter=64 channel=99
    13, 6, 2, -11, 12, 3, -8, -5, -1,
    -- filter=64 channel=100
    9, 6, 7, 0, -4, 7, -7, 7, 2,
    -- filter=64 channel=101
    2, 7, -6, 1, -3, 3, 4, 0, 5,
    -- filter=64 channel=102
    -1, 2, -2, 1, 0, 2, -2, -6, -5,
    -- filter=64 channel=103
    -1, -8, 0, -7, -7, 0, -7, -1, 4,
    -- filter=64 channel=104
    -11, -1, -7, -8, -9, 5, -7, -14, -5,
    -- filter=64 channel=105
    -2, 4, 2, 10, 6, 0, 5, -5, -5,
    -- filter=64 channel=106
    -1, -8, -8, 0, -4, -4, 2, -9, -10,
    -- filter=64 channel=107
    6, 0, 4, -3, 13, 7, -7, 3, 3,
    -- filter=64 channel=108
    8, 2, 3, 0, 9, 5, -2, 0, 4,
    -- filter=64 channel=109
    8, -4, 6, -3, -1, 14, -3, -5, 12,
    -- filter=64 channel=110
    4, 5, 2, 7, 6, 6, 2, 1, 0,
    -- filter=64 channel=111
    3, 5, 1, 5, 2, -5, 8, 2, 0,
    -- filter=64 channel=112
    2, -1, -4, -8, 11, -1, 4, -1, 10,
    -- filter=64 channel=113
    11, -2, -1, -7, 2, -3, 1, -9, 4,
    -- filter=64 channel=114
    -3, -8, 0, 2, 6, 14, 11, 5, 11,
    -- filter=64 channel=115
    0, 4, 4, -2, -2, 5, -3, -3, 5,
    -- filter=64 channel=116
    9, 8, 6, -5, -10, 7, 3, -15, -5,
    -- filter=64 channel=117
    0, 2, 3, -2, -2, -4, -4, 2, -5,
    -- filter=64 channel=118
    -1, -5, -5, 4, 5, 4, -4, 5, -5,
    -- filter=64 channel=119
    1, -5, 4, 0, 16, 6, 0, 8, 10,
    -- filter=64 channel=120
    5, -4, 3, -17, 5, 13, -6, -12, 12,
    -- filter=64 channel=121
    7, -4, 0, 3, -1, 5, -1, -8, -2,
    -- filter=64 channel=122
    -20, -25, -25, -21, -26, -9, -15, -16, -4,
    -- filter=64 channel=123
    -4, 1, 1, 5, 9, -3, -7, 1, 3,
    -- filter=64 channel=124
    -4, 5, 7, 7, 4, -2, -7, -6, 0,
    -- filter=64 channel=125
    -5, 5, -2, 1, -5, 9, 1, -10, 8,
    -- filter=64 channel=126
    5, 3, 0, 1, -6, 10, 2, -7, -1,
    -- filter=64 channel=127
    -3, 7, -2, 3, 0, -1, -5, 5, -2,
    -- filter=65 channel=0
    2, 11, 10, 9, 5, 0, -4, -10, -1,
    -- filter=65 channel=1
    6, 1, 9, -2, 0, 5, 0, 2, 6,
    -- filter=65 channel=2
    -6, 4, 8, -6, 0, -5, -1, 10, 5,
    -- filter=65 channel=3
    -2, -1, -14, 3, -8, -7, 3, 4, -11,
    -- filter=65 channel=4
    6, 0, -3, 6, 7, -4, 14, 13, 4,
    -- filter=65 channel=5
    9, 2, 8, 1, -3, 1, -8, -9, -3,
    -- filter=65 channel=6
    7, -3, 4, 11, 0, 0, 11, -1, -8,
    -- filter=65 channel=7
    5, 6, -6, -2, 1, -1, 6, -7, 2,
    -- filter=65 channel=8
    -9, 0, 14, -5, 9, 0, -6, 0, -1,
    -- filter=65 channel=9
    5, -7, 1, -4, -1, 9, -8, 2, 8,
    -- filter=65 channel=10
    0, -4, 3, -9, -5, 7, 2, 0, 6,
    -- filter=65 channel=11
    0, 0, 0, 11, -6, -12, 6, -5, 2,
    -- filter=65 channel=12
    0, 3, 9, -1, 3, 5, -5, 6, 4,
    -- filter=65 channel=13
    -9, -11, -3, -6, -5, 0, 0, -11, 6,
    -- filter=65 channel=14
    6, -1, 6, 1, 2, 3, -3, -5, 2,
    -- filter=65 channel=15
    -2, -4, 0, 4, -11, 3, 0, 0, 2,
    -- filter=65 channel=16
    1, 1, 0, -6, -12, -2, -9, 0, -3,
    -- filter=65 channel=17
    -2, 0, 2, 5, -7, 0, 0, -2, 7,
    -- filter=65 channel=18
    0, -9, 3, 7, -13, 5, 6, 0, 7,
    -- filter=65 channel=19
    -7, 2, 4, 4, 1, -7, 2, 2, -5,
    -- filter=65 channel=20
    15, -2, 7, 10, -5, -6, 1, 3, 1,
    -- filter=65 channel=21
    -7, -4, -5, -18, -7, 0, -20, -4, 0,
    -- filter=65 channel=22
    -4, -1, 9, 0, 2, 10, 4, -4, -4,
    -- filter=65 channel=23
    0, -8, 7, -15, -8, 10, -1, -2, 10,
    -- filter=65 channel=24
    -6, 1, -5, 6, 3, 0, 1, 5, -6,
    -- filter=65 channel=25
    -11, -13, 4, -5, -10, 11, 4, -1, 19,
    -- filter=65 channel=26
    -3, -2, 0, -4, 1, 8, -1, -3, 6,
    -- filter=65 channel=27
    -5, -11, 12, -11, -13, 14, 0, 4, 21,
    -- filter=65 channel=28
    7, 2, 0, -2, 2, -3, -2, -4, 4,
    -- filter=65 channel=29
    13, -1, -7, 18, -2, -3, 18, 1, -12,
    -- filter=65 channel=30
    0, -4, 10, 0, -6, 7, 0, 5, 6,
    -- filter=65 channel=31
    -13, -18, 14, -16, -4, 15, -19, 6, 16,
    -- filter=65 channel=32
    3, -9, -1, 4, -17, -1, 0, 3, 9,
    -- filter=65 channel=33
    -1, -5, -7, 0, -4, 8, -8, -5, 5,
    -- filter=65 channel=34
    -6, -4, 23, -16, 0, 17, -1, 1, 6,
    -- filter=65 channel=35
    -6, 3, -1, -5, -2, 1, 0, 1, 1,
    -- filter=65 channel=36
    2, 0, -3, -2, -7, 6, -5, -1, -3,
    -- filter=65 channel=37
    4, 6, 8, -4, 8, 9, -2, 4, -8,
    -- filter=65 channel=38
    -10, -5, 1, -11, -9, 5, -8, 0, 2,
    -- filter=65 channel=39
    -1, -6, -2, 7, 4, -4, 10, 3, 0,
    -- filter=65 channel=40
    0, 0, -6, 0, -4, -8, 7, 0, -5,
    -- filter=65 channel=41
    0, 2, -1, 0, -4, 9, 0, -6, 1,
    -- filter=65 channel=42
    5, 0, -6, -3, -5, -3, 0, 5, -4,
    -- filter=65 channel=43
    3, 0, 3, 0, 1, -7, 9, -1, -2,
    -- filter=65 channel=44
    -8, -3, 10, -1, -2, 12, -6, -7, -2,
    -- filter=65 channel=45
    1, 1, 1, 5, 2, -5, -4, 6, 5,
    -- filter=65 channel=46
    5, -5, -1, 1, -5, -6, -1, -2, 2,
    -- filter=65 channel=47
    -12, -16, 2, -6, -3, 0, -15, -9, 0,
    -- filter=65 channel=48
    0, -6, 10, -9, -10, 16, -7, 1, 17,
    -- filter=65 channel=49
    -5, 3, -2, 2, 2, 3, 12, 0, 2,
    -- filter=65 channel=50
    -10, -13, 0, -10, -9, 8, -1, 11, 11,
    -- filter=65 channel=51
    3, 1, 0, 5, 4, -7, 1, -1, 1,
    -- filter=65 channel=52
    -9, -7, 6, -4, -1, 8, 5, -1, 6,
    -- filter=65 channel=53
    -3, -7, 0, 8, -7, 3, 3, -3, 1,
    -- filter=65 channel=54
    -7, 6, -2, 1, -3, 6, -7, 6, -5,
    -- filter=65 channel=55
    3, -12, -5, 0, -10, 4, -2, -7, -1,
    -- filter=65 channel=56
    -7, 5, 16, 1, 11, 3, 4, -4, 0,
    -- filter=65 channel=57
    0, 0, -5, -7, 0, 1, 3, -3, 1,
    -- filter=65 channel=58
    9, 10, 9, -2, -3, 1, 0, 1, -8,
    -- filter=65 channel=59
    -3, -14, 0, -4, -15, 15, -7, -5, 4,
    -- filter=65 channel=60
    7, -3, -5, 0, 3, -5, 0, 5, -7,
    -- filter=65 channel=61
    -6, -7, -5, -2, -4, 4, -2, -3, -6,
    -- filter=65 channel=62
    5, -1, -1, 5, 2, 5, -6, 2, 5,
    -- filter=65 channel=63
    -3, 7, -1, 0, 2, 1, 3, -10, 0,
    -- filter=65 channel=64
    3, -3, -2, -2, 2, -5, 6, -2, 3,
    -- filter=65 channel=65
    -7, 7, 6, 0, -5, 4, 1, 4, 3,
    -- filter=65 channel=66
    -7, 7, 4, -10, -4, 2, 2, -5, 9,
    -- filter=65 channel=67
    -1, 4, -1, 0, -6, 3, 2, 5, 0,
    -- filter=65 channel=68
    2, -7, -7, 2, -1, 2, 8, -2, -5,
    -- filter=65 channel=69
    -1, 5, 0, 0, -2, 3, -6, 3, 4,
    -- filter=65 channel=70
    -3, -1, 14, -3, -6, 8, -10, 5, 7,
    -- filter=65 channel=71
    -6, -7, -11, 0, 1, -3, -7, -5, 1,
    -- filter=65 channel=72
    -10, -14, 2, -16, -10, 8, -13, 2, 7,
    -- filter=65 channel=73
    -5, -1, 9, -3, 2, 11, -1, 11, 0,
    -- filter=65 channel=74
    -13, -6, 27, -16, -4, 11, -10, 13, 4,
    -- filter=65 channel=75
    -7, 8, -3, 7, 4, 1, -8, 0, -4,
    -- filter=65 channel=76
    12, 0, -11, 3, -10, -10, 13, -10, -2,
    -- filter=65 channel=77
    -7, 4, 5, -6, -6, 0, -1, -1, -3,
    -- filter=65 channel=78
    0, -5, 9, -2, 3, -2, -1, 3, -4,
    -- filter=65 channel=79
    5, -19, 7, -4, -18, 5, 7, -11, 2,
    -- filter=65 channel=80
    -16, -17, -5, -13, -10, 8, -17, -2, 9,
    -- filter=65 channel=81
    0, -7, -3, -5, 7, 0, 3, 7, 2,
    -- filter=65 channel=82
    -5, 3, -4, 4, 6, 0, 0, -6, -7,
    -- filter=65 channel=83
    -8, 0, -7, 1, 3, -2, -1, -2, 7,
    -- filter=65 channel=84
    2, 0, 6, -2, 3, 0, 11, 0, 3,
    -- filter=65 channel=85
    -6, 3, -2, 6, -6, -1, -5, -2, 6,
    -- filter=65 channel=86
    5, -4, 13, 4, 0, 2, -3, -5, 7,
    -- filter=65 channel=87
    -4, 2, 8, -3, 3, 1, 5, -5, 4,
    -- filter=65 channel=88
    3, -6, 11, -10, 4, 3, -6, -3, 2,
    -- filter=65 channel=89
    -3, -11, -1, -11, -12, 8, -8, 1, 13,
    -- filter=65 channel=90
    -10, -2, 11, -5, 0, 6, -14, -2, 4,
    -- filter=65 channel=91
    1, -12, 10, -3, -8, 7, 6, 0, 16,
    -- filter=65 channel=92
    3, -4, -3, 2, 1, 6, 4, 0, 8,
    -- filter=65 channel=93
    0, 1, 8, -6, -1, 10, 0, 1, -1,
    -- filter=65 channel=94
    1, 3, 2, 0, 0, -2, 7, 0, 0,
    -- filter=65 channel=95
    0, 5, -6, 3, 5, 6, -4, -5, -5,
    -- filter=65 channel=96
    -5, 0, 3, -5, 5, 0, -1, 3, 0,
    -- filter=65 channel=97
    2, 2, -4, -5, -4, -9, -6, -1, -5,
    -- filter=65 channel=98
    -9, -18, 8, -9, -16, 13, -7, 2, 23,
    -- filter=65 channel=99
    -13, -14, 12, -20, -5, 18, -10, 11, 20,
    -- filter=65 channel=100
    -3, -3, 8, 2, 1, 6, 7, 0, 2,
    -- filter=65 channel=101
    2, -8, -7, -3, 5, -6, 8, 2, -8,
    -- filter=65 channel=102
    6, -4, 5, 5, 3, -3, -6, 0, 0,
    -- filter=65 channel=103
    -3, -14, -12, 0, -2, 4, -16, -1, 6,
    -- filter=65 channel=104
    -3, -11, 7, -7, -2, 10, -13, -2, 7,
    -- filter=65 channel=105
    7, -6, -7, 15, -8, -9, 11, -9, -4,
    -- filter=65 channel=106
    6, -2, -1, 7, -5, -10, 8, 0, -12,
    -- filter=65 channel=107
    6, 0, 5, 4, 5, 4, 7, -6, -7,
    -- filter=65 channel=108
    -4, 9, -3, -2, -5, -2, 4, -7, -2,
    -- filter=65 channel=109
    -2, -15, 15, -12, 0, 19, -5, 5, 19,
    -- filter=65 channel=110
    2, 1, 0, 1, -3, -5, -2, -10, 8,
    -- filter=65 channel=111
    -5, 4, -4, 8, -1, 3, 0, 2, 5,
    -- filter=65 channel=112
    -7, -5, 17, -14, 7, 16, -5, 10, 10,
    -- filter=65 channel=113
    -12, -7, -4, -11, 0, 6, 0, -3, 7,
    -- filter=65 channel=114
    6, -1, 7, 10, -2, 9, 15, 6, 4,
    -- filter=65 channel=115
    -1, -4, -1, 3, 5, -5, -1, -4, 2,
    -- filter=65 channel=116
    -5, -7, -4, -4, -13, 4, 3, 1, 11,
    -- filter=65 channel=117
    1, -2, -7, -7, 3, 0, -1, -5, 3,
    -- filter=65 channel=118
    3, 1, -5, 3, 5, -6, -6, 7, 2,
    -- filter=65 channel=119
    0, 0, 14, -3, 12, 12, -8, 6, 5,
    -- filter=65 channel=120
    -8, -10, 22, -17, -5, 15, 3, 10, 23,
    -- filter=65 channel=121
    -4, -5, -5, -5, 0, -2, -9, -3, 3,
    -- filter=65 channel=122
    -23, -13, -4, -20, -7, 0, -25, -19, 2,
    -- filter=65 channel=123
    -5, 3, 11, 0, -3, 1, -6, 5, -2,
    -- filter=65 channel=124
    10, -3, -3, 3, 3, 3, 9, -3, -6,
    -- filter=65 channel=125
    -16, -9, 4, -10, -10, 6, -9, 1, 13,
    -- filter=65 channel=126
    0, -4, -8, -5, -8, -4, -5, 2, 0,
    -- filter=65 channel=127
    1, -4, -6, -2, 4, -6, 0, -6, -1,
    -- filter=66 channel=0
    -6, 0, 11, -12, 3, 8, -1, 0, 9,
    -- filter=66 channel=1
    0, 0, 7, -10, -6, 2, 1, 7, 10,
    -- filter=66 channel=2
    1, 0, -3, -4, 0, -4, -6, 7, 7,
    -- filter=66 channel=3
    1, -2, -2, -4, -8, 5, -10, 0, 7,
    -- filter=66 channel=4
    -7, -12, -8, -8, 1, 9, 5, 3, 12,
    -- filter=66 channel=5
    1, 1, -5, -10, -11, 5, 2, -4, 0,
    -- filter=66 channel=6
    -2, -7, 2, -3, 4, 5, 1, 0, -6,
    -- filter=66 channel=7
    4, -6, -1, 3, 6, 6, 4, -7, -1,
    -- filter=66 channel=8
    1, 0, -2, -3, 3, -1, 3, -1, 9,
    -- filter=66 channel=9
    7, -3, -7, -3, -4, -4, 0, -3, 1,
    -- filter=66 channel=10
    0, 4, -11, 0, -3, -1, 8, 4, 5,
    -- filter=66 channel=11
    7, 3, -6, 6, -5, 5, -9, -3, 0,
    -- filter=66 channel=12
    -3, -3, 8, 7, -1, -7, 5, 2, -5,
    -- filter=66 channel=13
    -1, -1, -4, 0, -2, -4, -4, -2, -1,
    -- filter=66 channel=14
    -6, -3, -2, -2, -4, -2, 2, -5, 5,
    -- filter=66 channel=15
    -8, -5, 4, -3, 6, 0, -5, -5, 8,
    -- filter=66 channel=16
    0, 0, 2, -3, 5, -1, -1, 3, -2,
    -- filter=66 channel=17
    -3, 0, 0, 1, 5, -6, -5, -2, 0,
    -- filter=66 channel=18
    0, 6, 13, -1, 8, 11, -16, -3, 7,
    -- filter=66 channel=19
    0, -1, -7, -3, -1, 4, 2, 4, -4,
    -- filter=66 channel=20
    -3, 4, -8, -1, 2, 1, -10, -2, -3,
    -- filter=66 channel=21
    10, 3, -2, 7, -11, -7, 1, 2, -4,
    -- filter=66 channel=22
    -4, 0, 9, -1, 7, 8, -4, 0, 0,
    -- filter=66 channel=23
    7, -3, 1, 6, 1, -6, -7, 8, 6,
    -- filter=66 channel=24
    0, -1, -5, 1, -3, -3, 0, 0, -6,
    -- filter=66 channel=25
    5, 2, -2, -1, 3, 3, -6, 1, 2,
    -- filter=66 channel=26
    -5, -1, 3, -6, 0, -5, -2, -6, -4,
    -- filter=66 channel=27
    1, -6, 6, -9, 0, -1, -6, -3, 0,
    -- filter=66 channel=28
    0, 0, 4, 6, 5, -7, 3, 0, 1,
    -- filter=66 channel=29
    0, -7, 1, -7, -3, -3, -9, -10, -7,
    -- filter=66 channel=30
    -2, -3, 3, 0, -6, -2, -6, 5, 0,
    -- filter=66 channel=31
    6, -11, -6, 12, -9, -14, 11, 10, -1,
    -- filter=66 channel=32
    -1, 7, -2, -8, 1, 0, -10, -5, 8,
    -- filter=66 channel=33
    1, -1, 0, -9, -1, 7, -9, -4, 2,
    -- filter=66 channel=34
    7, 4, 9, 9, -2, 1, -1, 8, -6,
    -- filter=66 channel=35
    -7, 5, -7, 2, 6, 6, -3, 5, -2,
    -- filter=66 channel=36
    5, 2, -6, -2, -3, 1, 7, 2, 1,
    -- filter=66 channel=37
    -8, 5, 6, -4, -8, 6, -1, -6, 10,
    -- filter=66 channel=38
    4, -2, 5, -4, -5, 0, 0, 2, 6,
    -- filter=66 channel=39
    0, 2, 2, -6, 3, 2, -9, -4, -4,
    -- filter=66 channel=40
    3, 0, 3, 3, 2, -2, 2, 2, 5,
    -- filter=66 channel=41
    2, -4, -2, 8, 9, -8, 3, 3, 1,
    -- filter=66 channel=42
    -2, 4, 0, -6, 2, 3, 3, -3, -3,
    -- filter=66 channel=43
    -10, 1, 6, -3, 2, 5, -8, -8, 5,
    -- filter=66 channel=44
    6, -4, 7, 2, -2, -5, 4, 1, 0,
    -- filter=66 channel=45
    -2, 2, 7, 0, -4, -2, -7, -2, -6,
    -- filter=66 channel=46
    -3, 3, -4, 2, 0, -2, 0, -1, -1,
    -- filter=66 channel=47
    -2, 1, -2, -4, 1, -8, 11, 1, 0,
    -- filter=66 channel=48
    3, 3, -6, 1, -6, 1, 1, -4, 8,
    -- filter=66 channel=49
    0, -6, 6, -6, -6, 4, -4, 4, 8,
    -- filter=66 channel=50
    -1, -1, 0, -5, 1, -1, 7, 5, 4,
    -- filter=66 channel=51
    0, 2, 2, -6, -1, -5, 0, -3, 2,
    -- filter=66 channel=52
    -1, 0, 6, 1, -3, 4, 8, 5, 1,
    -- filter=66 channel=53
    8, 1, 4, 2, -2, 0, 1, -5, 0,
    -- filter=66 channel=54
    0, -2, 4, 1, 5, 2, -5, -3, 3,
    -- filter=66 channel=55
    2, 0, 4, -3, -1, -7, -3, 6, -6,
    -- filter=66 channel=56
    3, 0, 6, 5, 7, 3, 2, 0, 7,
    -- filter=66 channel=57
    4, 5, -1, 2, 0, -3, -2, 6, 0,
    -- filter=66 channel=58
    4, -5, -4, -6, 3, -6, -4, -8, -5,
    -- filter=66 channel=59
    6, 3, -4, 1, -1, -1, 8, 2, 0,
    -- filter=66 channel=60
    4, 6, 7, -3, -7, -2, -2, 5, 0,
    -- filter=66 channel=61
    2, 3, -5, 0, 0, -1, 3, 6, -3,
    -- filter=66 channel=62
    -5, -6, 4, -4, 3, 6, -4, 4, -2,
    -- filter=66 channel=63
    2, -6, 0, -5, -7, -7, 0, -3, 0,
    -- filter=66 channel=64
    2, 0, -1, 8, 0, -2, 7, 5, -6,
    -- filter=66 channel=65
    -2, 7, -4, 2, -1, 2, 0, 4, 6,
    -- filter=66 channel=66
    -2, 7, -2, 3, 1, 0, 7, 0, -2,
    -- filter=66 channel=67
    -1, -5, -3, 1, 0, -4, 0, 0, 3,
    -- filter=66 channel=68
    -5, 3, -6, 7, 2, 0, -2, 0, 5,
    -- filter=66 channel=69
    0, -5, 0, 2, -3, -4, 3, 0, 3,
    -- filter=66 channel=70
    1, -3, 7, -4, 4, 0, -3, 4, 2,
    -- filter=66 channel=71
    -1, 3, 2, -5, -5, -2, -1, 1, 6,
    -- filter=66 channel=72
    10, -3, -11, -1, -6, -14, 7, 7, -9,
    -- filter=66 channel=73
    -1, -4, 1, 3, -5, -4, -8, 1, -5,
    -- filter=66 channel=74
    5, -2, 7, -3, 3, 4, 0, 6, -4,
    -- filter=66 channel=75
    -9, 5, 5, 0, -6, 10, 0, 0, 12,
    -- filter=66 channel=76
    8, 0, 0, -1, 6, 5, -2, 1, 0,
    -- filter=66 channel=77
    5, -1, 7, -6, -5, 2, -6, -1, 3,
    -- filter=66 channel=78
    0, -5, -5, 1, -7, -8, -5, -3, 0,
    -- filter=66 channel=79
    -1, -1, 12, -9, 3, 14, -5, -4, 1,
    -- filter=66 channel=80
    0, -1, -5, -4, -5, -16, 5, -1, -1,
    -- filter=66 channel=81
    -4, 6, -6, 7, -5, -5, 0, 6, 0,
    -- filter=66 channel=82
    -6, 6, -2, -3, 0, 7, 4, -5, 0,
    -- filter=66 channel=83
    6, 0, 1, -8, 4, -6, 4, -3, 3,
    -- filter=66 channel=84
    -2, 5, 6, 0, 2, -1, 1, -3, 3,
    -- filter=66 channel=85
    2, 1, -3, -4, -6, -1, 3, -6, 4,
    -- filter=66 channel=86
    1, 7, 8, -1, -6, -4, 4, 4, -3,
    -- filter=66 channel=87
    -4, 0, 7, 0, 3, 8, 4, -5, -3,
    -- filter=66 channel=88
    3, 0, -6, 7, -1, -5, 8, 7, -7,
    -- filter=66 channel=89
    4, 5, -7, 8, -2, -8, 0, 0, 6,
    -- filter=66 channel=90
    1, 1, -9, 13, -3, -3, 0, 2, 4,
    -- filter=66 channel=91
    -5, 1, 4, -7, 8, 0, -7, 5, 10,
    -- filter=66 channel=92
    -5, -4, 0, 7, -3, 6, 4, 6, -1,
    -- filter=66 channel=93
    3, 2, 0, 3, -7, -7, 4, 2, 8,
    -- filter=66 channel=94
    0, 0, 5, 1, 2, 0, 2, 3, -1,
    -- filter=66 channel=95
    0, -2, 7, -4, -5, 4, -5, 4, 1,
    -- filter=66 channel=96
    -6, 0, 3, 0, 2, 3, -1, 0, 1,
    -- filter=66 channel=97
    -6, -2, -6, 6, -2, 1, -1, -5, -4,
    -- filter=66 channel=98
    1, -5, -4, -6, 3, -3, -9, 5, 6,
    -- filter=66 channel=99
    4, -11, -1, 3, -5, -11, 7, 0, -1,
    -- filter=66 channel=100
    5, -1, 5, 7, -2, -5, -3, -3, -3,
    -- filter=66 channel=101
    2, 1, -8, 0, 0, 3, 1, 0, 2,
    -- filter=66 channel=102
    -5, 0, -7, 0, 1, -3, 3, 0, -4,
    -- filter=66 channel=103
    6, 0, -5, -3, -13, -4, -4, -5, 0,
    -- filter=66 channel=104
    9, -3, -14, 5, 1, -17, 0, 7, -8,
    -- filter=66 channel=105
    -2, 5, -7, -6, 5, 0, -10, -6, -4,
    -- filter=66 channel=106
    -5, 8, 0, 6, 5, 1, -1, 1, -4,
    -- filter=66 channel=107
    -2, -6, 9, -2, -5, 1, -12, -1, 2,
    -- filter=66 channel=108
    -8, 0, -2, -3, 4, 4, 0, 2, -2,
    -- filter=66 channel=109
    0, 2, -4, 2, 4, 3, 0, 7, -1,
    -- filter=66 channel=110
    -3, -4, 1, 4, 3, -4, 9, 5, -7,
    -- filter=66 channel=111
    -4, -5, -5, -7, 7, -7, -5, 0, -1,
    -- filter=66 channel=112
    3, -8, -5, -2, 0, 0, -7, 0, 7,
    -- filter=66 channel=113
    0, 7, 3, 4, 0, -9, -4, -5, 3,
    -- filter=66 channel=114
    -8, -3, 14, -10, 2, 11, -19, 0, 3,
    -- filter=66 channel=115
    -3, 3, 0, -2, 5, -5, -1, 0, 3,
    -- filter=66 channel=116
    5, 0, -9, -4, -8, -4, 6, 6, -2,
    -- filter=66 channel=117
    1, 0, -4, 2, 1, 0, 4, 9, -6,
    -- filter=66 channel=118
    5, -3, -1, -6, 0, -2, 2, -6, 0,
    -- filter=66 channel=119
    3, -5, 2, 8, 4, 0, 0, 0, -4,
    -- filter=66 channel=120
    1, 0, 2, -9, -9, -1, -10, 0, 4,
    -- filter=66 channel=121
    9, -4, 3, 5, 2, -3, 1, -3, 6,
    -- filter=66 channel=122
    13, 3, -3, 10, -1, -15, 19, 11, 4,
    -- filter=66 channel=123
    8, 3, 3, -3, -2, 0, -3, -3, -1,
    -- filter=66 channel=124
    -1, 0, -3, -9, 5, 6, -7, -2, -8,
    -- filter=66 channel=125
    5, 1, 0, 3, -9, -9, 6, 1, -7,
    -- filter=66 channel=126
    1, -3, 0, 2, -3, -8, -8, -4, 2,
    -- filter=66 channel=127
    1, 0, 5, -6, 3, -3, 5, 1, -4,
    -- filter=67 channel=0
    -7, -12, 0, -4, -8, 6, 3, -7, 1,
    -- filter=67 channel=1
    -6, -1, 12, -6, -8, 5, -2, 2, 2,
    -- filter=67 channel=2
    -6, 0, -3, 3, -8, 0, 4, -7, 3,
    -- filter=67 channel=3
    -5, 0, -5, -2, -3, -1, -1, -8, -4,
    -- filter=67 channel=4
    5, -4, -3, -4, 0, -1, 4, -4, 0,
    -- filter=67 channel=5
    -7, -4, 5, -12, 2, 5, -3, -3, 2,
    -- filter=67 channel=6
    -2, -1, 2, 1, 3, 2, 3, -7, 4,
    -- filter=67 channel=7
    0, -2, 5, -7, 1, 0, 1, -5, -1,
    -- filter=67 channel=8
    3, 0, -6, -2, -7, 1, 0, 2, 5,
    -- filter=67 channel=9
    0, 5, 3, 0, 6, -4, 1, -6, -3,
    -- filter=67 channel=10
    6, 7, -5, 7, 8, -6, -1, 0, 0,
    -- filter=67 channel=11
    -3, 2, -9, 0, 5, 1, 3, -7, 0,
    -- filter=67 channel=12
    5, -6, 7, 5, -5, 2, 0, -1, -1,
    -- filter=67 channel=13
    3, -9, -10, 2, -1, 0, 5, 0, 0,
    -- filter=67 channel=14
    3, 6, 1, 4, -6, 0, 6, 3, -4,
    -- filter=67 channel=15
    -7, -15, -9, 4, -14, -6, 17, -4, -11,
    -- filter=67 channel=16
    -3, 16, 12, -10, -1, 7, -13, -3, 0,
    -- filter=67 channel=17
    -2, 2, 0, 4, 4, -3, -6, 0, 5,
    -- filter=67 channel=18
    -2, -21, -16, 12, -21, -5, 16, 3, -4,
    -- filter=67 channel=19
    -3, -4, -1, 2, 5, 0, -5, 2, -5,
    -- filter=67 channel=20
    0, -15, -13, 8, -11, 0, 3, 0, 0,
    -- filter=67 channel=21
    11, 14, 13, 7, 11, -1, -3, -7, -7,
    -- filter=67 channel=22
    -5, -10, 2, 0, -8, 1, -3, 1, 6,
    -- filter=67 channel=23
    -5, -12, -13, -5, -19, -14, 7, -11, -16,
    -- filter=67 channel=24
    -4, -4, 5, -7, 7, 1, 5, 2, 0,
    -- filter=67 channel=25
    9, 0, -7, 2, -6, 0, 14, 9, 7,
    -- filter=67 channel=26
    0, 5, 3, -3, 3, 5, -7, 4, 1,
    -- filter=67 channel=27
    1, -17, -11, 10, -6, -15, 15, -6, -11,
    -- filter=67 channel=28
    3, 3, -6, -2, -3, -7, 2, 1, 6,
    -- filter=67 channel=29
    -8, -12, -12, 8, -10, -11, 2, 0, -7,
    -- filter=67 channel=30
    -4, 4, 0, -4, -1, -9, -4, -4, -1,
    -- filter=67 channel=31
    0, 13, 1, 4, 2, -1, -11, -1, -12,
    -- filter=67 channel=32
    6, -8, -11, 9, -8, -14, 14, 2, -5,
    -- filter=67 channel=33
    5, -11, -8, -2, -13, -8, 13, 4, -10,
    -- filter=67 channel=34
    -1, -3, 0, -6, -14, -10, -4, -7, -5,
    -- filter=67 channel=35
    7, 5, 3, -5, 0, -6, -5, -3, -3,
    -- filter=67 channel=36
    3, 9, -4, 9, 0, 2, -10, -5, 1,
    -- filter=67 channel=37
    -7, 0, 2, -5, -11, 10, -7, -7, 10,
    -- filter=67 channel=38
    -8, -7, 1, 0, 1, -7, 7, 1, -3,
    -- filter=67 channel=39
    -3, -3, -2, -5, -2, -6, 8, -1, 0,
    -- filter=67 channel=40
    -4, 4, -7, 0, -1, 3, 5, -3, 5,
    -- filter=67 channel=41
    -3, -3, 11, 0, 0, 7, 10, 5, 16,
    -- filter=67 channel=42
    -6, -6, 6, -3, -5, -8, -2, -5, -4,
    -- filter=67 channel=43
    0, -5, -3, 0, -7, 0, 11, -2, -4,
    -- filter=67 channel=44
    -3, 0, 1, -1, -2, 4, -6, -1, 5,
    -- filter=67 channel=45
    -2, -6, 4, 1, -8, -7, 4, -1, -1,
    -- filter=67 channel=46
    2, 0, -5, 2, -1, 5, 4, 7, -5,
    -- filter=67 channel=47
    -1, 8, 18, -7, 10, 11, -10, 0, 0,
    -- filter=67 channel=48
    10, 11, 3, 6, 11, 0, 4, 5, 3,
    -- filter=67 channel=49
    -9, -6, 1, 4, -12, -6, 6, 4, -5,
    -- filter=67 channel=50
    4, -7, -10, 7, -8, -5, 10, 1, -11,
    -- filter=67 channel=51
    0, 0, -7, -3, -7, -4, 1, 0, -1,
    -- filter=67 channel=52
    -5, -6, -4, 0, -8, -9, 5, -9, 0,
    -- filter=67 channel=53
    -2, -1, -10, -2, 1, -1, 0, 1, -9,
    -- filter=67 channel=54
    7, -5, 2, 1, 4, 0, -3, -3, 2,
    -- filter=67 channel=55
    7, -13, -16, 5, -15, -5, 14, 4, -5,
    -- filter=67 channel=56
    3, -8, 3, 1, -8, 5, 2, 0, -5,
    -- filter=67 channel=57
    1, -3, 6, 0, -2, 0, -5, -6, 9,
    -- filter=67 channel=58
    -1, 0, 3, 0, -8, 2, -1, -5, 2,
    -- filter=67 channel=59
    5, 2, 0, 14, 8, 0, 0, -4, 0,
    -- filter=67 channel=60
    -5, 4, -3, -2, 1, -1, 6, -5, 1,
    -- filter=67 channel=61
    0, 3, -5, -5, 5, 6, -7, 4, 1,
    -- filter=67 channel=62
    -6, 5, 4, -1, -5, 1, 6, 3, 3,
    -- filter=67 channel=63
    -1, -2, 7, -8, 6, 11, -2, -4, 3,
    -- filter=67 channel=64
    7, -4, -2, 5, 0, -4, 6, -7, 4,
    -- filter=67 channel=65
    -6, -1, -3, -5, -5, 2, 7, 0, -5,
    -- filter=67 channel=66
    -1, 1, 0, 0, -4, 6, 0, -4, 10,
    -- filter=67 channel=67
    0, 5, -7, -4, -1, 5, 1, -1, -2,
    -- filter=67 channel=68
    -1, 6, 4, 3, -4, 6, 5, 2, 6,
    -- filter=67 channel=69
    4, 7, 7, -5, 1, 8, 3, 0, 2,
    -- filter=67 channel=70
    -8, -16, -9, 0, -9, -9, 6, 1, -2,
    -- filter=67 channel=71
    -1, 6, 6, -7, 1, -5, -1, -1, -4,
    -- filter=67 channel=72
    9, 7, -10, 11, 10, -9, 4, 7, -2,
    -- filter=67 channel=73
    -2, -15, -7, 2, -10, -9, 14, -3, -3,
    -- filter=67 channel=74
    -11, 0, 0, -11, -9, 0, 2, -2, -7,
    -- filter=67 channel=75
    -8, 0, 8, -11, -2, 4, 7, -6, -2,
    -- filter=67 channel=76
    5, -6, -13, 0, -5, -9, 9, -9, 1,
    -- filter=67 channel=77
    0, 3, 0, -3, -6, 2, 1, 4, -6,
    -- filter=67 channel=78
    1, 7, 0, -9, -6, -4, -12, 1, -7,
    -- filter=67 channel=79
    -7, -13, -12, 0, -24, -3, 20, -6, -2,
    -- filter=67 channel=80
    3, 13, -2, 13, 6, -8, 8, -3, -12,
    -- filter=67 channel=81
    0, 2, 2, -5, -7, -4, 6, 2, -6,
    -- filter=67 channel=82
    1, -3, -7, -4, -8, -6, -7, 2, -5,
    -- filter=67 channel=83
    3, 6, 0, 9, 11, -5, 2, -2, 3,
    -- filter=67 channel=84
    5, -13, -6, 10, -7, -1, 5, 0, -1,
    -- filter=67 channel=85
    2, -1, 2, -5, -2, -2, -4, 7, 7,
    -- filter=67 channel=86
    1, 0, -2, 1, -7, 1, -7, 0, 5,
    -- filter=67 channel=87
    -4, -2, 3, 0, -7, 2, 0, 0, -2,
    -- filter=67 channel=88
    11, 0, 2, 6, 10, -5, -1, 0, -2,
    -- filter=67 channel=89
    0, -10, -5, 10, -1, -11, 16, 1, -11,
    -- filter=67 channel=90
    -3, 0, -7, -3, 8, 7, -14, -8, -2,
    -- filter=67 channel=91
    0, -10, -12, 0, -13, -11, 10, -4, -5,
    -- filter=67 channel=92
    3, 2, -6, 4, 3, 5, -2, -8, -1,
    -- filter=67 channel=93
    1, 15, 11, -4, 9, -2, -1, -4, 0,
    -- filter=67 channel=94
    -1, 2, 5, 1, -5, 5, 1, -2, -6,
    -- filter=67 channel=95
    -1, -1, -2, 2, 3, 4, -7, -7, -7,
    -- filter=67 channel=96
    -4, 1, 5, 6, 3, 2, 6, 4, -5,
    -- filter=67 channel=97
    1, -2, 2, -4, 0, 1, 3, -4, 4,
    -- filter=67 channel=98
    -4, -3, 0, 10, 0, 0, 11, -7, -5,
    -- filter=67 channel=99
    2, -1, -11, 2, -10, -13, 6, -6, -11,
    -- filter=67 channel=100
    -4, -2, 4, 6, -2, -6, 4, 2, -6,
    -- filter=67 channel=101
    -6, 5, 9, 1, -10, 5, -7, -3, 5,
    -- filter=67 channel=102
    -6, 4, 5, 3, -4, 1, 0, 5, -4,
    -- filter=67 channel=103
    0, 10, 15, -4, 3, 13, -10, -1, 0,
    -- filter=67 channel=104
    6, 5, -2, 5, 11, -3, 0, 4, -1,
    -- filter=67 channel=105
    -2, -12, -4, 4, -3, -10, 5, 0, -3,
    -- filter=67 channel=106
    -1, -2, -1, 6, 0, 2, 5, -1, 1,
    -- filter=67 channel=107
    -10, -18, -16, -1, -15, 0, 1, -1, -9,
    -- filter=67 channel=108
    -4, 4, -2, -4, -2, 2, -1, 3, 3,
    -- filter=67 channel=109
    7, -4, -11, 4, 0, -2, 18, 6, -3,
    -- filter=67 channel=110
    3, 0, -10, 4, 0, -1, 1, -3, -5,
    -- filter=67 channel=111
    6, -4, 3, 8, -5, 1, 6, 0, 8,
    -- filter=67 channel=112
    -6, -2, 5, -4, -5, -9, -7, 2, -3,
    -- filter=67 channel=113
    2, 1, -8, 5, -1, -5, -1, -8, -10,
    -- filter=67 channel=114
    -9, -20, -10, -2, -15, -15, 10, 0, -7,
    -- filter=67 channel=115
    7, 2, 5, -4, -1, 0, 2, -7, 1,
    -- filter=67 channel=116
    6, 5, 0, 17, 7, 0, 8, 6, 3,
    -- filter=67 channel=117
    8, 7, 2, -5, -2, -5, -3, 4, -6,
    -- filter=67 channel=118
    -6, -5, 5, 0, 2, 3, 3, -7, -1,
    -- filter=67 channel=119
    -5, -10, -9, -9, -8, -6, 2, -9, -6,
    -- filter=67 channel=120
    2, -18, -10, 4, -12, -16, 3, -10, -5,
    -- filter=67 channel=121
    -1, -2, -1, 5, -5, 4, 0, -3, -5,
    -- filter=67 channel=122
    0, 32, 11, -12, 20, 17, -22, -2, -6,
    -- filter=67 channel=123
    -5, 6, 0, 1, -2, 3, 0, -7, 2,
    -- filter=67 channel=124
    -3, -2, -5, 3, -4, 3, -4, 2, 4,
    -- filter=67 channel=125
    7, 7, 1, 9, -2, -11, -3, 6, -4,
    -- filter=67 channel=126
    -2, -8, -3, -2, -5, 0, 15, 2, -4,
    -- filter=67 channel=127
    -3, -5, -2, -5, -3, -3, 3, 3, 0,
    -- filter=68 channel=0
    -5, 0, 2, 0, 5, 0, 1, -4, -4,
    -- filter=68 channel=1
    1, -1, 3, -7, 1, -1, -3, -4, 5,
    -- filter=68 channel=2
    2, -7, -5, -1, 4, -3, 5, 5, -1,
    -- filter=68 channel=3
    7, -3, -5, 1, 5, 8, -4, 3, -6,
    -- filter=68 channel=4
    -1, -6, -1, -2, 0, 3, -6, 5, 8,
    -- filter=68 channel=5
    2, -3, 2, 5, -6, 5, 6, 1, -7,
    -- filter=68 channel=6
    -2, 5, 6, 0, -2, 0, 3, 4, 1,
    -- filter=68 channel=7
    0, -3, 1, 2, 0, -3, 0, 6, 4,
    -- filter=68 channel=8
    4, -1, 1, 0, -7, 6, -2, 4, -2,
    -- filter=68 channel=9
    -2, 6, 3, 5, 0, -7, -5, -6, 0,
    -- filter=68 channel=10
    -2, 3, 2, 0, -3, 0, 0, -3, 4,
    -- filter=68 channel=11
    6, -5, -2, 7, 1, -5, -2, -4, -4,
    -- filter=68 channel=12
    3, -6, -2, -6, -6, -4, -5, 0, 0,
    -- filter=68 channel=13
    1, -6, -2, -5, 5, -5, -2, 3, 0,
    -- filter=68 channel=14
    -6, 3, 3, -1, -5, 0, -2, -5, -4,
    -- filter=68 channel=15
    -4, 0, -2, 0, 2, -7, -2, 0, 0,
    -- filter=68 channel=16
    4, -2, -2, 4, 5, -7, 4, -3, 1,
    -- filter=68 channel=17
    -2, -5, 5, 3, -4, 1, -7, 0, 6,
    -- filter=68 channel=18
    2, -7, -5, 0, 2, -3, 5, -5, -1,
    -- filter=68 channel=19
    6, -6, -4, 4, -5, 0, -6, -4, 3,
    -- filter=68 channel=20
    2, 6, 8, 1, 5, -5, 0, 4, 6,
    -- filter=68 channel=21
    -4, 1, 2, -1, 4, -2, -6, 0, 2,
    -- filter=68 channel=22
    3, -3, -1, 0, 3, 5, 0, 0, 1,
    -- filter=68 channel=23
    7, 8, 10, -2, -7, -5, 5, 5, -3,
    -- filter=68 channel=24
    1, -6, -2, 0, -4, 2, -6, -3, -1,
    -- filter=68 channel=25
    -4, -1, 0, 2, 5, -6, 4, 3, -3,
    -- filter=68 channel=26
    5, -1, -1, -2, -2, -2, -4, -1, -1,
    -- filter=68 channel=27
    4, 1, 3, -8, -5, 5, -6, -4, -2,
    -- filter=68 channel=28
    1, -1, -6, 3, -5, -2, -6, 1, 1,
    -- filter=68 channel=29
    -1, -4, 7, 2, -1, 3, 7, -2, 7,
    -- filter=68 channel=30
    -8, -7, 3, -2, 4, 3, -3, 0, -1,
    -- filter=68 channel=31
    6, 6, 9, 3, 1, 3, 5, -7, -6,
    -- filter=68 channel=32
    -6, 3, -4, -3, -6, -7, 6, -4, 0,
    -- filter=68 channel=33
    2, -6, -1, -4, -4, -4, 4, -4, -4,
    -- filter=68 channel=34
    -4, 3, 4, -1, -6, 0, -3, 1, 5,
    -- filter=68 channel=35
    2, -5, -1, 0, 3, 4, -1, 0, -1,
    -- filter=68 channel=36
    5, 4, 2, 2, -2, -5, -2, 6, 2,
    -- filter=68 channel=37
    1, -5, -2, -3, -2, 2, -2, -3, -2,
    -- filter=68 channel=38
    -1, 0, 0, 0, -5, 1, 0, 0, 5,
    -- filter=68 channel=39
    -3, 0, -1, 0, 3, 1, 7, 8, -6,
    -- filter=68 channel=40
    -1, 0, 7, -1, 6, -1, -2, 2, -5,
    -- filter=68 channel=41
    2, 0, -8, -5, -2, 0, 4, -2, -6,
    -- filter=68 channel=42
    -3, 0, -2, 3, -5, 3, 1, 6, -1,
    -- filter=68 channel=43
    -2, -5, 5, 1, -1, 0, 3, 0, 0,
    -- filter=68 channel=44
    -3, 1, 5, 6, -7, 0, 7, -2, 4,
    -- filter=68 channel=45
    -3, -5, -5, 5, 5, -2, 3, -1, -5,
    -- filter=68 channel=46
    -2, -4, 4, -1, -6, -1, -7, 0, -5,
    -- filter=68 channel=47
    -7, 1, 0, 1, -3, 2, -3, -3, 3,
    -- filter=68 channel=48
    -4, -7, 2, 2, 0, 5, 5, 0, -6,
    -- filter=68 channel=49
    -5, -8, 0, 6, 0, 0, -3, 4, 5,
    -- filter=68 channel=50
    1, -5, -3, 4, 2, 7, -4, -5, 3,
    -- filter=68 channel=51
    0, 6, 0, -6, -7, -5, 3, 3, -3,
    -- filter=68 channel=52
    8, 0, 1, 1, 0, -3, -3, -6, -3,
    -- filter=68 channel=53
    -5, 7, 7, 2, 7, 4, 0, 6, 3,
    -- filter=68 channel=54
    6, 5, 6, -7, 0, 4, 5, -2, 0,
    -- filter=68 channel=55
    -6, -5, -5, 2, 6, 5, 0, -1, 6,
    -- filter=68 channel=56
    4, -7, -1, -3, -4, -4, 6, -2, -1,
    -- filter=68 channel=57
    -4, -4, 1, 2, -6, -7, -2, -6, -1,
    -- filter=68 channel=58
    -3, 5, -3, 3, -2, 7, -6, 3, -4,
    -- filter=68 channel=59
    5, -1, 3, -5, -5, -6, 2, -7, -1,
    -- filter=68 channel=60
    6, 6, -7, 3, 5, 0, 0, 4, -6,
    -- filter=68 channel=61
    1, -5, -6, 4, 0, 2, 5, 4, 5,
    -- filter=68 channel=62
    -3, 7, -2, -6, 1, 5, -4, 6, 3,
    -- filter=68 channel=63
    4, 0, 2, 0, 5, -6, 3, 6, 5,
    -- filter=68 channel=64
    0, 0, -4, -2, 2, 4, 1, -6, 2,
    -- filter=68 channel=65
    1, 6, 7, 1, 0, 5, 1, 2, 2,
    -- filter=68 channel=66
    3, 7, 3, 0, -1, 5, -3, 4, 0,
    -- filter=68 channel=67
    4, 0, 4, -3, -3, 2, 7, 7, 1,
    -- filter=68 channel=68
    4, -3, 3, 3, 4, 1, 2, 0, -1,
    -- filter=68 channel=69
    6, -2, -2, 6, 5, -6, 1, -4, 5,
    -- filter=68 channel=70
    2, 0, -5, -5, 1, 3, -5, 1, -5,
    -- filter=68 channel=71
    0, -3, -4, -3, 4, -6, -7, -3, -4,
    -- filter=68 channel=72
    3, 4, -5, -5, -6, 4, 2, -5, 3,
    -- filter=68 channel=73
    0, 6, -2, -4, -2, 4, 1, 4, 1,
    -- filter=68 channel=74
    7, 0, -3, 6, -6, -6, 3, 3, 3,
    -- filter=68 channel=75
    -5, -1, 1, 5, -7, 3, 4, 0, -7,
    -- filter=68 channel=76
    1, 8, -3, 7, -3, 0, 3, 6, 2,
    -- filter=68 channel=77
    -6, -5, -5, 2, 5, -4, 3, 6, 6,
    -- filter=68 channel=78
    5, -2, -6, 7, -6, -6, 2, 3, 4,
    -- filter=68 channel=79
    -8, 0, -5, 0, 0, -8, -5, -5, 4,
    -- filter=68 channel=80
    2, 0, -5, 2, 3, -8, -2, 6, -5,
    -- filter=68 channel=81
    6, -7, -7, -4, -2, 1, -4, -6, -3,
    -- filter=68 channel=82
    -6, 7, -2, -6, 4, 0, 0, -1, 6,
    -- filter=68 channel=83
    -2, -6, 0, 0, -1, -5, 3, 5, 1,
    -- filter=68 channel=84
    -3, 0, 3, 4, 2, 7, -6, 3, 5,
    -- filter=68 channel=85
    0, 0, -6, -2, 5, -4, -6, -2, 1,
    -- filter=68 channel=86
    0, 3, -2, 4, 3, 7, -6, -7, -1,
    -- filter=68 channel=87
    -5, -4, 8, -2, -4, -4, 3, 6, 0,
    -- filter=68 channel=88
    0, 5, 8, 0, -3, 8, 3, 0, -6,
    -- filter=68 channel=89
    4, -6, 0, -3, -3, -6, 5, 6, -5,
    -- filter=68 channel=90
    4, 2, 0, 2, 0, 3, 0, -5, 0,
    -- filter=68 channel=91
    -2, -7, 3, -7, 3, -2, 7, -3, -6,
    -- filter=68 channel=92
    -1, -5, 7, -4, -7, 5, 1, 5, -1,
    -- filter=68 channel=93
    -3, -8, -1, 2, -2, -8, -2, 4, 6,
    -- filter=68 channel=94
    -5, -4, 4, -5, 6, -2, -5, -1, 4,
    -- filter=68 channel=95
    4, 5, 0, 5, 6, 2, -1, -1, 7,
    -- filter=68 channel=96
    -5, 0, 7, 0, -2, 6, -3, 0, 6,
    -- filter=68 channel=97
    2, -4, 7, 4, 6, 7, 4, 6, -3,
    -- filter=68 channel=98
    6, 1, 6, -5, 4, -7, -4, -3, -6,
    -- filter=68 channel=99
    6, 4, 8, -6, 2, -5, 0, -6, -6,
    -- filter=68 channel=100
    1, 0, -7, 0, 0, 2, -2, 4, -1,
    -- filter=68 channel=101
    0, -2, 1, 7, 7, 0, 4, 5, 5,
    -- filter=68 channel=102
    -5, -5, -6, -1, 3, 0, 7, 1, 5,
    -- filter=68 channel=103
    -5, 2, 0, -4, -6, 2, 1, -6, -7,
    -- filter=68 channel=104
    -4, -6, 7, -4, -7, 2, -3, 1, 4,
    -- filter=68 channel=105
    -5, -1, -4, -3, 3, -5, -6, 1, 5,
    -- filter=68 channel=106
    -6, 0, -3, -4, 6, -5, 4, 1, 1,
    -- filter=68 channel=107
    0, 4, 7, 0, 5, 0, 2, -4, 3,
    -- filter=68 channel=108
    -6, 2, 0, -6, -3, -1, -1, 0, 7,
    -- filter=68 channel=109
    1, 0, 3, -7, 0, -6, -1, -3, -4,
    -- filter=68 channel=110
    2, -4, 0, -3, -6, 5, -3, -6, 5,
    -- filter=68 channel=111
    -2, 1, -4, -2, 0, -1, -4, -6, 1,
    -- filter=68 channel=112
    -6, -4, -3, -3, 3, -1, -1, 0, -1,
    -- filter=68 channel=113
    -2, -1, 3, -4, -4, 4, -2, -1, -5,
    -- filter=68 channel=114
    -1, -8, 6, -2, -6, -4, 0, 2, 0,
    -- filter=68 channel=115
    -6, 2, -6, -3, 6, 4, 7, -3, -6,
    -- filter=68 channel=116
    5, 0, 1, 3, 0, 3, 4, -5, 8,
    -- filter=68 channel=117
    -3, -1, -4, -7, 5, 6, 0, 0, 1,
    -- filter=68 channel=118
    -5, 6, 4, 0, 0, 3, 5, 5, 7,
    -- filter=68 channel=119
    -6, 0, 4, -1, 0, 0, 2, -1, -5,
    -- filter=68 channel=120
    -7, -6, 7, -2, -7, -6, -1, 1, 7,
    -- filter=68 channel=121
    -3, 0, 6, -6, -3, -1, 3, 7, 0,
    -- filter=68 channel=122
    2, -6, 5, 4, 3, -6, 5, 2, 1,
    -- filter=68 channel=123
    6, -4, 7, 6, 0, 1, -1, -3, 0,
    -- filter=68 channel=124
    -6, 0, -4, -3, -6, -3, 0, -6, 0,
    -- filter=68 channel=125
    -2, 3, 4, -7, 0, 5, -5, -3, 4,
    -- filter=68 channel=126
    -7, 0, 5, 6, 5, -2, -8, 1, 1,
    -- filter=68 channel=127
    3, 5, 4, -5, 0, -5, 0, -2, -6,
    -- filter=69 channel=0
    -1, -5, 7, -2, 6, 6, -2, 8, 3,
    -- filter=69 channel=1
    -4, 6, 1, -1, 0, -3, 0, 0, -3,
    -- filter=69 channel=2
    -8, -7, 6, 2, 2, 0, 5, 0, -3,
    -- filter=69 channel=3
    -6, -3, 3, -7, -8, 1, 0, 6, 0,
    -- filter=69 channel=4
    -14, 5, -1, 2, 9, 5, 13, 0, 4,
    -- filter=69 channel=5
    1, 4, 6, 1, 2, 1, 2, -2, 4,
    -- filter=69 channel=6
    -3, -6, 0, -8, 2, -2, -1, 7, -6,
    -- filter=69 channel=7
    2, 7, 5, -4, -4, 0, -4, -4, -3,
    -- filter=69 channel=8
    -8, -5, -5, 8, 8, -7, 7, -7, 0,
    -- filter=69 channel=9
    -3, -4, 1, 7, 0, 2, -5, 5, -3,
    -- filter=69 channel=10
    0, -9, -2, -1, 2, 8, 2, 8, -2,
    -- filter=69 channel=11
    -9, -2, 2, -1, -5, 3, 8, 3, 0,
    -- filter=69 channel=12
    -5, -9, 10, -8, -4, 0, 3, 0, 1,
    -- filter=69 channel=13
    -2, -14, -5, -6, 0, -1, 0, 5, 2,
    -- filter=69 channel=14
    2, 1, 5, 4, 5, -3, -6, 0, -7,
    -- filter=69 channel=15
    -2, -8, 0, -6, -5, 0, 10, 1, 0,
    -- filter=69 channel=16
    3, 10, 0, 5, 3, -4, -2, -5, -1,
    -- filter=69 channel=17
    0, -4, -4, 6, -7, 4, -4, 4, 4,
    -- filter=69 channel=18
    -9, -11, 0, -6, -4, 4, 10, 14, -3,
    -- filter=69 channel=19
    -7, 6, 4, -3, -5, 7, 4, 2, -6,
    -- filter=69 channel=20
    -1, -3, 0, -16, -11, -2, 7, 0, 8,
    -- filter=69 channel=21
    2, 8, 3, -1, -2, 6, -2, -9, -7,
    -- filter=69 channel=22
    2, -6, -2, 2, -1, -6, 1, -1, 4,
    -- filter=69 channel=23
    -12, -13, 1, -20, -9, -5, 11, 0, -4,
    -- filter=69 channel=24
    4, 3, 7, -1, -5, -6, 0, -2, -2,
    -- filter=69 channel=25
    -2, 3, -4, -1, 7, 6, 1, 6, 3,
    -- filter=69 channel=26
    0, 0, 1, 5, 0, -6, -2, -1, 1,
    -- filter=69 channel=27
    -8, -8, 13, -6, 4, -4, 18, 0, 1,
    -- filter=69 channel=28
    -4, 2, 0, 0, -5, -6, -6, -2, -5,
    -- filter=69 channel=29
    -3, -3, 6, -2, -11, -4, 12, 10, 3,
    -- filter=69 channel=30
    -5, 0, 0, 0, 10, -1, 8, -1, -4,
    -- filter=69 channel=31
    0, 7, 10, -7, 5, -2, 5, 0, -8,
    -- filter=69 channel=32
    1, -11, -2, -16, -2, -2, 3, 10, -3,
    -- filter=69 channel=33
    -8, -11, 3, -3, 3, 4, 3, 3, -7,
    -- filter=69 channel=34
    0, -3, 6, 4, 5, 1, 2, 1, -8,
    -- filter=69 channel=35
    7, 0, 7, 0, -3, 3, -2, 4, 0,
    -- filter=69 channel=36
    -4, 0, -2, 0, 3, -3, 3, -6, 2,
    -- filter=69 channel=37
    -7, 5, 0, 9, 2, 5, 2, -9, -2,
    -- filter=69 channel=38
    1, 0, 1, -9, -7, 5, -5, -4, -6,
    -- filter=69 channel=39
    -8, 2, -7, 0, -8, 3, -2, -3, 3,
    -- filter=69 channel=40
    2, -4, 0, -6, -3, -1, -3, -1, -6,
    -- filter=69 channel=41
    9, -1, -1, -7, -2, -4, -6, 11, 0,
    -- filter=69 channel=42
    -1, 6, -4, -3, 0, -4, -3, -7, -6,
    -- filter=69 channel=43
    2, -7, 1, -13, 3, -7, 4, 0, -4,
    -- filter=69 channel=44
    -6, 0, 8, 6, 8, 6, 1, -2, -6,
    -- filter=69 channel=45
    0, 0, -8, 6, 0, -2, 1, -7, 6,
    -- filter=69 channel=46
    0, 0, 1, 6, 3, 2, 0, 5, 0,
    -- filter=69 channel=47
    5, -1, -6, 3, -3, 0, -15, -11, 0,
    -- filter=69 channel=48
    3, -1, 5, 6, 10, 6, 4, 2, 1,
    -- filter=69 channel=49
    -5, -2, -6, -5, 0, -3, 10, -1, -7,
    -- filter=69 channel=50
    -6, -6, -2, -8, 0, 4, 11, -5, -9,
    -- filter=69 channel=51
    6, -3, 0, 3, -4, 0, -1, -5, 1,
    -- filter=69 channel=52
    1, -2, -2, 4, -7, 4, 8, 3, -2,
    -- filter=69 channel=53
    -6, -2, 3, 0, -8, 6, 6, 1, 0,
    -- filter=69 channel=54
    7, -2, -6, -4, -6, -2, 3, 3, 4,
    -- filter=69 channel=55
    3, -16, 1, -7, -1, -4, 17, 15, 3,
    -- filter=69 channel=56
    -4, -2, 6, -4, -1, 0, 1, -5, 4,
    -- filter=69 channel=57
    -6, -5, 0, 1, -1, 5, 1, 0, 0,
    -- filter=69 channel=58
    -7, 6, 3, -4, -1, -1, -6, 3, 0,
    -- filter=69 channel=59
    9, -2, 1, 0, -4, 4, 6, -3, 3,
    -- filter=69 channel=60
    -6, 7, -3, -6, -3, 5, 5, 1, 3,
    -- filter=69 channel=61
    4, 4, -2, -3, 0, -1, 1, 2, -4,
    -- filter=69 channel=62
    7, -1, 7, 3, 3, -6, 1, 2, -1,
    -- filter=69 channel=63
    -2, 3, -1, 1, -5, 5, -7, -7, -4,
    -- filter=69 channel=64
    5, -6, 0, -1, -7, 3, -6, 6, 3,
    -- filter=69 channel=65
    0, -4, 0, 1, 5, 7, 6, 2, 1,
    -- filter=69 channel=66
    -2, 1, 3, -1, 1, -2, -1, 4, 1,
    -- filter=69 channel=67
    7, -6, 6, -4, 3, 3, 3, -3, 2,
    -- filter=69 channel=68
    3, 3, 2, 0, -3, -3, 0, 6, -2,
    -- filter=69 channel=69
    4, -6, -1, 2, 3, 2, -5, -4, -4,
    -- filter=69 channel=70
    -4, -3, 3, -5, 5, -7, 6, 6, -2,
    -- filter=69 channel=71
    0, -6, 2, -5, -3, 2, 0, 5, -4,
    -- filter=69 channel=72
    1, -5, -1, -8, -5, 3, -4, -6, 2,
    -- filter=69 channel=73
    -12, -2, -3, 0, -2, -4, 6, -2, -7,
    -- filter=69 channel=74
    -12, 9, 1, -2, 0, -6, 6, -7, -5,
    -- filter=69 channel=75
    1, -5, -9, -4, -9, 7, -9, 3, -2,
    -- filter=69 channel=76
    -8, -13, 3, -4, -4, 3, 10, 1, 8,
    -- filter=69 channel=77
    6, -5, 6, -6, -4, -3, -4, 1, -6,
    -- filter=69 channel=78
    -7, 4, -2, -4, 0, 4, 0, -4, -1,
    -- filter=69 channel=79
    -2, -16, 7, -12, -3, 11, 15, 6, -9,
    -- filter=69 channel=80
    12, 0, 7, 2, 0, 1, -2, -6, -1,
    -- filter=69 channel=81
    1, 2, 2, -2, 0, -1, 5, 6, 5,
    -- filter=69 channel=82
    6, 0, 1, 0, 3, -2, -5, -3, 2,
    -- filter=69 channel=83
    1, -1, 6, 9, -3, -2, -3, 2, -6,
    -- filter=69 channel=84
    -6, -8, 5, 0, -4, -5, 9, -4, -3,
    -- filter=69 channel=85
    -1, 4, 5, 0, -4, -6, 0, -6, 0,
    -- filter=69 channel=86
    0, 4, 5, -6, 8, 4, -6, 0, -6,
    -- filter=69 channel=87
    -1, 3, 5, -3, -6, 2, 8, 3, 0,
    -- filter=69 channel=88
    0, 8, 2, -5, 0, 0, 0, 0, 3,
    -- filter=69 channel=89
    -3, -9, 0, -11, 0, 7, 6, 15, -5,
    -- filter=69 channel=90
    2, 4, 3, 2, -4, 0, -6, 1, -5,
    -- filter=69 channel=91
    -7, -9, -2, -4, 5, -5, 4, -5, -9,
    -- filter=69 channel=92
    -1, -6, 1, 4, -1, 2, -4, -4, 2,
    -- filter=69 channel=93
    -1, 12, -4, 7, 9, 0, -3, -1, -1,
    -- filter=69 channel=94
    5, 3, 3, -6, 7, 6, 0, 4, -7,
    -- filter=69 channel=95
    -6, -5, -5, 0, 3, 0, 3, -4, 6,
    -- filter=69 channel=96
    -1, -5, -4, 2, 1, 0, 3, -2, 3,
    -- filter=69 channel=97
    7, 0, -6, -1, -7, -1, -6, -3, -7,
    -- filter=69 channel=98
    -5, -3, 11, -5, 5, 10, 11, -4, -6,
    -- filter=69 channel=99
    3, 2, 7, -7, 8, 7, 13, -1, 1,
    -- filter=69 channel=100
    4, -5, 4, 5, -1, 3, -2, -4, 8,
    -- filter=69 channel=101
    -9, -5, -6, -1, 9, -6, 9, 7, -2,
    -- filter=69 channel=102
    -1, 2, -6, -4, 6, 0, -2, -5, -4,
    -- filter=69 channel=103
    9, -3, -7, 3, 4, 5, -16, -10, -3,
    -- filter=69 channel=104
    1, 2, 9, 6, -2, 4, -3, -3, -5,
    -- filter=69 channel=105
    -7, -4, -2, -13, -5, 0, 0, 6, 7,
    -- filter=69 channel=106
    -2, -4, -1, -6, 0, 6, -5, -2, 0,
    -- filter=69 channel=107
    -2, -6, -1, -2, -3, 3, 7, 3, -6,
    -- filter=69 channel=108
    5, 0, 0, -4, -1, 8, 2, -5, -2,
    -- filter=69 channel=109
    -1, -9, 11, -8, 9, 8, 12, 3, -3,
    -- filter=69 channel=110
    2, 3, -2, -3, -9, 0, -1, -4, 5,
    -- filter=69 channel=111
    -1, 4, 0, 7, -1, -3, 4, 2, 2,
    -- filter=69 channel=112
    3, 4, 8, -4, 9, -8, -2, -7, -7,
    -- filter=69 channel=113
    -5, -7, -5, -10, -4, -1, -6, 5, 4,
    -- filter=69 channel=114
    -8, -15, 2, -15, 4, 0, 12, 6, -9,
    -- filter=69 channel=115
    0, -6, -5, 0, 7, 4, -7, -4, 0,
    -- filter=69 channel=116
    -8, 0, -2, -7, 5, 10, 5, 6, -7,
    -- filter=69 channel=117
    8, 0, -3, 1, 0, -3, 2, -1, 2,
    -- filter=69 channel=118
    -6, -2, -3, 4, 5, 0, 7, 0, -6,
    -- filter=69 channel=119
    -4, 2, 5, 0, 7, -6, 1, -4, 3,
    -- filter=69 channel=120
    -18, -2, 13, 0, 7, 2, 17, 2, -2,
    -- filter=69 channel=121
    8, 0, 5, -5, -7, 2, -2, 6, 4,
    -- filter=69 channel=122
    4, 6, 0, 3, 7, -4, -15, -21, -10,
    -- filter=69 channel=123
    3, 1, -1, 1, 3, 5, -5, 5, -2,
    -- filter=69 channel=124
    -6, -3, 2, -9, -5, -4, 2, 9, -4,
    -- filter=69 channel=125
    2, -4, 0, 2, 1, 4, 11, -3, 1,
    -- filter=69 channel=126
    -2, -3, 2, -7, -6, 2, 0, 13, 3,
    -- filter=69 channel=127
    9, 0, 2, -6, 4, 8, -5, 6, 0,
    -- filter=70 channel=0
    0, -1, 6, -4, 9, 5, -1, 3, -1,
    -- filter=70 channel=1
    -4, -7, 5, 0, 6, 3, 9, 8, -5,
    -- filter=70 channel=2
    -4, 6, 1, -6, -2, 0, 5, 0, 4,
    -- filter=70 channel=3
    8, -5, 5, 8, 3, 11, 4, -6, 2,
    -- filter=70 channel=4
    4, -5, -6, -4, 0, -2, 4, -1, 7,
    -- filter=70 channel=5
    0, -3, -3, 0, 2, -2, -3, -4, 2,
    -- filter=70 channel=6
    -4, 3, -6, 2, 0, 2, -2, 2, 0,
    -- filter=70 channel=7
    1, 5, -3, 0, -7, 4, 0, 5, 3,
    -- filter=70 channel=8
    1, 1, 5, -5, -4, -4, -4, -3, 4,
    -- filter=70 channel=9
    -3, 0, -1, -2, 2, 4, -4, -6, -3,
    -- filter=70 channel=10
    6, -4, 0, -5, -2, 3, -5, 3, -2,
    -- filter=70 channel=11
    3, -1, 2, -1, 0, -1, -1, 1, 1,
    -- filter=70 channel=12
    3, 5, -8, 2, -7, 0, -1, 7, 2,
    -- filter=70 channel=13
    -2, -5, 1, 4, -1, 1, 0, 0, -5,
    -- filter=70 channel=14
    5, 3, -2, 2, 2, 2, -2, -2, 0,
    -- filter=70 channel=15
    2, 6, 4, -4, -1, -4, -6, 0, -2,
    -- filter=70 channel=16
    -7, -2, 7, 4, 2, 0, 2, -2, 0,
    -- filter=70 channel=17
    -4, -4, 4, 3, 0, 3, 5, -3, 5,
    -- filter=70 channel=18
    -7, 5, -8, 0, -7, -2, 5, -5, -3,
    -- filter=70 channel=19
    -4, -5, 0, -3, 0, 4, -7, -4, -6,
    -- filter=70 channel=20
    -3, 0, -8, -3, 0, -6, 2, 3, 7,
    -- filter=70 channel=21
    0, 0, 4, 3, -5, -5, 1, 5, 5,
    -- filter=70 channel=22
    4, -5, -3, 0, -5, -2, -4, 1, 5,
    -- filter=70 channel=23
    0, 1, 5, -1, 2, 3, -3, -4, -7,
    -- filter=70 channel=24
    3, -4, 0, 0, -5, 6, -6, 2, -4,
    -- filter=70 channel=25
    3, -6, 5, 6, -5, 1, -8, -1, -5,
    -- filter=70 channel=26
    0, 2, 4, 1, 3, 0, 7, -4, 6,
    -- filter=70 channel=27
    -6, -8, -2, 0, -7, -6, 0, 1, 4,
    -- filter=70 channel=28
    0, -1, 1, 6, -5, -2, -1, 1, -4,
    -- filter=70 channel=29
    -2, -7, -4, -4, 4, 1, -3, -4, 6,
    -- filter=70 channel=30
    -1, -7, -2, 4, 6, -4, 0, 3, 0,
    -- filter=70 channel=31
    0, 6, -2, 0, -7, -5, -3, 5, -5,
    -- filter=70 channel=32
    -1, 1, -2, 0, 0, 4, 0, 0, -4,
    -- filter=70 channel=33
    -2, 1, 5, 0, 5, -5, 0, -5, -1,
    -- filter=70 channel=34
    -4, 0, 1, -2, 1, 5, -3, 7, 0,
    -- filter=70 channel=35
    0, 0, 1, -6, -6, -6, 4, -4, -4,
    -- filter=70 channel=36
    0, 5, 4, -4, 5, -6, 0, -3, -4,
    -- filter=70 channel=37
    -6, 3, 0, 4, 7, -2, 0, 7, 0,
    -- filter=70 channel=38
    -2, -6, -5, 0, 6, -1, -3, -6, 2,
    -- filter=70 channel=39
    6, 6, 6, 0, -5, 5, -2, -3, -4,
    -- filter=70 channel=40
    -6, 7, 3, 0, 7, 3, 0, 6, -1,
    -- filter=70 channel=41
    0, 8, 0, -4, 8, -9, 6, 10, -6,
    -- filter=70 channel=42
    1, -3, -3, -2, 6, 6, -2, 3, 5,
    -- filter=70 channel=43
    -1, 3, 5, 0, 2, 1, -2, -3, 5,
    -- filter=70 channel=44
    -8, 0, -4, 5, 5, 7, -2, 0, -6,
    -- filter=70 channel=45
    0, 0, -4, -3, -4, 4, 6, 7, -5,
    -- filter=70 channel=46
    -4, -2, -2, 0, 6, 4, -1, 6, 3,
    -- filter=70 channel=47
    2, 0, 2, 2, 6, 3, -1, -1, -3,
    -- filter=70 channel=48
    5, 1, -8, 6, -7, -7, 0, 5, -1,
    -- filter=70 channel=49
    -3, -1, -3, -4, -6, -3, 3, 4, 6,
    -- filter=70 channel=50
    4, 6, -6, 0, -8, -7, -7, 2, -1,
    -- filter=70 channel=51
    -7, 6, -3, -7, -5, 2, 1, 4, -4,
    -- filter=70 channel=52
    -5, 1, -3, 1, 4, -4, -2, -6, 2,
    -- filter=70 channel=53
    0, 2, -4, 2, 0, 2, 0, -7, 0,
    -- filter=70 channel=54
    4, -4, -2, 0, 7, -5, 0, -2, -5,
    -- filter=70 channel=55
    3, -1, 0, -4, 1, 1, -1, 2, -5,
    -- filter=70 channel=56
    3, 0, -4, 1, -6, 2, 0, -3, 6,
    -- filter=70 channel=57
    -5, 4, 3, 5, 2, -4, 3, 2, 2,
    -- filter=70 channel=58
    3, -3, 4, -6, -1, 5, 6, 0, -5,
    -- filter=70 channel=59
    -5, 6, -3, -5, 5, -6, -4, 4, 4,
    -- filter=70 channel=60
    -7, 4, -6, 2, -5, -2, -4, 2, 4,
    -- filter=70 channel=61
    -1, 6, 3, 5, 1, -4, -2, 2, -2,
    -- filter=70 channel=62
    1, 2, -2, 0, -1, 0, -3, 4, 6,
    -- filter=70 channel=63
    2, 2, -4, -3, 0, 0, -3, -5, -6,
    -- filter=70 channel=64
    5, -4, -4, 0, -5, 3, 7, -2, -6,
    -- filter=70 channel=65
    5, -5, -3, 7, -5, 4, -2, 7, 6,
    -- filter=70 channel=66
    0, 6, -6, 1, -3, -6, -3, -5, -6,
    -- filter=70 channel=67
    -6, 1, 5, -5, 0, 6, 6, -4, -1,
    -- filter=70 channel=68
    2, -3, 0, -5, -5, 0, 0, 3, -2,
    -- filter=70 channel=69
    4, 1, -2, -4, -4, -3, -1, 1, 2,
    -- filter=70 channel=70
    3, -2, 5, 2, -9, 0, -3, 0, 0,
    -- filter=70 channel=71
    2, 4, 0, -4, 0, 5, -2, 4, -2,
    -- filter=70 channel=72
    4, 2, -1, -5, -5, 0, 4, 1, 5,
    -- filter=70 channel=73
    -7, -3, 2, 5, -4, -4, 1, 6, 5,
    -- filter=70 channel=74
    7, -3, 7, 0, 0, -2, 0, -3, 0,
    -- filter=70 channel=75
    -1, 1, 6, 4, 10, -1, 8, 0, -1,
    -- filter=70 channel=76
    5, 2, -6, 5, -5, -5, 4, -1, -1,
    -- filter=70 channel=77
    5, 6, -7, 5, -3, -1, 0, 1, 1,
    -- filter=70 channel=78
    -6, -2, 4, 2, -3, 8, 6, -7, 4,
    -- filter=70 channel=79
    -5, 5, -7, -6, -3, -7, -8, 1, 6,
    -- filter=70 channel=80
    0, 0, 3, 0, -1, -8, -2, -6, 1,
    -- filter=70 channel=81
    -6, 5, -2, 7, -1, 2, -6, 6, 5,
    -- filter=70 channel=82
    -3, -5, 2, 1, 3, 6, -1, -1, 7,
    -- filter=70 channel=83
    -3, 0, -1, 1, 3, -5, -1, -4, 1,
    -- filter=70 channel=84
    -6, -3, 1, -6, -6, 6, 5, 2, -2,
    -- filter=70 channel=85
    -6, -3, 0, -3, -5, 4, -4, -3, -3,
    -- filter=70 channel=86
    2, -3, 2, -2, 1, 6, 0, -4, 0,
    -- filter=70 channel=87
    0, -6, -5, -7, 2, 1, 1, -4, 0,
    -- filter=70 channel=88
    -1, 6, 1, 1, -1, 0, -3, -1, 0,
    -- filter=70 channel=89
    -6, 4, 3, 6, -1, 0, 0, -8, 6,
    -- filter=70 channel=90
    1, 3, -4, -1, -3, 2, 0, -5, 5,
    -- filter=70 channel=91
    -2, -1, -2, -6, 0, -2, -3, -5, 4,
    -- filter=70 channel=92
    7, 3, 5, 0, -4, 6, 7, 0, -7,
    -- filter=70 channel=93
    -4, -2, -1, 0, 3, 1, 8, -4, 8,
    -- filter=70 channel=94
    1, 0, -4, 4, -1, -4, 7, -5, -6,
    -- filter=70 channel=95
    -2, 2, -2, -4, -5, 2, -4, 3, 0,
    -- filter=70 channel=96
    -4, 7, 0, 3, 6, 0, 4, 4, 7,
    -- filter=70 channel=97
    1, 4, 4, -6, 2, 0, 2, -3, 0,
    -- filter=70 channel=98
    -1, 3, 6, -3, -4, -2, -6, 4, 7,
    -- filter=70 channel=99
    -2, 7, 6, -3, -2, -5, -1, -4, 6,
    -- filter=70 channel=100
    3, 4, -6, -3, -4, -4, 5, 4, 5,
    -- filter=70 channel=101
    -7, -3, 3, -5, 0, 0, 8, -2, 5,
    -- filter=70 channel=102
    3, 2, 3, -5, 4, 6, 0, 1, -1,
    -- filter=70 channel=103
    2, 6, 0, 0, 8, -5, 1, 0, -5,
    -- filter=70 channel=104
    1, 0, 2, -4, -2, -7, -5, -7, 0,
    -- filter=70 channel=105
    0, 0, -6, 1, 4, 3, 5, 5, 4,
    -- filter=70 channel=106
    -3, 4, 2, 0, -6, -5, 0, -4, 2,
    -- filter=70 channel=107
    1, -2, -2, 3, -5, 5, 0, 3, 2,
    -- filter=70 channel=108
    7, -4, 1, -6, -4, -1, -6, 2, 5,
    -- filter=70 channel=109
    -8, 1, 3, -2, -1, -9, -8, -6, 8,
    -- filter=70 channel=110
    4, -1, -5, -1, -5, -6, -1, -5, 2,
    -- filter=70 channel=111
    -1, -6, 3, 7, 0, -3, 5, 7, -6,
    -- filter=70 channel=112
    0, -1, -6, -1, -7, 0, 5, 6, -3,
    -- filter=70 channel=113
    -4, 8, -2, -6, 6, 1, 2, -4, 2,
    -- filter=70 channel=114
    -4, -5, 0, 7, -7, 6, -2, -4, -1,
    -- filter=70 channel=115
    -3, -1, 5, 1, 1, -6, -7, 7, -1,
    -- filter=70 channel=116
    1, 4, 6, 4, -1, -4, 5, 6, 10,
    -- filter=70 channel=117
    1, 0, -5, -6, 2, 6, 5, 5, 0,
    -- filter=70 channel=118
    0, -1, -3, 0, -6, 5, 5, -5, 0,
    -- filter=70 channel=119
    0, 4, 1, 2, -6, -8, 3, 5, 1,
    -- filter=70 channel=120
    1, 2, -2, 6, -6, 0, 1, 10, 10,
    -- filter=70 channel=121
    6, 6, -3, -4, 2, -3, -7, -7, -4,
    -- filter=70 channel=122
    -5, 2, 1, -3, 8, 4, -1, -6, -4,
    -- filter=70 channel=123
    1, 3, 7, -3, 1, -1, 0, -3, 0,
    -- filter=70 channel=124
    3, -7, 5, 0, 3, -5, 1, -7, 6,
    -- filter=70 channel=125
    1, 2, -3, -1, 4, -7, -1, 3, -4,
    -- filter=70 channel=126
    2, 1, 4, 5, -5, 0, -4, -5, 3,
    -- filter=70 channel=127
    3, 5, 5, 2, 5, 0, -4, -2, 2,
    -- filter=71 channel=0
    1, 0, 7, 6, -4, -5, 2, -5, 0,
    -- filter=71 channel=1
    4, 7, 4, -1, -6, -4, 2, 4, -5,
    -- filter=71 channel=2
    -1, 3, 6, -5, 0, 0, -4, -5, 0,
    -- filter=71 channel=3
    7, -1, -4, -3, 5, -4, 0, -6, 3,
    -- filter=71 channel=4
    -2, 4, -1, 1, 0, 4, 0, 8, -6,
    -- filter=71 channel=5
    0, -5, -6, 2, -6, -5, 6, 2, 3,
    -- filter=71 channel=6
    -7, 0, -2, 0, -7, 1, 6, -1, -4,
    -- filter=71 channel=7
    -2, -5, -2, 6, -4, -5, -7, 3, -6,
    -- filter=71 channel=8
    4, 5, 1, 2, 0, -4, 4, -4, -3,
    -- filter=71 channel=9
    6, -1, -6, 5, 3, 0, 5, 1, -6,
    -- filter=71 channel=10
    7, 0, 6, 4, -7, 1, -7, -2, 0,
    -- filter=71 channel=11
    6, -3, 5, -2, 2, 0, 0, -2, 0,
    -- filter=71 channel=12
    -6, 5, -3, -5, -6, -3, -7, 6, -1,
    -- filter=71 channel=13
    3, 4, -3, 0, 4, 2, -5, -5, -4,
    -- filter=71 channel=14
    1, 0, 4, 1, -3, 1, -5, 4, 0,
    -- filter=71 channel=15
    3, 6, -2, 3, -4, -1, 4, -3, 2,
    -- filter=71 channel=16
    6, -3, -6, -6, 0, 0, 0, -2, -4,
    -- filter=71 channel=17
    1, 3, -2, -6, 0, -2, -5, 0, -4,
    -- filter=71 channel=18
    7, -4, -2, -5, 1, 1, 6, 0, -3,
    -- filter=71 channel=19
    -2, 3, -6, -2, 0, -4, 1, -5, 5,
    -- filter=71 channel=20
    0, 3, 2, -6, 0, -7, 2, 6, -1,
    -- filter=71 channel=21
    -6, 4, 4, -5, 0, -4, 7, 4, 2,
    -- filter=71 channel=22
    -5, 0, -3, 3, 1, 0, -2, -4, -7,
    -- filter=71 channel=23
    5, 5, 2, -5, -6, -1, -1, 6, -2,
    -- filter=71 channel=24
    5, 4, -4, -3, 2, -5, -5, 3, 5,
    -- filter=71 channel=25
    4, 2, 6, 4, 4, -1, -5, 1, -4,
    -- filter=71 channel=26
    0, -4, 4, -5, -4, -4, 4, 2, 7,
    -- filter=71 channel=27
    -2, 1, -5, -7, -8, 2, -4, 5, 1,
    -- filter=71 channel=28
    5, -2, 0, 1, 3, -4, 1, 2, 0,
    -- filter=71 channel=29
    4, 2, 3, -6, -7, 0, 0, -4, 2,
    -- filter=71 channel=30
    -3, 6, 0, -6, -2, 6, 2, 7, 6,
    -- filter=71 channel=31
    0, -7, 0, 1, -6, 5, 0, 5, 1,
    -- filter=71 channel=32
    -6, 0, 3, -1, 2, -5, 2, -1, 0,
    -- filter=71 channel=33
    6, 4, 3, 0, -4, -5, -7, -4, -2,
    -- filter=71 channel=34
    4, -3, -6, -1, -4, -3, 4, -2, 5,
    -- filter=71 channel=35
    5, -2, 2, 0, 1, -6, 0, -4, 2,
    -- filter=71 channel=36
    -6, 1, 7, -3, 0, -2, -3, 0, 1,
    -- filter=71 channel=37
    0, -6, 3, -6, -7, 5, 4, -4, -5,
    -- filter=71 channel=38
    -4, -2, 4, -6, -4, -6, 2, -5, 0,
    -- filter=71 channel=39
    5, 7, 0, 2, 2, -4, 0, -6, 4,
    -- filter=71 channel=40
    -1, 7, -2, -3, -6, -3, -6, -3, 3,
    -- filter=71 channel=41
    6, -3, 3, 2, -2, 4, 1, -8, -1,
    -- filter=71 channel=42
    3, 1, 7, -3, 1, 0, -6, 5, -6,
    -- filter=71 channel=43
    -7, 5, 4, 6, 1, 2, -3, -2, 1,
    -- filter=71 channel=44
    4, 2, -1, -1, 2, 4, -1, 0, -4,
    -- filter=71 channel=45
    0, -3, 5, -1, 2, 3, 5, 0, 4,
    -- filter=71 channel=46
    1, 3, 6, 6, 4, -1, 0, 3, 0,
    -- filter=71 channel=47
    6, 7, 7, -1, 0, 0, -5, -2, -6,
    -- filter=71 channel=48
    -2, -3, -3, -3, 0, -4, 7, 1, -4,
    -- filter=71 channel=49
    -6, 2, -5, -6, -3, 0, 0, 3, -6,
    -- filter=71 channel=50
    -5, -3, -2, 6, 4, -2, -3, -1, 0,
    -- filter=71 channel=51
    2, 5, -2, 6, 1, 1, 6, 4, -4,
    -- filter=71 channel=52
    -6, -6, -1, -6, -3, -3, 1, 6, -4,
    -- filter=71 channel=53
    5, -5, 3, -4, 0, 0, -1, -5, 4,
    -- filter=71 channel=54
    -6, 3, 3, 7, -6, 3, 6, 0, 4,
    -- filter=71 channel=55
    5, 1, -5, 1, -3, -1, -1, 2, -7,
    -- filter=71 channel=56
    -5, -2, -1, -2, 0, -7, 0, 1, 3,
    -- filter=71 channel=57
    -6, -7, -6, 5, 0, 6, -1, -4, 7,
    -- filter=71 channel=58
    -7, 0, 7, 2, -4, 3, -5, 2, 5,
    -- filter=71 channel=59
    7, 1, 6, 4, 6, -6, -2, -4, -6,
    -- filter=71 channel=60
    7, 7, -3, 4, 4, -1, 5, 1, -4,
    -- filter=71 channel=61
    3, 5, 5, -5, 0, 4, 5, -3, 6,
    -- filter=71 channel=62
    5, 3, -5, 0, 7, -5, -2, 2, 1,
    -- filter=71 channel=63
    4, 4, 3, 6, 6, -2, 2, 3, 0,
    -- filter=71 channel=64
    2, -1, -4, 5, -4, 3, -1, 0, 3,
    -- filter=71 channel=65
    -7, 3, 5, 1, -2, 1, 0, 5, -4,
    -- filter=71 channel=66
    3, 5, 5, 4, -2, -2, -3, 6, -2,
    -- filter=71 channel=67
    -5, 6, -1, 5, 5, 7, 0, -7, -1,
    -- filter=71 channel=68
    5, -6, 3, 0, 0, 3, -1, 0, -1,
    -- filter=71 channel=69
    -5, -5, -2, -4, -5, -7, -4, -3, -7,
    -- filter=71 channel=70
    -5, 3, 1, -3, 0, -3, -5, 6, -1,
    -- filter=71 channel=71
    5, 7, -4, -3, 0, 5, 3, -2, -4,
    -- filter=71 channel=72
    0, -3, 1, -3, 5, -2, -6, -4, -3,
    -- filter=71 channel=73
    -3, 0, -2, -2, -1, -5, -6, -7, 2,
    -- filter=71 channel=74
    3, -2, 2, -2, 1, 6, 6, 3, -5,
    -- filter=71 channel=75
    -1, 0, -2, 3, 3, 0, 2, -5, -6,
    -- filter=71 channel=76
    -5, 0, 0, -2, 6, 1, -1, -1, 3,
    -- filter=71 channel=77
    -3, -3, 0, 2, 5, 0, 5, -6, -3,
    -- filter=71 channel=78
    2, 0, 6, -3, 0, 4, -1, -2, -5,
    -- filter=71 channel=79
    2, -5, -1, -3, -2, -2, -2, 3, 0,
    -- filter=71 channel=80
    -3, 4, 0, -6, 5, -3, -1, 1, -4,
    -- filter=71 channel=81
    -4, 1, 2, 5, -6, -4, 0, 3, 4,
    -- filter=71 channel=82
    5, -3, 3, -3, -6, 1, -1, 1, -2,
    -- filter=71 channel=83
    0, 0, -5, -3, -4, -6, 1, -5, 1,
    -- filter=71 channel=84
    -3, -2, -7, -1, -7, -4, 7, -4, -5,
    -- filter=71 channel=85
    6, -4, 0, -7, 0, -3, -1, 0, 6,
    -- filter=71 channel=86
    0, -2, 2, -6, -4, 0, 6, -7, -1,
    -- filter=71 channel=87
    -4, 0, 0, -6, 6, -6, 5, 7, 0,
    -- filter=71 channel=88
    -2, 1, -1, -7, 0, -7, 1, 1, 1,
    -- filter=71 channel=89
    -4, -7, -8, -6, 5, 0, -4, 5, -5,
    -- filter=71 channel=90
    -7, 2, 7, 0, -2, 1, 3, 1, -1,
    -- filter=71 channel=91
    -4, -6, -2, 3, 6, -5, -2, 5, -2,
    -- filter=71 channel=92
    -6, 0, 5, 6, 2, -1, -5, -2, 0,
    -- filter=71 channel=93
    -5, -7, -3, -6, 7, 1, 4, -2, -7,
    -- filter=71 channel=94
    -6, 3, 2, 4, -1, -6, 0, -2, 1,
    -- filter=71 channel=95
    -5, -5, 4, 5, -1, 3, 1, -1, -4,
    -- filter=71 channel=96
    0, 0, -3, 2, 5, 1, -1, -4, -1,
    -- filter=71 channel=97
    5, 4, -6, -3, 5, -3, 1, 3, 5,
    -- filter=71 channel=98
    4, 4, 0, -7, 5, -1, 5, -4, 2,
    -- filter=71 channel=99
    2, -2, 2, 0, -7, -6, 2, 6, -6,
    -- filter=71 channel=100
    -6, -5, 4, 4, 2, 1, -1, 3, 2,
    -- filter=71 channel=101
    6, -2, 1, -2, -5, -6, 5, 0, 2,
    -- filter=71 channel=102
    -1, 0, -2, -1, -1, -2, 2, -5, 4,
    -- filter=71 channel=103
    0, 0, -3, 1, 5, 4, -1, 3, -3,
    -- filter=71 channel=104
    -4, 3, 4, -1, -5, 0, 4, 5, -1,
    -- filter=71 channel=105
    6, 6, 0, 5, -5, -6, -3, -4, 1,
    -- filter=71 channel=106
    3, -3, 7, 3, 5, -6, 6, -2, 1,
    -- filter=71 channel=107
    -1, 6, -6, 0, -2, -4, -4, 5, 3,
    -- filter=71 channel=108
    0, 2, 0, -5, -5, -1, -1, 1, -7,
    -- filter=71 channel=109
    -3, 1, 3, -6, 0, 0, 0, -3, -4,
    -- filter=71 channel=110
    1, 5, -7, 6, -5, -4, 2, 0, -6,
    -- filter=71 channel=111
    -4, 5, 0, 4, 2, -2, 5, 2, 2,
    -- filter=71 channel=112
    0, 6, 3, -1, 3, -2, -2, -3, 0,
    -- filter=71 channel=113
    -2, 6, 1, 0, -3, 4, 5, 6, 0,
    -- filter=71 channel=114
    2, 5, 0, -7, -1, 2, -3, -1, 0,
    -- filter=71 channel=115
    -5, 3, 5, -3, 0, -3, -4, -3, 6,
    -- filter=71 channel=116
    4, -5, 3, -4, 2, 4, 2, -3, 6,
    -- filter=71 channel=117
    -4, 0, -3, -3, 0, -2, 4, 0, 4,
    -- filter=71 channel=118
    7, -6, -5, -1, 0, -2, -3, -2, -2,
    -- filter=71 channel=119
    0, 7, -2, 5, 3, -3, 5, 4, 6,
    -- filter=71 channel=120
    -5, -8, -7, -3, -5, 2, 2, 5, -4,
    -- filter=71 channel=121
    1, -3, -3, -4, -5, 5, -4, 2, 1,
    -- filter=71 channel=122
    -6, 1, -6, 0, 1, 0, 1, -4, -1,
    -- filter=71 channel=123
    0, 3, 3, 6, 2, -3, -4, -2, -3,
    -- filter=71 channel=124
    2, -1, 5, 1, 5, 6, 0, 0, 6,
    -- filter=71 channel=125
    -3, -2, 1, -7, -5, -1, 1, 0, -1,
    -- filter=71 channel=126
    5, -6, 4, 4, -1, 3, 2, 0, -3,
    -- filter=71 channel=127
    0, -4, 5, 0, -3, -4, 4, 2, -5,
    -- filter=72 channel=0
    0, 6, -6, 3, 6, 4, 3, -5, -2,
    -- filter=72 channel=1
    -4, 0, 4, 9, -13, -11, 8, 22, 0,
    -- filter=72 channel=2
    0, 12, 6, 4, -5, -9, -2, 13, -3,
    -- filter=72 channel=3
    24, 14, -8, 12, 48, 18, 17, -1, -1,
    -- filter=72 channel=4
    13, 33, 18, 23, 10, -3, 19, 51, 4,
    -- filter=72 channel=5
    8, -1, -14, 1, 6, 8, -6, -13, 1,
    -- filter=72 channel=6
    2, 2, 4, 5, -2, 0, 6, 0, 5,
    -- filter=72 channel=7
    5, -1, 2, 0, 4, 0, 3, 0, -3,
    -- filter=72 channel=8
    3, -4, -7, 2, 5, 7, -1, 0, -1,
    -- filter=72 channel=9
    2, 15, 6, -10, -5, 0, 2, 7, 0,
    -- filter=72 channel=10
    5, 10, 4, -6, -10, 9, 6, -11, -9,
    -- filter=72 channel=11
    2, 3, 4, -9, 2, -1, -4, 1, -9,
    -- filter=72 channel=12
    2, -7, 10, 5, -9, -3, -11, 0, 10,
    -- filter=72 channel=13
    3, 16, 0, -11, -29, -1, 11, 9, -1,
    -- filter=72 channel=14
    -2, -4, -3, 6, 4, 0, -2, 3, 0,
    -- filter=72 channel=15
    1, 5, -1, -15, -14, 13, 6, 0, -13,
    -- filter=72 channel=16
    2, 6, 3, -1, -4, 9, 8, -5, 0,
    -- filter=72 channel=17
    -7, -5, 0, -1, 1, -5, -3, 0, 1,
    -- filter=72 channel=18
    -6, 3, 2, -5, -37, -2, 4, 5, -3,
    -- filter=72 channel=19
    0, -3, -7, 2, -2, 4, -5, 0, 1,
    -- filter=72 channel=20
    -3, 2, -10, -4, -3, 7, 0, -7, 3,
    -- filter=72 channel=21
    -5, 4, 1, -18, -18, 6, 11, -5, -10,
    -- filter=72 channel=22
    9, 1, -8, -9, 5, 15, 3, -11, -4,
    -- filter=72 channel=23
    28, 18, -19, -41, 6, 21, 38, -25, -2,
    -- filter=72 channel=24
    4, -5, 0, 1, 0, 1, 7, -4, 5,
    -- filter=72 channel=25
    1, 25, 3, -21, -46, 1, 21, 15, -15,
    -- filter=72 channel=26
    4, 0, -6, 8, -10, -6, -3, 12, -3,
    -- filter=72 channel=27
    6, 18, -6, -51, -47, 13, 38, 16, -13,
    -- filter=72 channel=28
    6, -4, -3, 0, 4, -7, 4, 0, -5,
    -- filter=72 channel=29
    -7, -2, 0, 8, -1, 12, -5, 2, 2,
    -- filter=72 channel=30
    3, 6, 6, -19, -27, 1, 21, 20, -2,
    -- filter=72 channel=31
    17, 30, -2, -42, -29, 19, 27, -11, -11,
    -- filter=72 channel=32
    0, 23, 4, -19, -26, 13, 25, 3, -10,
    -- filter=72 channel=33
    6, 16, -4, -22, -12, 17, 15, -5, -15,
    -- filter=72 channel=34
    24, -10, -10, -24, 16, 12, -2, -22, 0,
    -- filter=72 channel=35
    -5, 4, -2, -6, 4, 1, -3, -3, -1,
    -- filter=72 channel=36
    2, 1, 11, -3, -19, -12, 9, 1, 0,
    -- filter=72 channel=37
    -3, -2, 0, 4, -15, 3, 0, 9, -1,
    -- filter=72 channel=38
    15, 13, -10, -12, -12, 10, 16, -4, -4,
    -- filter=72 channel=39
    2, 6, -6, -3, -7, 3, -4, 5, -3,
    -- filter=72 channel=40
    -7, 0, -11, 0, 3, 7, -2, -5, -6,
    -- filter=72 channel=41
    -18, 2, 8, 37, -33, -19, 1, 26, -12,
    -- filter=72 channel=42
    -7, -2, 0, -10, -2, -8, 3, 0, -6,
    -- filter=72 channel=43
    8, 2, -9, 3, 23, 9, 2, -11, -5,
    -- filter=72 channel=44
    10, 7, -1, -18, -9, 4, 0, -2, 5,
    -- filter=72 channel=45
    5, -1, 2, -1, -2, -2, 6, 1, -6,
    -- filter=72 channel=46
    -2, -3, -1, 10, 4, -10, 0, 6, 2,
    -- filter=72 channel=47
    4, 11, -4, -20, -16, 4, 14, 2, 2,
    -- filter=72 channel=48
    3, 15, 10, -24, -44, -7, 22, 26, -3,
    -- filter=72 channel=49
    -14, 13, 8, 2, -21, -8, 15, 25, -1,
    -- filter=72 channel=50
    9, 17, -2, -31, -15, 7, 9, -2, -3,
    -- filter=72 channel=51
    0, -6, 0, -6, -2, -1, -5, -1, 6,
    -- filter=72 channel=52
    4, 6, -8, -5, 7, 5, 1, -12, 0,
    -- filter=72 channel=53
    0, 2, 3, 0, -9, 2, 4, 5, -4,
    -- filter=72 channel=54
    -5, 4, 4, 4, 7, -6, 2, 5, 2,
    -- filter=72 channel=55
    -3, 13, 7, -17, -22, 15, 7, -8, -6,
    -- filter=72 channel=56
    9, 0, -6, -18, -2, 2, -4, -10, -1,
    -- filter=72 channel=57
    -5, 8, 12, 20, 1, -3, 9, 9, 0,
    -- filter=72 channel=58
    9, -7, -3, 0, 6, -4, 7, -2, -3,
    -- filter=72 channel=59
    -2, 15, 11, -18, -34, 1, 9, 6, -13,
    -- filter=72 channel=60
    -5, -7, -7, 4, 0, -4, -3, 2, 0,
    -- filter=72 channel=61
    6, 0, 6, 0, 0, -6, 8, -2, -2,
    -- filter=72 channel=62
    4, -5, -2, -4, 8, 4, -1, -7, 5,
    -- filter=72 channel=63
    -2, -3, -5, -6, 5, -4, -9, 4, 7,
    -- filter=72 channel=64
    -8, 9, -3, 1, -8, 6, -4, -5, 3,
    -- filter=72 channel=65
    -7, 0, 3, 0, -1, 2, -3, 0, -3,
    -- filter=72 channel=66
    -8, -1, 4, 13, -22, -5, -1, 1, -2,
    -- filter=72 channel=67
    0, 3, -1, -1, 1, -1, -2, 4, -3,
    -- filter=72 channel=68
    -5, 5, 5, 0, -11, -2, 5, 13, -5,
    -- filter=72 channel=69
    -2, 0, -3, -3, 0, 2, -8, -4, 5,
    -- filter=72 channel=70
    2, 10, -10, -17, -12, 18, 9, 3, -9,
    -- filter=72 channel=71
    10, 4, -3, 3, 12, 13, 2, -15, 0,
    -- filter=72 channel=72
    -4, 14, 2, -26, -30, 0, 20, 0, 0,
    -- filter=72 channel=73
    -2, 11, 15, -8, -16, -7, 4, 17, 8,
    -- filter=72 channel=74
    6, 7, -8, -22, -10, 13, 8, -12, -14,
    -- filter=72 channel=75
    10, 5, -21, -8, -4, 10, 7, -10, -13,
    -- filter=72 channel=76
    1, 4, 0, -6, -5, -1, 0, -11, -10,
    -- filter=72 channel=77
    0, -7, -5, 2, -1, 5, 2, 6, 6,
    -- filter=72 channel=78
    2, 3, 1, -7, -2, -5, -5, -9, 7,
    -- filter=72 channel=79
    -5, 22, -10, -29, -28, 13, 24, 5, -15,
    -- filter=72 channel=80
    6, 33, 13, -38, -47, 0, 27, 12, -15,
    -- filter=72 channel=81
    -4, 1, 2, 4, 6, 1, -5, 1, -6,
    -- filter=72 channel=82
    5, -4, -6, 0, 9, 5, 5, -10, 0,
    -- filter=72 channel=83
    -2, 5, 8, -1, -18, 0, 4, 13, -3,
    -- filter=72 channel=84
    -8, 8, -1, -8, -30, -3, 13, 19, 2,
    -- filter=72 channel=85
    -1, 3, 4, -1, -3, 1, 6, 4, 5,
    -- filter=72 channel=86
    4, 5, -11, 2, 1, 10, 4, -12, 0,
    -- filter=72 channel=87
    11, 0, -1, -11, 7, -1, 5, -5, 0,
    -- filter=72 channel=88
    2, 6, 5, -12, -12, -4, -4, -8, 1,
    -- filter=72 channel=89
    3, 13, 0, -28, -19, 6, 16, -3, -4,
    -- filter=72 channel=90
    17, 3, -8, -9, 18, 13, -5, -24, 3,
    -- filter=72 channel=91
    -6, 21, 8, -19, -40, 6, 26, 24, -5,
    -- filter=72 channel=92
    6, -3, 0, 2, 18, -1, 6, -5, 1,
    -- filter=72 channel=93
    -2, 9, 7, -6, -30, -9, 4, 22, 5,
    -- filter=72 channel=94
    -1, -2, -1, 1, 3, 5, 5, -4, -4,
    -- filter=72 channel=95
    10, -1, 3, 5, 5, 0, 4, -3, 0,
    -- filter=72 channel=96
    4, 3, 4, -6, -12, -1, -3, -3, 2,
    -- filter=72 channel=97
    13, 1, -2, 3, 21, 4, 7, -8, 0,
    -- filter=72 channel=98
    13, 19, 4, -27, -23, 0, 20, 1, -12,
    -- filter=72 channel=99
    19, 24, -4, -29, -10, 5, 16, -13, -11,
    -- filter=72 channel=100
    -2, -9, 6, 1, 2, -6, 1, 2, 1,
    -- filter=72 channel=101
    6, 23, 7, 25, 16, 0, 9, 22, 1,
    -- filter=72 channel=102
    5, 0, 5, 4, 3, -6, 0, -7, -1,
    -- filter=72 channel=103
    3, 11, 0, -13, 7, 13, 3, -15, 2,
    -- filter=72 channel=104
    6, 10, 7, -12, -35, 4, 17, 8, -4,
    -- filter=72 channel=105
    -2, 0, 1, 9, 9, 6, -6, 2, -3,
    -- filter=72 channel=106
    1, -4, -5, -4, 4, 0, 0, 5, 4,
    -- filter=72 channel=107
    12, -4, -13, -1, 12, 2, -2, 2, -2,
    -- filter=72 channel=108
    -9, 0, -4, 11, 0, 0, -1, 10, -5,
    -- filter=72 channel=109
    2, 23, 0, -32, -47, -3, 21, 12, -7,
    -- filter=72 channel=110
    0, 10, -5, -10, -5, 14, 15, -8, 1,
    -- filter=72 channel=111
    -6, 7, 2, 7, -2, -2, 2, 6, -2,
    -- filter=72 channel=112
    8, 9, -4, -26, 4, 2, 7, -10, -11,
    -- filter=72 channel=113
    18, 13, -12, -26, 7, 8, 12, -11, -3,
    -- filter=72 channel=114
    -2, 9, 2, -5, -37, 3, 20, 24, 6,
    -- filter=72 channel=115
    0, -2, -4, -4, 0, 0, 5, 0, -5,
    -- filter=72 channel=116
    -10, 35, 18, -8, -49, -8, 23, 21, 2,
    -- filter=72 channel=117
    -4, 6, 3, -10, -10, 4, 12, 11, -1,
    -- filter=72 channel=118
    4, 5, 4, 4, -8, -3, 6, -6, 2,
    -- filter=72 channel=119
    2, -8, -9, -26, 0, 0, -6, -19, 6,
    -- filter=72 channel=120
    2, 3, 0, -27, -17, 6, 9, 3, 1,
    -- filter=72 channel=121
    -3, 2, 0, 0, -6, -4, 7, -3, -6,
    -- filter=72 channel=122
    7, 24, 14, -17, -29, 2, 11, -5, -7,
    -- filter=72 channel=123
    9, 6, -5, -9, 20, 11, 8, -12, -3,
    -- filter=72 channel=124
    -4, 0, 0, -5, 10, 11, -4, -4, -1,
    -- filter=72 channel=125
    -1, 25, 10, -21, -41, -4, 12, 7, -8,
    -- filter=72 channel=126
    -5, 0, -9, -1, -1, 8, -2, -4, 1,
    -- filter=72 channel=127
    -5, -9, -5, 4, 0, -11, -7, -3, 1,
    -- filter=73 channel=0
    -14, -1, 4, -13, -14, 5, 1, 5, 14,
    -- filter=73 channel=1
    -8, 3, 4, -5, -10, 10, 10, 6, 9,
    -- filter=73 channel=2
    -2, -3, 0, -3, 5, -4, 6, 2, 6,
    -- filter=73 channel=3
    5, 4, -4, 1, -7, -10, 7, 7, 2,
    -- filter=73 channel=4
    -5, -4, 4, 0, 9, -6, 18, 8, -4,
    -- filter=73 channel=5
    0, 4, 4, -12, -10, 8, 4, 12, 0,
    -- filter=73 channel=6
    5, 7, 10, 8, 10, 4, 5, 1, -9,
    -- filter=73 channel=7
    -4, 5, -1, 1, -2, 6, -3, 7, 3,
    -- filter=73 channel=8
    1, -5, 9, -1, 15, 1, 10, 5, 7,
    -- filter=73 channel=9
    0, -10, 2, -12, -7, -1, 4, 4, 0,
    -- filter=73 channel=10
    -1, -3, -10, 0, -15, 1, -7, -3, 12,
    -- filter=73 channel=11
    4, 6, 5, 7, 2, -7, 3, -5, -10,
    -- filter=73 channel=12
    3, -3, 13, 1, -3, 17, 7, 8, 2,
    -- filter=73 channel=13
    0, 2, -11, 0, -19, 3, -8, 3, 0,
    -- filter=73 channel=14
    3, 6, -4, 3, 7, -5, -6, -1, -1,
    -- filter=73 channel=15
    -5, -4, -3, 4, -6, -5, 5, -2, -7,
    -- filter=73 channel=16
    7, -5, 11, -9, -11, 5, 1, 4, 2,
    -- filter=73 channel=17
    5, 2, -1, 4, -3, 0, 2, 6, 6,
    -- filter=73 channel=18
    -1, 3, -10, 3, -5, 1, 0, 2, 5,
    -- filter=73 channel=19
    -4, -1, -5, -6, 1, 7, -5, -4, -1,
    -- filter=73 channel=20
    10, 10, 3, 5, 13, 0, -1, -15, -6,
    -- filter=73 channel=21
    0, -12, 3, -5, -15, 10, -6, 3, 12,
    -- filter=73 channel=22
    1, 1, 3, 1, 1, 1, -6, 7, -11,
    -- filter=73 channel=23
    7, -12, -7, -10, -12, 2, 2, -1, -5,
    -- filter=73 channel=24
    2, -1, 3, -5, -1, -1, 1, -2, -4,
    -- filter=73 channel=25
    -8, -14, 7, -16, -19, 10, 0, 5, 14,
    -- filter=73 channel=26
    -4, 4, 6, -4, -1, 6, 0, -2, 0,
    -- filter=73 channel=27
    -10, -30, 11, -26, -17, 25, 3, 16, 7,
    -- filter=73 channel=28
    0, -4, 2, 1, 7, -4, -2, 2, 5,
    -- filter=73 channel=29
    11, 5, -4, 11, 7, 9, -2, -9, -13,
    -- filter=73 channel=30
    -4, -10, 11, -18, -7, 8, 1, 7, 9,
    -- filter=73 channel=31
    -3, -26, -6, -16, -18, 14, -8, 11, 12,
    -- filter=73 channel=32
    7, -11, 7, 0, -18, 7, -5, 3, 0,
    -- filter=73 channel=33
    6, -2, -15, -15, -16, 0, 2, 0, 10,
    -- filter=73 channel=34
    0, 0, 15, -14, 3, 4, 8, 7, -1,
    -- filter=73 channel=35
    1, 3, -4, 4, -3, -2, -7, -6, 0,
    -- filter=73 channel=36
    5, -9, 4, 2, 2, 5, -6, 3, -8,
    -- filter=73 channel=37
    -14, -5, 10, -10, 3, 13, -5, 8, 4,
    -- filter=73 channel=38
    2, -8, 2, -11, -13, 10, 3, 0, 1,
    -- filter=73 channel=39
    6, 1, -3, 2, 0, 6, -2, -10, -10,
    -- filter=73 channel=40
    4, 8, -4, 8, -8, -6, -3, -9, -9,
    -- filter=73 channel=41
    -3, 0, -1, 2, -3, -9, -4, 5, 5,
    -- filter=73 channel=42
    -8, -5, -4, -1, -5, 5, 1, 8, -5,
    -- filter=73 channel=43
    5, 0, -13, -2, -5, 0, 2, 0, -4,
    -- filter=73 channel=44
    -7, -15, 3, -13, 1, 14, 5, 19, 10,
    -- filter=73 channel=45
    0, 5, 0, 0, 4, 0, 1, -1, -6,
    -- filter=73 channel=46
    -8, -2, 4, -2, -3, -5, -2, 3, 4,
    -- filter=73 channel=47
    0, -3, 0, -4, -5, 7, 0, 16, 14,
    -- filter=73 channel=48
    -7, -24, 0, -17, -1, 15, 6, 14, 12,
    -- filter=73 channel=49
    5, 1, 5, 2, 12, 4, 9, 9, -4,
    -- filter=73 channel=50
    -3, -18, -3, -15, -11, 3, 4, 5, 3,
    -- filter=73 channel=51
    1, 4, 2, 6, -2, 4, -1, -5, -1,
    -- filter=73 channel=52
    0, -7, 4, 3, 10, 10, 1, 0, -9,
    -- filter=73 channel=53
    -1, -1, 3, -4, 6, 8, -8, 5, 1,
    -- filter=73 channel=54
    0, 6, 0, 0, -4, 3, -7, -5, 3,
    -- filter=73 channel=55
    6, 0, -7, -2, -9, 2, -3, 0, 3,
    -- filter=73 channel=56
    -2, 4, 9, 1, 9, 10, -2, 6, 3,
    -- filter=73 channel=57
    0, -6, -7, -8, -1, 0, -2, -4, 2,
    -- filter=73 channel=58
    2, 8, -2, -3, -3, 7, -1, 1, 6,
    -- filter=73 channel=59
    -5, -16, -5, -11, -23, 4, -5, 1, 5,
    -- filter=73 channel=60
    2, 6, 2, -5, -4, -5, 0, 0, -1,
    -- filter=73 channel=61
    5, -1, 5, -3, 0, -2, 3, 0, -5,
    -- filter=73 channel=62
    -5, -4, -6, -2, 6, 0, -3, 0, 3,
    -- filter=73 channel=63
    0, 3, 7, -4, 6, -3, 1, -1, -2,
    -- filter=73 channel=64
    0, 0, 1, 1, 7, 2, 4, 3, -3,
    -- filter=73 channel=65
    5, 5, 5, -5, -6, -6, -6, 0, 5,
    -- filter=73 channel=66
    0, -2, 10, -1, -7, 4, -2, 7, 0,
    -- filter=73 channel=67
    -9, 4, 3, 5, 1, 5, 5, -2, 3,
    -- filter=73 channel=68
    1, 4, 4, 5, 1, 4, 4, 0, -2,
    -- filter=73 channel=69
    6, 2, -4, -4, 1, -1, -4, 4, -2,
    -- filter=73 channel=70
    0, -21, -4, -16, -11, 6, 6, 4, 1,
    -- filter=73 channel=71
    -3, 6, -8, 6, -4, -10, 0, -5, 3,
    -- filter=73 channel=72
    2, -13, -3, -7, -12, 3, -3, 1, 13,
    -- filter=73 channel=73
    0, -4, 11, -7, 5, 3, -1, 11, 2,
    -- filter=73 channel=74
    0, -17, 12, -19, 7, 14, 7, 7, -2,
    -- filter=73 channel=75
    -1, -1, -6, -12, -11, -3, -1, 0, 20,
    -- filter=73 channel=76
    9, 9, -2, 14, -4, -7, -6, -11, -3,
    -- filter=73 channel=77
    6, 6, -2, 6, 2, 0, -6, 3, 3,
    -- filter=73 channel=78
    -4, 4, 3, -10, -7, 2, 2, 8, -3,
    -- filter=73 channel=79
    0, -12, -6, 1, -20, 6, 0, 4, 0,
    -- filter=73 channel=80
    0, -15, -1, -9, -29, 12, -8, 7, 17,
    -- filter=73 channel=81
    2, -2, -3, -6, -7, -2, 4, 0, 7,
    -- filter=73 channel=82
    2, -6, -7, 4, 3, -4, 5, 3, 3,
    -- filter=73 channel=83
    -2, -1, -5, -8, -1, 3, 4, -2, 1,
    -- filter=73 channel=84
    6, -9, 5, -4, -3, 5, 6, 7, 2,
    -- filter=73 channel=85
    0, -3, 7, 5, 5, 6, -2, 4, -1,
    -- filter=73 channel=86
    5, 0, 7, 1, 0, 0, 7, 8, 1,
    -- filter=73 channel=87
    6, 9, 3, 8, 7, 6, 2, 2, -10,
    -- filter=73 channel=88
    -1, -5, 9, -9, 7, 11, 2, -4, -5,
    -- filter=73 channel=89
    7, -6, -7, -4, -19, 2, -10, 0, 12,
    -- filter=73 channel=90
    -2, -6, 7, 0, 7, 6, -3, 1, 3,
    -- filter=73 channel=91
    -6, -19, 2, -13, -4, 10, 7, 1, -7,
    -- filter=73 channel=92
    -4, 0, -8, 0, 2, 1, 3, -2, 6,
    -- filter=73 channel=93
    -14, -4, 11, -11, -6, 14, 10, 13, 13,
    -- filter=73 channel=94
    2, 4, -3, 7, 6, -6, -1, -3, -3,
    -- filter=73 channel=95
    -4, 2, 0, 8, -6, 2, 6, 7, 6,
    -- filter=73 channel=96
    -2, 0, 0, 0, -9, -7, 3, 3, 5,
    -- filter=73 channel=97
    -3, 5, -9, 2, -12, -9, -3, 5, 1,
    -- filter=73 channel=98
    3, -6, -7, -18, -17, 23, -3, 8, 18,
    -- filter=73 channel=99
    2, -13, 0, -9, -4, 19, -5, 14, -4,
    -- filter=73 channel=100
    -5, 7, 7, 0, 5, -4, 2, -2, -3,
    -- filter=73 channel=101
    2, 2, 7, -3, 13, 4, 5, 5, -6,
    -- filter=73 channel=102
    -3, -2, 0, 3, -7, -6, 2, 4, -3,
    -- filter=73 channel=103
    7, -5, 0, -13, -23, 7, 6, 1, 23,
    -- filter=73 channel=104
    1, -16, -4, -5, -7, 12, -8, 3, 8,
    -- filter=73 channel=105
    1, 8, -4, 9, 12, -4, -4, -8, -12,
    -- filter=73 channel=106
    0, -1, 3, 9, 0, 2, 0, -6, -7,
    -- filter=73 channel=107
    0, -2, 8, -5, 7, 0, -4, -8, -16,
    -- filter=73 channel=108
    -1, 11, 6, 7, -4, -5, 5, 3, -3,
    -- filter=73 channel=109
    2, -14, 10, -20, -8, 15, -7, 12, 0,
    -- filter=73 channel=110
    -1, -9, 1, -5, -14, 2, -6, 6, 1,
    -- filter=73 channel=111
    -1, 1, -1, 6, -3, 6, 2, 4, -5,
    -- filter=73 channel=112
    -5, -6, 11, -14, 0, 5, -3, 6, 1,
    -- filter=73 channel=113
    -4, 1, -6, -5, -18, 3, 0, 6, 3,
    -- filter=73 channel=114
    2, -10, 4, -10, 0, 17, 6, 16, 3,
    -- filter=73 channel=115
    2, -4, -3, 0, 1, -5, -4, -5, -2,
    -- filter=73 channel=116
    -4, -15, -5, -3, -13, 8, 4, 7, 0,
    -- filter=73 channel=117
    6, -4, -7, 5, -5, -6, 0, -4, -3,
    -- filter=73 channel=118
    5, 6, 0, 1, 1, -2, -2, 7, 3,
    -- filter=73 channel=119
    -3, -3, 26, -21, 20, 7, 6, 4, 0,
    -- filter=73 channel=120
    -5, -26, 16, -24, 10, 29, 2, 16, 5,
    -- filter=73 channel=121
    5, 2, -3, 0, -10, 5, -2, 6, 8,
    -- filter=73 channel=122
    4, -9, 11, -12, -2, 17, 3, 9, 23,
    -- filter=73 channel=123
    -9, 0, 8, -9, 0, -2, -3, 4, -2,
    -- filter=73 channel=124
    10, 1, 2, 1, -1, 0, 2, 0, 2,
    -- filter=73 channel=125
    5, -26, 4, -9, -5, 15, -7, 6, 11,
    -- filter=73 channel=126
    0, 1, -1, 6, -11, 4, 0, 2, 14,
    -- filter=73 channel=127
    4, -3, -1, 5, 4, -3, -3, 6, -3,
    -- filter=74 channel=0
    17, 17, 7, 8, 5, 10, -10, -9, -1,
    -- filter=74 channel=1
    4, 11, 5, 5, 6, 4, -6, 2, -6,
    -- filter=74 channel=2
    2, -4, -2, -4, 5, 0, -5, -4, -5,
    -- filter=74 channel=3
    1, 7, -5, 0, 1, 1, -3, -1, -7,
    -- filter=74 channel=4
    9, 3, 15, -5, 0, 8, -6, -6, -3,
    -- filter=74 channel=5
    -4, -9, -13, -2, 3, 0, -5, 2, 1,
    -- filter=74 channel=6
    3, 6, 0, -4, 1, -1, 4, 0, -13,
    -- filter=74 channel=7
    -5, -7, 6, 0, -6, 6, 0, 6, 3,
    -- filter=74 channel=8
    6, 2, 0, -4, 7, 5, 4, 4, -7,
    -- filter=74 channel=9
    -1, 0, -9, -4, 7, 9, 4, 1, -3,
    -- filter=74 channel=10
    -13, -12, -16, -8, -12, 5, 3, -2, 8,
    -- filter=74 channel=11
    -1, 8, 0, -2, -6, 3, -5, -6, -8,
    -- filter=74 channel=12
    3, -9, 5, 5, -11, 2, -5, 1, -7,
    -- filter=74 channel=13
    -3, 7, -3, 0, -5, 2, -2, -8, -9,
    -- filter=74 channel=14
    -1, 3, 0, 0, 1, 2, 3, -4, -7,
    -- filter=74 channel=15
    4, 11, 7, 0, 4, -1, 0, -8, -14,
    -- filter=74 channel=16
    -7, -4, -2, -7, 3, 0, -1, 1, 3,
    -- filter=74 channel=17
    3, 5, -4, -1, -3, 5, 6, 0, -6,
    -- filter=74 channel=18
    13, 8, 1, 0, 0, -2, -1, -12, -11,
    -- filter=74 channel=19
    2, 2, -3, -6, 0, 7, -5, 6, -3,
    -- filter=74 channel=20
    8, 6, 9, 4, 1, 7, -1, -11, -12,
    -- filter=74 channel=21
    -2, -14, -9, -5, 9, 13, 8, 9, 24,
    -- filter=74 channel=22
    -3, 6, -4, 1, 6, 0, 0, -7, -12,
    -- filter=74 channel=23
    -3, -5, -5, 7, -6, 7, -4, -6, -8,
    -- filter=74 channel=24
    2, -6, -7, -1, 3, 6, 1, -7, 4,
    -- filter=74 channel=25
    8, 1, -13, -7, 7, 0, -5, -5, -9,
    -- filter=74 channel=26
    -8, -3, 0, -2, -5, 8, 5, -1, 3,
    -- filter=74 channel=27
    11, 0, -11, -3, 2, 5, 1, -6, 2,
    -- filter=74 channel=28
    3, 2, 1, -4, 6, 1, 5, 6, -2,
    -- filter=74 channel=29
    7, 13, 14, -2, 6, 4, -8, -8, -15,
    -- filter=74 channel=30
    8, 4, -5, -6, 12, 13, -5, -4, 4,
    -- filter=74 channel=31
    -4, -21, -23, -12, 2, 12, 0, 7, 28,
    -- filter=74 channel=32
    8, 1, -4, 8, 5, 6, 6, -15, -19,
    -- filter=74 channel=33
    0, -10, -1, 3, 8, -4, -5, 0, 0,
    -- filter=74 channel=34
    -2, 1, 1, 0, -4, -4, -3, -9, -7,
    -- filter=74 channel=35
    -1, 4, -2, 1, -2, 0, 2, 5, 6,
    -- filter=74 channel=36
    5, -2, 2, -5, -3, 0, 6, 2, 13,
    -- filter=74 channel=37
    11, 0, 6, 0, 13, 10, 3, 8, 2,
    -- filter=74 channel=38
    -1, 0, -7, 2, 3, -1, -6, -5, 5,
    -- filter=74 channel=39
    8, 11, 0, 7, 1, 6, -3, -5, 3,
    -- filter=74 channel=40
    9, 10, 11, 7, 8, 1, 11, 6, 2,
    -- filter=74 channel=41
    1, 4, 8, -7, -18, -17, -2, -12, -21,
    -- filter=74 channel=42
    8, 4, 0, 2, 0, 2, -5, 2, -1,
    -- filter=74 channel=43
    7, -3, -3, -5, -6, 0, -8, -8, -2,
    -- filter=74 channel=44
    4, -13, -12, 3, 4, 14, -3, 6, 14,
    -- filter=74 channel=45
    -2, 11, -3, 8, 0, 11, 5, 3, 9,
    -- filter=74 channel=46
    3, -2, 0, -2, -1, -4, -4, 5, -6,
    -- filter=74 channel=47
    -1, -7, -9, -7, 10, 6, -9, 15, 13,
    -- filter=74 channel=48
    -3, -14, -10, 0, 0, 11, -6, 1, 0,
    -- filter=74 channel=49
    2, 6, 13, 3, 5, 0, 0, -7, -7,
    -- filter=74 channel=50
    -3, -8, -10, -1, 0, 3, 1, 8, 2,
    -- filter=74 channel=51
    -1, 4, -1, -6, 3, -3, 6, 5, 1,
    -- filter=74 channel=52
    8, 6, 5, 0, 2, 2, 11, 2, -9,
    -- filter=74 channel=53
    -7, 1, 8, -2, -5, 6, 5, -9, -4,
    -- filter=74 channel=54
    -1, -4, -1, -2, 3, 5, -7, 6, -7,
    -- filter=74 channel=55
    2, -1, 5, 3, -5, -7, 1, -9, -11,
    -- filter=74 channel=56
    6, -5, 3, 3, 3, -9, 5, 1, -9,
    -- filter=74 channel=57
    3, -1, 6, -2, 0, -5, -5, 0, -1,
    -- filter=74 channel=58
    2, 1, 4, -6, 8, -4, 1, -4, 5,
    -- filter=74 channel=59
    1, -2, -8, -7, 0, 6, 0, 1, 7,
    -- filter=74 channel=60
    -5, -1, 2, -3, 5, 4, 2, 1, -6,
    -- filter=74 channel=61
    2, 5, 5, -6, 3, 4, 1, 0, -1,
    -- filter=74 channel=62
    -3, 1, -6, 2, -4, 0, 2, -6, -7,
    -- filter=74 channel=63
    -5, -4, -1, 4, 7, 4, 3, -3, 0,
    -- filter=74 channel=64
    -2, -1, -1, 5, 4, 4, 7, -4, 8,
    -- filter=74 channel=65
    -7, 1, 2, -2, 0, 5, -1, -3, 2,
    -- filter=74 channel=66
    0, -1, -3, 4, -3, -3, 6, -7, -10,
    -- filter=74 channel=67
    4, -5, 3, 0, -6, -4, 6, 0, 6,
    -- filter=74 channel=68
    0, 0, 1, -4, 0, 8, -1, 2, 2,
    -- filter=74 channel=69
    -7, -7, 2, -4, -4, 0, -5, 3, 3,
    -- filter=74 channel=70
    2, 4, -3, 5, 7, 8, 0, 0, -6,
    -- filter=74 channel=71
    0, 2, 1, 0, -3, 2, 1, -3, -1,
    -- filter=74 channel=72
    -3, -11, -9, 0, -8, 2, 3, 7, 7,
    -- filter=74 channel=73
    1, -4, 3, -3, 1, 8, 1, 1, -6,
    -- filter=74 channel=74
    6, -7, -8, 0, 0, 4, 1, 3, 7,
    -- filter=74 channel=75
    14, 6, -3, 0, 2, 0, -7, 3, -5,
    -- filter=74 channel=76
    12, 18, 18, 1, -1, 6, 6, -9, -4,
    -- filter=74 channel=77
    -4, 3, 0, 6, -5, 3, -6, 1, -4,
    -- filter=74 channel=78
    1, -9, -9, -3, -7, 5, 4, -2, -4,
    -- filter=74 channel=79
    14, 4, -1, 0, -1, 6, 6, -7, -20,
    -- filter=74 channel=80
    -2, -24, -23, -5, -1, 6, 5, 3, 15,
    -- filter=74 channel=81
    -2, -3, -2, -2, -2, -2, -2, 0, -7,
    -- filter=74 channel=82
    -2, -7, -4, 5, 4, 7, 4, -3, 9,
    -- filter=74 channel=83
    1, -1, 0, 2, 1, 4, -7, 0, 9,
    -- filter=74 channel=84
    0, 3, 6, 4, 6, 3, -4, -5, -11,
    -- filter=74 channel=85
    -3, 7, 5, 7, 5, -5, -2, -3, 0,
    -- filter=74 channel=86
    7, 4, 6, 6, -2, 4, 2, -4, -2,
    -- filter=74 channel=87
    1, 1, 9, 0, -3, -4, -1, -9, -6,
    -- filter=74 channel=88
    1, 0, 6, 2, 1, 9, 11, 0, 11,
    -- filter=74 channel=89
    -13, 0, -8, -7, -10, -4, 5, -3, 0,
    -- filter=74 channel=90
    0, -2, 6, 3, 6, 2, 5, 10, 17,
    -- filter=74 channel=91
    1, 4, 11, 1, 0, 9, 8, 2, -2,
    -- filter=74 channel=92
    7, -4, -3, 2, -1, -3, 5, 3, -4,
    -- filter=74 channel=93
    2, -2, -10, -15, 2, 5, 3, -5, 7,
    -- filter=74 channel=94
    -4, -5, 0, -2, 2, 3, 0, -5, 6,
    -- filter=74 channel=95
    5, 0, 0, 1, -3, -1, 4, -4, -7,
    -- filter=74 channel=96
    2, -6, -1, 7, 3, -6, 0, 6, -1,
    -- filter=74 channel=97
    3, -3, -7, 5, 10, 0, -7, 4, -3,
    -- filter=74 channel=98
    -9, -7, -21, -7, 4, 4, 2, -1, -8,
    -- filter=74 channel=99
    -7, -15, -18, -3, -2, 0, 7, -9, 1,
    -- filter=74 channel=100
    4, 2, 2, 5, -8, -2, -5, -4, -4,
    -- filter=74 channel=101
    8, 1, 7, -1, 3, 11, -4, -5, -7,
    -- filter=74 channel=102
    5, 0, -2, -1, 3, -3, 1, -3, 5,
    -- filter=74 channel=103
    -8, -11, -19, -9, 8, 1, -7, 11, 9,
    -- filter=74 channel=104
    -2, -15, -8, -9, 0, 11, 0, 4, 12,
    -- filter=74 channel=105
    3, 2, 12, -7, -1, 2, 2, -8, -14,
    -- filter=74 channel=106
    6, 10, 0, 4, 6, -4, -3, 8, 0,
    -- filter=74 channel=107
    11, 16, 17, 12, 8, 0, -5, -2, -8,
    -- filter=74 channel=108
    7, 6, 6, 0, 5, 0, 0, 1, -8,
    -- filter=74 channel=109
    1, -7, -11, 1, 0, 7, 0, -1, -7,
    -- filter=74 channel=110
    -6, -2, -1, -10, -7, 5, -8, -4, 6,
    -- filter=74 channel=111
    2, 7, 7, 2, 6, -3, 7, 2, -5,
    -- filter=74 channel=112
    -2, -4, -4, -7, -5, -2, 6, -8, -4,
    -- filter=74 channel=113
    -8, -9, -11, -1, -3, 4, -3, 4, 5,
    -- filter=74 channel=114
    6, 12, 7, 3, -3, 4, -13, -20, -19,
    -- filter=74 channel=115
    -6, -3, 5, -6, -1, 2, 0, -2, 2,
    -- filter=74 channel=116
    -3, -11, -9, -4, -5, 8, 7, -5, -3,
    -- filter=74 channel=117
    6, -5, 3, 2, -3, 1, 2, 7, 0,
    -- filter=74 channel=118
    6, 5, -2, 0, 1, 0, 2, 1, -5,
    -- filter=74 channel=119
    -9, -4, -7, -7, 2, -9, 8, -7, -6,
    -- filter=74 channel=120
    3, -6, 5, -3, -1, -1, -1, -7, -6,
    -- filter=74 channel=121
    -10, -4, 0, -5, -1, 2, 2, 2, -3,
    -- filter=74 channel=122
    -13, -13, -15, 2, 10, 16, 4, 22, 36,
    -- filter=74 channel=123
    0, -5, 3, 1, 2, 3, 0, 3, 1,
    -- filter=74 channel=124
    -5, 3, 5, 4, -1, -3, 4, -12, -13,
    -- filter=74 channel=125
    -10, -6, -17, -6, 3, 9, 4, 4, 7,
    -- filter=74 channel=126
    -2, -7, -3, -5, 4, 3, -3, -9, -6,
    -- filter=74 channel=127
    -2, -2, -3, -7, -7, -6, 6, 0, 4,
    -- filter=75 channel=0
    3, 13, -11, 14, 12, -14, 4, -1, -12,
    -- filter=75 channel=1
    11, 6, 4, 14, 2, -15, -6, -5, -9,
    -- filter=75 channel=2
    0, 4, -3, 0, -6, 4, -2, 3, -3,
    -- filter=75 channel=3
    9, 3, -2, -1, 9, 2, -2, 2, 5,
    -- filter=75 channel=4
    -5, 6, -1, 1, 2, -2, -5, -4, -4,
    -- filter=75 channel=5
    -1, 4, -7, 9, 0, -9, 1, -4, -8,
    -- filter=75 channel=6
    4, 1, -2, -9, 2, -4, -3, 1, 1,
    -- filter=75 channel=7
    3, 0, 6, 4, -7, -4, -5, -6, 3,
    -- filter=75 channel=8
    -6, 1, -1, -5, 1, -1, 1, 2, 5,
    -- filter=75 channel=9
    5, 5, -1, -1, 5, -5, -8, 6, -7,
    -- filter=75 channel=10
    2, 3, -4, -11, -9, -1, -1, -8, 0,
    -- filter=75 channel=11
    -9, -3, -1, -2, 1, -5, -12, -10, -3,
    -- filter=75 channel=12
    0, 0, -6, 5, -2, -3, -3, -8, 0,
    -- filter=75 channel=13
    10, 3, 3, 0, -3, 9, -7, -5, 4,
    -- filter=75 channel=14
    -5, 3, 1, -2, 4, 5, -2, 5, -1,
    -- filter=75 channel=15
    5, 5, 4, 0, 0, 1, -8, 0, 1,
    -- filter=75 channel=16
    4, 1, -3, 6, 9, 2, 6, -2, -2,
    -- filter=75 channel=17
    0, 3, 4, -1, -6, 0, 3, -5, 3,
    -- filter=75 channel=18
    9, 12, 5, -1, -4, -3, -8, -7, -4,
    -- filter=75 channel=19
    0, 3, 1, -3, 0, -3, 2, -5, 5,
    -- filter=75 channel=20
    -12, -8, -11, -15, -12, 0, -13, -14, -11,
    -- filter=75 channel=21
    -4, 1, -5, 0, 0, 7, -1, -5, 8,
    -- filter=75 channel=22
    4, -2, -8, 5, 1, 0, 1, 2, -1,
    -- filter=75 channel=23
    12, 12, 3, -5, 3, 7, -17, -2, 7,
    -- filter=75 channel=24
    -5, 2, -8, 5, -4, -7, -3, -5, -4,
    -- filter=75 channel=25
    0, 1, 6, -2, -6, 1, -1, 0, -5,
    -- filter=75 channel=26
    0, -3, -3, 3, 4, 0, 4, -1, 2,
    -- filter=75 channel=27
    7, 9, 8, 1, -1, 4, -6, -7, -1,
    -- filter=75 channel=28
    6, -3, -4, 1, 2, -2, -6, 0, 6,
    -- filter=75 channel=29
    1, -9, -9, -5, -5, -13, -6, -15, -11,
    -- filter=75 channel=30
    1, -1, -8, 0, 0, -4, -5, 4, -9,
    -- filter=75 channel=31
    0, -4, 11, -5, 10, 16, -1, 0, 15,
    -- filter=75 channel=32
    12, 13, -2, -4, -6, 3, -6, -15, -10,
    -- filter=75 channel=33
    14, 14, 7, 1, 8, 9, 0, -1, -4,
    -- filter=75 channel=34
    0, 9, -3, -7, 9, -8, -6, -7, 4,
    -- filter=75 channel=35
    6, 5, -5, 6, -6, -1, -3, 5, 0,
    -- filter=75 channel=36
    -13, 2, -1, -4, -8, 10, 5, 0, 7,
    -- filter=75 channel=37
    11, 3, 3, 3, 12, -9, -4, 9, -2,
    -- filter=75 channel=38
    1, -4, -7, -6, 4, 7, 2, 4, 1,
    -- filter=75 channel=39
    0, -6, -5, 2, -7, 3, -5, -2, 0,
    -- filter=75 channel=40
    5, -1, -3, -4, -8, 7, -4, -7, 1,
    -- filter=75 channel=41
    12, 13, -2, -9, -10, -3, -5, -14, -10,
    -- filter=75 channel=42
    4, -1, 0, 7, 9, 1, 5, 7, 0,
    -- filter=75 channel=43
    9, 2, 0, 1, -7, -5, -3, -9, -8,
    -- filter=75 channel=44
    4, 6, 5, 3, 9, -5, 1, 2, 5,
    -- filter=75 channel=45
    0, 6, -7, 2, -3, 0, 6, 1, -2,
    -- filter=75 channel=46
    -1, 8, 3, -3, 3, -3, -4, 0, 5,
    -- filter=75 channel=47
    10, -6, -10, 2, 0, 8, 12, 7, 0,
    -- filter=75 channel=48
    1, 1, 3, 6, 5, 0, 1, -2, 7,
    -- filter=75 channel=49
    0, 4, 7, -9, 3, -6, -13, -11, -3,
    -- filter=75 channel=50
    5, 11, 9, -3, 11, 4, -10, -3, -3,
    -- filter=75 channel=51
    -4, 6, -2, 5, 4, -5, -6, 0, 3,
    -- filter=75 channel=52
    0, 7, -4, -3, -5, 0, 0, 0, 2,
    -- filter=75 channel=53
    -7, -4, 1, -9, -8, -5, -1, -10, -4,
    -- filter=75 channel=54
    4, 4, -1, 3, -4, -6, 1, 3, -4,
    -- filter=75 channel=55
    -3, -3, -3, -17, -5, -3, -6, -3, -9,
    -- filter=75 channel=56
    -4, 5, 2, -6, -3, -7, 2, -5, 2,
    -- filter=75 channel=57
    5, 6, 5, 5, 1, -4, 3, -4, -8,
    -- filter=75 channel=58
    -2, -2, -1, 0, -3, -4, 3, 6, -12,
    -- filter=75 channel=59
    1, -3, 0, 1, 4, 6, -7, -6, -2,
    -- filter=75 channel=60
    -2, 3, 1, -3, 0, -6, 7, 4, 7,
    -- filter=75 channel=61
    -5, -6, 5, -2, -6, -6, 1, -2, -5,
    -- filter=75 channel=62
    -3, 0, -6, 0, 1, 0, 5, -3, 0,
    -- filter=75 channel=63
    -7, -11, -16, 2, -6, -11, -7, 0, -5,
    -- filter=75 channel=64
    -7, 2, 6, -4, -1, 5, 3, 0, 1,
    -- filter=75 channel=65
    7, -6, -6, -1, -2, 2, -4, -1, 6,
    -- filter=75 channel=66
    8, 8, 4, 6, -8, -6, -6, -2, -2,
    -- filter=75 channel=67
    4, 0, -6, 4, 1, -5, -2, -1, -3,
    -- filter=75 channel=68
    -2, -2, 0, -8, 6, 1, -6, 1, -6,
    -- filter=75 channel=69
    6, -4, 2, -5, -3, -6, 1, 2, -6,
    -- filter=75 channel=70
    7, 16, 2, -1, 7, 12, -11, 5, 4,
    -- filter=75 channel=71
    12, 4, -2, 6, 3, 0, -2, 0, 10,
    -- filter=75 channel=72
    2, -8, 10, -2, -4, 15, -2, 1, 9,
    -- filter=75 channel=73
    2, -1, 8, -7, -9, 1, -5, -11, 2,
    -- filter=75 channel=74
    10, 4, 3, -6, 3, -1, -7, 1, 1,
    -- filter=75 channel=75
    20, 6, -12, 11, 12, -8, 6, 2, -6,
    -- filter=75 channel=76
    -10, 1, -9, -14, -15, -9, -4, -11, -8,
    -- filter=75 channel=77
    7, -2, 4, 4, -2, -3, -2, 4, -6,
    -- filter=75 channel=78
    0, -2, -10, 5, 0, -4, 1, 3, -7,
    -- filter=75 channel=79
    15, 7, 8, -7, 1, -5, -10, -3, -2,
    -- filter=75 channel=80
    4, 1, -2, 6, -4, 15, 3, -4, 9,
    -- filter=75 channel=81
    0, 7, 6, -2, -1, -6, -2, 5, 6,
    -- filter=75 channel=82
    6, 7, 0, 2, -6, 5, 5, 5, 0,
    -- filter=75 channel=83
    -3, -4, 0, -4, 0, 5, -8, -7, -2,
    -- filter=75 channel=84
    -4, 10, 5, -11, -9, -6, -1, -7, -6,
    -- filter=75 channel=85
    -2, 0, -4, -1, -4, -1, 0, 0, -5,
    -- filter=75 channel=86
    -5, 4, -8, 6, 0, -2, 5, -1, -9,
    -- filter=75 channel=87
    2, 5, -8, -12, -2, -10, -4, -8, -2,
    -- filter=75 channel=88
    -7, 1, -5, 0, 2, 5, -4, 8, 6,
    -- filter=75 channel=89
    9, 7, 13, -10, -12, 13, -1, 0, 4,
    -- filter=75 channel=90
    -6, -1, 0, 1, 6, 3, -7, 4, 6,
    -- filter=75 channel=91
    7, 1, 5, -7, -3, -2, -2, 0, -3,
    -- filter=75 channel=92
    -1, -3, -2, 0, -5, 3, -2, 7, -3,
    -- filter=75 channel=93
    0, -4, -8, -1, 4, -5, -4, 4, 3,
    -- filter=75 channel=94
    -6, -3, 3, 7, 0, -3, -2, 5, 1,
    -- filter=75 channel=95
    1, -1, 0, -1, -2, -1, 2, 3, 0,
    -- filter=75 channel=96
    0, 0, -3, -6, -6, -5, 1, -3, 7,
    -- filter=75 channel=97
    3, 8, 2, 6, 1, 3, 1, 0, 8,
    -- filter=75 channel=98
    4, 3, 1, -6, -6, 7, -4, -8, 0,
    -- filter=75 channel=99
    -6, -7, 0, -5, -2, 9, -8, -12, 2,
    -- filter=75 channel=100
    0, -3, 7, -8, 1, -3, -4, -4, 0,
    -- filter=75 channel=101
    -4, 6, 8, 4, -5, -6, 2, -8, -3,
    -- filter=75 channel=102
    -4, -7, -5, -3, 1, 0, 6, 5, 2,
    -- filter=75 channel=103
    10, 3, 0, 11, 2, 3, 3, 11, 0,
    -- filter=75 channel=104
    -9, 2, -4, 2, 5, 11, -3, -6, 0,
    -- filter=75 channel=105
    0, -9, 1, -3, -7, -11, 1, -1, -11,
    -- filter=75 channel=106
    -6, 0, -4, -5, -2, -3, -3, 4, 1,
    -- filter=75 channel=107
    -2, -4, -5, -4, -12, -9, -4, -1, -3,
    -- filter=75 channel=108
    -3, -3, 0, 5, -11, 0, -4, -9, -6,
    -- filter=75 channel=109
    3, 7, -1, -3, 0, -6, -9, -5, 0,
    -- filter=75 channel=110
    -7, 4, 9, 0, -5, 0, 1, -5, -2,
    -- filter=75 channel=111
    -2, 0, 0, -6, 4, -9, 0, 0, -2,
    -- filter=75 channel=112
    3, 8, -5, 4, 0, -1, -3, 3, 2,
    -- filter=75 channel=113
    11, 9, 6, 7, 8, 1, -5, -3, 1,
    -- filter=75 channel=114
    12, 2, 0, -3, -8, -7, -16, -6, -15,
    -- filter=75 channel=115
    -7, 5, -2, 4, -3, 0, -2, -5, -7,
    -- filter=75 channel=116
    1, -9, -1, -8, -13, 1, -11, -5, 3,
    -- filter=75 channel=117
    -1, 0, -3, -1, -4, 0, -5, -6, 8,
    -- filter=75 channel=118
    4, 1, -1, 6, 0, -5, 5, 4, -7,
    -- filter=75 channel=119
    -1, 6, -3, -7, 6, 3, -6, -3, -5,
    -- filter=75 channel=120
    -5, 3, 2, -16, 1, -9, -17, -12, -5,
    -- filter=75 channel=121
    -1, 8, -5, -8, 0, 10, -6, -3, 3,
    -- filter=75 channel=122
    -4, -6, -9, 15, 10, 3, 14, 4, 5,
    -- filter=75 channel=123
    -5, 11, -5, -5, 0, 7, -1, 5, 1,
    -- filter=75 channel=124
    3, 0, 0, -2, -5, 0, 0, 1, -1,
    -- filter=75 channel=125
    -6, -7, -2, -11, -8, 6, -12, -7, 8,
    -- filter=75 channel=126
    11, 1, -5, 0, 2, 8, 2, -4, 0,
    -- filter=75 channel=127
    3, 0, 0, -1, 0, -2, -6, 1, 0,
    -- filter=76 channel=0
    5, 1, 4, 0, 5, -4, -2, 0, 2,
    -- filter=76 channel=1
    1, 5, -6, -3, 0, 0, -2, 6, -5,
    -- filter=76 channel=2
    3, -4, -4, -1, 0, -7, -7, 1, 4,
    -- filter=76 channel=3
    -1, -1, 7, -7, -3, 0, 0, 8, 0,
    -- filter=76 channel=4
    2, -7, 6, -4, 3, 2, -4, 0, 5,
    -- filter=76 channel=5
    0, 7, -2, 4, 2, 5, 1, 4, 7,
    -- filter=76 channel=6
    3, -3, -2, 7, -1, -5, 6, -5, -6,
    -- filter=76 channel=7
    1, 1, 3, 4, -2, 4, -1, -1, -6,
    -- filter=76 channel=8
    0, 1, -5, 6, -3, -7, -5, -2, -7,
    -- filter=76 channel=9
    -7, -2, 3, -1, -6, 0, -2, -6, -7,
    -- filter=76 channel=10
    3, -5, 4, -4, -8, -2, 7, 6, -5,
    -- filter=76 channel=11
    6, 7, -6, -2, 3, 6, -5, 7, -4,
    -- filter=76 channel=12
    5, 6, -3, 0, -1, -4, 3, 2, 6,
    -- filter=76 channel=13
    4, 0, -4, 1, 0, -4, 2, 5, -5,
    -- filter=76 channel=14
    0, 4, -6, 3, 6, 0, 6, 0, 7,
    -- filter=76 channel=15
    5, -6, -3, -5, 0, 1, 4, 2, -7,
    -- filter=76 channel=16
    -4, -7, -6, 0, 4, -3, -4, -1, 0,
    -- filter=76 channel=17
    -7, -6, 6, 2, 1, 0, -1, 6, 4,
    -- filter=76 channel=18
    9, -4, 3, 5, -7, -3, 0, -1, 1,
    -- filter=76 channel=19
    -1, 0, 3, 4, -2, -2, 6, -6, 2,
    -- filter=76 channel=20
    -4, 1, 0, 8, 5, -5, -2, -5, 4,
    -- filter=76 channel=21
    -3, 4, 0, 4, -4, 6, 5, -2, -4,
    -- filter=76 channel=22
    0, 2, -5, 2, -4, -1, -3, 6, -6,
    -- filter=76 channel=23
    3, -5, 0, 0, -2, -1, 6, 0, -4,
    -- filter=76 channel=24
    -3, 0, 1, 1, -4, -2, 1, 7, -6,
    -- filter=76 channel=25
    1, 0, 4, -6, 0, -3, -3, 3, -3,
    -- filter=76 channel=26
    -3, 2, 1, -6, 5, 6, 0, -2, 0,
    -- filter=76 channel=27
    -7, -6, 3, 2, -3, -4, 1, -3, -2,
    -- filter=76 channel=28
    4, -5, -5, 3, 7, 1, 3, 3, 3,
    -- filter=76 channel=29
    -4, 1, -3, 0, -2, -1, -4, -2, 1,
    -- filter=76 channel=30
    2, -2, 1, 0, 0, 6, 4, 1, 0,
    -- filter=76 channel=31
    -4, -6, 3, -6, -1, -8, 6, -5, -5,
    -- filter=76 channel=32
    3, 0, 0, -5, 4, -3, -6, 4, 0,
    -- filter=76 channel=33
    0, -3, -8, -2, 3, -4, 1, 3, 7,
    -- filter=76 channel=34
    -6, 6, -2, -1, 6, -5, 3, 2, 1,
    -- filter=76 channel=35
    -5, 1, 0, -5, 6, -3, 0, -6, 1,
    -- filter=76 channel=36
    -4, -4, 6, 4, 3, 4, 5, 6, 2,
    -- filter=76 channel=37
    5, -6, 2, -3, 2, -4, -6, 5, -6,
    -- filter=76 channel=38
    -4, 5, 5, -2, 0, 6, -4, 0, -6,
    -- filter=76 channel=39
    2, -6, 3, 1, -4, -5, 2, 1, 0,
    -- filter=76 channel=40
    3, 3, 0, 4, 4, 6, 5, -5, -5,
    -- filter=76 channel=41
    6, 3, -2, -1, 8, 7, -3, 3, 7,
    -- filter=76 channel=42
    3, -7, 4, 2, -1, -7, 2, 0, -4,
    -- filter=76 channel=43
    8, 0, -2, 0, 0, 2, 6, 2, 6,
    -- filter=76 channel=44
    -8, -4, -6, -5, 2, -6, -4, -2, -4,
    -- filter=76 channel=45
    7, -5, 2, -6, -2, -5, 7, -1, 3,
    -- filter=76 channel=46
    0, 5, -1, 0, -3, -2, 7, 5, -5,
    -- filter=76 channel=47
    2, 0, -6, 5, -7, -5, -3, -4, -4,
    -- filter=76 channel=48
    -6, 2, 0, -1, 5, -7, 2, -4, 5,
    -- filter=76 channel=49
    -3, -2, 2, 1, -3, 2, 5, 3, 4,
    -- filter=76 channel=50
    -5, -7, 0, -3, 0, 4, 0, -6, -4,
    -- filter=76 channel=51
    0, 1, 5, -6, -1, 6, 7, 0, 4,
    -- filter=76 channel=52
    4, -6, -4, 5, 1, 0, 0, 0, -7,
    -- filter=76 channel=53
    1, 5, -5, 6, 0, 1, -2, 0, 0,
    -- filter=76 channel=54
    0, 3, -7, 2, 7, 3, -5, -2, -5,
    -- filter=76 channel=55
    6, 0, -3, 0, 0, 3, 3, -5, 3,
    -- filter=76 channel=56
    -1, -3, 3, 5, 4, -1, -3, -6, 0,
    -- filter=76 channel=57
    5, 0, 5, -2, 5, 6, 0, 3, 2,
    -- filter=76 channel=58
    0, -2, -2, 5, 0, -2, -4, 0, -3,
    -- filter=76 channel=59
    -5, 0, 2, -4, -8, -3, -1, 0, -3,
    -- filter=76 channel=60
    0, 4, -6, -4, -5, 0, -1, -1, -3,
    -- filter=76 channel=61
    -4, 7, -6, -2, -5, -1, 2, 6, -2,
    -- filter=76 channel=62
    1, 4, 2, 2, 1, 5, 7, -1, 0,
    -- filter=76 channel=63
    4, 7, -2, 0, 8, 6, -3, 0, 1,
    -- filter=76 channel=64
    0, -1, 0, 0, 3, -5, 6, -2, 3,
    -- filter=76 channel=65
    -5, -1, -4, -4, 7, -6, -6, 0, 7,
    -- filter=76 channel=66
    7, -6, 5, 0, 5, -3, -1, 6, 7,
    -- filter=76 channel=67
    -6, -4, 5, 4, 5, 2, 5, 4, -4,
    -- filter=76 channel=68
    2, -2, 5, 7, -5, 0, 2, -4, 7,
    -- filter=76 channel=69
    5, -4, 3, 0, 0, 0, 6, -3, -2,
    -- filter=76 channel=70
    -6, -4, 1, 3, 6, 2, 5, 4, 0,
    -- filter=76 channel=71
    0, 0, 0, 0, 0, -1, 7, 0, 6,
    -- filter=76 channel=72
    2, 0, -2, 6, 0, -1, 4, -7, 5,
    -- filter=76 channel=73
    -6, 0, 1, 6, 6, -2, -6, 0, -2,
    -- filter=76 channel=74
    -5, -6, 1, -5, 3, -6, -9, -1, 0,
    -- filter=76 channel=75
    5, -1, 1, 6, 0, 5, -2, -4, -3,
    -- filter=76 channel=76
    -3, 1, -1, 7, -6, -7, 0, 8, 8,
    -- filter=76 channel=77
    5, 2, -1, -2, 6, 4, -2, 6, -3,
    -- filter=76 channel=78
    -5, 7, -5, -3, -6, -3, 1, 5, -6,
    -- filter=76 channel=79
    7, 4, -8, 6, -7, -4, 8, -2, 4,
    -- filter=76 channel=80
    -4, -1, -1, 0, -8, -7, -6, -9, 2,
    -- filter=76 channel=81
    -7, 5, 0, -1, 6, 2, 6, 6, 0,
    -- filter=76 channel=82
    0, -2, 6, 6, 0, -1, 6, 3, -7,
    -- filter=76 channel=83
    -3, 0, -7, -4, 6, 1, 5, -6, 2,
    -- filter=76 channel=84
    0, 5, -3, -2, 7, -3, 4, -4, -1,
    -- filter=76 channel=85
    -6, -4, -5, 5, 5, -3, -5, 6, 3,
    -- filter=76 channel=86
    1, -5, -2, -6, -4, -6, 3, 0, 1,
    -- filter=76 channel=87
    -2, 3, 1, 0, -3, 0, 0, -4, 4,
    -- filter=76 channel=88
    -4, 4, -3, -5, -3, -4, 6, -3, 3,
    -- filter=76 channel=89
    3, -5, -5, 6, -5, 0, 7, 1, -1,
    -- filter=76 channel=90
    5, 8, 6, -5, 4, 5, 7, 1, -6,
    -- filter=76 channel=91
    2, -8, -5, -4, -2, 2, -2, -4, -4,
    -- filter=76 channel=92
    5, -5, 0, 0, -2, -7, 1, 6, 0,
    -- filter=76 channel=93
    -8, 0, 5, 6, -5, 2, 3, 0, -4,
    -- filter=76 channel=94
    -4, 3, 4, 0, 5, -6, 3, 7, 4,
    -- filter=76 channel=95
    -4, -6, -4, 1, 0, 1, -3, 6, 1,
    -- filter=76 channel=96
    -4, 7, -6, 0, -3, -3, 2, -5, -3,
    -- filter=76 channel=97
    -4, 2, -4, -6, 5, -6, 0, 3, -1,
    -- filter=76 channel=98
    -1, -5, 0, 5, -8, -6, 0, 0, -8,
    -- filter=76 channel=99
    -8, 1, -4, -4, -4, 0, 6, 5, 4,
    -- filter=76 channel=100
    -4, 3, 2, 7, -2, 2, 6, -3, 2,
    -- filter=76 channel=101
    -5, -5, 6, -4, 6, -2, 5, -3, -1,
    -- filter=76 channel=102
    6, -6, -2, -6, -3, 0, 5, -4, -3,
    -- filter=76 channel=103
    -6, -8, 6, 3, 2, 0, 0, -4, 2,
    -- filter=76 channel=104
    -7, -2, -2, 5, -3, -2, 5, -8, 0,
    -- filter=76 channel=105
    -2, -5, 2, -4, -3, -2, 3, 5, -5,
    -- filter=76 channel=106
    2, 2, -1, -5, -2, -5, 0, 5, -1,
    -- filter=76 channel=107
    -1, 1, 3, 0, -1, 7, -3, -5, 4,
    -- filter=76 channel=108
    -2, -5, -4, 3, 6, -3, 5, 0, 4,
    -- filter=76 channel=109
    -3, 4, -5, 0, 0, -1, -3, -2, 5,
    -- filter=76 channel=110
    3, -5, -7, -7, 6, -5, 5, 3, 2,
    -- filter=76 channel=111
    6, 5, -6, -4, 4, 6, 1, 0, 7,
    -- filter=76 channel=112
    3, 1, -6, 4, -4, 0, -2, 0, -1,
    -- filter=76 channel=113
    -6, -7, 0, -5, 0, 0, 6, 2, -6,
    -- filter=76 channel=114
    3, -5, 6, 5, 1, -5, -2, 5, 4,
    -- filter=76 channel=115
    6, 2, 5, 6, 6, 0, 1, 0, 6,
    -- filter=76 channel=116
    4, -7, 4, 2, 1, 1, 0, 5, 2,
    -- filter=76 channel=117
    5, 6, 6, 6, -7, 0, 0, 1, 6,
    -- filter=76 channel=118
    -3, 6, 1, -4, 0, 3, 2, -4, -5,
    -- filter=76 channel=119
    -2, -3, 4, 1, 4, 3, 1, -1, -1,
    -- filter=76 channel=120
    -10, -6, 3, -2, -1, 2, 1, 3, -6,
    -- filter=76 channel=121
    -6, -3, -2, -5, -3, 1, 5, -2, 6,
    -- filter=76 channel=122
    -6, 3, 2, 0, -2, -1, 0, -1, 6,
    -- filter=76 channel=123
    -4, 4, 0, -4, -3, -7, 5, -3, 5,
    -- filter=76 channel=124
    6, -3, 1, -5, 2, 0, 3, 3, -5,
    -- filter=76 channel=125
    -7, -8, -1, 0, -5, 2, -6, -1, 1,
    -- filter=76 channel=126
    -4, 1, -2, 0, -5, 1, 7, 2, 3,
    -- filter=76 channel=127
    -4, 0, 1, -5, 5, -1, 4, 5, 4,
    -- filter=77 channel=0
    0, 0, -7, 4, -11, -4, 3, -4, -11,
    -- filter=77 channel=1
    -5, -3, -10, 2, -6, -4, -7, -8, -1,
    -- filter=77 channel=2
    -5, 7, -5, -5, -2, 5, 0, 1, -2,
    -- filter=77 channel=3
    -2, 0, 0, -1, -8, -1, -7, -3, 0,
    -- filter=77 channel=4
    -11, 4, 0, -4, 0, 0, -4, 5, 10,
    -- filter=77 channel=5
    9, -6, -6, 11, 0, -5, 11, 0, -7,
    -- filter=77 channel=6
    -8, -7, -4, 2, 1, 2, -2, -7, -2,
    -- filter=77 channel=7
    4, 0, 0, -3, -1, 1, 5, 0, 3,
    -- filter=77 channel=8
    0, -4, -4, 5, 7, 2, 1, 4, -2,
    -- filter=77 channel=9
    -6, 2, -4, 4, 0, -1, -4, 7, 0,
    -- filter=77 channel=10
    -9, 8, 1, -10, 0, -1, -14, 0, 5,
    -- filter=77 channel=11
    0, 0, 4, -10, 2, -1, -9, -5, -3,
    -- filter=77 channel=12
    -8, -5, 3, 6, 0, 2, 0, 6, -3,
    -- filter=77 channel=13
    -8, 2, 7, -17, -1, -4, -8, -6, -1,
    -- filter=77 channel=14
    -4, 7, -1, 3, -1, 3, 6, -3, -6,
    -- filter=77 channel=15
    0, -4, -5, -13, -4, 3, -6, -6, 2,
    -- filter=77 channel=16
    4, 1, 3, 3, 10, 5, -1, 5, 0,
    -- filter=77 channel=17
    3, 5, 2, -3, -1, 6, 6, 0, -2,
    -- filter=77 channel=18
    -14, -9, 2, -15, -4, -8, -14, -6, -1,
    -- filter=77 channel=19
    -5, -1, -2, -6, -4, -6, -3, -3, -4,
    -- filter=77 channel=20
    -1, -6, 2, -9, 0, 0, -3, -9, 2,
    -- filter=77 channel=21
    -6, 3, -5, 5, 18, -7, 3, 14, 0,
    -- filter=77 channel=22
    3, -9, 5, -6, 0, 6, -2, -7, -1,
    -- filter=77 channel=23
    -8, 3, 5, -16, -7, 9, -8, 0, 4,
    -- filter=77 channel=24
    0, -6, -4, -3, -3, -2, 2, -6, 1,
    -- filter=77 channel=25
    -14, 2, 1, -12, -4, 0, -4, 0, 6,
    -- filter=77 channel=26
    6, 5, 0, 1, 4, -6, 10, 0, -1,
    -- filter=77 channel=27
    -4, -5, 1, -15, -8, 3, -4, -11, 8,
    -- filter=77 channel=28
    -7, 5, -1, 4, 0, -3, 5, 0, 1,
    -- filter=77 channel=29
    -3, 0, 5, -10, -9, 4, 1, -3, -3,
    -- filter=77 channel=30
    -2, -6, 0, -8, -4, 3, 0, 0, 6,
    -- filter=77 channel=31
    2, 17, 2, 1, 19, -6, -2, 5, 7,
    -- filter=77 channel=32
    -2, 3, 5, -15, -7, 1, -10, -14, 2,
    -- filter=77 channel=33
    -8, 5, -4, -4, 2, 0, -6, -2, -7,
    -- filter=77 channel=34
    7, 4, 6, 5, 3, 0, 7, -1, 4,
    -- filter=77 channel=35
    4, 2, 1, 5, 0, -3, -4, -5, -4,
    -- filter=77 channel=36
    3, 9, 6, 2, 0, -1, -6, -1, -7,
    -- filter=77 channel=37
    -4, 0, -10, 5, -5, -5, -4, -1, -2,
    -- filter=77 channel=38
    -1, -4, 7, -7, 2, -5, -4, 6, 2,
    -- filter=77 channel=39
    4, 5, 5, 1, 4, -7, -5, 5, 1,
    -- filter=77 channel=40
    0, 3, 7, -7, 3, -1, 2, -6, 1,
    -- filter=77 channel=41
    -11, 2, 2, -11, 0, 0, -13, -5, -3,
    -- filter=77 channel=42
    -6, 2, -1, 0, 6, -7, 3, -7, 2,
    -- filter=77 channel=43
    -10, -4, 8, -1, -7, -3, 4, -5, -4,
    -- filter=77 channel=44
    -2, -3, -1, -4, 2, -1, 3, -1, 1,
    -- filter=77 channel=45
    2, -4, -1, 0, -1, 0, -4, -4, -7,
    -- filter=77 channel=46
    0, 4, 1, 0, 5, 4, 0, -7, -2,
    -- filter=77 channel=47
    2, 12, -9, 6, 18, -1, -2, 11, 1,
    -- filter=77 channel=48
    -7, -2, -8, -6, 8, -4, -8, 0, -3,
    -- filter=77 channel=49
    -4, 2, -4, -14, -8, -2, -13, -3, -1,
    -- filter=77 channel=50
    -2, 5, -4, -5, 1, 0, 0, 0, -6,
    -- filter=77 channel=51
    -6, 0, 3, 5, 5, 5, -2, -7, -5,
    -- filter=77 channel=52
    0, -1, -3, -5, 6, 9, 3, -4, 4,
    -- filter=77 channel=53
    0, 6, 7, 0, -7, 6, 0, 3, 7,
    -- filter=77 channel=54
    0, -5, -3, -5, 4, 0, 0, 3, -5,
    -- filter=77 channel=55
    -4, 3, 3, -8, -3, 6, -10, 0, -4,
    -- filter=77 channel=56
    -2, 2, 5, 1, 8, 7, 6, 1, 7,
    -- filter=77 channel=57
    1, -2, -3, 5, 0, 6, -3, -1, -5,
    -- filter=77 channel=58
    2, -7, -6, 5, 0, 3, -2, 6, 1,
    -- filter=77 channel=59
    -3, 9, 0, -2, 2, -8, -6, -1, -7,
    -- filter=77 channel=60
    -6, 1, 0, 2, -1, -3, 7, -1, -5,
    -- filter=77 channel=61
    0, -3, 7, 1, 2, 1, 3, 0, -6,
    -- filter=77 channel=62
    3, 4, -6, 2, 2, 3, 4, 0, -4,
    -- filter=77 channel=63
    5, 8, 3, 13, 9, -5, 0, 5, 7,
    -- filter=77 channel=64
    6, 1, -3, 7, 5, 0, -4, 0, 2,
    -- filter=77 channel=65
    -5, -6, 0, 6, -6, -3, 5, 1, 5,
    -- filter=77 channel=66
    -9, 1, 8, 6, 4, 4, -5, 0, 1,
    -- filter=77 channel=67
    -5, 2, 5, 0, 0, -2, -3, 4, -6,
    -- filter=77 channel=68
    -6, -6, -3, 0, -7, 3, -8, 0, -5,
    -- filter=77 channel=69
    5, 2, -6, 5, -5, -5, -5, -2, 0,
    -- filter=77 channel=70
    -3, -9, 10, -11, -6, 9, -13, -9, 1,
    -- filter=77 channel=71
    6, 1, 3, 0, 3, 0, 6, 4, -7,
    -- filter=77 channel=72
    -4, 2, -5, -6, 9, -7, -12, -1, 3,
    -- filter=77 channel=73
    -13, -7, -3, -12, 2, -5, -4, -8, -4,
    -- filter=77 channel=74
    0, -2, 10, 9, -2, 6, -1, 0, 7,
    -- filter=77 channel=75
    1, 0, 0, -4, 1, 2, -7, 6, -3,
    -- filter=77 channel=76
    -8, -7, 1, -6, 3, 8, -5, -7, -8,
    -- filter=77 channel=77
    0, -4, 6, 3, -5, -1, -3, 5, 2,
    -- filter=77 channel=78
    8, 10, 5, -1, 11, -5, -4, 4, 5,
    -- filter=77 channel=79
    -11, -10, 1, -27, -10, -1, -20, -11, 3,
    -- filter=77 channel=80
    -12, 3, 1, 2, 19, -2, 1, 15, 2,
    -- filter=77 channel=81
    -4, 7, -4, 1, 0, 4, 0, -1, -6,
    -- filter=77 channel=82
    -2, -6, 5, -7, 2, -5, 0, 0, -6,
    -- filter=77 channel=83
    0, -3, 6, -4, 4, -7, -1, 0, 5,
    -- filter=77 channel=84
    -10, 3, 7, -4, -2, 6, -9, -9, -2,
    -- filter=77 channel=85
    4, 0, -4, 0, -7, 4, 0, 3, 4,
    -- filter=77 channel=86
    0, 1, 0, -3, -7, 8, 5, 1, 4,
    -- filter=77 channel=87
    2, 0, 0, 1, 2, 8, 3, 0, -3,
    -- filter=77 channel=88
    -5, -1, -6, 9, 11, -3, 8, 5, 1,
    -- filter=77 channel=89
    -11, 4, -5, -19, -6, -6, -10, -1, 0,
    -- filter=77 channel=90
    2, 5, 7, 10, 13, 4, -4, 13, 2,
    -- filter=77 channel=91
    -15, -2, 3, -8, -11, -1, -11, -3, 0,
    -- filter=77 channel=92
    6, 4, 9, 3, -2, 0, -4, -4, 5,
    -- filter=77 channel=93
    -5, 2, -5, 6, 5, -11, -2, 1, 0,
    -- filter=77 channel=94
    -2, 0, -3, -4, -4, -1, -4, 5, -1,
    -- filter=77 channel=95
    -7, -2, -5, -7, 5, 3, -5, 6, 5,
    -- filter=77 channel=96
    -5, 3, -5, -7, -7, -3, 0, -7, 0,
    -- filter=77 channel=97
    5, 1, 3, -1, 9, 3, -2, 0, 4,
    -- filter=77 channel=98
    -4, 0, -2, -14, 3, -7, -12, 2, 2,
    -- filter=77 channel=99
    7, 11, 3, 4, 9, -2, -4, 6, 6,
    -- filter=77 channel=100
    -5, 0, -1, -2, -4, 5, -7, 0, 4,
    -- filter=77 channel=101
    -3, 3, 5, 0, 0, -3, 5, -7, -2,
    -- filter=77 channel=102
    1, 7, 1, 5, 2, -4, -4, -5, 0,
    -- filter=77 channel=103
    2, 0, -2, 11, 20, -7, 2, 9, 0,
    -- filter=77 channel=104
    0, 4, 1, 1, 16, -5, -8, 7, -5,
    -- filter=77 channel=105
    0, 4, 1, -8, 1, -4, -8, 0, -4,
    -- filter=77 channel=106
    -9, -3, 1, -4, -1, -8, -3, -3, 2,
    -- filter=77 channel=107
    -6, -4, -5, -2, -3, 7, -8, -4, -3,
    -- filter=77 channel=108
    -7, -4, 6, -1, -7, 3, 4, 6, -7,
    -- filter=77 channel=109
    -16, 5, -1, -9, -3, -5, -3, -3, 2,
    -- filter=77 channel=110
    0, 10, 1, -2, 9, 4, -7, 1, -6,
    -- filter=77 channel=111
    -8, -3, -5, 4, -6, -6, 0, 0, -5,
    -- filter=77 channel=112
    0, 0, -1, 2, -3, -1, 0, -1, 9,
    -- filter=77 channel=113
    -4, 2, 1, 0, 1, -1, 2, 9, -4,
    -- filter=77 channel=114
    -9, -5, -9, -15, -14, -7, -12, -7, 0,
    -- filter=77 channel=115
    0, -2, -2, 4, 6, 7, 3, 6, 3,
    -- filter=77 channel=116
    -13, -1, 2, -16, 2, -7, -14, -8, -2,
    -- filter=77 channel=117
    2, -5, -3, -10, 6, 3, -9, 0, 0,
    -- filter=77 channel=118
    -2, 3, -2, 5, 2, -1, -4, -3, 2,
    -- filter=77 channel=119
    7, -3, 6, 14, 0, 10, 9, 9, 5,
    -- filter=77 channel=120
    -10, 2, 8, -10, -3, -2, -6, -7, 4,
    -- filter=77 channel=121
    2, 7, -1, -2, 1, 4, 1, -1, 0,
    -- filter=77 channel=122
    8, 15, -7, 8, 31, -13, -2, 23, 0,
    -- filter=77 channel=123
    -2, -5, 10, 5, 6, -3, -1, 2, 7,
    -- filter=77 channel=124
    -4, 4, 7, -5, -3, 2, -7, 0, 4,
    -- filter=77 channel=125
    -3, 5, 3, -8, 9, 4, -16, 2, 6,
    -- filter=77 channel=126
    -4, -5, -5, -9, -6, 1, -5, 2, -6,
    -- filter=77 channel=127
    -7, 0, 3, -3, -3, 7, 0, 1, -5,
    -- filter=78 channel=0
    0, -18, -30, 10, -4, -25, 16, -1, -13,
    -- filter=78 channel=1
    2, -21, -22, 5, -18, -14, 14, 11, -10,
    -- filter=78 channel=2
    1, -1, 2, -5, 4, -2, -2, -3, 0,
    -- filter=78 channel=3
    -4, -13, 1, -1, -13, -1, 1, -4, -9,
    -- filter=78 channel=4
    0, -2, -8, 1, -20, -8, -3, -8, -7,
    -- filter=78 channel=5
    6, -10, -12, 5, 3, -6, 4, 3, -3,
    -- filter=78 channel=6
    -1, 8, 0, -5, 13, 10, 1, -7, 0,
    -- filter=78 channel=7
    2, -5, -3, -3, 1, -5, -2, 2, -2,
    -- filter=78 channel=8
    3, -4, 1, -4, 3, 4, 1, 0, 0,
    -- filter=78 channel=9
    4, -2, -5, 0, -2, -5, 0, -1, 4,
    -- filter=78 channel=10
    8, -5, 9, 1, 6, 0, -7, -6, 5,
    -- filter=78 channel=11
    -17, 7, 16, -2, 15, 24, -6, -12, -7,
    -- filter=78 channel=12
    0, -1, 4, 6, 3, -7, 3, 5, -3,
    -- filter=78 channel=13
    -8, 8, 0, -1, 3, 5, -4, -6, 2,
    -- filter=78 channel=14
    -5, 2, 3, 0, -1, 0, -4, 6, 7,
    -- filter=78 channel=15
    -6, 8, 13, -18, 4, 5, 0, 0, -16,
    -- filter=78 channel=16
    1, -2, -5, 10, 0, -13, 3, -5, 2,
    -- filter=78 channel=17
    -4, 5, -4, 5, -2, -7, 4, 0, 1,
    -- filter=78 channel=18
    -6, 5, 16, -7, 5, 12, -5, -1, -13,
    -- filter=78 channel=19
    3, 5, -1, 7, 2, 0, -2, -3, -4,
    -- filter=78 channel=20
    -13, 24, 37, -20, 25, 26, -19, -17, -6,
    -- filter=78 channel=21
    0, 0, -12, 10, -4, 2, 8, 6, 8,
    -- filter=78 channel=22
    -3, -8, 0, -6, -3, -2, 3, -4, -10,
    -- filter=78 channel=23
    -18, 15, 5, -11, 3, 5, -2, 0, -5,
    -- filter=78 channel=24
    -5, 0, -6, -2, -1, 3, -2, -6, 1,
    -- filter=78 channel=25
    5, -7, -5, 5, -8, -1, 3, 7, -2,
    -- filter=78 channel=26
    5, 3, -12, 0, 3, -6, 9, -3, -7,
    -- filter=78 channel=27
    0, -4, -1, 9, -7, 2, 0, 2, 2,
    -- filter=78 channel=28
    -1, -5, -1, 2, -5, 4, 0, -6, 7,
    -- filter=78 channel=29
    -9, 20, 38, -20, 26, 33, -23, -6, -2,
    -- filter=78 channel=30
    -4, -13, -2, -1, 1, -5, 7, 4, 1,
    -- filter=78 channel=31
    12, 8, 2, 0, -10, -7, 3, 10, 11,
    -- filter=78 channel=32
    -11, 0, 0, -10, 0, 6, -6, -9, -3,
    -- filter=78 channel=33
    1, -1, -4, -5, -5, -9, 4, -2, -4,
    -- filter=78 channel=34
    5, 10, 4, 5, 4, 5, 15, 3, -1,
    -- filter=78 channel=35
    -6, 6, 0, 4, 4, 1, -3, -5, 5,
    -- filter=78 channel=36
    3, 9, 12, 6, 0, 4, -1, 4, 5,
    -- filter=78 channel=37
    -6, -16, -23, 17, -6, -22, 10, 4, -6,
    -- filter=78 channel=38
    1, -3, 1, -3, 4, -4, -4, 0, -5,
    -- filter=78 channel=39
    -6, 12, 20, -1, 6, 6, -1, -9, -2,
    -- filter=78 channel=40
    1, 10, 4, -5, 5, 11, -10, -6, 0,
    -- filter=78 channel=41
    18, 7, 0, 1, 7, -11, 10, 23, 3,
    -- filter=78 channel=42
    8, 4, -10, 4, -8, -7, 7, -1, 8,
    -- filter=78 channel=43
    -4, -4, -3, -4, -6, -2, 0, 0, -10,
    -- filter=78 channel=44
    2, -14, -21, 12, -11, -8, 8, 1, 9,
    -- filter=78 channel=45
    4, 7, -5, -7, -2, 7, -1, 0, -4,
    -- filter=78 channel=46
    3, 5, -4, -2, -6, -8, 0, 5, 3,
    -- filter=78 channel=47
    6, -15, -13, 0, -9, -8, 3, 4, 7,
    -- filter=78 channel=48
    8, -17, -11, 6, -11, -11, 3, 0, 5,
    -- filter=78 channel=49
    -12, 9, 2, 0, 1, -4, -6, -7, -8,
    -- filter=78 channel=50
    3, -9, 4, 4, -8, 3, 8, 3, -5,
    -- filter=78 channel=51
    1, -1, 6, 7, -1, -3, -5, 1, -7,
    -- filter=78 channel=52
    -9, 5, 5, 3, 0, 5, -1, -1, 0,
    -- filter=78 channel=53
    -7, 14, 18, -8, 3, 14, -7, -5, -5,
    -- filter=78 channel=54
    -4, 0, 1, 0, -1, 3, 3, 5, -1,
    -- filter=78 channel=55
    -18, 20, 30, -8, 16, 15, -17, -11, 0,
    -- filter=78 channel=56
    4, -3, 3, 1, -6, 0, 1, -3, -7,
    -- filter=78 channel=57
    9, -5, 2, -2, -6, -3, 0, -5, 2,
    -- filter=78 channel=58
    7, -2, 1, 1, -4, -6, -2, 6, 1,
    -- filter=78 channel=59
    7, -6, -8, 1, -7, -3, -2, 10, 0,
    -- filter=78 channel=60
    -4, -3, 1, 6, -3, -1, 2, 2, 5,
    -- filter=78 channel=61
    -3, 0, 0, -2, 1, 9, -7, -7, 3,
    -- filter=78 channel=62
    -5, -3, -2, -5, 0, 2, -1, -5, 2,
    -- filter=78 channel=63
    7, 3, -6, 8, 4, 1, 1, 2, 0,
    -- filter=78 channel=64
    -5, 7, 3, -1, 2, 2, -6, -3, -4,
    -- filter=78 channel=65
    -5, -6, 7, 0, 4, 2, 2, 2, -6,
    -- filter=78 channel=66
    10, 1, 5, 12, 3, -5, -1, 9, 3,
    -- filter=78 channel=67
    -4, -2, -5, 0, -1, 0, -2, 6, 4,
    -- filter=78 channel=68
    3, 2, 4, -2, 3, -1, 6, -6, 5,
    -- filter=78 channel=69
    4, 0, 5, 1, 2, 1, -4, -3, 0,
    -- filter=78 channel=70
    -7, -5, 0, -4, 0, -7, 1, 0, -12,
    -- filter=78 channel=71
    4, -6, 0, 0, -8, -9, 0, 2, -2,
    -- filter=78 channel=72
    0, 0, 7, 7, 1, 1, 4, 7, 12,
    -- filter=78 channel=73
    -3, 9, 4, -3, 2, 5, 0, -5, 1,
    -- filter=78 channel=74
    4, 5, -2, 0, 6, 5, 4, 3, 0,
    -- filter=78 channel=75
    13, -16, -26, 6, -17, -19, 15, 13, -12,
    -- filter=78 channel=76
    -8, 24, 32, -16, 16, 24, -11, 0, -9,
    -- filter=78 channel=77
    -6, -5, 0, -6, 4, 5, 5, -1, 7,
    -- filter=78 channel=78
    8, -1, -5, 3, 10, -4, 7, 11, 5,
    -- filter=78 channel=79
    -2, 7, 1, -1, 11, 2, 3, 3, -7,
    -- filter=78 channel=80
    3, 0, 0, -2, -5, 2, -1, 6, 13,
    -- filter=78 channel=81
    -3, -1, -2, 4, -2, 3, -6, -5, 2,
    -- filter=78 channel=82
    2, 4, 3, -6, -4, -7, 4, 1, 2,
    -- filter=78 channel=83
    2, -4, -6, 0, -8, 0, -1, -6, -6,
    -- filter=78 channel=84
    -3, 8, 5, -9, 11, 4, -2, -9, -1,
    -- filter=78 channel=85
    7, 0, -5, 0, 6, 4, 1, -2, 0,
    -- filter=78 channel=86
    -2, 0, 0, 8, -4, 1, 5, 6, 0,
    -- filter=78 channel=87
    -2, 4, 10, 0, 9, 3, -6, 2, -3,
    -- filter=78 channel=88
    1, 8, -1, -7, -1, 0, -5, 4, 5,
    -- filter=78 channel=89
    -5, 1, 13, 2, 3, 6, -4, 0, -1,
    -- filter=78 channel=90
    1, 0, 0, -5, -1, 2, 2, 5, 0,
    -- filter=78 channel=91
    -7, -2, 9, 5, -3, 3, -4, -4, -6,
    -- filter=78 channel=92
    -5, 5, -5, -6, -6, -6, 0, -5, -5,
    -- filter=78 channel=93
    1, -21, -24, 8, -18, -12, 10, -2, -1,
    -- filter=78 channel=94
    2, -2, 2, -3, 6, 6, 5, -1, 2,
    -- filter=78 channel=95
    6, -6, -1, 1, 2, 2, 6, -6, -6,
    -- filter=78 channel=96
    6, 0, 4, 6, 4, -2, -4, -3, 6,
    -- filter=78 channel=97
    7, -6, 3, 5, -11, -2, 6, -2, -8,
    -- filter=78 channel=98
    1, -2, -3, -1, -3, -11, 3, 3, -3,
    -- filter=78 channel=99
    3, 14, 7, -10, 12, 4, -13, 4, -2,
    -- filter=78 channel=100
    0, 5, -5, 2, 2, -6, 7, 6, -4,
    -- filter=78 channel=101
    2, -11, 6, 3, -16, -2, 0, -5, 4,
    -- filter=78 channel=102
    -2, 4, 3, -6, 3, 1, 1, 6, -3,
    -- filter=78 channel=103
    -2, -9, -11, -2, -12, -15, 6, -3, 4,
    -- filter=78 channel=104
    6, 3, -7, 1, -8, -5, -2, 5, 1,
    -- filter=78 channel=105
    -15, 8, 14, -3, 20, 22, -7, -1, 4,
    -- filter=78 channel=106
    -4, 9, 12, -6, 3, 7, -2, -9, -9,
    -- filter=78 channel=107
    -11, 13, 11, -7, 8, -2, -4, -8, -15,
    -- filter=78 channel=108
    1, 0, -8, 8, -1, -5, 8, -2, 4,
    -- filter=78 channel=109
    -7, 1, 3, -5, 7, -3, 1, -6, 3,
    -- filter=78 channel=110
    8, 8, -4, 2, -3, 5, -3, 0, 7,
    -- filter=78 channel=111
    -7, -5, 8, -7, -4, -4, 8, 6, 0,
    -- filter=78 channel=112
    -2, -4, -6, -5, 0, -10, 6, 2, -5,
    -- filter=78 channel=113
    3, -7, -2, 1, -6, -2, -2, 4, 4,
    -- filter=78 channel=114
    -4, 5, 3, 2, 6, -10, 7, -1, -18,
    -- filter=78 channel=115
    0, -2, 0, -6, -6, 5, 2, -1, 4,
    -- filter=78 channel=116
    -7, 2, 4, 4, 5, -2, 1, -2, -1,
    -- filter=78 channel=117
    -2, 5, -7, -1, 7, -5, -4, 5, 1,
    -- filter=78 channel=118
    7, 6, 5, 3, 7, 0, 7, 4, 4,
    -- filter=78 channel=119
    7, -1, -2, 7, 9, 2, 4, 2, 1,
    -- filter=78 channel=120
    -19, 4, 12, -11, -3, -1, 0, -9, -15,
    -- filter=78 channel=121
    -1, -4, 5, 1, -4, -1, 0, -6, 3,
    -- filter=78 channel=122
    1, -25, -17, 4, -13, -17, 13, 11, 3,
    -- filter=78 channel=123
    -6, -1, 0, 6, -4, -6, 9, 6, -4,
    -- filter=78 channel=124
    -8, 10, 19, -2, 0, 15, -12, -7, -8,
    -- filter=78 channel=125
    -3, 3, 6, 1, 3, 0, 1, 7, 3,
    -- filter=78 channel=126
    2, -4, 3, -4, 5, 0, 7, -6, -8,
    -- filter=78 channel=127
    4, -5, -4, 5, 4, -1, 2, 9, -6,
    -- filter=79 channel=0
    -21, -3, -7, -23, 13, 15, -14, 0, 16,
    -- filter=79 channel=1
    -23, 4, 8, -21, 4, 14, -7, -2, 19,
    -- filter=79 channel=2
    -1, 2, -5, -5, -4, 0, -2, 4, -5,
    -- filter=79 channel=3
    -1, -3, 1, -13, -5, -4, 0, -10, -3,
    -- filter=79 channel=4
    -4, -6, -3, 1, -4, 1, -7, -4, -10,
    -- filter=79 channel=5
    -10, 11, 3, -14, 16, 10, -9, 20, 16,
    -- filter=79 channel=6
    7, -2, 0, 1, 0, -7, 7, -8, -7,
    -- filter=79 channel=7
    5, 0, 0, 6, 6, -1, -3, 4, 4,
    -- filter=79 channel=8
    -4, -6, 7, -2, 0, 0, 0, -3, 6,
    -- filter=79 channel=9
    3, 6, 2, -11, 11, 7, 1, 2, 1,
    -- filter=79 channel=10
    0, 5, 2, 6, 0, 0, 1, -1, 3,
    -- filter=79 channel=11
    4, -2, 9, 10, -16, -6, 6, -1, 1,
    -- filter=79 channel=12
    -2, 5, 7, 0, -2, 0, 1, 0, 0,
    -- filter=79 channel=13
    5, 0, 7, 11, -20, -4, 4, -8, -7,
    -- filter=79 channel=14
    6, 5, -4, 4, -3, 7, 5, -1, -5,
    -- filter=79 channel=15
    13, -8, -8, 10, -17, -13, 9, -6, -1,
    -- filter=79 channel=16
    -8, 3, 0, -7, 8, -4, -14, 13, 7,
    -- filter=79 channel=17
    1, -2, -1, -2, 1, -5, 6, 4, -2,
    -- filter=79 channel=18
    10, -11, -6, 4, -16, -7, 3, -7, 0,
    -- filter=79 channel=19
    -5, 5, 6, 0, 0, 0, -2, 3, -6,
    -- filter=79 channel=20
    26, -10, -6, 24, -9, -20, 11, -2, -8,
    -- filter=79 channel=21
    -1, 13, -2, 0, 21, -6, -11, 6, -1,
    -- filter=79 channel=22
    3, 1, 3, -2, 0, 2, 0, 7, 6,
    -- filter=79 channel=23
    8, -9, 4, 3, -1, -14, 12, 6, 0,
    -- filter=79 channel=24
    2, -2, 2, 0, 5, 0, 5, 1, -3,
    -- filter=79 channel=25
    -3, 3, -6, 0, 6, 2, -10, 6, -2,
    -- filter=79 channel=26
    -6, 5, 2, -11, 1, 1, -5, 0, 8,
    -- filter=79 channel=27
    -8, 4, 0, -11, 11, 1, -10, 4, 13,
    -- filter=79 channel=28
    -4, 2, 1, -5, -2, 2, 0, -2, 5,
    -- filter=79 channel=29
    23, -5, 6, 13, -11, -10, 14, -6, -4,
    -- filter=79 channel=30
    -14, 8, 8, -12, 0, 5, -9, 3, 8,
    -- filter=79 channel=31
    -2, 12, -3, -4, 14, -15, -16, 3, 0,
    -- filter=79 channel=32
    10, 0, 6, 4, -8, 3, 4, 0, -1,
    -- filter=79 channel=33
    1, 0, 6, -2, 7, 6, -11, -2, 2,
    -- filter=79 channel=34
    0, 9, 6, -3, 23, -7, 2, 19, 4,
    -- filter=79 channel=35
    1, 0, 3, 0, 5, 1, -5, -2, 1,
    -- filter=79 channel=36
    5, 3, -10, 1, 0, -9, -1, 0, -15,
    -- filter=79 channel=37
    -17, 0, 4, -25, 8, 20, -18, 10, 18,
    -- filter=79 channel=38
    -1, 7, -4, -4, 8, -2, 4, 3, -5,
    -- filter=79 channel=39
    7, -5, 4, 12, -4, 2, 10, -8, -10,
    -- filter=79 channel=40
    2, -8, 0, 1, -4, -13, 3, 0, -10,
    -- filter=79 channel=41
    4, -8, 11, 3, -16, 11, 0, 0, -5,
    -- filter=79 channel=42
    -9, -1, 10, -8, 3, 5, -10, -6, 11,
    -- filter=79 channel=43
    9, -11, 0, -5, -7, -1, -4, 1, 6,
    -- filter=79 channel=44
    -19, 2, 0, -26, 9, 10, -16, 9, 11,
    -- filter=79 channel=45
    0, -4, -3, -3, -1, 1, -2, -3, 1,
    -- filter=79 channel=46
    6, -4, -7, 4, 2, 1, -6, 1, -6,
    -- filter=79 channel=47
    -7, 9, -8, -13, 16, 12, -19, 11, 1,
    -- filter=79 channel=48
    -9, -3, 7, -17, 5, -1, -13, 5, 4,
    -- filter=79 channel=49
    1, -13, -6, -4, -7, -5, 1, -13, 4,
    -- filter=79 channel=50
    3, -6, 6, -10, 2, -6, 4, 2, -1,
    -- filter=79 channel=51
    5, 0, -1, 1, -5, 3, 7, -3, 7,
    -- filter=79 channel=52
    7, -3, 0, 6, 6, -6, -2, 3, -9,
    -- filter=79 channel=53
    1, 0, 6, 5, -7, -10, 11, 1, -7,
    -- filter=79 channel=54
    6, -5, -2, -2, -4, -2, 5, -5, 4,
    -- filter=79 channel=55
    15, -9, -8, 21, -17, -19, 14, -11, -13,
    -- filter=79 channel=56
    1, 6, -3, -1, 11, -4, 0, 0, -7,
    -- filter=79 channel=57
    -3, -8, -6, 5, 1, 5, 0, -1, -7,
    -- filter=79 channel=58
    -8, 7, 0, -11, 10, 5, -5, 2, 4,
    -- filter=79 channel=59
    -7, 3, -4, -2, 2, 4, -4, 3, 4,
    -- filter=79 channel=60
    -4, -2, 3, -4, 2, 0, -4, -3, 3,
    -- filter=79 channel=61
    5, -2, 4, 11, 2, -3, 3, 8, 0,
    -- filter=79 channel=62
    5, 4, 3, -5, 1, 5, -3, 0, 6,
    -- filter=79 channel=63
    -3, 7, 4, -3, 7, 10, -9, 11, 10,
    -- filter=79 channel=64
    1, -8, -7, 4, -1, -6, -3, -1, -9,
    -- filter=79 channel=65
    1, 4, 2, 2, 3, -6, -6, 6, -5,
    -- filter=79 channel=66
    4, -2, 7, 10, -4, 6, 1, -6, -3,
    -- filter=79 channel=67
    -2, 0, 0, -4, 2, -3, 3, -2, -5,
    -- filter=79 channel=68
    2, -3, -2, 2, -11, 2, -4, -10, -2,
    -- filter=79 channel=69
    0, -2, 2, -2, -2, 7, -3, -6, -5,
    -- filter=79 channel=70
    -6, 4, 5, 1, -11, 4, -4, -10, 0,
    -- filter=79 channel=71
    6, -8, -4, 4, -6, -6, -6, -1, 0,
    -- filter=79 channel=72
    10, 5, -9, 0, -4, -4, -1, -8, -1,
    -- filter=79 channel=73
    -2, -6, 3, 6, -8, -7, 10, 0, -10,
    -- filter=79 channel=74
    1, 0, -3, 1, 16, -6, 0, 0, -1,
    -- filter=79 channel=75
    -19, 5, -3, -16, 18, 29, -10, 0, 23,
    -- filter=79 channel=76
    14, -6, -7, 18, -15, -19, 20, -4, -9,
    -- filter=79 channel=77
    -4, -4, 0, 4, 3, -3, 4, 3, -1,
    -- filter=79 channel=78
    -3, 8, 2, -14, 5, 9, -12, 8, 6,
    -- filter=79 channel=79
    3, -8, -1, 4, -13, 1, 2, -11, 3,
    -- filter=79 channel=80
    -4, 7, 1, -3, 4, 2, -16, -4, -1,
    -- filter=79 channel=81
    4, -5, 3, 4, 1, -4, 7, -4, -4,
    -- filter=79 channel=82
    3, 1, 2, 2, -7, 1, -2, 4, -6,
    -- filter=79 channel=83
    -1, 6, 3, -8, 5, -5, -10, 8, 6,
    -- filter=79 channel=84
    -3, -2, 1, -2, -11, 7, 3, -5, 2,
    -- filter=79 channel=85
    -2, 0, 0, 1, -1, 1, 0, 1, 2,
    -- filter=79 channel=86
    1, 9, 5, -8, 4, 0, -4, -2, 12,
    -- filter=79 channel=87
    12, 1, 7, 3, -1, -1, 6, -3, -3,
    -- filter=79 channel=88
    -2, 3, -1, 0, 8, -9, 0, -1, -16,
    -- filter=79 channel=89
    12, -15, 0, 13, -11, -5, 11, -13, -10,
    -- filter=79 channel=90
    -3, 0, -6, -3, 4, -4, 4, -8, -15,
    -- filter=79 channel=91
    -8, 0, 7, -2, -6, 7, 6, -6, 3,
    -- filter=79 channel=92
    0, -4, 6, 5, 3, -1, 0, 3, 1,
    -- filter=79 channel=93
    -13, 3, 7, -19, 17, 12, -18, 5, 14,
    -- filter=79 channel=94
    2, -4, 4, 3, 2, 7, 2, 3, 7,
    -- filter=79 channel=95
    5, 4, 7, 1, -1, 3, 2, -1, 0,
    -- filter=79 channel=96
    -5, 0, 3, 4, -3, 6, -4, -3, 8,
    -- filter=79 channel=97
    -3, 4, -1, -2, -7, -2, -5, 0, 7,
    -- filter=79 channel=98
    -8, 5, 5, -14, -6, 9, 0, -3, 8,
    -- filter=79 channel=99
    13, 13, 0, 12, 13, -3, 12, 11, 0,
    -- filter=79 channel=100
    0, -2, 8, -2, 0, -4, 1, -4, 5,
    -- filter=79 channel=101
    -1, -1, 5, -7, -12, -6, -1, -5, -5,
    -- filter=79 channel=102
    1, 7, -4, -4, 5, 4, 2, 0, 6,
    -- filter=79 channel=103
    -12, 12, -12, -12, 15, 6, -15, 12, 5,
    -- filter=79 channel=104
    -3, 7, 1, -6, 10, -1, -8, 1, 0,
    -- filter=79 channel=105
    19, -3, -2, 5, -11, -8, 11, 5, 0,
    -- filter=79 channel=106
    4, 3, -2, 7, -12, -4, 3, -7, -7,
    -- filter=79 channel=107
    10, -8, -3, 5, -17, -9, 3, -1, -5,
    -- filter=79 channel=108
    0, 5, 0, 6, 1, -4, 2, 6, -3,
    -- filter=79 channel=109
    6, 9, -3, -4, 5, 3, -2, 8, -2,
    -- filter=79 channel=110
    3, 0, 0, 0, -6, -2, 0, -2, 8,
    -- filter=79 channel=111
    0, 6, -8, 4, 4, -6, 7, 7, -1,
    -- filter=79 channel=112
    -10, -3, -1, -8, 13, 5, -8, 10, 1,
    -- filter=79 channel=113
    0, 5, -5, -7, 3, -2, 1, 0, 9,
    -- filter=79 channel=114
    0, -2, -7, -2, 1, 3, -3, 0, 12,
    -- filter=79 channel=115
    1, 2, -3, -1, 0, -1, -3, 5, -2,
    -- filter=79 channel=116
    -3, 3, -5, 5, -6, -8, 3, 2, -8,
    -- filter=79 channel=117
    -5, 4, -3, 0, -2, -4, 7, -5, -9,
    -- filter=79 channel=118
    -2, -5, -1, -3, 1, -4, 0, -3, 0,
    -- filter=79 channel=119
    7, 12, 0, 9, 20, -6, 1, 16, -5,
    -- filter=79 channel=120
    6, -4, 7, -3, 4, -4, 0, -2, 1,
    -- filter=79 channel=121
    8, 5, 1, 10, -6, 0, 4, 0, 3,
    -- filter=79 channel=122
    -12, 25, -5, -19, 36, -2, -26, 18, -7,
    -- filter=79 channel=123
    -2, -4, -3, -4, 7, -3, 6, 8, 0,
    -- filter=79 channel=124
    6, 5, -2, 7, -9, -8, 7, -1, -4,
    -- filter=79 channel=125
    -2, -1, -6, 0, 8, 1, -4, 2, -1,
    -- filter=79 channel=126
    4, -12, -2, 3, -13, 4, 6, -7, 3,
    -- filter=79 channel=127
    6, 1, -6, 3, -7, -2, 4, -3, 0,
    -- filter=80 channel=0
    -9, 11, -2, -19, 13, 8, -12, 11, -3,
    -- filter=80 channel=1
    -6, 7, -6, -6, 25, -11, -2, 16, -7,
    -- filter=80 channel=2
    -2, 0, 4, 7, 1, 6, 0, 0, 2,
    -- filter=80 channel=3
    -2, 0, -1, 0, 6, 3, 2, 3, -2,
    -- filter=80 channel=4
    6, 0, 4, 5, 3, 0, -4, 7, 7,
    -- filter=80 channel=5
    1, 15, -9, 5, 24, -6, 4, 20, -3,
    -- filter=80 channel=6
    -5, -6, 8, -1, 3, -1, 0, 6, -1,
    -- filter=80 channel=7
    -5, 6, 7, 0, -3, -6, 4, -7, -4,
    -- filter=80 channel=8
    1, -6, 11, -4, 5, 11, 1, -7, 2,
    -- filter=80 channel=9
    -1, 0, 5, 0, -1, 4, -1, -6, -7,
    -- filter=80 channel=10
    0, 4, -1, 1, 3, -7, 0, -5, 0,
    -- filter=80 channel=11
    4, -1, 0, 1, -12, 9, 0, -7, 12,
    -- filter=80 channel=12
    -1, 3, 0, 0, 10, -3, 2, 6, -1,
    -- filter=80 channel=13
    0, 0, 5, -9, 1, 3, 0, 1, -8,
    -- filter=80 channel=14
    4, -3, 2, 5, 2, 0, -1, -5, 3,
    -- filter=80 channel=15
    0, 0, 2, 4, -7, 6, -1, 0, 1,
    -- filter=80 channel=16
    5, 8, -6, 6, 12, -11, -6, 9, -4,
    -- filter=80 channel=17
    6, 1, -3, 3, -5, -1, 5, -3, -5,
    -- filter=80 channel=18
    4, 1, 5, -6, 0, -2, -2, -1, 6,
    -- filter=80 channel=19
    -1, -4, 6, 1, 3, -6, -6, -6, 6,
    -- filter=80 channel=20
    3, -9, 7, 0, -16, 13, 1, -6, 12,
    -- filter=80 channel=21
    -4, 5, -7, 4, 1, -14, 6, 5, -14,
    -- filter=80 channel=22
    1, 3, 2, 0, 6, -3, 4, 5, -3,
    -- filter=80 channel=23
    1, -3, 12, 3, -16, 11, 7, -18, 24,
    -- filter=80 channel=24
    -3, 2, 4, -7, -5, 2, 3, 2, 0,
    -- filter=80 channel=25
    -4, -3, -12, 3, 11, -7, 6, -1, -4,
    -- filter=80 channel=26
    4, 6, -7, -4, 4, -5, 0, 2, -6,
    -- filter=80 channel=27
    4, -7, -1, 4, -16, 6, 4, -11, 11,
    -- filter=80 channel=28
    5, -4, 2, 2, 5, 1, -3, 6, -5,
    -- filter=80 channel=29
    0, -1, 6, 0, -12, 15, 5, -2, 14,
    -- filter=80 channel=30
    -5, -4, -6, 6, 0, 5, 2, 0, -1,
    -- filter=80 channel=31
    9, -8, 3, 11, -8, 7, 4, -12, -3,
    -- filter=80 channel=32
    -7, -6, 4, 5, 2, -1, 8, 3, 6,
    -- filter=80 channel=33
    -6, -6, 3, -2, -1, -4, -5, -10, 5,
    -- filter=80 channel=34
    -8, -11, 6, -8, -3, 17, 3, -6, 16,
    -- filter=80 channel=35
    0, 2, 3, -2, 1, 7, 6, -6, -1,
    -- filter=80 channel=36
    3, 5, -3, -7, -2, -3, -1, -6, 0,
    -- filter=80 channel=37
    -3, 0, -12, -6, 21, -1, -7, 6, 3,
    -- filter=80 channel=38
    -2, 0, -3, 9, -1, -6, -2, -4, 6,
    -- filter=80 channel=39
    -5, 0, -1, 0, -1, -2, 8, 5, 0,
    -- filter=80 channel=40
    5, 3, 6, -4, -4, 3, -5, 2, 8,
    -- filter=80 channel=41
    3, 10, -7, -13, 6, -11, -9, 8, -14,
    -- filter=80 channel=42
    -9, 0, -3, -2, 8, 0, -5, 9, -4,
    -- filter=80 channel=43
    2, 2, -2, 0, 1, 2, -1, 6, 8,
    -- filter=80 channel=44
    3, 10, -10, -3, 10, -7, -8, 0, 0,
    -- filter=80 channel=45
    7, 0, -5, 0, 6, -6, 0, 3, -7,
    -- filter=80 channel=46
    -1, -2, 0, -4, 1, 0, -6, 4, -7,
    -- filter=80 channel=47
    -1, 7, -15, 6, 23, -8, 7, 6, -6,
    -- filter=80 channel=48
    3, -1, -6, 11, 4, -5, -2, 2, -5,
    -- filter=80 channel=49
    -4, 2, 8, -1, -4, 9, 0, 0, 9,
    -- filter=80 channel=50
    1, -9, -6, 1, -14, 3, 0, -13, -3,
    -- filter=80 channel=51
    0, -4, -4, 6, -2, -7, 0, 1, 0,
    -- filter=80 channel=52
    1, -8, 6, -3, 0, 1, -1, -4, 11,
    -- filter=80 channel=53
    2, -6, 3, 7, -3, 9, 4, 4, 6,
    -- filter=80 channel=54
    -4, 5, -6, -4, 3, 5, 1, 4, -3,
    -- filter=80 channel=55
    -2, -5, 1, -5, -20, -1, 5, -7, 3,
    -- filter=80 channel=56
    7, -6, 0, 6, -6, -3, -5, -6, 3,
    -- filter=80 channel=57
    -7, -5, 0, 2, 4, -1, 0, 0, 1,
    -- filter=80 channel=58
    -1, 0, -5, -4, 11, 6, -5, 17, 2,
    -- filter=80 channel=59
    2, 4, -11, 7, 0, -13, 2, -2, -15,
    -- filter=80 channel=60
    0, 3, -4, 0, 5, 0, -2, 2, 4,
    -- filter=80 channel=61
    5, 5, 7, 0, 0, 10, -7, 0, 2,
    -- filter=80 channel=62
    2, -4, 7, 7, -7, -2, 3, 0, 0,
    -- filter=80 channel=63
    -4, 11, -4, 2, 10, 3, 1, 4, 3,
    -- filter=80 channel=64
    4, -7, -3, 0, -8, 1, -2, -5, -2,
    -- filter=80 channel=65
    -6, 0, -6, -7, 2, 4, -7, 3, 1,
    -- filter=80 channel=66
    -9, -1, 2, -10, 6, 3, -8, 4, -9,
    -- filter=80 channel=67
    -6, 3, 6, 0, -1, -4, 6, -5, 7,
    -- filter=80 channel=68
    1, 1, 0, 5, -8, 0, -1, -3, -2,
    -- filter=80 channel=69
    -5, 7, -6, -2, 10, 1, -1, 2, -5,
    -- filter=80 channel=70
    0, -6, 3, -2, -14, 14, 0, -13, 5,
    -- filter=80 channel=71
    0, 1, -3, 0, 1, 0, 4, -8, 4,
    -- filter=80 channel=72
    -4, 4, 6, 8, -10, -4, 2, -1, 0,
    -- filter=80 channel=73
    -1, -7, 0, 6, -10, 7, -4, -4, 6,
    -- filter=80 channel=74
    1, -4, 1, 7, -17, 8, -4, -12, 13,
    -- filter=80 channel=75
    -12, 12, -14, -13, 32, -4, -10, 9, -6,
    -- filter=80 channel=76
    -4, -5, 10, -1, -9, 4, -4, -3, 2,
    -- filter=80 channel=77
    1, -4, -5, -4, -4, 4, 4, 6, -6,
    -- filter=80 channel=78
    -4, 9, 0, -2, 1, 2, 0, 0, 9,
    -- filter=80 channel=79
    -1, -4, -6, -9, -11, 6, 4, -1, 9,
    -- filter=80 channel=80
    -5, 4, -10, 7, 7, -3, 2, -5, -15,
    -- filter=80 channel=81
    3, -6, -6, 3, 1, -3, 1, -7, 0,
    -- filter=80 channel=82
    3, 5, 1, -3, 2, -3, 2, -1, -2,
    -- filter=80 channel=83
    4, -6, -1, 7, -6, 0, 6, -3, -4,
    -- filter=80 channel=84
    -7, 1, 10, -3, -1, 7, 0, -3, 9,
    -- filter=80 channel=85
    3, 1, -2, 1, 6, 4, -2, 7, -4,
    -- filter=80 channel=86
    -4, 6, 1, -1, 4, 9, -3, 0, 9,
    -- filter=80 channel=87
    -2, 2, 6, -6, 2, 6, 4, -6, 1,
    -- filter=80 channel=88
    6, 4, -1, 6, -2, 4, -7, 0, 2,
    -- filter=80 channel=89
    3, 0, -2, -8, -5, -6, -5, -10, -2,
    -- filter=80 channel=90
    -1, 2, -1, 0, -2, 0, -2, -9, 7,
    -- filter=80 channel=91
    -6, -2, 1, 2, -11, 6, 1, -7, 10,
    -- filter=80 channel=92
    2, 2, 6, -7, 1, 2, 2, -7, 10,
    -- filter=80 channel=93
    -10, 10, -3, -5, 19, 3, -1, 14, -4,
    -- filter=80 channel=94
    0, 4, 2, -6, -2, -1, -3, 4, -2,
    -- filter=80 channel=95
    -3, 0, 1, -2, -1, 6, -4, 3, -5,
    -- filter=80 channel=96
    4, 3, -8, 0, 4, 5, -7, -2, -8,
    -- filter=80 channel=97
    -7, -7, -7, -5, 0, -3, -6, -6, 6,
    -- filter=80 channel=98
    2, -1, -4, -1, 5, 1, 8, -5, -5,
    -- filter=80 channel=99
    -2, -9, 12, 6, -14, 13, -1, -15, 17,
    -- filter=80 channel=100
    6, 3, 1, 3, 5, -3, 1, 2, -3,
    -- filter=80 channel=101
    2, 0, -3, 6, 2, -5, 1, 3, 0,
    -- filter=80 channel=102
    2, -2, 3, 0, 5, -1, -2, 0, -4,
    -- filter=80 channel=103
    -5, 9, -6, 12, 14, -10, -1, 2, -12,
    -- filter=80 channel=104
    0, -5, -3, 4, -2, 0, 10, -4, -10,
    -- filter=80 channel=105
    7, 4, 6, -6, -11, 0, 5, -8, 8,
    -- filter=80 channel=106
    -3, -2, 6, -2, -9, -4, -3, -8, 0,
    -- filter=80 channel=107
    1, -7, 10, -4, 0, 9, 2, 1, 10,
    -- filter=80 channel=108
    3, 0, -2, -8, 5, 4, 0, 9, 4,
    -- filter=80 channel=109
    6, -2, 0, 12, -5, 2, 4, -10, 4,
    -- filter=80 channel=110
    -3, -5, 10, 0, -4, 11, -1, 1, 10,
    -- filter=80 channel=111
    0, 0, -2, 4, 6, 1, 5, 0, -8,
    -- filter=80 channel=112
    4, -8, 0, 2, 1, 6, -3, 0, 6,
    -- filter=80 channel=113
    -2, -9, -5, -1, -10, 2, -1, 1, 1,
    -- filter=80 channel=114
    -3, 0, 2, -5, 5, 3, 3, 5, 11,
    -- filter=80 channel=115
    2, 7, -4, -7, -4, 0, 2, 2, 0,
    -- filter=80 channel=116
    3, 5, -5, 3, -1, -1, 11, -9, -4,
    -- filter=80 channel=117
    -3, 7, 4, -6, 5, 0, -1, -5, 0,
    -- filter=80 channel=118
    1, 4, -2, 0, -4, -3, 0, -3, 3,
    -- filter=80 channel=119
    7, -6, 8, 7, -7, 0, 4, -2, 6,
    -- filter=80 channel=120
    -2, -9, 13, 9, -23, 17, 12, -20, 14,
    -- filter=80 channel=121
    0, 2, -4, -1, -2, -5, 6, 4, 2,
    -- filter=80 channel=122
    0, 12, -18, 3, 19, -11, 4, 5, -14,
    -- filter=80 channel=123
    5, 0, 4, -4, 2, 0, 1, -2, 10,
    -- filter=80 channel=124
    3, 4, 0, -3, -7, 8, -4, -5, -1,
    -- filter=80 channel=125
    8, 0, -2, 10, -13, -2, 3, -12, 3,
    -- filter=80 channel=126
    -4, -3, 1, 2, 10, -6, 6, -4, 0,
    -- filter=80 channel=127
    -2, -2, -2, 0, 0, -5, 2, 5, 5,
    -- filter=81 channel=0
    7, 11, 8, 10, 15, 7, 2, 18, 9,
    -- filter=81 channel=1
    5, 2, 6, 7, 4, 0, 7, 12, 12,
    -- filter=81 channel=2
    -2, 5, 1, -1, 0, 4, 9, 5, 4,
    -- filter=81 channel=3
    7, 13, 0, -10, -7, 1, 2, 4, -2,
    -- filter=81 channel=4
    1, 1, 3, 8, 1, 1, 13, 13, 12,
    -- filter=81 channel=5
    3, -4, 8, 8, 0, 5, -1, 3, 11,
    -- filter=81 channel=6
    4, 0, 4, 7, 16, 8, 0, 11, 1,
    -- filter=81 channel=7
    -6, -3, 0, 0, -5, -6, 7, 1, -2,
    -- filter=81 channel=8
    1, 0, -4, -6, -4, 6, 2, 6, 3,
    -- filter=81 channel=9
    -8, 0, 3, -6, 0, -10, 1, -1, -9,
    -- filter=81 channel=10
    0, -5, 3, -3, -9, 2, 4, -13, -3,
    -- filter=81 channel=11
    -7, 11, 8, 9, 3, -4, 5, 6, -1,
    -- filter=81 channel=12
    10, 5, 2, 7, 2, 0, -1, -6, 9,
    -- filter=81 channel=13
    -1, -7, 5, -1, -11, -2, 3, 4, -2,
    -- filter=81 channel=14
    -4, 0, -3, 1, 0, -6, -3, -2, -1,
    -- filter=81 channel=15
    -11, -2, -4, 5, -2, -11, 3, 6, -9,
    -- filter=81 channel=16
    0, -1, 4, -1, -8, 9, 2, 3, 3,
    -- filter=81 channel=17
    -2, -2, -6, -5, -6, 3, 2, 0, -5,
    -- filter=81 channel=18
    -1, 1, 3, 10, -1, -6, 8, 13, -10,
    -- filter=81 channel=19
    -2, -1, 2, -3, 4, -4, 0, 5, 0,
    -- filter=81 channel=20
    -6, 6, 14, 15, 22, 6, 0, 16, 0,
    -- filter=81 channel=21
    -8, -4, -3, 0, -11, 2, -4, -6, 1,
    -- filter=81 channel=22
    1, 2, -5, -5, 8, 3, 6, -1, -1,
    -- filter=81 channel=23
    -3, 5, -5, -2, -11, -12, 0, -9, -18,
    -- filter=81 channel=24
    5, -6, -2, -4, 5, 8, -2, 0, 7,
    -- filter=81 channel=25
    -11, -2, 0, 0, -13, -14, -3, 0, -9,
    -- filter=81 channel=26
    7, -1, -5, 1, -3, 6, 8, 3, 6,
    -- filter=81 channel=27
    -15, -7, -20, -11, -27, -23, 3, -13, -26,
    -- filter=81 channel=28
    6, -7, -3, 7, 0, -5, -6, -6, 6,
    -- filter=81 channel=29
    1, 9, -1, 10, 9, -1, -2, 13, -1,
    -- filter=81 channel=30
    -7, 1, 0, 0, -4, 0, 0, -6, 0,
    -- filter=81 channel=31
    -11, -12, -4, -2, -12, -3, -1, -7, -15,
    -- filter=81 channel=32
    -7, -8, -3, 0, -7, -5, 12, 5, -8,
    -- filter=81 channel=33
    -12, -9, -2, -2, -13, -2, -4, -5, -6,
    -- filter=81 channel=34
    5, 0, -2, -1, -2, -1, -1, -3, 0,
    -- filter=81 channel=35
    1, 6, -1, -1, 0, 6, -4, -4, 5,
    -- filter=81 channel=36
    1, 2, 6, 4, 0, 7, 3, 9, 4,
    -- filter=81 channel=37
    5, -3, -7, -3, -1, 0, 4, 0, 13,
    -- filter=81 channel=38
    -6, 0, -6, -2, -12, -6, 5, -8, -7,
    -- filter=81 channel=39
    -1, 1, -2, 9, 7, 0, 5, 8, 2,
    -- filter=81 channel=40
    -8, 3, 7, -1, 4, 0, -2, 7, -7,
    -- filter=81 channel=41
    4, -5, 0, 19, 3, 10, 20, 10, 18,
    -- filter=81 channel=42
    5, 0, 4, -7, 0, 2, -6, 4, 3,
    -- filter=81 channel=43
    -4, 11, 12, 0, 2, 0, 3, 5, 4,
    -- filter=81 channel=44
    -10, -3, -9, -9, -13, 0, 5, -5, 0,
    -- filter=81 channel=45
    2, 0, 7, 2, 8, 8, 0, 4, 3,
    -- filter=81 channel=46
    -2, 2, 3, -4, 8, 3, 9, 6, 0,
    -- filter=81 channel=47
    -9, -14, -1, -11, -8, -7, -5, -4, -12,
    -- filter=81 channel=48
    -12, -11, -6, -4, -15, -20, 9, -4, -4,
    -- filter=81 channel=49
    -3, -5, -3, 7, 6, -6, -1, 6, -4,
    -- filter=81 channel=50
    -6, -4, -1, -13, -19, -16, -5, -12, -7,
    -- filter=81 channel=51
    6, -3, 2, 2, 0, 2, 6, -5, -6,
    -- filter=81 channel=52
    0, -4, 4, 4, 5, 0, 4, -2, 1,
    -- filter=81 channel=53
    0, 4, -5, 4, 5, 0, 1, -4, 2,
    -- filter=81 channel=54
    7, 4, -3, 0, 0, -4, 4, -4, -6,
    -- filter=81 channel=55
    -5, 4, 0, 10, 8, -10, 3, 2, -9,
    -- filter=81 channel=56
    0, 0, -4, -2, -4, -1, -4, -2, 2,
    -- filter=81 channel=57
    0, -6, 2, 5, 6, -4, 4, -2, 1,
    -- filter=81 channel=58
    7, 11, -3, 1, 7, 9, -1, 5, 12,
    -- filter=81 channel=59
    -13, -7, -7, 0, -18, -18, 7, -2, -11,
    -- filter=81 channel=60
    -1, -4, 2, -1, 4, 2, -6, 5, 4,
    -- filter=81 channel=61
    -4, -2, 1, 5, -2, 9, 0, 1, 10,
    -- filter=81 channel=62
    -1, 2, 5, -6, -5, 0, 1, -2, 1,
    -- filter=81 channel=63
    2, -4, 3, 6, 5, 7, 0, 11, 14,
    -- filter=81 channel=64
    5, -3, 2, 2, 4, 0, 2, 0, 3,
    -- filter=81 channel=65
    5, -1, -4, -2, -6, -1, -2, 1, -3,
    -- filter=81 channel=66
    5, -1, 0, 3, 0, 8, 7, -2, 4,
    -- filter=81 channel=67
    -2, -3, 6, 0, 8, -3, -4, 8, 6,
    -- filter=81 channel=68
    -3, -5, 2, -4, -3, -3, 0, 5, 10,
    -- filter=81 channel=69
    -2, -3, 2, -4, 0, 2, -3, -2, 9,
    -- filter=81 channel=70
    -12, -10, -8, -9, -11, -18, 2, 0, -20,
    -- filter=81 channel=71
    0, 5, 4, 4, -7, 4, -4, 3, 4,
    -- filter=81 channel=72
    -7, -13, 0, -7, -3, -1, -4, -4, -8,
    -- filter=81 channel=73
    1, -5, -3, 2, 1, -10, 6, 3, -7,
    -- filter=81 channel=74
    -5, -4, -6, 5, -11, -2, 1, -13, 1,
    -- filter=81 channel=75
    0, 1, 10, 1, 0, 8, 4, 9, 14,
    -- filter=81 channel=76
    3, 12, 7, 14, 12, 10, 10, 10, 5,
    -- filter=81 channel=77
    6, 1, -5, 0, 3, -3, 0, 1, 3,
    -- filter=81 channel=78
    3, -7, 0, 6, 0, 6, 6, 2, 4,
    -- filter=81 channel=79
    -4, -2, -8, 7, -6, -20, 10, 3, -3,
    -- filter=81 channel=80
    -7, -6, -7, -10, -16, -16, 2, -14, -5,
    -- filter=81 channel=81
    -3, 0, -1, -6, -1, 5, 3, 7, -4,
    -- filter=81 channel=82
    -6, 1, -1, 5, -2, 6, -3, 5, 6,
    -- filter=81 channel=83
    -3, -6, -1, -8, 0, -5, -5, 2, 4,
    -- filter=81 channel=84
    -1, 0, 0, 10, 9, -6, 10, 13, 0,
    -- filter=81 channel=85
    -2, 1, -6, -3, 2, 0, -1, 7, -7,
    -- filter=81 channel=86
    11, -2, 1, 2, 8, -2, 10, 8, 1,
    -- filter=81 channel=87
    7, 0, 1, 15, 11, 13, 3, 7, 11,
    -- filter=81 channel=88
    4, 10, 8, 7, -1, 1, 2, 0, 2,
    -- filter=81 channel=89
    -6, -3, -6, -6, -4, -13, -3, -4, -12,
    -- filter=81 channel=90
    1, -5, 4, 4, -1, 4, 9, -5, 2,
    -- filter=81 channel=91
    -12, -12, -7, 1, -7, -21, 8, -7, -14,
    -- filter=81 channel=92
    -4, 7, 2, -2, 2, 2, 1, -1, -2,
    -- filter=81 channel=93
    -9, -12, -4, -10, -6, -9, 6, 1, 6,
    -- filter=81 channel=94
    6, -1, -7, 0, -3, 4, 4, -2, -3,
    -- filter=81 channel=95
    -7, -1, 6, -2, -4, -6, -3, 1, -4,
    -- filter=81 channel=96
    -2, 2, -5, -5, -1, 4, 5, 1, 3,
    -- filter=81 channel=97
    0, 6, 3, -5, -2, 2, 0, -2, -3,
    -- filter=81 channel=98
    -5, 0, -7, -13, -11, -21, -6, -13, -7,
    -- filter=81 channel=99
    -2, -6, 1, -8, -14, -6, 7, 0, -13,
    -- filter=81 channel=100
    3, -5, -8, 9, -5, 6, 5, 1, 1,
    -- filter=81 channel=101
    6, 2, -6, 1, 0, -5, 7, 9, 0,
    -- filter=81 channel=102
    -5, 3, 3, -4, -3, -5, -2, -6, 0,
    -- filter=81 channel=103
    -9, -3, -5, -11, -15, 1, -3, -12, -7,
    -- filter=81 channel=104
    -9, -10, 1, -9, -6, -11, 4, -8, -8,
    -- filter=81 channel=105
    0, 4, 3, 3, 4, 6, 2, 9, 7,
    -- filter=81 channel=106
    8, 10, 4, 8, 2, 5, -2, 5, 8,
    -- filter=81 channel=107
    1, 9, 4, 7, 9, 11, 4, 8, 5,
    -- filter=81 channel=108
    7, 1, 9, 13, 13, 7, 0, 1, 3,
    -- filter=81 channel=109
    -9, -11, -11, -2, -9, -24, 5, 1, -7,
    -- filter=81 channel=110
    6, -7, 8, 4, -7, 7, -3, -3, -3,
    -- filter=81 channel=111
    5, -3, 4, 8, 7, 3, 6, -3, 5,
    -- filter=81 channel=112
    -7, -2, -11, -12, -12, -7, 1, 1, -13,
    -- filter=81 channel=113
    -3, -10, 2, 0, -9, -4, 0, -7, -6,
    -- filter=81 channel=114
    -3, 0, -4, 7, 17, 5, 3, 16, 14,
    -- filter=81 channel=115
    1, 7, -3, -1, -4, 6, 6, 3, 0,
    -- filter=81 channel=116
    0, -8, -5, 1, -2, -19, 5, 5, -6,
    -- filter=81 channel=117
    5, -7, 4, 3, -6, -1, 6, 2, -8,
    -- filter=81 channel=118
    -4, -1, -5, 0, 0, -1, 3, 7, 3,
    -- filter=81 channel=119
    6, -2, -7, 4, -3, -7, -2, 4, -3,
    -- filter=81 channel=120
    -12, -8, -16, -11, -12, -13, 2, -9, -14,
    -- filter=81 channel=121
    3, -1, -3, -5, 0, -7, 0, -7, -5,
    -- filter=81 channel=122
    -3, -18, -10, -4, -10, -1, 4, -9, -11,
    -- filter=81 channel=123
    -5, -5, -3, 6, 3, 2, -6, -4, -1,
    -- filter=81 channel=124
    -5, 6, 0, 4, 0, -2, -3, -4, 7,
    -- filter=81 channel=125
    -3, -4, -7, -3, -15, -8, 6, 2, -7,
    -- filter=81 channel=126
    1, 3, 1, 2, -1, 0, 0, -3, -2,
    -- filter=81 channel=127
    -2, -3, -6, 7, -6, 4, 2, -3, 8,
    -- filter=82 channel=0
    -3, 5, 5, 0, -4, -9, -8, -5, -6,
    -- filter=82 channel=1
    6, 9, 0, -5, -7, -1, -5, -3, -12,
    -- filter=82 channel=2
    -9, -7, -9, 0, 3, 3, -2, -4, -3,
    -- filter=82 channel=3
    2, -1, 4, -11, 1, -3, -6, -9, -6,
    -- filter=82 channel=4
    -9, -10, -3, -8, -14, -9, -7, 0, -10,
    -- filter=82 channel=5
    2, -5, -1, -7, -8, 3, -2, -15, -1,
    -- filter=82 channel=6
    -12, 2, -7, -1, 7, -4, -4, 3, -2,
    -- filter=82 channel=7
    -6, -3, -4, 6, 0, 7, -4, -7, 4,
    -- filter=82 channel=8
    -4, 3, -1, 9, -4, 0, 5, 4, -1,
    -- filter=82 channel=9
    5, 0, -5, -4, -7, 5, -7, 1, 1,
    -- filter=82 channel=10
    0, 3, 9, 1, 7, -1, 11, 6, 2,
    -- filter=82 channel=11
    -9, -4, -6, 0, 3, -4, 3, 7, 11,
    -- filter=82 channel=12
    1, 3, 5, 10, 4, 2, 12, 3, 2,
    -- filter=82 channel=13
    0, 5, -6, -7, 15, -1, 14, 15, -5,
    -- filter=82 channel=14
    1, 5, 6, 0, 0, 0, 0, -1, -4,
    -- filter=82 channel=15
    -6, -5, 4, -12, -2, 3, -7, 9, 11,
    -- filter=82 channel=16
    3, 9, -2, -4, -6, -3, -6, -12, -11,
    -- filter=82 channel=17
    -4, 7, 4, 1, 4, 0, 5, 6, 0,
    -- filter=82 channel=18
    -10, -8, 3, -8, 11, 1, -4, 2, 6,
    -- filter=82 channel=19
    -2, -7, 3, 0, -4, 0, -3, -4, 4,
    -- filter=82 channel=20
    -13, -19, -11, -15, -3, 1, 0, 19, 8,
    -- filter=82 channel=21
    4, 3, 11, 2, -4, -1, -9, -5, -12,
    -- filter=82 channel=22
    1, 0, 7, -5, -4, 6, 0, 2, 6,
    -- filter=82 channel=23
    -2, -6, 3, -3, 9, 9, 7, 12, 18,
    -- filter=82 channel=24
    -1, 6, 5, 0, 4, 6, 6, 6, 0,
    -- filter=82 channel=25
    -7, 10, -4, 7, 0, 3, 9, 1, -1,
    -- filter=82 channel=26
    0, 6, 2, -4, -9, -3, -6, -6, 3,
    -- filter=82 channel=27
    -4, 12, 1, 4, 0, 8, 0, -11, -2,
    -- filter=82 channel=28
    0, 1, 4, -3, -5, -1, 6, 3, -1,
    -- filter=82 channel=29
    -11, -19, -8, -14, 5, -6, -9, 6, 9,
    -- filter=82 channel=30
    1, -6, -3, 0, -10, 4, 0, -14, -6,
    -- filter=82 channel=31
    4, 5, 4, 4, -2, 4, 0, -14, 1,
    -- filter=82 channel=32
    -11, 1, 6, -2, 9, 5, 5, 8, 1,
    -- filter=82 channel=33
    -6, 12, 5, 2, 3, 5, 4, -3, -3,
    -- filter=82 channel=34
    4, 2, 2, -2, 3, 7, 3, 0, 12,
    -- filter=82 channel=35
    4, 0, 3, 4, -6, -2, -4, -4, 7,
    -- filter=82 channel=36
    5, -7, -5, 5, 9, -1, -1, -6, 5,
    -- filter=82 channel=37
    6, 4, 5, -2, -3, -10, -10, -11, -12,
    -- filter=82 channel=38
    4, 2, 3, -4, 3, 6, 1, -9, -2,
    -- filter=82 channel=39
    -4, -1, -7, -10, -2, 5, 2, 7, 3,
    -- filter=82 channel=40
    -3, -7, -2, -1, 7, -4, 4, 9, -1,
    -- filter=82 channel=41
    4, 3, 5, 2, 24, -4, 9, 14, -9,
    -- filter=82 channel=42
    0, -5, 2, -3, -7, -8, 3, 0, -2,
    -- filter=82 channel=43
    2, 5, -4, -11, 7, -1, -6, 8, 5,
    -- filter=82 channel=44
    -1, 13, 2, -4, -9, -7, -8, -12, -9,
    -- filter=82 channel=45
    -2, -10, -9, 2, -5, 3, 0, -5, 7,
    -- filter=82 channel=46
    8, -4, 3, 0, -1, 3, -1, -3, 3,
    -- filter=82 channel=47
    13, 2, 4, -5, -9, 3, -8, -16, -2,
    -- filter=82 channel=48
    8, 0, 9, 1, -10, 3, -9, -12, -4,
    -- filter=82 channel=49
    -8, -2, -10, 0, -8, 1, -9, -7, 3,
    -- filter=82 channel=50
    4, 6, 8, -7, 0, -1, -4, -5, 0,
    -- filter=82 channel=51
    2, -2, 0, -5, 4, 2, -5, -3, 1,
    -- filter=82 channel=52
    -4, 2, -4, 0, 7, 8, 4, -1, 8,
    -- filter=82 channel=53
    -12, -11, -6, 1, -3, -3, 4, 2, 6,
    -- filter=82 channel=54
    -3, 6, 4, -3, -1, 1, 3, 4, -3,
    -- filter=82 channel=55
    -8, 4, -6, -9, 16, -1, 3, 8, 16,
    -- filter=82 channel=56
    3, 5, 2, 9, -1, -5, 0, 5, -5,
    -- filter=82 channel=57
    0, 5, -6, -8, 3, -1, -4, -5, -1,
    -- filter=82 channel=58
    -8, -2, 0, -9, -5, -5, -1, -10, -1,
    -- filter=82 channel=59
    10, 6, 1, -1, 0, 1, 2, -5, -3,
    -- filter=82 channel=60
    3, -3, 4, 3, 4, 0, 2, -1, -3,
    -- filter=82 channel=61
    -5, -2, -7, -2, 7, -4, 8, 5, 7,
    -- filter=82 channel=62
    -4, -6, -5, 2, 0, 0, 0, 1, 4,
    -- filter=82 channel=63
    -3, -7, -5, -1, -3, 2, -8, -7, -6,
    -- filter=82 channel=64
    -1, 2, 1, 3, 8, -2, 0, 4, 1,
    -- filter=82 channel=65
    3, -3, -1, -4, 1, 0, -2, 6, 3,
    -- filter=82 channel=66
    0, 11, -6, 9, 14, -4, 6, 1, -8,
    -- filter=82 channel=67
    5, -5, -2, -3, 5, -6, 1, -5, 3,
    -- filter=82 channel=68
    -2, -1, -8, 4, -3, -8, -2, -6, -9,
    -- filter=82 channel=69
    0, 3, 0, 0, 7, -5, 6, 6, 5,
    -- filter=82 channel=70
    -4, 10, -1, 0, -2, 0, 0, 0, 0,
    -- filter=82 channel=71
    -2, 4, 0, -4, -5, 0, -4, -3, -6,
    -- filter=82 channel=72
    9, -2, 2, 0, -1, 0, -1, 3, -2,
    -- filter=82 channel=73
    -11, -4, 0, 5, 0, -2, 0, -7, 2,
    -- filter=82 channel=74
    -1, 5, -5, 6, 2, 11, -1, 5, -2,
    -- filter=82 channel=75
    0, 3, 10, -4, 2, -6, -6, -9, -10,
    -- filter=82 channel=76
    -7, -12, -10, -3, 12, -9, -3, 20, 0,
    -- filter=82 channel=77
    -6, 0, -4, 1, 7, 2, 1, 5, 2,
    -- filter=82 channel=78
    4, 4, 5, 4, -7, 6, -7, 1, 4,
    -- filter=82 channel=79
    -4, 4, 2, -7, 6, 0, 4, 13, 0,
    -- filter=82 channel=80
    12, 0, 6, 0, -5, 4, -3, -13, -3,
    -- filter=82 channel=81
    4, 2, -1, -7, 7, -4, -3, -5, 4,
    -- filter=82 channel=82
    6, 2, 5, 5, 4, 6, 3, -4, 6,
    -- filter=82 channel=83
    2, -6, -1, -5, 1, -3, -3, 0, -5,
    -- filter=82 channel=84
    -2, 4, -9, -9, 0, 0, -6, 5, 1,
    -- filter=82 channel=85
    -1, -2, 0, 6, -4, -1, 1, 2, -4,
    -- filter=82 channel=86
    5, 10, 6, -5, 7, 1, -2, 8, 4,
    -- filter=82 channel=87
    -8, 6, -6, -3, 0, 0, -1, 10, 4,
    -- filter=82 channel=88
    3, 0, 0, 3, 8, -5, 7, 7, 7,
    -- filter=82 channel=89
    3, -2, 0, 1, 16, -8, 14, 7, 1,
    -- filter=82 channel=90
    7, 8, -6, 0, -3, -7, 7, -3, 6,
    -- filter=82 channel=91
    -13, 0, -3, -7, -1, 0, 3, -5, 7,
    -- filter=82 channel=92
    0, 1, 2, 5, -7, -1, -2, -5, 3,
    -- filter=82 channel=93
    2, 10, 2, 4, -7, -3, -4, -19, -2,
    -- filter=82 channel=94
    1, -4, -5, -1, 1, -1, 0, 2, 4,
    -- filter=82 channel=95
    6, -3, 5, -6, 5, 2, 8, 7, 0,
    -- filter=82 channel=96
    1, 0, 4, -1, 5, -7, 3, -1, 1,
    -- filter=82 channel=97
    -1, -5, -1, 0, 3, -5, -9, 2, 4,
    -- filter=82 channel=98
    -6, 6, 0, -2, 0, -2, 4, 2, -1,
    -- filter=82 channel=99
    -7, 7, -7, 14, 13, -2, 7, -2, 12,
    -- filter=82 channel=100
    5, 0, 0, -5, 9, 1, 5, -3, -6,
    -- filter=82 channel=101
    0, -4, -10, -2, 0, 0, -5, -2, -1,
    -- filter=82 channel=102
    -6, -6, -3, 7, -2, -4, 5, 3, -4,
    -- filter=82 channel=103
    12, 0, 3, -5, -16, -1, -8, -14, -1,
    -- filter=82 channel=104
    0, 0, 6, 3, 3, 9, 3, -11, 5,
    -- filter=82 channel=105
    -6, -4, -8, -6, 8, -2, 2, 13, 8,
    -- filter=82 channel=106
    -8, -9, -10, -7, -3, 1, -1, -2, 3,
    -- filter=82 channel=107
    -10, -4, -12, -3, 2, 0, 0, 1, 12,
    -- filter=82 channel=108
    -8, -5, 4, -6, 0, 3, 5, 9, 3,
    -- filter=82 channel=109
    -10, 1, 5, 2, 6, 0, 2, -5, 9,
    -- filter=82 channel=110
    -1, 1, 9, 9, 0, -5, 4, 1, 0,
    -- filter=82 channel=111
    1, 6, -1, -1, 0, 0, -5, 3, 1,
    -- filter=82 channel=112
    -6, 10, 5, -2, -9, 0, 1, -4, -2,
    -- filter=82 channel=113
    9, 10, 8, -2, 5, 0, -4, 1, -1,
    -- filter=82 channel=114
    -15, -1, -3, -10, 2, -8, -8, -6, -8,
    -- filter=82 channel=115
    3, -3, 6, -3, -5, 3, 3, 3, -3,
    -- filter=82 channel=116
    -6, 0, -5, 0, 6, 5, 2, 4, 5,
    -- filter=82 channel=117
    6, -6, 0, -3, 0, -6, 7, 7, -8,
    -- filter=82 channel=118
    -2, 2, 3, 0, -4, -3, 2, -3, 2,
    -- filter=82 channel=119
    6, 5, 6, 11, 4, 0, 0, 4, -2,
    -- filter=82 channel=120
    -14, 7, -5, 0, 7, 4, -1, 0, 12,
    -- filter=82 channel=121
    11, 3, -4, 3, 12, -5, 5, 0, 2,
    -- filter=82 channel=122
    17, 15, 4, 8, -5, -3, -5, -23, -6,
    -- filter=82 channel=123
    -6, 0, -3, -6, -4, 5, -5, 6, 2,
    -- filter=82 channel=124
    -7, -1, -9, -6, 5, 4, 5, 5, 0,
    -- filter=82 channel=125
    -3, 7, -5, 5, -1, 8, 0, -9, -2,
    -- filter=82 channel=126
    5, 1, 7, 3, 3, 1, 4, 3, 1,
    -- filter=82 channel=127
    1, 0, 4, -6, 1, 5, -5, 0, 2,
    -- filter=83 channel=0
    -19, -11, -19, -22, -28, -15, -11, -12, -5,
    -- filter=83 channel=1
    -21, -26, -10, -12, -17, -9, -10, -9, -9,
    -- filter=83 channel=2
    2, 9, 0, -4, -3, 5, 6, -2, 2,
    -- filter=83 channel=3
    -5, -9, 0, -13, -14, -15, -6, -5, -6,
    -- filter=83 channel=4
    0, 0, -7, 1, 3, 8, 6, 4, 1,
    -- filter=83 channel=5
    -16, -13, -5, -13, -18, -5, -14, 0, -4,
    -- filter=83 channel=6
    4, 8, 0, -7, -8, -6, 4, -7, -3,
    -- filter=83 channel=7
    0, -3, 2, -3, 4, -5, -1, 1, -6,
    -- filter=83 channel=8
    5, 7, -5, 7, -4, 3, 0, -1, -2,
    -- filter=83 channel=9
    1, 6, 0, 2, -3, -1, -2, 8, 0,
    -- filter=83 channel=10
    4, -4, -7, 8, 2, -4, 5, -2, 9,
    -- filter=83 channel=11
    3, 12, 3, 9, 11, 0, -5, -1, -5,
    -- filter=83 channel=12
    5, 1, 3, -2, 0, 4, 1, -2, -7,
    -- filter=83 channel=13
    1, -7, 2, -4, -4, 0, 12, -6, -1,
    -- filter=83 channel=14
    -2, 5, 5, 0, -2, -6, -3, 6, 4,
    -- filter=83 channel=15
    -11, -3, -9, -6, -7, -9, -3, -4, -5,
    -- filter=83 channel=16
    0, 0, -4, -13, -13, -8, -6, -2, -4,
    -- filter=83 channel=17
    -4, -1, 5, 5, -3, -2, -4, 1, -6,
    -- filter=83 channel=18
    -17, -12, -7, -1, -5, -9, 8, -3, 4,
    -- filter=83 channel=19
    -2, 5, -2, 3, 0, -2, 7, 0, -1,
    -- filter=83 channel=20
    -3, 7, 15, 2, 6, 2, -13, 0, -11,
    -- filter=83 channel=21
    -6, -3, 7, -3, -6, 9, 1, 5, 2,
    -- filter=83 channel=22
    -2, -6, -12, 0, -6, -4, -8, 3, 4,
    -- filter=83 channel=23
    -12, 0, -13, -2, 4, 4, -2, 6, -6,
    -- filter=83 channel=24
    -3, 0, -6, -4, -1, 2, 4, -5, -6,
    -- filter=83 channel=25
    -9, -13, -1, 2, -1, 3, 1, 13, 15,
    -- filter=83 channel=26
    3, -9, 0, -2, 0, 5, -8, -2, -5,
    -- filter=83 channel=27
    -17, -14, -14, -8, -7, 5, 11, 12, 17,
    -- filter=83 channel=28
    -7, 4, 1, 1, 6, 0, -5, -4, 3,
    -- filter=83 channel=29
    3, 15, 10, -2, 12, 2, -8, -3, 1,
    -- filter=83 channel=30
    -1, 0, 0, -2, -9, 2, -3, -2, 5,
    -- filter=83 channel=31
    2, 2, 1, 10, 0, 3, 2, 0, 9,
    -- filter=83 channel=32
    -13, -5, -14, -3, 4, -1, 0, -2, -5,
    -- filter=83 channel=33
    -14, -11, -7, -2, -5, -1, 4, -5, 9,
    -- filter=83 channel=34
    -1, 2, 6, -7, -3, 0, -9, -6, 6,
    -- filter=83 channel=35
    6, -2, -2, -6, 6, 0, -7, 0, 0,
    -- filter=83 channel=36
    5, 14, 15, 3, 11, 4, -6, 3, -6,
    -- filter=83 channel=37
    -23, -19, -8, -16, -17, -16, -7, -11, 1,
    -- filter=83 channel=38
    -8, 0, 5, -1, -5, -4, 8, 3, 0,
    -- filter=83 channel=39
    -1, -1, 10, 7, 10, 8, 0, -2, 0,
    -- filter=83 channel=40
    -3, 7, 2, -2, 0, -6, -3, -2, -11,
    -- filter=83 channel=41
    -6, 13, 0, 7, 12, -8, 3, 1, 6,
    -- filter=83 channel=42
    -2, -7, -3, 1, -10, 0, 4, 6, 3,
    -- filter=83 channel=43
    -8, -1, -10, -10, -9, -7, -11, -2, -3,
    -- filter=83 channel=44
    -3, -19, -3, -4, -15, 3, -1, -1, 1,
    -- filter=83 channel=45
    3, -3, 1, 3, 0, -2, -3, -8, 5,
    -- filter=83 channel=46
    2, 0, 0, 0, 1, -10, -6, -7, -4,
    -- filter=83 channel=47
    -8, -6, 0, -11, -20, 0, -9, -8, 0,
    -- filter=83 channel=48
    0, 0, -3, 0, -4, 10, 7, 8, 16,
    -- filter=83 channel=49
    -8, -1, -2, 8, 6, 2, 4, 5, 6,
    -- filter=83 channel=50
    -6, -7, -3, -3, 7, 0, 11, -1, 4,
    -- filter=83 channel=51
    0, 7, -4, 1, 3, 0, 1, 5, 0,
    -- filter=83 channel=52
    -6, 1, 0, 2, -2, 0, 2, -2, 0,
    -- filter=83 channel=53
    -2, 2, 7, 5, 0, 9, 2, 2, 3,
    -- filter=83 channel=54
    7, 3, -6, 0, -5, -5, -6, 1, 3,
    -- filter=83 channel=55
    1, 0, 2, 7, 5, -4, 1, 8, 2,
    -- filter=83 channel=56
    0, 2, -5, 7, 5, 5, 3, 2, -5,
    -- filter=83 channel=57
    2, 0, 1, 0, 0, 0, 4, -6, -6,
    -- filter=83 channel=58
    -11, -7, -9, -8, -12, -3, 0, -8, -8,
    -- filter=83 channel=59
    -3, -8, 1, 7, 5, 5, 11, 5, 8,
    -- filter=83 channel=60
    -1, 1, -4, 4, -5, 5, -6, -3, -2,
    -- filter=83 channel=61
    9, 10, 0, 5, 5, 0, -5, 1, 0,
    -- filter=83 channel=62
    -2, 0, -4, -7, 6, -4, -5, -7, -1,
    -- filter=83 channel=63
    -6, 1, 5, -4, 2, -1, -10, 2, -4,
    -- filter=83 channel=64
    -3, 0, -3, 0, 2, 7, 4, 0, 2,
    -- filter=83 channel=65
    6, -1, 1, -3, 0, 4, 0, 3, 2,
    -- filter=83 channel=66
    -2, 7, 8, 2, 9, -3, 1, 0, 0,
    -- filter=83 channel=67
    1, -6, -6, -5, 5, 3, -3, 0, -6,
    -- filter=83 channel=68
    3, 3, 5, 7, -2, 1, 2, -1, -4,
    -- filter=83 channel=69
    7, 7, 6, 0, 4, 1, 1, -1, 4,
    -- filter=83 channel=70
    -9, -16, -12, 1, -2, -3, 9, 1, -4,
    -- filter=83 channel=71
    1, -4, 3, -9, -2, 2, -10, -2, 2,
    -- filter=83 channel=72
    -1, 6, -2, 8, 2, 2, 15, 2, 6,
    -- filter=83 channel=73
    -3, 3, -5, 11, -1, 9, 1, 11, 5,
    -- filter=83 channel=74
    -1, 2, -9, 5, 8, 2, -5, 8, 0,
    -- filter=83 channel=75
    -21, -18, -18, -25, -25, -19, -11, -1, 2,
    -- filter=83 channel=76
    4, 10, 10, -2, 1, 2, -5, -3, -10,
    -- filter=83 channel=77
    -6, 5, -4, -4, 0, 0, 0, 6, -6,
    -- filter=83 channel=78
    -5, 0, -4, 0, 2, 0, -5, -3, 7,
    -- filter=83 channel=79
    -15, -9, -9, -10, -14, -13, 8, 2, -4,
    -- filter=83 channel=80
    0, -5, 0, 5, 8, 6, 11, 10, 12,
    -- filter=83 channel=81
    3, -7, -3, 3, -6, 6, 6, -1, -7,
    -- filter=83 channel=82
    3, -4, -3, 0, 1, 2, -8, 0, -8,
    -- filter=83 channel=83
    -5, 3, -3, -3, 9, 10, 3, 4, 3,
    -- filter=83 channel=84
    -9, 0, -4, 8, 7, -2, 0, 3, 0,
    -- filter=83 channel=85
    -6, 5, 5, -1, 3, -1, -2, 7, 2,
    -- filter=83 channel=86
    0, -10, -4, -8, -1, -3, 0, -4, -2,
    -- filter=83 channel=87
    -2, 0, 3, 2, 9, -2, -5, -3, 0,
    -- filter=83 channel=88
    1, 9, 5, 8, 3, 3, -6, 1, 0,
    -- filter=83 channel=89
    -7, -11, 2, 10, -2, 3, 10, 8, 8,
    -- filter=83 channel=90
    0, 7, -3, 2, 11, 7, 0, 1, -3,
    -- filter=83 channel=91
    0, 4, 2, 8, 4, 5, 4, 9, 0,
    -- filter=83 channel=92
    -3, -7, -2, -7, 1, -6, 1, 0, 6,
    -- filter=83 channel=93
    -9, -21, -17, -10, -21, -10, 0, 0, -6,
    -- filter=83 channel=94
    -4, -4, -3, -4, -1, 0, 4, 4, -4,
    -- filter=83 channel=95
    -1, -2, -6, 1, 0, -5, -7, 2, 3,
    -- filter=83 channel=96
    -5, 2, -7, 7, -6, 0, -5, 6, -2,
    -- filter=83 channel=97
    -6, -9, -7, -6, -4, -9, 2, -2, -7,
    -- filter=83 channel=98
    -11, -11, 1, 8, 0, -2, 14, 9, 12,
    -- filter=83 channel=99
    11, 4, 6, 16, 20, 12, 7, 12, 10,
    -- filter=83 channel=100
    0, 7, 2, -3, 5, 2, 6, 9, 2,
    -- filter=83 channel=101
    0, -5, 7, 6, -5, 0, -3, 0, -2,
    -- filter=83 channel=102
    -3, 0, 3, 1, 6, 1, 3, 1, -1,
    -- filter=83 channel=103
    -9, -11, 1, -19, -9, -11, -14, -2, 2,
    -- filter=83 channel=104
    6, 2, 1, 0, 13, 4, 6, 11, 13,
    -- filter=83 channel=105
    -4, 0, 4, -7, 6, -8, 1, -13, -1,
    -- filter=83 channel=106
    -6, 4, 3, 9, 9, 5, 3, -6, 1,
    -- filter=83 channel=107
    -15, 2, -9, -8, -4, -2, -14, -1, -9,
    -- filter=83 channel=108
    3, -6, 2, -6, -7, -3, 2, -3, -4,
    -- filter=83 channel=109
    -8, -3, -10, 4, 12, 3, 17, 15, 16,
    -- filter=83 channel=110
    0, 1, -6, 2, -2, 3, 7, 6, 5,
    -- filter=83 channel=111
    -5, -6, -5, -5, -4, -5, -5, 0, -5,
    -- filter=83 channel=112
    -1, -2, -5, 0, 1, 6, 2, -2, 9,
    -- filter=83 channel=113
    1, -1, -10, -1, -1, -9, 6, -2, 0,
    -- filter=83 channel=114
    -11, -12, -15, -16, -11, -6, 0, -2, -4,
    -- filter=83 channel=115
    4, -3, -4, 1, 1, 7, 7, -6, 7,
    -- filter=83 channel=116
    1, 1, 5, 15, 11, 6, 15, 3, 15,
    -- filter=83 channel=117
    1, 2, -2, 0, -3, -4, -2, 3, 0,
    -- filter=83 channel=118
    1, 3, -2, 6, -3, -4, 0, 5, -1,
    -- filter=83 channel=119
    0, -4, 5, 4, 5, 4, 3, 7, -3,
    -- filter=83 channel=120
    -4, -1, -6, 0, 11, 10, 8, 8, 12,
    -- filter=83 channel=121
    -5, -6, 1, 3, 3, 4, 9, -7, -3,
    -- filter=83 channel=122
    -13, -14, 2, -18, -16, -8, -19, -15, 7,
    -- filter=83 channel=123
    6, -6, -1, -7, 4, -3, -1, -2, -5,
    -- filter=83 channel=124
    -9, -2, -3, 4, -8, 4, -9, -6, -10,
    -- filter=83 channel=125
    1, -3, 2, 5, 17, 16, 7, 10, 17,
    -- filter=83 channel=126
    1, 0, 3, -3, -1, 2, 2, 0, -3,
    -- filter=83 channel=127
    -3, 4, -5, -3, 1, 0, 7, -5, 2,
    -- filter=84 channel=0
    2, 0, 5, 6, 6, 2, 4, -4, -2,
    -- filter=84 channel=1
    -6, -2, 0, 7, -5, 2, 0, -6, 4,
    -- filter=84 channel=2
    -1, 2, 0, -1, 3, 7, -6, -3, 6,
    -- filter=84 channel=3
    -7, 2, -3, -7, -4, 6, -2, 1, 4,
    -- filter=84 channel=4
    6, 2, 0, 0, 3, -5, 4, 0, -7,
    -- filter=84 channel=5
    1, -3, 2, 3, -7, -4, 0, -4, -1,
    -- filter=84 channel=6
    -5, 0, 4, -3, -7, 7, -1, 0, -6,
    -- filter=84 channel=7
    6, 3, -7, -1, 0, -6, 6, 3, 4,
    -- filter=84 channel=8
    -5, 0, 7, 0, 5, -2, 5, 5, 1,
    -- filter=84 channel=9
    0, -2, -1, 0, -2, -1, -1, -2, 5,
    -- filter=84 channel=10
    -6, 1, 0, -1, -1, 2, 6, -2, 5,
    -- filter=84 channel=11
    -5, 4, 4, 1, 2, 6, 0, 2, 6,
    -- filter=84 channel=12
    6, 0, -4, 0, -1, 0, -1, 0, 3,
    -- filter=84 channel=13
    5, -3, 0, 3, -4, 1, -6, -2, 0,
    -- filter=84 channel=14
    2, 7, 4, 6, 1, 3, 6, 0, 5,
    -- filter=84 channel=15
    -7, 2, -7, 0, -5, -2, -1, -1, 3,
    -- filter=84 channel=16
    2, -5, 1, 1, -4, -2, 6, -1, -3,
    -- filter=84 channel=17
    3, 5, -3, 4, 3, -1, -1, 2, 0,
    -- filter=84 channel=18
    0, 3, -2, 2, 0, -3, 0, 0, 5,
    -- filter=84 channel=19
    6, 5, 0, 0, 0, 1, -3, -6, -6,
    -- filter=84 channel=20
    0, 1, -6, 0, 0, 5, -7, -4, 0,
    -- filter=84 channel=21
    6, 4, 6, 5, 1, 2, -6, -1, -6,
    -- filter=84 channel=22
    0, 3, -5, -4, 2, -2, -2, -3, 1,
    -- filter=84 channel=23
    1, 0, -4, 2, 0, 3, -2, 5, 5,
    -- filter=84 channel=24
    -2, 4, 0, -3, 4, 4, -4, -2, -4,
    -- filter=84 channel=25
    -6, -5, 0, 0, 5, 1, -6, 0, 1,
    -- filter=84 channel=26
    4, -1, -4, -6, 4, -4, 1, -6, 2,
    -- filter=84 channel=27
    -2, 1, 0, 3, 2, 4, -5, 2, 5,
    -- filter=84 channel=28
    -7, -1, -6, 2, 1, 7, -1, 5, 7,
    -- filter=84 channel=29
    1, 1, -6, -4, -1, 2, 1, -5, -4,
    -- filter=84 channel=30
    1, -7, 2, 5, -2, -2, 6, -2, -5,
    -- filter=84 channel=31
    -8, -2, -2, 4, 1, -2, 5, -4, -3,
    -- filter=84 channel=32
    3, 0, -7, -4, -1, 2, 0, 6, 4,
    -- filter=84 channel=33
    1, 0, -3, 3, -2, 2, 1, -4, 7,
    -- filter=84 channel=34
    -3, 1, 0, 2, 5, 0, 7, -5, 1,
    -- filter=84 channel=35
    -2, 0, 0, 3, 3, -5, -4, -3, -2,
    -- filter=84 channel=36
    -3, 0, -3, -1, 7, 0, -5, -1, -6,
    -- filter=84 channel=37
    2, -6, 4, -3, 0, -4, 5, 4, 0,
    -- filter=84 channel=38
    1, -1, 1, -4, -4, 5, -4, 6, -1,
    -- filter=84 channel=39
    0, 2, 3, -2, 3, 4, 6, -5, -7,
    -- filter=84 channel=40
    -5, -2, 7, -3, 0, -5, -4, -6, 3,
    -- filter=84 channel=41
    1, -5, 0, 0, -5, -5, 5, 1, 2,
    -- filter=84 channel=42
    0, -3, -1, 6, -2, -7, -7, -6, 4,
    -- filter=84 channel=43
    -5, 5, -6, 3, -2, 4, -2, 0, -1,
    -- filter=84 channel=44
    -4, -6, 6, -6, -4, 6, 2, -4, -7,
    -- filter=84 channel=45
    -7, -7, -6, 2, -4, 6, 3, 2, 6,
    -- filter=84 channel=46
    -2, 5, 7, 4, -7, 3, -6, -1, -1,
    -- filter=84 channel=47
    0, 4, -2, 3, 1, -1, 5, -6, 4,
    -- filter=84 channel=48
    4, 5, -6, -4, -4, 5, 7, -5, -5,
    -- filter=84 channel=49
    -1, 5, 3, -7, 4, 3, 3, -6, 3,
    -- filter=84 channel=50
    -7, -4, 4, 1, -5, 7, -6, -3, -3,
    -- filter=84 channel=51
    0, 5, -2, -4, 2, -1, 4, 0, 5,
    -- filter=84 channel=52
    6, 5, 5, 0, 2, 3, 5, 4, -5,
    -- filter=84 channel=53
    1, 3, -7, -4, -5, -4, 3, -5, 5,
    -- filter=84 channel=54
    -1, 1, 1, -5, 1, -7, 0, -2, 1,
    -- filter=84 channel=55
    0, -1, 2, -2, 0, 1, -3, -1, 2,
    -- filter=84 channel=56
    6, 3, -5, 4, -2, 7, 4, 0, -6,
    -- filter=84 channel=57
    7, -2, -4, -5, 0, 5, 5, -2, 7,
    -- filter=84 channel=58
    -3, -5, -6, 2, 1, -4, -7, 1, 4,
    -- filter=84 channel=59
    5, -5, 3, 6, 2, -3, 2, 0, -4,
    -- filter=84 channel=60
    2, 4, 4, 0, 2, 6, 0, -4, 6,
    -- filter=84 channel=61
    5, 0, 5, -5, 6, -4, -2, 3, 3,
    -- filter=84 channel=62
    -1, 3, -1, 6, -1, 4, -5, 0, 0,
    -- filter=84 channel=63
    -5, -7, -4, -6, -3, 0, 1, 6, -2,
    -- filter=84 channel=64
    4, -2, -1, 4, 0, -1, -7, 4, -4,
    -- filter=84 channel=65
    -2, -5, 0, 1, -1, 4, 4, 0, 5,
    -- filter=84 channel=66
    -6, 1, -2, -5, 4, -3, 6, 7, 6,
    -- filter=84 channel=67
    0, 7, 4, 2, 1, 4, -1, 0, -5,
    -- filter=84 channel=68
    1, 1, -1, -7, -3, 7, -6, -1, 0,
    -- filter=84 channel=69
    0, 3, 5, -5, 7, -1, -3, 6, 0,
    -- filter=84 channel=70
    3, -4, -6, 3, 0, 2, -7, 4, -4,
    -- filter=84 channel=71
    0, 0, -7, -7, -2, 4, -6, 6, -2,
    -- filter=84 channel=72
    1, -7, 5, 3, 7, 6, -4, 1, 1,
    -- filter=84 channel=73
    3, -6, 0, 4, 5, -5, -1, 7, -2,
    -- filter=84 channel=74
    3, 5, -7, 2, 3, 1, -1, -1, -4,
    -- filter=84 channel=75
    4, 6, -3, 3, -3, -2, 6, -6, 5,
    -- filter=84 channel=76
    -5, -6, -7, -6, 1, -3, 3, 0, 2,
    -- filter=84 channel=77
    -5, -2, 6, -1, 0, -2, -1, 0, 6,
    -- filter=84 channel=78
    -5, 3, -2, -7, 3, 4, -3, 2, -4,
    -- filter=84 channel=79
    -2, -2, -6, -4, 6, 2, -4, -1, -1,
    -- filter=84 channel=80
    -4, -6, -5, -8, 3, 0, 1, -6, 2,
    -- filter=84 channel=81
    -1, -2, 6, 0, -1, -7, -2, -3, -2,
    -- filter=84 channel=82
    2, 4, 6, -5, 3, -3, -7, -7, 6,
    -- filter=84 channel=83
    -5, 0, -6, 0, -1, -3, -2, 1, 5,
    -- filter=84 channel=84
    -1, 4, 4, -4, -4, 4, 0, -1, 1,
    -- filter=84 channel=85
    5, -4, 5, 0, -7, 0, -6, -6, -3,
    -- filter=84 channel=86
    -7, 5, 0, 5, 4, 1, -4, 0, 2,
    -- filter=84 channel=87
    1, 4, -2, -4, -3, -6, 1, -1, 4,
    -- filter=84 channel=88
    2, 5, 1, 1, 4, -6, 0, -6, -3,
    -- filter=84 channel=89
    -4, 2, 1, -5, -2, 2, 1, 3, 5,
    -- filter=84 channel=90
    -4, -4, -4, 5, -5, 4, 0, 0, 1,
    -- filter=84 channel=91
    -6, -6, 0, -7, 4, 0, -2, 0, -6,
    -- filter=84 channel=92
    0, 6, -6, 6, 0, -5, 2, 4, 3,
    -- filter=84 channel=93
    0, 2, -3, 4, 2, 2, -1, -4, -5,
    -- filter=84 channel=94
    -5, -2, 5, 0, 6, 5, 0, -4, 2,
    -- filter=84 channel=95
    -7, -5, 2, 4, -4, -5, 6, 3, 1,
    -- filter=84 channel=96
    2, -3, 5, -6, 5, -3, 6, -5, 6,
    -- filter=84 channel=97
    5, 3, -7, 2, 5, -1, -3, -3, 3,
    -- filter=84 channel=98
    2, -5, 1, -2, 6, -6, 3, -6, -5,
    -- filter=84 channel=99
    0, -3, 4, -3, -5, -4, -6, 5, -2,
    -- filter=84 channel=100
    -2, 0, 2, -2, 6, 0, 7, 1, -1,
    -- filter=84 channel=101
    0, 1, 7, 1, 0, 1, -2, -7, 6,
    -- filter=84 channel=102
    5, 7, -5, -6, -3, -2, -5, 0, -4,
    -- filter=84 channel=103
    4, 5, -1, 3, -6, -2, -5, -2, -5,
    -- filter=84 channel=104
    -6, 2, -1, 0, 5, 6, 4, 0, -3,
    -- filter=84 channel=105
    -5, -3, -6, -7, -5, 5, 1, -4, -1,
    -- filter=84 channel=106
    6, 6, -7, -6, 1, 1, -6, -5, -1,
    -- filter=84 channel=107
    5, 0, -1, -6, -6, -5, 1, -1, 5,
    -- filter=84 channel=108
    -2, -3, 1, -5, 2, 4, -3, -3, 5,
    -- filter=84 channel=109
    1, 5, 4, 5, -1, 0, -6, -4, 4,
    -- filter=84 channel=110
    3, 5, 1, -5, -7, -4, 6, 0, 6,
    -- filter=84 channel=111
    2, 3, -3, 4, 7, -2, -1, -7, -1,
    -- filter=84 channel=112
    1, -7, 0, -6, -2, 1, 5, 0, -7,
    -- filter=84 channel=113
    3, 0, -2, 4, -2, 1, -2, 7, 4,
    -- filter=84 channel=114
    -1, -1, 4, -7, 1, -4, -4, 4, -3,
    -- filter=84 channel=115
    -3, -4, 2, 0, 0, -7, 6, 3, -2,
    -- filter=84 channel=116
    -1, -6, -1, -1, 1, -5, 1, 6, -2,
    -- filter=84 channel=117
    2, 0, 5, 5, -6, -3, 7, 0, 0,
    -- filter=84 channel=118
    2, -6, -3, 1, -3, 3, 5, 0, -1,
    -- filter=84 channel=119
    3, 4, -2, 0, 4, -5, 0, 0, 1,
    -- filter=84 channel=120
    -1, -7, -2, -5, 7, -1, 0, -2, 3,
    -- filter=84 channel=121
    2, -1, 0, 4, -4, -1, 4, -1, 3,
    -- filter=84 channel=122
    1, -6, 1, -3, -4, 0, 2, -7, -3,
    -- filter=84 channel=123
    -6, -1, 5, -2, -4, 4, 4, 1, 3,
    -- filter=84 channel=124
    -4, 4, 1, -6, 7, 3, 4, -6, 2,
    -- filter=84 channel=125
    -7, -1, -6, -1, -3, -4, -3, 2, -2,
    -- filter=84 channel=126
    2, 6, -8, 0, -6, -6, -6, 6, -6,
    -- filter=84 channel=127
    2, 6, -1, -1, 3, 2, -2, -5, 0,
    -- filter=85 channel=0
    2, 0, -6, 7, -18, -19, 8, -1, -1,
    -- filter=85 channel=1
    10, -13, -5, 8, -14, -11, 17, -12, -1,
    -- filter=85 channel=2
    4, -4, 6, 2, -5, 4, 3, -3, 1,
    -- filter=85 channel=3
    2, 0, -5, 2, 2, 2, -6, -1, -11,
    -- filter=85 channel=4
    -1, 0, 6, -2, -7, 3, -6, -7, 0,
    -- filter=85 channel=5
    18, -4, 3, 6, -1, 1, -1, -11, 4,
    -- filter=85 channel=6
    -7, -3, 3, -6, 12, -6, -1, 12, -1,
    -- filter=85 channel=7
    4, 0, -4, 2, 0, 0, 5, -6, 0,
    -- filter=85 channel=8
    2, 0, -1, -7, 2, -9, -2, 12, -7,
    -- filter=85 channel=9
    0, 3, 4, -9, -5, 6, -1, -5, 6,
    -- filter=85 channel=10
    3, 11, 5, -13, 0, 3, -3, -4, 4,
    -- filter=85 channel=11
    -8, 8, 3, -6, 0, -3, -13, -2, -6,
    -- filter=85 channel=12
    3, 2, -1, 12, 7, -11, 6, 4, -12,
    -- filter=85 channel=13
    0, 12, -6, -7, 10, 2, 10, -1, 3,
    -- filter=85 channel=14
    4, 6, 5, -7, 4, 7, -5, 7, -3,
    -- filter=85 channel=15
    -8, 11, -2, -4, 6, 3, -14, 11, -6,
    -- filter=85 channel=16
    6, -1, -7, -3, 0, 7, 0, -3, 7,
    -- filter=85 channel=17
    0, 6, 2, 2, -2, -6, 4, 7, -6,
    -- filter=85 channel=18
    -6, 13, -6, -12, 12, -3, -7, 1, -6,
    -- filter=85 channel=19
    -1, -5, 2, -7, 3, -2, -6, 0, -2,
    -- filter=85 channel=20
    -8, 7, -2, -4, 10, -10, -4, 15, 2,
    -- filter=85 channel=21
    -4, -3, -2, 0, -2, 10, 0, 1, 12,
    -- filter=85 channel=22
    1, 8, 2, -1, 5, -1, -4, 7, 3,
    -- filter=85 channel=23
    -5, 7, -9, -18, 24, -14, -18, 19, -8,
    -- filter=85 channel=24
    0, 1, -7, -5, -4, 2, 5, 2, -2,
    -- filter=85 channel=25
    2, 5, 0, -8, 2, 0, -2, 2, 4,
    -- filter=85 channel=26
    8, -2, 1, -4, -4, 2, 2, -8, 0,
    -- filter=85 channel=27
    -4, 2, -4, -13, 9, -9, -18, 11, 4,
    -- filter=85 channel=28
    0, 0, -4, 7, 1, -1, -6, -5, 5,
    -- filter=85 channel=29
    -4, 13, 5, -9, 20, -4, -4, 4, 2,
    -- filter=85 channel=30
    -1, 2, 4, 1, 2, -2, -8, 0, 0,
    -- filter=85 channel=31
    4, -1, -11, -30, 2, -1, -25, 3, 12,
    -- filter=85 channel=32
    -5, 14, 0, -11, 14, -10, 2, 11, 3,
    -- filter=85 channel=33
    -5, 7, 1, -12, 1, -8, 2, 6, -3,
    -- filter=85 channel=34
    11, 6, -1, 5, 31, -12, 1, 29, -5,
    -- filter=85 channel=35
    -1, 1, 4, 0, 0, 1, -6, -2, 0,
    -- filter=85 channel=36
    -6, -2, -5, -10, 0, 4, -3, 1, 3,
    -- filter=85 channel=37
    13, -12, -5, 4, -11, -8, 12, -6, -5,
    -- filter=85 channel=38
    -2, 0, 2, -8, 10, 2, -12, 4, 4,
    -- filter=85 channel=39
    2, 8, -4, -4, 11, -8, -10, 2, -3,
    -- filter=85 channel=40
    0, 1, -8, -6, -3, 4, -9, 0, 3,
    -- filter=85 channel=41
    -9, 5, 5, 18, 0, -6, 19, 9, 5,
    -- filter=85 channel=42
    -1, -8, -2, -1, -8, 4, 3, -8, 0,
    -- filter=85 channel=43
    -2, 9, -7, -7, 8, -7, -7, 0, 0,
    -- filter=85 channel=44
    1, -3, -3, 2, -4, -1, 2, -3, 1,
    -- filter=85 channel=45
    7, 2, 2, 3, -3, 0, 0, -6, 5,
    -- filter=85 channel=46
    0, -4, 0, 0, 6, 0, -3, -4, -4,
    -- filter=85 channel=47
    5, 0, 2, 0, -3, 5, 6, -16, 6,
    -- filter=85 channel=48
    -5, 3, 6, 0, 1, 7, -9, -10, 4,
    -- filter=85 channel=49
    -12, 1, -7, -11, 4, -7, 0, 4, 1,
    -- filter=85 channel=50
    3, 4, -1, -7, 6, 1, -14, 3, 6,
    -- filter=85 channel=51
    -4, 1, 7, -2, -5, 1, -6, -1, -1,
    -- filter=85 channel=52
    0, 13, -4, -9, 10, -1, -2, 19, -1,
    -- filter=85 channel=53
    -1, 8, 0, 1, 9, 3, 0, 8, -6,
    -- filter=85 channel=54
    5, 4, 1, -1, -6, -5, -7, 6, -1,
    -- filter=85 channel=55
    -10, 11, -2, -10, 20, -8, -12, 12, -4,
    -- filter=85 channel=56
    -2, -2, 0, -5, 1, -7, 2, 12, 0,
    -- filter=85 channel=57
    5, 0, 0, 4, -3, -4, -2, -5, 6,
    -- filter=85 channel=58
    13, -8, -3, 10, -10, -3, 5, 3, 5,
    -- filter=85 channel=59
    3, 7, -1, -3, 4, 12, 4, 0, 15,
    -- filter=85 channel=60
    -3, 3, 6, -6, -7, 3, 6, 4, -5,
    -- filter=85 channel=61
    -5, 9, -1, -1, 13, 2, -6, 10, -2,
    -- filter=85 channel=62
    6, 6, -4, -1, -4, 3, 0, -3, -2,
    -- filter=85 channel=63
    2, -2, 4, 1, -2, -4, 7, -4, -5,
    -- filter=85 channel=64
    -1, 0, 4, 2, 4, 1, -7, -4, -4,
    -- filter=85 channel=65
    5, 4, 2, 6, 0, -5, 4, -4, -5,
    -- filter=85 channel=66
    9, 5, -3, 10, 8, -2, 19, 7, 0,
    -- filter=85 channel=67
    6, -7, 2, -4, -3, 5, 0, -2, -2,
    -- filter=85 channel=68
    -7, 3, 4, 0, -6, -1, -8, 0, -6,
    -- filter=85 channel=69
    0, -3, -8, 8, -3, -3, -2, 6, 1,
    -- filter=85 channel=70
    6, 12, -3, -8, 17, 1, -13, 2, -11,
    -- filter=85 channel=71
    7, -4, 5, 0, 4, 1, 0, 0, -8,
    -- filter=85 channel=72
    3, 1, -8, -3, 3, 4, -2, 5, 2,
    -- filter=85 channel=73
    -8, 2, 3, -3, 14, 0, -2, 6, -2,
    -- filter=85 channel=74
    2, 11, -12, -10, 15, -13, -14, 17, -2,
    -- filter=85 channel=75
    11, -7, 2, 11, -12, -4, 16, -17, -5,
    -- filter=85 channel=76
    0, 3, -6, -10, 9, 0, -14, 10, 1,
    -- filter=85 channel=77
    0, -3, -4, -1, 0, 2, 7, -2, -4,
    -- filter=85 channel=78
    10, -3, -3, 0, 6, -5, -1, 6, -2,
    -- filter=85 channel=79
    -3, 11, -2, -15, 11, -9, 7, 11, -4,
    -- filter=85 channel=80
    8, 5, 0, -14, -3, 6, -8, -13, 12,
    -- filter=85 channel=81
    -3, 5, -4, 5, -4, 5, 6, 7, -2,
    -- filter=85 channel=82
    8, -5, 5, 4, -4, 0, 1, -4, 0,
    -- filter=85 channel=83
    1, 1, -5, 0, -7, 0, -1, 1, 5,
    -- filter=85 channel=84
    -4, 8, -11, -8, 11, -8, -3, 4, 1,
    -- filter=85 channel=85
    0, -1, -5, -4, -3, -6, 3, -6, -3,
    -- filter=85 channel=86
    3, 2, -9, 3, 3, -16, 6, 3, -2,
    -- filter=85 channel=87
    -6, 12, -3, -3, 11, -4, 1, 13, 0,
    -- filter=85 channel=88
    -9, 1, -4, -11, 0, 2, -1, 4, 1,
    -- filter=85 channel=89
    -2, 6, 8, -9, 6, 5, -9, -3, 0,
    -- filter=85 channel=90
    6, -4, 0, -6, 12, -2, -8, 10, -2,
    -- filter=85 channel=91
    -9, 10, -2, -19, 18, -5, -16, 12, 5,
    -- filter=85 channel=92
    5, 0, -6, -6, 11, 6, 5, 10, 5,
    -- filter=85 channel=93
    4, 2, 5, 2, -10, 5, 0, -8, 11,
    -- filter=85 channel=94
    1, 2, 1, -6, -2, 1, 6, -6, 0,
    -- filter=85 channel=95
    3, -6, -5, -3, 4, -7, 5, -3, -2,
    -- filter=85 channel=96
    3, 0, 2, -1, 4, -1, -1, -1, 3,
    -- filter=85 channel=97
    5, -1, 5, 1, 3, -9, -6, -7, 5,
    -- filter=85 channel=98
    0, 4, -2, -18, 9, -7, -5, 1, 7,
    -- filter=85 channel=99
    0, 7, -7, -21, 26, -9, -10, 28, -1,
    -- filter=85 channel=100
    6, -2, -4, 7, 7, 4, 11, 5, 0,
    -- filter=85 channel=101
    -7, -7, -5, 5, -2, 0, -1, -7, 4,
    -- filter=85 channel=102
    0, -6, -1, 6, 7, 0, -3, 0, 7,
    -- filter=85 channel=103
    1, -2, 0, 4, 1, 0, -6, -13, 8,
    -- filter=85 channel=104
    4, 3, -6, -15, -3, 8, -2, -3, 7,
    -- filter=85 channel=105
    5, 14, 1, -6, 12, -3, -9, 13, 3,
    -- filter=85 channel=106
    -4, -6, -5, -2, 5, 7, -10, -2, 5,
    -- filter=85 channel=107
    -6, 6, -1, 2, 16, -6, 0, 15, -11,
    -- filter=85 channel=108
    0, 1, 0, 1, 1, 6, 4, 5, 7,
    -- filter=85 channel=109
    -10, 13, -2, -14, 16, 0, -2, 11, 6,
    -- filter=85 channel=110
    8, 7, 0, -4, 2, 5, -9, 11, 0,
    -- filter=85 channel=111
    0, 2, 3, -4, 0, 6, -1, 4, 5,
    -- filter=85 channel=112
    -4, 4, -5, -5, 1, -6, 0, -1, 0,
    -- filter=85 channel=113
    -5, 0, 0, -10, 2, -2, -3, 4, 1,
    -- filter=85 channel=114
    4, 10, -2, 0, 13, -14, 7, 11, -8,
    -- filter=85 channel=115
    0, 0, 2, -6, 0, 3, -1, 8, -5,
    -- filter=85 channel=116
    -14, 10, -3, -16, 9, 9, -9, 3, 16,
    -- filter=85 channel=117
    -7, 2, 1, -6, -5, -1, -1, -2, -2,
    -- filter=85 channel=118
    -4, -3, 5, -2, 0, -2, 1, -6, 5,
    -- filter=85 channel=119
    -4, 8, 0, -3, 18, 0, -2, 15, -3,
    -- filter=85 channel=120
    -9, 9, -10, -25, 17, -6, -18, 25, -11,
    -- filter=85 channel=121
    2, -4, -5, -8, 0, 7, -4, 1, -1,
    -- filter=85 channel=122
    3, -1, -1, -7, -9, 0, -7, -7, 11,
    -- filter=85 channel=123
    7, 8, 5, -2, 16, 4, -3, 9, -6,
    -- filter=85 channel=124
    7, 11, -1, 3, 11, 0, -2, 4, 3,
    -- filter=85 channel=125
    1, -2, -6, -17, 5, 0, -12, 12, 6,
    -- filter=85 channel=126
    1, 6, 7, 2, 0, -3, -2, -9, 7,
    -- filter=85 channel=127
    -3, 4, -2, 5, -2, -6, 10, -3, -1,
    -- filter=86 channel=0
    -4, -4, -1, 3, -3, 8, 1, -1, -1,
    -- filter=86 channel=1
    0, 5, -3, 8, 5, -4, 8, -1, -3,
    -- filter=86 channel=2
    -1, 1, -2, 5, 7, -5, -1, 3, -3,
    -- filter=86 channel=3
    -2, 3, -1, 0, 7, -6, 3, 1, 0,
    -- filter=86 channel=4
    2, -1, -2, 5, 1, 0, -5, 5, -6,
    -- filter=86 channel=5
    -5, -2, 5, 0, 7, 4, -6, 6, 0,
    -- filter=86 channel=6
    0, 5, -4, 0, -2, -5, -3, -6, 0,
    -- filter=86 channel=7
    -3, -4, 0, 5, 0, -6, 6, -2, 4,
    -- filter=86 channel=8
    -4, -5, 3, 1, 6, 2, -5, -6, 0,
    -- filter=86 channel=9
    5, 2, 6, 2, -6, -2, -1, 3, 0,
    -- filter=86 channel=10
    2, 5, -6, -7, -3, -7, 0, 4, 2,
    -- filter=86 channel=11
    -1, 5, 1, -5, 5, 1, -3, -2, -3,
    -- filter=86 channel=12
    -6, -7, -5, -4, 1, -7, 0, 4, -1,
    -- filter=86 channel=13
    0, -6, -2, -2, 4, 0, 3, 0, -8,
    -- filter=86 channel=14
    -7, 0, -1, -6, -5, -3, 0, 4, 4,
    -- filter=86 channel=15
    -7, -8, -1, 4, 3, 5, -5, -1, 0,
    -- filter=86 channel=16
    -5, 8, 0, 6, 0, -4, 5, -2, -4,
    -- filter=86 channel=17
    -3, 0, -1, -2, -5, -3, -4, 6, -5,
    -- filter=86 channel=18
    -3, 1, 0, 6, 0, 0, -2, -2, -6,
    -- filter=86 channel=19
    -6, 6, 7, -6, 4, 1, 3, 0, 5,
    -- filter=86 channel=20
    0, -1, 3, 6, 1, 5, 8, 8, -1,
    -- filter=86 channel=21
    3, 6, 1, 4, 0, 0, -3, 2, -2,
    -- filter=86 channel=22
    1, 3, -6, 3, 5, 4, -6, 2, 5,
    -- filter=86 channel=23
    4, 4, -7, 0, 2, 1, -8, -2, 0,
    -- filter=86 channel=24
    0, -4, -4, -6, 7, 2, 4, 5, -5,
    -- filter=86 channel=25
    -4, -7, 0, 4, -3, 0, -6, 0, -7,
    -- filter=86 channel=26
    1, -2, 6, -6, 1, -5, -3, 2, 0,
    -- filter=86 channel=27
    -8, 0, 2, -6, -1, -8, -5, -2, 0,
    -- filter=86 channel=28
    -7, 5, 5, -5, 5, -7, 1, -3, -7,
    -- filter=86 channel=29
    -4, 5, 6, -1, 3, -2, 6, 0, -4,
    -- filter=86 channel=30
    -1, -7, 4, 1, 0, 5, 6, -3, 1,
    -- filter=86 channel=31
    -3, -4, -4, -4, -3, -7, -6, -7, 1,
    -- filter=86 channel=32
    -8, 5, -7, -1, 5, -1, -7, -4, -5,
    -- filter=86 channel=33
    3, -7, -8, -9, -8, -3, -7, -5, -5,
    -- filter=86 channel=34
    5, 6, 2, -6, -2, 6, 2, -7, 0,
    -- filter=86 channel=35
    1, -5, -6, -6, -3, -2, -1, -2, 7,
    -- filter=86 channel=36
    -3, -4, 7, 5, 3, -4, 7, -6, 6,
    -- filter=86 channel=37
    -1, 0, 2, -4, -6, 3, -1, -1, 8,
    -- filter=86 channel=38
    2, -5, -5, 0, 0, -4, -3, 3, -7,
    -- filter=86 channel=39
    6, 0, 0, 4, 1, 3, -4, -4, 6,
    -- filter=86 channel=40
    -5, -4, -4, 0, 2, 5, 0, -5, 0,
    -- filter=86 channel=41
    11, -6, -8, 9, 1, 3, 6, -5, 1,
    -- filter=86 channel=42
    2, 0, 6, -4, -1, 5, 0, 6, 5,
    -- filter=86 channel=43
    6, 0, 2, 0, -3, 5, 3, 4, -7,
    -- filter=86 channel=44
    0, -6, 0, 5, -3, 8, -3, -4, 0,
    -- filter=86 channel=45
    -3, -4, 7, -3, 0, -3, 0, -5, -2,
    -- filter=86 channel=46
    7, 5, 6, -4, 5, 2, 5, 0, 0,
    -- filter=86 channel=47
    6, 0, 2, 4, 3, 6, -5, 3, 2,
    -- filter=86 channel=48
    4, -2, -4, 1, -8, 4, 4, -4, 2,
    -- filter=86 channel=49
    5, -6, -6, 3, -2, -5, -1, 4, -4,
    -- filter=86 channel=50
    -8, -3, 3, -5, -7, -1, 4, -5, -2,
    -- filter=86 channel=51
    3, 3, -4, -1, -1, -2, -5, 1, -5,
    -- filter=86 channel=52
    -1, 1, -4, 0, 5, 0, 7, -2, 6,
    -- filter=86 channel=53
    -3, 3, -2, -1, 1, -4, 6, 7, -1,
    -- filter=86 channel=54
    -3, 3, 0, 4, -7, -4, -1, -1, 4,
    -- filter=86 channel=55
    2, 2, -1, 0, 4, -5, 0, -3, -1,
    -- filter=86 channel=56
    1, -3, -2, 5, 3, 0, 2, -3, 0,
    -- filter=86 channel=57
    2, -6, -2, 1, -4, -6, -5, 4, 0,
    -- filter=86 channel=58
    -1, 0, 0, -4, 4, 5, 4, -4, 8,
    -- filter=86 channel=59
    -7, -9, -8, -3, -1, -6, -6, -5, -4,
    -- filter=86 channel=60
    1, 0, -7, -4, -5, 0, 3, -4, -4,
    -- filter=86 channel=61
    -6, 2, 7, 0, 7, 6, -6, 4, -5,
    -- filter=86 channel=62
    7, -1, 0, -1, 1, -4, -3, -1, -3,
    -- filter=86 channel=63
    -1, -2, -5, 4, -2, 8, 1, 6, 5,
    -- filter=86 channel=64
    -1, -7, -2, 5, -6, 6, 3, 6, 4,
    -- filter=86 channel=65
    -2, 3, -3, -6, 6, -5, -2, -1, -6,
    -- filter=86 channel=66
    0, -7, -2, 6, -1, -3, -1, -7, 4,
    -- filter=86 channel=67
    -3, 0, 0, 7, -2, 7, 7, 4, -4,
    -- filter=86 channel=68
    6, -3, -4, -6, -3, -1, -3, -4, 7,
    -- filter=86 channel=69
    -5, -6, 1, -1, 5, -5, -3, 4, 0,
    -- filter=86 channel=70
    -9, -5, 1, -10, 2, 5, 1, 1, -2,
    -- filter=86 channel=71
    -5, 2, 5, -2, 1, -5, -4, -7, -4,
    -- filter=86 channel=72
    -7, 2, -2, -7, 1, -7, 7, 3, 6,
    -- filter=86 channel=73
    2, -6, -2, 5, 1, 0, -3, -7, 1,
    -- filter=86 channel=74
    0, -9, -4, -2, 2, 2, 4, 1, -5,
    -- filter=86 channel=75
    5, 2, 0, 5, 0, 0, 1, -7, -4,
    -- filter=86 channel=76
    0, -5, -3, 0, 2, 6, 6, 6, 5,
    -- filter=86 channel=77
    2, 6, -5, 2, -5, 5, -4, -5, 4,
    -- filter=86 channel=78
    -1, -6, 0, -3, 3, 8, -1, 3, 6,
    -- filter=86 channel=79
    3, 0, -1, 2, -9, -8, -4, -5, -1,
    -- filter=86 channel=80
    -3, 0, -5, -1, 1, 0, 6, 4, 6,
    -- filter=86 channel=81
    3, 5, -6, 0, -2, 0, 5, 4, 3,
    -- filter=86 channel=82
    6, 3, 0, -1, 2, 0, 3, -5, 2,
    -- filter=86 channel=83
    -7, -6, 6, 4, 0, 2, 6, 1, -4,
    -- filter=86 channel=84
    4, -7, 5, -6, 1, 3, -6, 2, 2,
    -- filter=86 channel=85
    -1, -1, -2, -5, 6, 7, 2, 0, -6,
    -- filter=86 channel=86
    6, -1, 3, 0, 5, 5, 0, 4, -3,
    -- filter=86 channel=87
    2, 6, 6, 5, 6, 0, 3, 0, -2,
    -- filter=86 channel=88
    -4, 1, 4, 0, -6, 2, 5, 2, 2,
    -- filter=86 channel=89
    -8, -1, -2, 3, -8, -5, 2, -9, -6,
    -- filter=86 channel=90
    -6, 6, -2, 7, 1, -3, 0, 0, 4,
    -- filter=86 channel=91
    -3, 0, -2, -8, 2, -7, -1, 3, -8,
    -- filter=86 channel=92
    2, 4, -6, 0, -4, 3, -1, 0, -5,
    -- filter=86 channel=93
    2, 4, 1, -4, -5, 6, 1, 2, -7,
    -- filter=86 channel=94
    -5, -4, 2, 0, -5, -5, -3, -5, 3,
    -- filter=86 channel=95
    -4, 4, 3, 0, -2, 2, -7, 1, 0,
    -- filter=86 channel=96
    4, -4, 0, -1, -5, -5, -5, 5, -1,
    -- filter=86 channel=97
    4, 5, 2, 2, 6, 0, 6, 5, 2,
    -- filter=86 channel=98
    0, 5, 3, -5, 5, -2, -3, -4, -1,
    -- filter=86 channel=99
    -5, -1, 1, -2, 0, 5, 0, -5, 0,
    -- filter=86 channel=100
    6, -6, 0, 6, -7, 2, 2, 0, 0,
    -- filter=86 channel=101
    -5, -5, 7, 3, 1, 3, 5, -5, 0,
    -- filter=86 channel=102
    5, -3, -5, -5, -5, 1, 2, -1, -3,
    -- filter=86 channel=103
    3, -7, -7, -7, -1, 1, -3, -1, -2,
    -- filter=86 channel=104
    -5, -7, -7, 2, -1, -7, 5, 3, -3,
    -- filter=86 channel=105
    6, 5, -3, 1, 0, 1, 5, 6, -1,
    -- filter=86 channel=106
    -4, 0, 0, 4, 4, 7, 7, 0, 2,
    -- filter=86 channel=107
    4, 4, -5, 1, -4, 0, 7, 7, 0,
    -- filter=86 channel=108
    2, -2, -2, 8, -4, 2, 5, 5, -1,
    -- filter=86 channel=109
    0, -8, 0, 1, 1, 3, 0, 0, -8,
    -- filter=86 channel=110
    0, -3, -1, 0, -5, -2, 4, 2, -7,
    -- filter=86 channel=111
    -3, -5, 0, -2, -6, 6, -2, -6, 5,
    -- filter=86 channel=112
    -8, -7, -6, 0, 2, -2, -2, -7, 4,
    -- filter=86 channel=113
    -5, 1, 3, 5, -3, 2, -6, -3, 4,
    -- filter=86 channel=114
    -7, -6, -4, -1, -6, -5, 6, -6, -2,
    -- filter=86 channel=115
    -6, -5, -6, 4, 6, 3, 3, 7, 6,
    -- filter=86 channel=116
    3, -3, -7, -5, -4, -8, 0, -6, -1,
    -- filter=86 channel=117
    2, -4, -2, 7, -7, 0, -1, 5, 4,
    -- filter=86 channel=118
    -2, 0, -6, -1, 3, 3, 0, 6, -4,
    -- filter=86 channel=119
    3, 1, 1, 0, -1, 6, 1, 2, 3,
    -- filter=86 channel=120
    0, -2, 3, -6, 2, -2, 0, 1, -7,
    -- filter=86 channel=121
    -3, 0, 4, 7, -1, 4, 4, -2, -1,
    -- filter=86 channel=122
    1, -3, -1, -6, 6, 1, 0, 5, 2,
    -- filter=86 channel=123
    -7, 2, -7, -7, 0, -4, 2, 6, 5,
    -- filter=86 channel=124
    -5, -1, -1, 4, 3, -6, -3, 1, -6,
    -- filter=86 channel=125
    3, 3, 3, -1, -4, -2, 5, 3, -5,
    -- filter=86 channel=126
    -4, -7, 3, 6, 1, 1, 9, -3, 1,
    -- filter=86 channel=127
    -5, -6, 4, 2, -5, -3, 0, 5, -1,
    -- filter=87 channel=0
    -12, -22, -20, -12, -18, -10, -2, -5, 0,
    -- filter=87 channel=1
    -2, -16, 1, -16, -21, -7, -6, -14, -3,
    -- filter=87 channel=2
    6, 9, 0, -4, 1, 2, -2, 5, -2,
    -- filter=87 channel=3
    -9, -15, -13, -8, -3, -3, 0, -4, -1,
    -- filter=87 channel=4
    -5, -2, -4, -12, -10, -4, -2, -4, 1,
    -- filter=87 channel=5
    -11, -16, -8, -16, -6, 2, -8, -6, 1,
    -- filter=87 channel=6
    2, 0, 0, 0, -8, -9, 0, 4, -3,
    -- filter=87 channel=7
    6, -2, 2, 1, 7, 4, 6, -6, 0,
    -- filter=87 channel=8
    1, -4, -1, -1, 3, 3, -4, 4, -5,
    -- filter=87 channel=9
    1, 0, 4, 1, 6, 2, -3, 0, 0,
    -- filter=87 channel=10
    -6, -5, 0, 0, 8, 11, 6, -2, 2,
    -- filter=87 channel=11
    -1, 0, 5, -3, 15, 12, 1, 3, 13,
    -- filter=87 channel=12
    5, -13, 2, 6, 1, -3, -4, -6, -2,
    -- filter=87 channel=13
    5, -5, -5, 7, 6, 7, 4, -1, 1,
    -- filter=87 channel=14
    3, -1, 4, 3, -2, -7, -7, 2, -5,
    -- filter=87 channel=15
    -7, -7, -8, 4, 5, 1, 7, -1, 0,
    -- filter=87 channel=16
    -1, -8, 0, -2, -5, -4, -8, -9, 0,
    -- filter=87 channel=17
    0, 6, 0, -6, 6, -2, -1, -2, 3,
    -- filter=87 channel=18
    -8, -16, -20, 1, -6, 2, 0, -2, 3,
    -- filter=87 channel=19
    0, 4, 7, 0, -5, 4, 2, -4, 4,
    -- filter=87 channel=20
    8, 3, 0, 5, 7, 16, 3, 7, 14,
    -- filter=87 channel=21
    2, -1, 15, 1, -1, 14, -8, 3, 8,
    -- filter=87 channel=22
    -1, -6, -3, 7, -3, -4, 1, -3, -8,
    -- filter=87 channel=23
    0, -23, -18, 3, 6, 0, 14, 16, 0,
    -- filter=87 channel=24
    1, 2, 0, 1, 4, -6, -6, 1, -2,
    -- filter=87 channel=25
    0, -11, -7, 0, -3, 5, -9, -7, -6,
    -- filter=87 channel=26
    2, -1, 10, -9, 0, -1, 0, 5, 2,
    -- filter=87 channel=27
    -9, -13, -17, 3, 5, 3, -6, 4, -3,
    -- filter=87 channel=28
    0, 2, 2, 2, -4, 7, -2, 6, -4,
    -- filter=87 channel=29
    3, 1, -7, 2, 15, 0, 2, 11, 15,
    -- filter=87 channel=30
    -10, -6, -9, -2, 1, 3, -2, -9, 7,
    -- filter=87 channel=31
    -2, 5, 0, 5, 11, 19, -9, 7, 7,
    -- filter=87 channel=32
    1, -18, -18, 8, -2, 2, -2, -9, 6,
    -- filter=87 channel=33
    -7, -14, -11, -5, -8, -1, -2, -4, 6,
    -- filter=87 channel=34
    6, -13, -4, 7, -11, -4, -1, -2, 2,
    -- filter=87 channel=35
    1, -6, 0, 1, 5, -7, -7, -2, 0,
    -- filter=87 channel=36
    2, 15, 10, 11, 3, 3, 4, 2, 0,
    -- filter=87 channel=37
    -16, -17, 1, -16, -21, 0, -8, -15, 2,
    -- filter=87 channel=38
    -7, -3, 4, 5, 0, 4, 5, 2, 9,
    -- filter=87 channel=39
    8, 7, 7, 9, 6, 4, 2, 2, 8,
    -- filter=87 channel=40
    1, 6, 5, 7, 8, -3, 4, 9, 10,
    -- filter=87 channel=41
    5, 7, -11, 0, -8, -9, 10, -14, 0,
    -- filter=87 channel=42
    0, -3, 2, 0, 0, 0, 0, 3, -3,
    -- filter=87 channel=43
    -9, -17, -5, 5, -4, -1, 12, 3, -5,
    -- filter=87 channel=44
    -12, -4, -3, -9, -12, 0, -8, -2, 4,
    -- filter=87 channel=45
    0, -2, -3, 5, 1, 3, 7, 0, 4,
    -- filter=87 channel=46
    3, 2, -9, 0, -7, -1, 2, -9, -2,
    -- filter=87 channel=47
    -12, -7, -4, -16, 2, 6, -11, -3, 0,
    -- filter=87 channel=48
    -1, -7, 6, 0, 7, 10, -10, 1, 4,
    -- filter=87 channel=49
    2, -2, -9, 8, 5, -1, -4, -3, 0,
    -- filter=87 channel=50
    1, -6, 0, 9, 10, 6, -5, 3, -3,
    -- filter=87 channel=51
    3, 3, -4, -1, 7, -5, -4, 6, -5,
    -- filter=87 channel=52
    4, -13, -5, 1, -3, -1, 10, -6, -3,
    -- filter=87 channel=53
    -2, -8, -7, 6, 3, 9, 0, 0, 3,
    -- filter=87 channel=54
    -4, 5, 5, 5, -5, 0, 6, 2, 5,
    -- filter=87 channel=55
    0, -14, -15, 5, 14, 0, 7, 5, 9,
    -- filter=87 channel=56
    -6, -3, -3, 0, 5, -5, 2, 1, -4,
    -- filter=87 channel=57
    6, 6, 0, -3, 4, -6, 7, -5, -1,
    -- filter=87 channel=58
    3, 0, -2, -7, -2, -5, -7, -1, 4,
    -- filter=87 channel=59
    0, -5, 4, -7, 12, 13, 2, -1, -2,
    -- filter=87 channel=60
    4, 1, 0, 1, -5, 6, -3, -2, -5,
    -- filter=87 channel=61
    6, -3, 11, -1, 0, 2, -1, 3, 4,
    -- filter=87 channel=62
    -2, -1, 2, 4, -7, -2, 4, 8, 1,
    -- filter=87 channel=63
    3, -6, 3, -2, 2, 6, 0, -5, 5,
    -- filter=87 channel=64
    -3, 1, 4, 8, 8, 6, 0, 0, 8,
    -- filter=87 channel=65
    -3, -1, 0, 0, -4, 2, 4, -5, 4,
    -- filter=87 channel=66
    6, -5, -4, 13, -11, 1, -2, 0, -3,
    -- filter=87 channel=67
    4, 0, -5, 4, 3, -2, -4, 4, 5,
    -- filter=87 channel=68
    -6, 4, 7, -2, 0, 8, -6, 4, 6,
    -- filter=87 channel=69
    3, 2, 6, 6, -7, 2, 6, 0, -2,
    -- filter=87 channel=70
    2, -14, -18, -1, -3, 0, 0, -3, -6,
    -- filter=87 channel=71
    -7, -9, -9, 3, 0, 1, 6, 3, 1,
    -- filter=87 channel=72
    0, 6, 1, 1, 18, 11, -3, 7, 11,
    -- filter=87 channel=73
    1, -11, -3, -2, 1, 9, 3, 1, 5,
    -- filter=87 channel=74
    4, -11, 0, 15, -5, 4, 1, 4, 3,
    -- filter=87 channel=75
    -8, -24, -17, -15, -14, -12, -10, -12, -6,
    -- filter=87 channel=76
    -4, -1, -6, 2, 3, 0, 7, 11, 12,
    -- filter=87 channel=77
    -1, -5, 3, 4, -2, 1, -2, -2, -3,
    -- filter=87 channel=78
    0, -1, -3, -2, 6, 7, -4, 2, 3,
    -- filter=87 channel=79
    -9, -22, -17, -4, -4, 5, -4, -2, 5,
    -- filter=87 channel=80
    1, 0, 6, 0, 18, 15, -6, 0, 3,
    -- filter=87 channel=81
    1, -5, -4, 3, -6, 5, 7, 5, 2,
    -- filter=87 channel=82
    -2, -6, -5, -5, 4, -1, -1, 3, 7,
    -- filter=87 channel=83
    5, 10, 3, 5, 14, 9, -7, 5, 0,
    -- filter=87 channel=84
    -3, -2, -6, 5, 6, 7, 0, 3, -7,
    -- filter=87 channel=85
    6, -4, 4, -2, -1, 0, -3, -7, 5,
    -- filter=87 channel=86
    -2, -5, -4, 6, -7, 0, -5, -3, 3,
    -- filter=87 channel=87
    0, 0, 2, 11, 0, 0, 3, 2, 3,
    -- filter=87 channel=88
    9, 10, 13, 12, 11, 12, 10, 11, 1,
    -- filter=87 channel=89
    -4, -15, -10, 4, 10, 9, 5, 7, 0,
    -- filter=87 channel=90
    8, -4, 1, -3, 3, -1, -1, 6, 0,
    -- filter=87 channel=91
    7, -7, -7, 13, 4, 10, -3, 3, -6,
    -- filter=87 channel=92
    4, -3, -10, -3, -6, -7, 2, 4, 6,
    -- filter=87 channel=93
    -18, -5, 6, -17, -2, -6, -9, -7, -6,
    -- filter=87 channel=94
    3, -5, -5, 6, 0, -5, -7, 0, 3,
    -- filter=87 channel=95
    -6, -5, -2, 0, -4, 0, -3, 3, 0,
    -- filter=87 channel=96
    -6, -3, 6, -1, -3, -6, 3, 6, -3,
    -- filter=87 channel=97
    -6, -9, -3, 0, -10, -9, -7, 8, 8,
    -- filter=87 channel=98
    0, -8, -8, -4, 7, 8, -2, -7, -3,
    -- filter=87 channel=99
    5, -9, 4, 11, 17, 14, -2, 17, 0,
    -- filter=87 channel=100
    -1, -5, 3, 7, -4, 2, -4, 1, -7,
    -- filter=87 channel=101
    -1, -1, 3, -2, -6, 7, 0, -3, 8,
    -- filter=87 channel=102
    6, -4, 6, -3, -1, 1, 3, -5, -6,
    -- filter=87 channel=103
    -18, -17, 2, -20, -10, 6, -10, -9, 6,
    -- filter=87 channel=104
    -4, -3, 4, 4, 16, 19, -3, -3, 12,
    -- filter=87 channel=105
    -5, -3, -9, 8, 0, -3, 2, 11, 5,
    -- filter=87 channel=106
    -4, -2, -1, 0, 3, 2, 9, -2, -4,
    -- filter=87 channel=107
    -3, -13, -9, 8, -12, 0, 10, 1, 1,
    -- filter=87 channel=108
    -6, -7, 3, -5, 4, 4, 6, -2, 2,
    -- filter=87 channel=109
    -7, -19, -5, 6, 8, 5, 4, 2, 0,
    -- filter=87 channel=110
    -3, -5, -9, 0, 7, 0, -5, 3, 0,
    -- filter=87 channel=111
    4, 6, -1, 4, -4, -3, -1, -1, 6,
    -- filter=87 channel=112
    -2, -7, -10, 6, -6, 5, 2, 0, -4,
    -- filter=87 channel=113
    0, -12, -7, -6, -8, 0, 0, 11, -4,
    -- filter=87 channel=114
    -5, -17, -15, 7, -15, -8, 7, -7, -8,
    -- filter=87 channel=115
    1, -5, 4, 6, 1, 6, 5, -3, -4,
    -- filter=87 channel=116
    5, 2, 5, 10, 4, 5, -5, -5, 0,
    -- filter=87 channel=117
    -3, 2, -3, -3, 1, 2, 3, -3, -5,
    -- filter=87 channel=118
    3, 6, -5, -4, -2, -2, 0, 6, -6,
    -- filter=87 channel=119
    4, -1, -2, 10, -1, -6, -2, -2, 0,
    -- filter=87 channel=120
    -6, -2, -4, 21, 4, 2, 7, 1, 5,
    -- filter=87 channel=121
    3, 0, -4, 7, -1, 6, 6, -7, -6,
    -- filter=87 channel=122
    -20, 2, 12, -20, 3, 5, -20, 0, 0,
    -- filter=87 channel=123
    4, -10, -9, 6, -5, -2, -5, 2, 2,
    -- filter=87 channel=124
    4, 4, -9, -4, 5, 8, -1, -4, -1,
    -- filter=87 channel=125
    -6, 1, -2, 4, 12, 10, 0, 9, 5,
    -- filter=87 channel=126
    -6, -8, -13, -3, 0, -4, -2, 4, 11,
    -- filter=87 channel=127
    -5, -3, 6, 0, -5, -5, 2, -7, 1,
    -- filter=88 channel=0
    -3, -11, -9, -4, -2, -8, 16, 13, 11,
    -- filter=88 channel=1
    -11, -8, 0, 0, 3, 3, 16, 13, 5,
    -- filter=88 channel=2
    6, 2, -3, 5, 3, 0, 2, -7, -6,
    -- filter=88 channel=3
    0, -5, -8, -6, -4, -5, 7, 1, 5,
    -- filter=88 channel=4
    6, -6, -11, 0, -2, -4, 0, -4, 6,
    -- filter=88 channel=5
    -17, -18, -9, -8, -10, 0, 10, 11, 11,
    -- filter=88 channel=6
    7, 7, -4, 11, -1, -7, -4, -12, -7,
    -- filter=88 channel=7
    -1, -1, 0, -6, 2, -3, 4, 0, 3,
    -- filter=88 channel=8
    3, -3, -6, -4, 0, -3, 2, 1, 3,
    -- filter=88 channel=9
    -6, -8, -2, 6, 8, 0, 4, -1, 3,
    -- filter=88 channel=10
    -10, 3, 7, 3, 5, 5, 0, -6, -4,
    -- filter=88 channel=11
    16, 6, 7, 7, 4, -9, -12, -12, -11,
    -- filter=88 channel=12
    -1, -1, -3, -8, -6, -5, -9, -11, 5,
    -- filter=88 channel=13
    1, 8, 4, 1, 5, -5, -9, -7, -4,
    -- filter=88 channel=14
    1, -2, 2, -1, 3, -3, 1, 6, 7,
    -- filter=88 channel=15
    3, 10, -3, 10, 2, 0, -4, -17, -8,
    -- filter=88 channel=16
    -12, -10, -9, -10, -7, 7, 7, 4, 1,
    -- filter=88 channel=17
    5, 1, 0, 5, 3, -5, -1, -6, -6,
    -- filter=88 channel=18
    10, 23, -2, 14, 6, -6, -2, -16, -8,
    -- filter=88 channel=19
    0, -6, 6, 5, -5, 1, -3, 7, 7,
    -- filter=88 channel=20
    18, 19, -4, 6, 1, -12, -11, -21, -15,
    -- filter=88 channel=21
    -5, -13, 1, 3, 0, 7, 6, 9, 8,
    -- filter=88 channel=22
    1, 1, -6, 6, 7, -6, 5, 5, -5,
    -- filter=88 channel=23
    -1, 15, 4, 5, -1, -8, -7, -7, -12,
    -- filter=88 channel=24
    -3, 2, -2, -1, -2, 2, 0, -6, -6,
    -- filter=88 channel=25
    -17, 6, 0, 5, 5, 2, 6, 6, -1,
    -- filter=88 channel=26
    -10, -11, -10, 0, 1, -1, -8, 3, -5,
    -- filter=88 channel=27
    0, 14, 0, 6, 13, 4, 3, -8, -2,
    -- filter=88 channel=28
    -4, 0, 1, -2, 5, 5, -2, 2, 4,
    -- filter=88 channel=29
    19, 8, -3, 15, 0, -13, -10, -22, -10,
    -- filter=88 channel=30
    -9, 0, 0, -4, 1, 0, 0, 4, 0,
    -- filter=88 channel=31
    -1, 1, 0, 2, -2, 5, -5, 8, 13,
    -- filter=88 channel=32
    -1, 10, -2, 6, 6, -5, -4, -6, -16,
    -- filter=88 channel=33
    -12, 0, -4, -2, 13, 3, -2, 0, -1,
    -- filter=88 channel=34
    -8, -6, 0, -3, -3, -8, -11, -2, -3,
    -- filter=88 channel=35
    -1, -7, -2, -4, -4, 3, 0, -1, 6,
    -- filter=88 channel=36
    0, 3, -1, -1, 2, -2, -7, -14, -3,
    -- filter=88 channel=37
    -4, -13, -4, 1, 0, 0, 8, 18, 6,
    -- filter=88 channel=38
    -7, -3, -5, -3, 2, 8, 1, -1, 4,
    -- filter=88 channel=39
    12, 1, -4, 7, 0, 1, 0, -4, -13,
    -- filter=88 channel=40
    5, 3, 4, 9, 1, -7, -7, -3, -7,
    -- filter=88 channel=41
    -2, -15, 1, -21, -10, -6, -4, -10, 0,
    -- filter=88 channel=42
    4, -1, -7, -1, 0, 4, 2, 1, -1,
    -- filter=88 channel=43
    0, -5, -3, -5, -2, -8, -1, -6, -10,
    -- filter=88 channel=44
    -5, -15, -4, -9, 0, 3, 5, 8, 15,
    -- filter=88 channel=45
    5, 3, 3, 0, 6, 1, 7, 2, 3,
    -- filter=88 channel=46
    -1, 5, 5, -5, -3, 3, 3, -6, -4,
    -- filter=88 channel=47
    -15, -12, 0, -11, -2, 8, 10, 6, 7,
    -- filter=88 channel=48
    -3, -8, 2, 1, 0, -2, 3, -4, 4,
    -- filter=88 channel=49
    11, 13, 4, 13, -4, 0, -4, -9, -10,
    -- filter=88 channel=50
    -4, -1, 0, 5, 4, -2, 0, 9, 1,
    -- filter=88 channel=51
    -2, 0, 2, 2, -3, -5, 1, 4, 0,
    -- filter=88 channel=52
    6, -3, 1, -8, -6, -7, -6, -13, -4,
    -- filter=88 channel=53
    6, 10, 0, 0, 5, -7, -9, -13, -9,
    -- filter=88 channel=54
    -4, 0, 5, 6, 1, 6, 0, 2, -4,
    -- filter=88 channel=55
    10, 19, 2, 5, 10, 0, -19, -22, -15,
    -- filter=88 channel=56
    6, -10, -7, -3, -9, 3, -6, -1, -2,
    -- filter=88 channel=57
    -5, 3, 3, 3, 1, -7, -5, -5, 4,
    -- filter=88 channel=58
    3, -16, 0, -6, 1, 2, 0, 2, 9,
    -- filter=88 channel=59
    -14, -1, 9, 4, 0, 7, -1, -1, 10,
    -- filter=88 channel=60
    2, 5, -4, -2, 6, -6, 6, 5, 1,
    -- filter=88 channel=61
    1, 3, -4, -3, 1, 5, 0, -5, -4,
    -- filter=88 channel=62
    -1, -4, -2, 7, -6, 1, -4, 4, 3,
    -- filter=88 channel=63
    -3, -15, -6, -6, -3, 4, -4, 6, 6,
    -- filter=88 channel=64
    7, -2, 2, -5, -8, 4, 0, 2, 0,
    -- filter=88 channel=65
    -6, -7, 6, -4, 5, -2, 7, 0, -5,
    -- filter=88 channel=66
    -6, -9, 4, -15, -1, -4, -11, -12, 0,
    -- filter=88 channel=67
    3, 1, 0, 0, 5, -5, -6, -5, 2,
    -- filter=88 channel=68
    4, 7, 0, 8, 1, 0, -1, -5, -7,
    -- filter=88 channel=69
    -6, 0, -3, 5, 5, 3, -5, -2, 0,
    -- filter=88 channel=70
    3, 5, 0, -3, 4, 0, 4, -2, -1,
    -- filter=88 channel=71
    -5, -7, -5, -1, 5, -6, 10, 4, 1,
    -- filter=88 channel=72
    -3, 2, -3, -6, 9, 7, -7, 1, 2,
    -- filter=88 channel=73
    3, 12, 3, 5, 0, 0, -12, -14, -3,
    -- filter=88 channel=74
    4, 4, 7, -6, -6, -3, -3, -6, 3,
    -- filter=88 channel=75
    -18, -6, -2, -11, 0, 2, 13, 10, 14,
    -- filter=88 channel=76
    11, 20, -4, 4, -2, -5, -9, -14, -19,
    -- filter=88 channel=77
    -3, 3, -4, -6, -7, 5, -1, -6, 6,
    -- filter=88 channel=78
    -7, 0, 1, 6, -7, 5, -2, 5, 3,
    -- filter=88 channel=79
    9, 14, 5, 1, 15, -6, -5, -11, -15,
    -- filter=88 channel=80
    -13, -3, -4, -7, 3, 8, -1, 5, 15,
    -- filter=88 channel=81
    1, -1, -7, -4, -2, -3, 1, -7, 7,
    -- filter=88 channel=82
    5, -7, 1, -2, 2, 1, 8, -3, 1,
    -- filter=88 channel=83
    2, 2, 0, -2, 5, 3, -3, 0, -7,
    -- filter=88 channel=84
    4, 2, 5, 8, -6, -2, -10, -5, -12,
    -- filter=88 channel=85
    1, 0, -3, 0, -4, -2, 4, -4, 3,
    -- filter=88 channel=86
    -2, -3, -8, 3, -12, -3, 0, -5, 8,
    -- filter=88 channel=87
    7, 0, 1, 2, -6, 1, -5, -9, -5,
    -- filter=88 channel=88
    -4, -4, 5, -4, 4, 10, -1, -11, 6,
    -- filter=88 channel=89
    -6, 7, 8, 9, 12, 2, 2, -4, -6,
    -- filter=88 channel=90
    2, -6, 5, -9, -5, 5, -6, -2, 6,
    -- filter=88 channel=91
    8, 4, 3, 2, 1, -5, -1, -13, -2,
    -- filter=88 channel=92
    -1, -3, 3, -6, -2, 1, 1, 4, -2,
    -- filter=88 channel=93
    -14, -11, -3, 4, -7, 1, 8, 7, 7,
    -- filter=88 channel=94
    5, -3, 1, -1, 6, 0, -6, -6, 6,
    -- filter=88 channel=95
    -3, 7, -1, 0, -4, 2, -2, -6, -8,
    -- filter=88 channel=96
    -1, 2, 7, 3, -5, 0, 0, 3, -5,
    -- filter=88 channel=97
    -3, -3, -5, -2, -3, -4, 9, 10, -1,
    -- filter=88 channel=98
    -8, -2, 3, 7, 2, 2, 1, 4, -2,
    -- filter=88 channel=99
    6, 5, 5, -3, 5, 10, -22, -11, -1,
    -- filter=88 channel=100
    -2, -4, -3, -6, -5, -3, -9, -6, -5,
    -- filter=88 channel=101
    -2, -5, -4, -5, 3, 0, 0, 1, 4,
    -- filter=88 channel=102
    4, 1, -5, -6, 2, 1, 0, -6, 5,
    -- filter=88 channel=103
    -10, -17, -4, 0, -3, 9, 14, 22, 15,
    -- filter=88 channel=104
    -15, -2, -3, -4, -2, 8, 5, -4, 1,
    -- filter=88 channel=105
    7, 13, -5, 1, 0, -10, -5, -18, -9,
    -- filter=88 channel=106
    -2, 1, 4, 5, 0, 2, -8, -9, -6,
    -- filter=88 channel=107
    14, 11, 4, 14, 3, -12, -4, -14, -9,
    -- filter=88 channel=108
    -5, -5, -3, -11, -6, -5, -1, 0, -7,
    -- filter=88 channel=109
    -6, 9, 3, -2, 10, -2, 0, -15, -11,
    -- filter=88 channel=110
    -5, 0, -5, -2, 5, 0, -10, 2, 9,
    -- filter=88 channel=111
    2, -4, 2, -9, 0, -5, -6, 3, -5,
    -- filter=88 channel=112
    -9, -5, 5, 3, 0, -5, 7, 2, 7,
    -- filter=88 channel=113
    -7, 5, -2, -5, -1, 9, 0, 0, 2,
    -- filter=88 channel=114
    -2, 3, 0, 6, 4, -12, 1, -19, -9,
    -- filter=88 channel=115
    -3, 0, 6, -1, 2, -6, -4, 6, -4,
    -- filter=88 channel=116
    5, 8, -4, 10, 0, 0, -4, -14, -6,
    -- filter=88 channel=117
    -3, 4, 2, 6, -4, -2, 5, 2, 0,
    -- filter=88 channel=118
    2, -3, 6, -4, -1, -5, -6, -6, -4,
    -- filter=88 channel=119
    -3, -12, -4, 0, -9, -6, -1, -9, -5,
    -- filter=88 channel=120
    14, 12, -4, 3, 2, -3, -17, -18, -1,
    -- filter=88 channel=121
    -5, -8, 10, -9, 0, 4, -7, -5, -3,
    -- filter=88 channel=122
    -21, -32, -8, -13, -5, 20, 6, 22, 28,
    -- filter=88 channel=123
    3, -2, 0, -8, -10, 3, 4, 3, -9,
    -- filter=88 channel=124
    12, 1, 4, 5, -2, -7, -4, -11, -4,
    -- filter=88 channel=125
    -7, -3, 7, 4, 10, 8, -13, -4, 3,
    -- filter=88 channel=126
    2, -3, 8, -4, 4, 0, 0, -6, 5,
    -- filter=88 channel=127
    2, -8, -1, 1, 4, 4, 0, -8, -1,
    -- filter=89 channel=0
    15, 14, -1, 12, 2, -1, -8, -6, -14,
    -- filter=89 channel=1
    12, 5, -1, 7, 7, -5, -5, -1, -2,
    -- filter=89 channel=2
    -3, 2, 1, 6, 13, 10, -5, 5, -5,
    -- filter=89 channel=3
    -1, 28, 17, 1, 0, -2, 14, 8, -1,
    -- filter=89 channel=4
    3, 10, 12, 25, 35, 9, 3, 12, 4,
    -- filter=89 channel=5
    12, 10, 4, 11, -3, 4, -9, 7, 3,
    -- filter=89 channel=6
    7, 13, -1, -2, 7, -4, -6, -12, -11,
    -- filter=89 channel=7
    -1, 3, -5, -5, -5, 3, 4, -4, 3,
    -- filter=89 channel=8
    7, -4, 8, -5, 0, 4, -7, 5, -4,
    -- filter=89 channel=9
    -6, 2, -1, -7, -2, -2, 5, 11, 6,
    -- filter=89 channel=10
    -11, -7, 7, 1, -11, -7, 12, 11, 5,
    -- filter=89 channel=11
    -5, 12, 7, 1, 8, 5, -3, -3, -1,
    -- filter=89 channel=12
    -5, 3, 5, 4, 0, -5, 0, -10, 6,
    -- filter=89 channel=13
    -10, -4, 10, 0, -13, -4, 0, 0, 1,
    -- filter=89 channel=14
    7, -6, -2, 1, 1, -4, 6, 0, -2,
    -- filter=89 channel=15
    6, 6, 18, 4, -1, 3, -1, -10, -1,
    -- filter=89 channel=16
    -1, -5, 1, 0, 0, -10, 3, 8, 7,
    -- filter=89 channel=17
    4, 0, 0, -2, 7, -2, 1, -3, -5,
    -- filter=89 channel=18
    4, -1, 0, 3, -7, 3, -12, -1, -13,
    -- filter=89 channel=19
    4, 0, -4, 5, 1, 4, 1, -7, -1,
    -- filter=89 channel=20
    -6, 14, 10, 0, 7, 14, -10, -15, -15,
    -- filter=89 channel=21
    -7, -16, -13, -10, -16, -6, 4, 13, 12,
    -- filter=89 channel=22
    5, 11, 4, 2, -8, -7, -8, 0, -5,
    -- filter=89 channel=23
    -11, 17, 10, -15, -11, 6, 7, 1, -1,
    -- filter=89 channel=24
    -4, -5, 7, 5, -2, 1, -3, -6, -5,
    -- filter=89 channel=25
    -4, -7, -9, 10, -8, -10, 10, 13, 3,
    -- filter=89 channel=26
    -8, 2, -12, 6, 3, -3, 5, 0, 0,
    -- filter=89 channel=27
    -7, -2, 5, 0, -5, -9, 6, 5, -11,
    -- filter=89 channel=28
    -6, -5, -6, -2, -6, 0, 5, 5, -7,
    -- filter=89 channel=29
    0, 15, 13, 3, 13, 12, -15, -18, -7,
    -- filter=89 channel=30
    -5, 2, -3, 6, 5, -2, 7, -1, 3,
    -- filter=89 channel=31
    -22, -22, -8, -7, -21, -5, 25, 25, 15,
    -- filter=89 channel=32
    6, -3, 7, 1, 0, -2, -4, 2, -6,
    -- filter=89 channel=33
    -8, -1, 0, -3, -22, -14, -2, 4, 2,
    -- filter=89 channel=34
    0, 11, 3, -7, -11, 4, 9, -3, -5,
    -- filter=89 channel=35
    0, 0, -1, 0, -2, -7, 4, -4, -5,
    -- filter=89 channel=36
    -10, -10, -6, 5, 0, 4, 7, 1, 5,
    -- filter=89 channel=37
    -1, -9, -10, 11, 0, 3, -10, 2, 0,
    -- filter=89 channel=38
    0, -1, -6, -4, -12, -4, 13, 12, -5,
    -- filter=89 channel=39
    -1, 0, 7, -1, 3, 0, -10, 0, -5,
    -- filter=89 channel=40
    -1, -1, 8, -5, -3, -2, -7, -2, 0,
    -- filter=89 channel=41
    6, -9, 4, 18, -5, -11, -3, -8, -6,
    -- filter=89 channel=42
    1, -2, -3, 5, 0, -1, 0, -4, -4,
    -- filter=89 channel=43
    8, 20, 15, -4, 2, 6, -1, -11, -10,
    -- filter=89 channel=44
    -5, -3, 1, -3, -1, 3, 4, 2, -4,
    -- filter=89 channel=45
    0, 0, 1, 1, -1, 5, -2, -1, -5,
    -- filter=89 channel=46
    -2, -5, -4, -2, 4, 3, -6, -5, 3,
    -- filter=89 channel=47
    -6, -13, -1, -5, -1, -6, 0, 8, 4,
    -- filter=89 channel=48
    -4, -23, -16, 3, 8, 5, 5, 8, 7,
    -- filter=89 channel=49
    3, -5, 11, 9, 17, 6, -7, -3, 1,
    -- filter=89 channel=50
    -13, -2, -3, 0, -14, -1, 8, 6, -1,
    -- filter=89 channel=51
    -5, 2, 0, 7, 0, -4, 6, 2, 0,
    -- filter=89 channel=52
    7, 8, 9, 0, -4, 0, -3, -11, -3,
    -- filter=89 channel=53
    -5, 10, 2, -4, 5, 10, 2, 0, -1,
    -- filter=89 channel=54
    5, 0, 0, 2, 7, 4, -3, 3, 4,
    -- filter=89 channel=55
    1, 3, 2, -2, 0, 0, -3, 1, -1,
    -- filter=89 channel=56
    1, 0, 0, -2, 5, 1, 4, 0, -2,
    -- filter=89 channel=57
    6, -3, 4, 4, 5, -4, -4, -5, -2,
    -- filter=89 channel=58
    9, 11, 3, 6, 7, 3, -3, -8, -3,
    -- filter=89 channel=59
    -18, -15, 0, -9, -8, -8, 14, 5, 7,
    -- filter=89 channel=60
    -6, -2, 0, 4, -6, 4, 6, -4, 1,
    -- filter=89 channel=61
    1, 1, 3, 0, 0, 6, 5, 1, -3,
    -- filter=89 channel=62
    4, -4, -1, 4, -3, -6, 7, 7, 5,
    -- filter=89 channel=63
    3, 6, -4, 7, 7, 3, -2, -4, -2,
    -- filter=89 channel=64
    -8, -3, -2, 4, 0, 6, -4, 2, -3,
    -- filter=89 channel=65
    -2, -2, -4, -5, 1, 0, 0, 4, 3,
    -- filter=89 channel=66
    9, -6, -5, -1, -10, -2, -2, 1, 0,
    -- filter=89 channel=67
    0, 6, 6, 0, -6, -6, 4, -4, -2,
    -- filter=89 channel=68
    4, 5, 5, 0, 12, 9, -1, -6, -6,
    -- filter=89 channel=69
    -4, -3, -7, -5, 3, 0, 6, 0, 6,
    -- filter=89 channel=70
    2, -4, 9, 0, -10, 0, 4, -5, -7,
    -- filter=89 channel=71
    -1, 0, 9, -8, -8, -6, 3, 4, 6,
    -- filter=89 channel=72
    -7, -16, -6, -10, -19, 0, 19, 22, 7,
    -- filter=89 channel=73
    3, -2, 2, 0, -1, 3, 4, 0, -5,
    -- filter=89 channel=74
    0, -3, 6, -12, 0, -6, 2, -1, -1,
    -- filter=89 channel=75
    7, 12, 3, 11, -2, -11, -6, 9, 4,
    -- filter=89 channel=76
    5, 11, 3, -6, 2, -4, -3, -13, -14,
    -- filter=89 channel=77
    2, 3, -6, 4, 6, 1, 0, -7, 0,
    -- filter=89 channel=78
    1, -4, 0, 2, 0, 9, 7, -4, -5,
    -- filter=89 channel=79
    -2, 3, 3, 0, -14, -11, -8, 0, -15,
    -- filter=89 channel=80
    -15, -16, -2, -8, -10, -16, 18, 23, 7,
    -- filter=89 channel=81
    0, 6, 5, 0, 5, -6, -5, 0, -2,
    -- filter=89 channel=82
    -3, -2, 3, -3, 3, 1, -4, 0, 4,
    -- filter=89 channel=83
    -1, -17, -11, 6, 10, -6, 7, 0, 8,
    -- filter=89 channel=84
    -3, 3, 9, 2, 10, 6, -9, -2, -1,
    -- filter=89 channel=85
    -3, 0, 1, 4, 1, -4, 0, -1, -1,
    -- filter=89 channel=86
    3, 1, 4, 0, -4, -3, 1, -7, -3,
    -- filter=89 channel=87
    3, 9, 7, -1, 2, 3, -6, -1, -1,
    -- filter=89 channel=88
    -2, -8, -1, -9, -6, -1, 10, 0, -2,
    -- filter=89 channel=89
    -3, 0, 0, -1, -19, -5, 7, 11, 3,
    -- filter=89 channel=90
    -7, 1, 9, 0, 0, -2, 10, 2, 0,
    -- filter=89 channel=91
    -11, -2, 5, -2, 0, 0, 6, 1, 3,
    -- filter=89 channel=92
    0, 12, 10, 0, -3, 2, 3, 3, -5,
    -- filter=89 channel=93
    0, -13, -2, 11, 9, 5, 5, 6, 0,
    -- filter=89 channel=94
    -3, -2, 1, 3, -2, 7, -3, -3, 0,
    -- filter=89 channel=95
    -4, 8, 0, 2, 1, 3, 3, 2, 3,
    -- filter=89 channel=96
    2, 0, -4, 0, -2, -3, 3, -2, 5,
    -- filter=89 channel=97
    -4, 15, 8, -7, -3, 7, 10, 2, -2,
    -- filter=89 channel=98
    -12, -9, -6, -9, -13, -3, 0, 16, 8,
    -- filter=89 channel=99
    -3, -10, 7, -10, -6, -3, 12, 5, -2,
    -- filter=89 channel=100
    5, 6, -2, 2, -3, 3, -3, 0, 2,
    -- filter=89 channel=101
    9, -2, 8, 10, 22, 18, 7, 10, -5,
    -- filter=89 channel=102
    1, -5, -2, -4, -2, -4, 6, 0, -1,
    -- filter=89 channel=103
    -4, 1, -3, -2, -5, -3, 12, 22, 4,
    -- filter=89 channel=104
    -16, -26, -6, -4, -6, -11, 8, 16, 15,
    -- filter=89 channel=105
    0, 15, 6, -5, 5, -2, 0, -5, -12,
    -- filter=89 channel=106
    4, 1, -4, 2, 7, -2, 1, 1, -7,
    -- filter=89 channel=107
    7, 14, 10, 4, 9, 12, -4, -6, -18,
    -- filter=89 channel=108
    13, 7, 0, 12, 5, -1, 1, 4, -2,
    -- filter=89 channel=109
    -6, -17, 5, -4, -11, -7, -3, 7, -1,
    -- filter=89 channel=110
    2, -6, 3, 0, -5, -5, 6, 3, 7,
    -- filter=89 channel=111
    -2, -1, -5, -3, 6, 4, -5, 6, -1,
    -- filter=89 channel=112
    -3, -7, -2, -7, -6, -1, 2, 2, -5,
    -- filter=89 channel=113
    1, 5, 5, -9, -19, -3, 12, 4, -5,
    -- filter=89 channel=114
    8, 11, 6, 20, 5, 2, -9, -21, -12,
    -- filter=89 channel=115
    -6, 3, -7, -6, -2, 0, -3, -2, -7,
    -- filter=89 channel=116
    -7, -18, 0, 3, 0, -5, 5, 11, 0,
    -- filter=89 channel=117
    -1, 0, 5, 0, -3, 0, 7, 6, 7,
    -- filter=89 channel=118
    2, 6, -1, 2, 3, -6, -5, 1, 1,
    -- filter=89 channel=119
    1, 2, 9, -4, 0, 6, -2, -8, 1,
    -- filter=89 channel=120
    -7, 0, 12, 0, 3, 11, 3, -8, -12,
    -- filter=89 channel=121
    0, -1, 1, 0, -12, -10, 1, 3, 1,
    -- filter=89 channel=122
    -16, -19, -3, -12, -11, -12, 5, 16, 5,
    -- filter=89 channel=123
    -6, -1, 3, -2, 3, 7, 1, -6, -6,
    -- filter=89 channel=124
    -2, 0, 0, -1, 0, 7, -9, -13, -7,
    -- filter=89 channel=125
    -12, -19, 0, 4, -13, -2, 16, 14, 7,
    -- filter=89 channel=126
    -5, 0, 0, -9, -6, 1, 8, 9, -4,
    -- filter=89 channel=127
    7, 4, -2, 7, -6, -2, -2, -6, 1,
    -- filter=90 channel=0
    -10, -22, -3, -16, -27, -14, -13, -19, 1,
    -- filter=90 channel=1
    0, -6, -11, -11, -17, -4, -18, -15, 8,
    -- filter=90 channel=2
    -5, 3, -2, 2, 2, 3, -2, -6, 0,
    -- filter=90 channel=3
    -7, -10, -8, -3, -1, -13, 0, 8, -2,
    -- filter=90 channel=4
    -3, 7, 5, -14, -6, -10, -10, -16, -7,
    -- filter=90 channel=5
    -12, -9, -4, -2, -18, 0, -6, -9, 1,
    -- filter=90 channel=6
    2, 1, -1, 0, 1, 1, -1, -3, -13,
    -- filter=90 channel=7
    -5, -2, 1, 6, 4, -4, 6, -5, 6,
    -- filter=90 channel=8
    2, 6, -4, -8, -8, 0, -9, -12, -1,
    -- filter=90 channel=9
    -3, -2, 0, 6, 2, 1, -5, 5, -3,
    -- filter=90 channel=10
    -6, -6, 2, 1, 14, 0, -1, 0, 1,
    -- filter=90 channel=11
    0, 3, 7, -3, 4, -1, 3, -9, -8,
    -- filter=90 channel=12
    0, -10, 0, 1, -10, 2, -4, -5, -1,
    -- filter=90 channel=13
    7, 0, -2, -5, -2, -2, -1, -12, -7,
    -- filter=90 channel=14
    3, -6, 0, 2, 2, -3, 6, 6, 4,
    -- filter=90 channel=15
    10, 4, -1, -4, -1, 4, -7, -13, -9,
    -- filter=90 channel=16
    -5, -1, -11, 0, 4, -7, 3, 0, 9,
    -- filter=90 channel=17
    -4, -6, -4, -4, -3, 2, 6, -3, 0,
    -- filter=90 channel=18
    5, 0, 2, -2, -5, -2, -19, -17, -17,
    -- filter=90 channel=19
    -4, 0, 1, -3, 3, 2, -6, -1, 7,
    -- filter=90 channel=20
    0, 0, -2, 2, -5, 3, -1, -8, -21,
    -- filter=90 channel=21
    -2, -4, -10, -1, 1, 6, 1, 8, 4,
    -- filter=90 channel=22
    8, 0, -6, -2, -5, 0, 0, -6, -9,
    -- filter=90 channel=23
    8, 7, -3, 16, 12, 4, 2, 5, 1,
    -- filter=90 channel=24
    -4, -5, 0, 1, 6, -6, 0, 4, -4,
    -- filter=90 channel=25
    6, -8, 11, 5, -4, 0, -2, -4, 6,
    -- filter=90 channel=26
    -11, 2, -9, -9, -9, -6, 0, -10, 0,
    -- filter=90 channel=27
    10, 3, 6, -3, 12, 10, -14, -11, -1,
    -- filter=90 channel=28
    6, 6, -1, 5, 6, 3, 3, 2, 0,
    -- filter=90 channel=29
    6, 12, -1, -2, -4, 1, -9, -5, -20,
    -- filter=90 channel=30
    -3, -8, -2, 0, 2, 5, 1, -10, 4,
    -- filter=90 channel=31
    -11, -7, -10, 12, 24, 16, 9, 18, 11,
    -- filter=90 channel=32
    17, 1, 3, -2, -11, 7, -14, -9, -4,
    -- filter=90 channel=33
    8, -9, 6, 4, 0, 13, -7, 0, 5,
    -- filter=90 channel=34
    4, -8, 10, -4, -3, -10, -7, -4, 8,
    -- filter=90 channel=35
    -4, -2, 6, 5, 1, -5, 3, -6, 1,
    -- filter=90 channel=36
    4, 2, -4, -1, 10, -4, 6, -4, -7,
    -- filter=90 channel=37
    -11, -19, -9, -8, -16, -1, -15, -8, 0,
    -- filter=90 channel=38
    -1, -7, 0, 0, 0, 10, 7, 6, -2,
    -- filter=90 channel=39
    -4, -2, -6, -1, 6, 0, -3, -10, 0,
    -- filter=90 channel=40
    -8, 2, 7, -5, 4, -3, 0, -2, -4,
    -- filter=90 channel=41
    0, 4, 3, -9, -14, -7, -7, -18, -16,
    -- filter=90 channel=42
    -2, -2, 0, -2, 4, -8, 0, -1, -7,
    -- filter=90 channel=43
    1, -5, -1, 3, -4, -3, -7, -11, -4,
    -- filter=90 channel=44
    -6, -8, -4, -12, -5, 0, -3, -2, 5,
    -- filter=90 channel=45
    -5, 6, -4, 0, -9, 3, -2, 0, 6,
    -- filter=90 channel=46
    5, 0, 4, 3, -9, -4, 1, -6, -2,
    -- filter=90 channel=47
    -17, -7, -6, -4, 7, 8, 2, 7, 19,
    -- filter=90 channel=48
    3, -5, -3, -10, 7, 0, -11, -2, 3,
    -- filter=90 channel=49
    9, 0, 13, -7, -8, 4, -13, -4, -13,
    -- filter=90 channel=50
    7, -1, -2, 9, 13, 6, 2, 6, 0,
    -- filter=90 channel=51
    3, -1, 3, 0, 7, 4, 0, 3, 3,
    -- filter=90 channel=52
    0, 3, 6, 3, -2, -2, 0, -12, 2,
    -- filter=90 channel=53
    -5, 5, -2, 9, -4, 0, 0, -4, -1,
    -- filter=90 channel=54
    6, 3, 7, 7, -2, -6, 1, -3, 0,
    -- filter=90 channel=55
    10, 9, 5, -1, 0, 8, -4, -1, -7,
    -- filter=90 channel=56
    -1, -5, 1, -5, -1, -2, -6, -8, 0,
    -- filter=90 channel=57
    1, -1, -4, 0, 0, -1, -6, -5, -7,
    -- filter=90 channel=58
    -6, -5, -3, -7, -11, -12, -4, -2, -7,
    -- filter=90 channel=59
    -1, -8, 4, -7, 6, 6, 0, -3, 3,
    -- filter=90 channel=60
    -1, 3, -7, -5, 5, 6, 1, 5, -2,
    -- filter=90 channel=61
    4, -2, -4, -3, -10, -4, -3, -10, -1,
    -- filter=90 channel=62
    3, 0, 6, 0, -2, 5, 0, -4, -6,
    -- filter=90 channel=63
    -8, 2, -10, -2, -7, -3, 0, 2, -3,
    -- filter=90 channel=64
    -3, 4, 5, -4, 4, -8, 3, 6, 3,
    -- filter=90 channel=65
    0, -4, -3, -1, -5, 0, -6, 3, -6,
    -- filter=90 channel=66
    -3, -5, 5, -7, -9, -1, 1, -5, 4,
    -- filter=90 channel=67
    4, 5, -4, -7, -6, -7, -1, -2, -3,
    -- filter=90 channel=68
    -1, 7, 5, -4, 3, -7, 2, 0, -1,
    -- filter=90 channel=69
    -7, 2, 6, -4, -6, -6, -3, 3, -6,
    -- filter=90 channel=70
    14, 4, 5, 9, 0, 5, 0, -6, 0,
    -- filter=90 channel=71
    0, 3, 1, 0, 6, 0, 5, 10, 6,
    -- filter=90 channel=72
    0, -6, 0, 1, 24, 5, 1, 11, 9,
    -- filter=90 channel=73
    3, 6, 2, 3, 1, -2, -7, -13, 0,
    -- filter=90 channel=74
    0, 0, 3, 10, 0, 1, 2, -7, 2,
    -- filter=90 channel=75
    -2, -9, -9, -11, -11, -6, -16, -9, 2,
    -- filter=90 channel=76
    2, 6, 5, 2, -6, -4, -3, -15, -12,
    -- filter=90 channel=77
    -2, 2, 3, 0, -1, -3, -6, 3, 2,
    -- filter=90 channel=78
    -8, -1, -8, 2, 5, 1, -8, 3, 7,
    -- filter=90 channel=79
    12, -5, 8, -7, -6, 6, -6, -25, -4,
    -- filter=90 channel=80
    0, -10, -1, 1, 16, 0, 2, 7, 7,
    -- filter=90 channel=81
    0, 0, 5, -6, -1, -6, 1, -6, 6,
    -- filter=90 channel=82
    -2, 1, 0, 3, 5, -2, -4, 8, -6,
    -- filter=90 channel=83
    -2, 4, 4, -7, 0, -3, -12, 0, -4,
    -- filter=90 channel=84
    8, 1, 12, 2, -3, 7, -5, -10, -9,
    -- filter=90 channel=85
    2, -3, 3, 0, -5, 3, 5, 2, -3,
    -- filter=90 channel=86
    -2, -12, 0, -7, -7, -3, 0, -1, -4,
    -- filter=90 channel=87
    7, -4, 5, -4, -1, 4, 0, -3, 0,
    -- filter=90 channel=88
    2, 2, 6, -1, 5, 2, 4, 1, 5,
    -- filter=90 channel=89
    13, -2, 0, 3, 4, 6, 6, 1, 5,
    -- filter=90 channel=90
    -8, -2, 0, -4, -3, -2, 5, 0, 10,
    -- filter=90 channel=91
    10, 1, 5, 1, 7, 10, -2, -5, -5,
    -- filter=90 channel=92
    -1, 1, 6, 6, -5, 1, 2, -5, 1,
    -- filter=90 channel=93
    -5, -10, -11, -9, -1, 1, -1, -15, -4,
    -- filter=90 channel=94
    -2, 5, 0, 0, 0, -7, -6, -6, -7,
    -- filter=90 channel=95
    0, -2, 2, -7, -5, 4, 1, -3, 5,
    -- filter=90 channel=96
    -5, -4, 5, -3, 0, 2, 0, 2, 4,
    -- filter=90 channel=97
    -3, -1, -4, 6, -3, -4, 2, 6, 0,
    -- filter=90 channel=98
    0, 2, 4, 2, 3, 13, -11, 0, 4,
    -- filter=90 channel=99
    -3, 6, -4, 10, 16, 14, 6, 5, 6,
    -- filter=90 channel=100
    4, 0, -1, 0, -1, -5, -3, 3, 0,
    -- filter=90 channel=101
    2, -4, 4, 1, -2, -1, -5, -12, 0,
    -- filter=90 channel=102
    5, -3, 1, 0, 4, 0, 3, -3, -4,
    -- filter=90 channel=103
    -7, -4, -7, -2, 6, 5, 0, 6, 17,
    -- filter=90 channel=104
    -7, -6, -5, 3, 15, 3, -2, 2, 2,
    -- filter=90 channel=105
    -2, 3, 0, 0, -5, -5, -6, -12, -15,
    -- filter=90 channel=106
    -3, 7, -2, -4, 6, -10, 5, 0, 0,
    -- filter=90 channel=107
    4, 0, 2, 1, -12, -9, -6, -18, -6,
    -- filter=90 channel=108
    3, -5, -1, -10, -4, -3, 0, -2, -1,
    -- filter=90 channel=109
    9, -1, 12, -3, 0, 16, -14, -13, 0,
    -- filter=90 channel=110
    -2, 2, 1, 5, 9, -3, 8, 0, -5,
    -- filter=90 channel=111
    2, 3, -3, 1, -1, 3, -1, -1, 2,
    -- filter=90 channel=112
    6, 2, -2, 4, 1, 9, -6, 0, 2,
    -- filter=90 channel=113
    7, 3, -4, 0, 6, 0, 4, 0, 14,
    -- filter=90 channel=114
    19, 3, -2, -12, -18, -3, -21, -33, -13,
    -- filter=90 channel=115
    0, 4, 5, -4, 3, 4, 1, 6, 0,
    -- filter=90 channel=116
    2, 9, 1, 6, 7, 0, -2, -12, -16,
    -- filter=90 channel=117
    1, 0, 5, -6, 6, 7, 7, -6, 3,
    -- filter=90 channel=118
    -7, 0, 3, 0, -7, -4, 0, -4, -4,
    -- filter=90 channel=119
    -10, 0, 3, 1, -8, 0, -10, -1, 5,
    -- filter=90 channel=120
    12, 0, 15, 8, 11, 13, -19, -18, -11,
    -- filter=90 channel=121
    3, 4, -2, 2, -8, 6, 3, -7, -6,
    -- filter=90 channel=122
    -15, -9, -12, -7, 8, 10, -1, 10, 17,
    -- filter=90 channel=123
    5, 1, 5, 2, -2, 0, 4, 2, 5,
    -- filter=90 channel=124
    -3, 4, -3, -3, -3, -3, -5, -4, -3,
    -- filter=90 channel=125
    6, 1, 8, -3, 8, 10, 0, -8, 2,
    -- filter=90 channel=126
    0, -6, 7, 4, 2, -1, -3, 0, -5,
    -- filter=90 channel=127
    0, 3, 6, 2, -8, -5, -8, 4, 0,
    -- filter=91 channel=0
    1, -9, 0, 15, -2, -2, 8, -2, -2,
    -- filter=91 channel=1
    6, 0, -2, 5, -8, 0, -6, -3, 8,
    -- filter=91 channel=2
    8, 2, -7, 2, -7, 3, 4, 6, -4,
    -- filter=91 channel=3
    -2, -5, -1, -4, -13, -7, 7, -9, 1,
    -- filter=91 channel=4
    14, 9, 2, -11, -14, -2, -7, -15, -8,
    -- filter=91 channel=5
    2, -3, -8, -5, 0, -1, 5, -3, 3,
    -- filter=91 channel=6
    -3, 6, 3, -4, -1, 2, -4, 2, 1,
    -- filter=91 channel=7
    4, -3, -2, 0, 3, 5, -5, -7, -3,
    -- filter=91 channel=8
    -3, -8, 1, -2, -12, -4, -2, 0, -1,
    -- filter=91 channel=9
    4, -2, -5, 0, 0, -6, 0, -1, -4,
    -- filter=91 channel=10
    0, -8, -3, 5, -3, 1, 5, -5, -5,
    -- filter=91 channel=11
    -2, 1, 2, 1, 6, -2, 8, -3, 3,
    -- filter=91 channel=12
    -6, -7, 10, -7, -17, 8, -7, -11, -3,
    -- filter=91 channel=13
    -7, -12, -10, 7, -2, 7, 3, -9, 5,
    -- filter=91 channel=14
    3, 6, -7, -4, 5, 2, 0, 5, 4,
    -- filter=91 channel=15
    -6, 2, -10, 11, 6, -5, 5, 2, -7,
    -- filter=91 channel=16
    -10, -10, 1, 3, 3, 4, 5, -2, 5,
    -- filter=91 channel=17
    -5, 0, -6, 4, -5, 1, -5, -1, -3,
    -- filter=91 channel=18
    9, -4, 1, 8, 4, 7, 12, 2, 7,
    -- filter=91 channel=19
    -6, -5, 1, 1, -5, -1, -4, 6, 1,
    -- filter=91 channel=20
    0, 6, 2, 4, -4, -10, 0, 5, 3,
    -- filter=91 channel=21
    -5, -5, -5, 3, 6, 0, 3, 7, 2,
    -- filter=91 channel=22
    1, -10, 0, 5, 0, 4, -1, 1, -4,
    -- filter=91 channel=23
    -15, -14, -21, -8, -5, -2, 3, 2, -9,
    -- filter=91 channel=24
    3, 0, 5, 4, 3, -3, -6, 2, -6,
    -- filter=91 channel=25
    2, -9, -3, 4, 2, 11, -4, 0, 9,
    -- filter=91 channel=26
    -3, -5, 7, -2, 5, -2, 1, -5, 5,
    -- filter=91 channel=27
    4, 0, -8, 17, -2, -3, 0, -1, 1,
    -- filter=91 channel=28
    -2, -6, -1, 2, -1, 4, -3, 6, 5,
    -- filter=91 channel=29
    -3, 3, -8, 3, 0, -7, 3, 7, -10,
    -- filter=91 channel=30
    0, -5, -2, 8, -2, 6, 2, 7, -4,
    -- filter=91 channel=31
    -20, -7, -19, 12, 7, -1, 7, 14, -3,
    -- filter=91 channel=32
    7, -12, -6, 9, -8, 2, 4, -5, 3,
    -- filter=91 channel=33
    2, -18, -4, 9, 1, 2, 3, 2, 5,
    -- filter=91 channel=34
    -12, -24, 4, -18, -21, -16, -13, -22, -13,
    -- filter=91 channel=35
    6, 0, 4, -1, 0, 5, -2, -2, -3,
    -- filter=91 channel=36
    -5, -3, -5, -8, -9, -7, -8, -5, 0,
    -- filter=91 channel=37
    9, 1, -2, 7, -9, -7, -5, -1, -5,
    -- filter=91 channel=38
    1, 0, -4, 6, 3, -1, 0, 1, 0,
    -- filter=91 channel=39
    4, 8, 2, 0, -2, -7, 1, 2, 0,
    -- filter=91 channel=40
    -9, 1, -3, -1, 5, -1, 0, -4, -1,
    -- filter=91 channel=41
    10, -13, 6, -6, -27, 10, 0, -25, 2,
    -- filter=91 channel=42
    3, 0, -8, 10, 2, 5, 8, 1, -8,
    -- filter=91 channel=43
    -3, -12, -8, -10, -5, -11, -1, -8, -9,
    -- filter=91 channel=44
    5, -8, -5, 5, -7, 2, 5, 4, -2,
    -- filter=91 channel=45
    7, 0, 6, -1, 2, 0, 7, 8, -1,
    -- filter=91 channel=46
    0, 3, -5, -4, 0, -1, -6, 1, -7,
    -- filter=91 channel=47
    -9, -14, 0, 0, 2, 12, 2, 8, 5,
    -- filter=91 channel=48
    1, -1, -1, 13, 1, 6, -3, 7, 6,
    -- filter=91 channel=49
    12, 0, -6, 7, 3, -2, 5, 0, -1,
    -- filter=91 channel=50
    -6, -4, -5, 4, 3, 7, 1, 4, -6,
    -- filter=91 channel=51
    -6, 0, 0, 0, 4, -3, 4, -1, -2,
    -- filter=91 channel=52
    -1, -1, -1, -2, -11, -9, -3, 0, -7,
    -- filter=91 channel=53
    1, 6, -7, -4, -4, 4, 0, -3, 3,
    -- filter=91 channel=54
    2, -5, 1, 6, -6, 6, -2, 0, -4,
    -- filter=91 channel=55
    -6, -4, -12, 4, -5, 0, 1, 5, -9,
    -- filter=91 channel=56
    -13, -13, -9, -5, -12, -4, -1, -7, 5,
    -- filter=91 channel=57
    0, -7, 7, -9, -7, 3, 2, -7, 6,
    -- filter=91 channel=58
    -5, -2, 0, -7, -2, -10, 0, -1, -2,
    -- filter=91 channel=59
    5, -2, 1, 10, 11, 13, 5, 8, 0,
    -- filter=91 channel=60
    3, -4, 0, 5, -7, -2, -2, -4, 1,
    -- filter=91 channel=61
    -9, -11, 3, 1, -12, 1, 1, -4, -2,
    -- filter=91 channel=62
    0, -3, 2, -7, 5, -5, 8, 4, 0,
    -- filter=91 channel=63
    8, 0, 0, 5, 0, -9, 6, -1, -3,
    -- filter=91 channel=64
    1, 0, 0, -1, 1, -6, 0, 0, 0,
    -- filter=91 channel=65
    0, -6, 1, 1, 0, 2, 2, -6, -5,
    -- filter=91 channel=66
    0, -14, 9, 0, -14, 0, -3, -9, 6,
    -- filter=91 channel=67
    -5, 5, -5, -6, 0, -6, -5, -3, -4,
    -- filter=91 channel=68
    1, -2, -2, 3, -2, 0, 3, -4, 6,
    -- filter=91 channel=69
    -4, -2, 4, 7, -3, 5, 6, -3, 5,
    -- filter=91 channel=70
    -8, -3, -15, 0, 0, -8, -2, 4, -8,
    -- filter=91 channel=71
    -4, -10, -5, -9, 4, -6, -4, 4, -5,
    -- filter=91 channel=72
    -10, -4, -3, 7, 15, 8, 3, 11, -5,
    -- filter=91 channel=73
    9, 4, -7, 4, 5, 5, -4, 4, -4,
    -- filter=91 channel=74
    -2, -4, 0, 1, -6, 3, -12, 0, 3,
    -- filter=91 channel=75
    1, -23, -16, 10, -8, -2, 3, 0, -4,
    -- filter=91 channel=76
    -3, 4, -2, 5, 2, -7, 10, -6, -3,
    -- filter=91 channel=77
    2, -6, -2, 5, -2, 2, 4, 1, 1,
    -- filter=91 channel=78
    0, 1, -1, 2, 0, -4, 1, 7, -5,
    -- filter=91 channel=79
    2, -8, -9, 7, 3, 0, 4, -3, 6,
    -- filter=91 channel=80
    1, -2, -13, 11, 15, 6, 14, 6, 4,
    -- filter=91 channel=81
    0, -4, 7, 0, 5, 7, 0, 7, -1,
    -- filter=91 channel=82
    0, -1, -5, 0, 7, -3, -4, -2, -1,
    -- filter=91 channel=83
    -5, 0, 0, 7, 10, -4, 4, 1, -6,
    -- filter=91 channel=84
    -2, 1, -7, 8, -5, 5, -6, -1, 0,
    -- filter=91 channel=85
    6, 2, 6, 1, -2, 1, -3, 0, 2,
    -- filter=91 channel=86
    -9, -6, 2, 0, -16, 3, 0, -11, -1,
    -- filter=91 channel=87
    -7, -7, 0, 0, -13, 0, -6, -6, -6,
    -- filter=91 channel=88
    -8, -5, 0, 0, -7, -10, -8, 6, -9,
    -- filter=91 channel=89
    0, -16, -1, 4, 12, 7, 1, 6, -4,
    -- filter=91 channel=90
    -18, -8, 0, -15, -13, -6, -6, 0, -8,
    -- filter=91 channel=91
    9, 0, 0, 9, -4, -1, -7, -5, -8,
    -- filter=91 channel=92
    -8, -6, -3, -2, -3, -6, 0, 0, -6,
    -- filter=91 channel=93
    10, 2, 0, 3, 0, 2, 8, 9, -4,
    -- filter=91 channel=94
    2, -5, 0, -4, -4, 6, -4, -1, 2,
    -- filter=91 channel=95
    0, 2, 1, -1, -3, 4, 3, -8, -2,
    -- filter=91 channel=96
    9, 0, 0, 0, -2, 1, -1, -4, -5,
    -- filter=91 channel=97
    -11, -2, 0, 2, 5, -7, 1, 1, -3,
    -- filter=91 channel=98
    1, -13, -9, 5, 14, 10, 6, -1, 9,
    -- filter=91 channel=99
    -20, -5, -16, -2, 0, -2, -2, 4, -8,
    -- filter=91 channel=100
    3, -5, 2, 0, -4, 3, 1, 3, 2,
    -- filter=91 channel=101
    1, 7, -2, 0, -14, -8, -7, -4, -9,
    -- filter=91 channel=102
    5, -7, -3, -6, -5, 2, 0, -3, -6,
    -- filter=91 channel=103
    -12, -14, -10, 12, 7, 8, 14, 2, 13,
    -- filter=91 channel=104
    0, 0, -3, 5, 6, 3, 4, 6, -2,
    -- filter=91 channel=105
    3, 7, 4, -1, -5, 2, -4, 0, 3,
    -- filter=91 channel=106
    -2, 0, -7, -4, -2, -5, 6, 3, -7,
    -- filter=91 channel=107
    7, -4, 6, 6, 1, -9, 5, 1, -7,
    -- filter=91 channel=108
    2, -9, 5, -8, -6, -5, -4, -8, 1,
    -- filter=91 channel=109
    -5, -6, -8, 11, 8, -3, 2, 1, 7,
    -- filter=91 channel=110
    -13, -4, 0, 1, 2, -3, 3, -5, -6,
    -- filter=91 channel=111
    2, -1, -4, 4, 3, 2, -3, 2, -2,
    -- filter=91 channel=112
    3, -5, -5, -2, -2, 0, 5, 0, -5,
    -- filter=91 channel=113
    -5, -5, -3, 2, 3, -7, -1, 0, 1,
    -- filter=91 channel=114
    11, -4, 0, 15, 5, 4, 0, 0, -2,
    -- filter=91 channel=115
    0, -1, -5, -4, 0, 0, 1, -2, 4,
    -- filter=91 channel=116
    9, 7, 0, 12, 2, 2, 3, -1, 0,
    -- filter=91 channel=117
    3, -3, -6, -5, -4, 8, 0, -6, 0,
    -- filter=91 channel=118
    1, 3, 6, 6, -2, 7, -6, 7, 6,
    -- filter=91 channel=119
    -12, -19, 2, -18, -16, -4, -10, -5, -8,
    -- filter=91 channel=120
    -8, -4, -10, 6, 9, -5, -5, 3, -9,
    -- filter=91 channel=121
    -2, -14, -2, 4, -7, 2, 8, -3, -2,
    -- filter=91 channel=122
    -15, -16, 0, 3, 4, 12, 12, 8, 18,
    -- filter=91 channel=123
    -3, -3, 2, -14, -5, -4, -10, -3, -4,
    -- filter=91 channel=124
    0, 3, 0, 3, -7, -6, -1, 5, -2,
    -- filter=91 channel=125
    -10, 2, -9, 8, 6, 6, 6, 0, 8,
    -- filter=91 channel=126
    3, -14, 0, 8, -4, 0, 10, 3, 9,
    -- filter=91 channel=127
    2, -2, 2, -1, -6, 4, 0, -1, -2,
    -- filter=92 channel=0
    -4, -7, 3, -1, 4, 9, 1, 1, 2,
    -- filter=92 channel=1
    0, 1, 1, -7, 0, 13, 3, 2, -2,
    -- filter=92 channel=2
    6, -2, 5, -3, -1, 4, -3, 0, 4,
    -- filter=92 channel=3
    -3, -5, 0, -2, -6, -4, -3, 8, 5,
    -- filter=92 channel=4
    0, 9, -4, -8, 1, -8, -4, 4, 9,
    -- filter=92 channel=5
    -9, 4, 7, -6, 2, 3, 1, 4, 1,
    -- filter=92 channel=6
    -3, -8, 4, -7, -10, 1, 3, -1, -6,
    -- filter=92 channel=7
    -6, -2, 1, -6, -4, -3, 5, 6, 0,
    -- filter=92 channel=8
    -2, 2, -3, -5, 3, -1, 4, 2, 2,
    -- filter=92 channel=9
    -1, 7, 5, 5, 6, 0, 1, 6, 2,
    -- filter=92 channel=10
    2, -4, -2, -7, -5, 0, 4, -8, -6,
    -- filter=92 channel=11
    1, -10, -3, -10, -5, 3, -5, -9, -11,
    -- filter=92 channel=12
    3, -3, 0, 5, 2, 6, -1, -5, -1,
    -- filter=92 channel=13
    -5, -14, -5, -7, 2, 2, 0, -2, 2,
    -- filter=92 channel=14
    4, -2, 5, -2, 0, 3, -5, -3, -7,
    -- filter=92 channel=15
    -11, -8, -3, -1, 0, 4, -11, 2, 7,
    -- filter=92 channel=16
    -2, -5, -1, 5, 7, 4, -2, 3, 4,
    -- filter=92 channel=17
    0, 7, -1, 0, 1, 6, -4, 7, -2,
    -- filter=92 channel=18
    -14, -17, 2, -7, -4, 0, -12, -4, 4,
    -- filter=92 channel=19
    4, -2, 3, -6, 0, 6, 6, -6, 6,
    -- filter=92 channel=20
    -4, -13, 0, -8, -2, -13, -12, -3, -4,
    -- filter=92 channel=21
    0, -6, -1, 1, 0, -4, -1, -6, -12,
    -- filter=92 channel=22
    -1, 0, 5, -6, -1, 0, -7, 2, -3,
    -- filter=92 channel=23
    -6, -9, 2, 1, -11, 0, -11, 1, -6,
    -- filter=92 channel=24
    6, 1, 1, 4, 1, 5, 6, -2, 0,
    -- filter=92 channel=25
    -2, -2, 6, -3, 1, 2, 4, 5, 11,
    -- filter=92 channel=26
    0, 3, -2, 4, -7, -4, 5, -8, 1,
    -- filter=92 channel=27
    -4, -5, 7, -3, 10, 19, -2, 1, 8,
    -- filter=92 channel=28
    -1, 2, 6, 6, -1, -5, -6, -2, 6,
    -- filter=92 channel=29
    -10, -9, 0, -4, -7, -9, -13, -12, -12,
    -- filter=92 channel=30
    0, -2, 7, -1, 10, 5, 7, 7, 2,
    -- filter=92 channel=31
    -8, -12, 0, 0, 5, -3, 3, -3, -3,
    -- filter=92 channel=32
    -10, -3, 6, -2, 3, 1, 4, 5, 13,
    -- filter=92 channel=33
    -7, -14, 1, -4, 8, 2, 1, 8, 13,
    -- filter=92 channel=34
    0, -2, 5, 2, 0, 0, 0, 5, 1,
    -- filter=92 channel=35
    6, -2, 0, 0, 0, -6, -2, -3, 4,
    -- filter=92 channel=36
    5, -12, -12, -10, -11, -1, -2, -8, -14,
    -- filter=92 channel=37
    -8, -5, 2, 6, 7, 14, 10, 9, 6,
    -- filter=92 channel=38
    0, 2, -3, 7, 2, -3, -5, 1, -4,
    -- filter=92 channel=39
    -9, 0, -9, 4, -1, -6, -7, -10, -3,
    -- filter=92 channel=40
    0, -1, -3, -9, -4, 1, -8, 0, -6,
    -- filter=92 channel=41
    1, -17, -8, -9, -11, 2, -3, -15, 0,
    -- filter=92 channel=42
    -9, -1, -3, -4, -2, 0, -3, 2, 0,
    -- filter=92 channel=43
    -3, -13, -3, -4, -8, -1, -6, 7, -4,
    -- filter=92 channel=44
    2, -2, 4, 0, 6, 13, 0, 0, 5,
    -- filter=92 channel=45
    0, -1, 2, -4, 0, 1, 0, 3, 0,
    -- filter=92 channel=46
    -3, -2, -4, -5, -6, 0, -6, 2, -2,
    -- filter=92 channel=47
    -5, -4, -3, 8, 11, 4, 3, -2, 5,
    -- filter=92 channel=48
    -5, 0, 0, 1, 5, 11, 7, 0, 3,
    -- filter=92 channel=49
    -6, 0, 0, -5, 3, -4, -5, -3, 9,
    -- filter=92 channel=50
    -4, 6, 7, -2, 2, 5, -2, -3, 0,
    -- filter=92 channel=51
    -2, 0, -6, -3, 6, -3, -5, -5, 4,
    -- filter=92 channel=52
    2, 0, 0, -2, -1, -8, 1, -7, -6,
    -- filter=92 channel=53
    -5, 0, 2, -2, -4, -5, -2, -1, -3,
    -- filter=92 channel=54
    6, 5, -3, 2, 0, 2, 4, -3, 0,
    -- filter=92 channel=55
    -11, -16, -4, -11, -9, -8, -12, -9, -6,
    -- filter=92 channel=56
    5, -2, -4, -3, -5, 0, 7, 3, -5,
    -- filter=92 channel=57
    -4, -4, -2, -7, -8, 0, 6, 0, 6,
    -- filter=92 channel=58
    -8, 3, 0, 2, 3, 6, -4, 4, 3,
    -- filter=92 channel=59
    -5, 0, -2, 5, 5, -2, 5, 5, 0,
    -- filter=92 channel=60
    -3, -4, 1, 2, 2, 0, -2, 4, 3,
    -- filter=92 channel=61
    0, -8, -4, 0, 0, -7, -2, 1, -3,
    -- filter=92 channel=62
    4, -3, 0, -5, -6, -6, 5, 4, -6,
    -- filter=92 channel=63
    -7, 4, -5, 0, 0, -8, -1, -3, -6,
    -- filter=92 channel=64
    2, -10, -8, -8, -7, -8, -2, 2, -3,
    -- filter=92 channel=65
    0, -3, -5, 1, -2, 6, -6, -3, -4,
    -- filter=92 channel=66
    -3, -9, 0, 0, -11, -2, 1, -5, -1,
    -- filter=92 channel=67
    -4, -2, -4, 0, 5, -7, -1, 2, 0,
    -- filter=92 channel=68
    5, 5, -10, 0, -7, -9, -7, -5, 1,
    -- filter=92 channel=69
    0, -8, -1, 1, -4, -3, -3, -5, 6,
    -- filter=92 channel=70
    -13, -4, 2, 3, 3, 0, -1, 8, 10,
    -- filter=92 channel=71
    -2, -9, -5, -5, -10, -7, 0, 4, 4,
    -- filter=92 channel=72
    0, 0, 0, -1, 2, 2, -12, -2, -9,
    -- filter=92 channel=73
    -9, -5, 3, 0, -1, -2, -8, 0, 0,
    -- filter=92 channel=74
    0, 9, 10, 6, 8, 8, 0, 7, 8,
    -- filter=92 channel=75
    -14, -14, 3, 1, -2, 4, 0, 1, 6,
    -- filter=92 channel=76
    0, -7, -9, -1, -2, -8, -1, -2, 0,
    -- filter=92 channel=77
    -2, -4, 1, 1, -2, -6, 2, 3, -1,
    -- filter=92 channel=78
    0, -4, 4, 5, 7, -1, 2, -5, 1,
    -- filter=92 channel=79
    -6, -12, 1, -4, -5, 13, -9, -7, 9,
    -- filter=92 channel=80
    -2, -10, 5, 3, 9, 7, -2, -4, 3,
    -- filter=92 channel=81
    -5, -1, -2, -1, 6, -7, 0, 0, -1,
    -- filter=92 channel=82
    -1, -8, 5, -7, 1, 5, 5, -4, -3,
    -- filter=92 channel=83
    3, -4, 0, 5, 3, 0, 1, 7, 3,
    -- filter=92 channel=84
    -10, -7, 7, 6, 0, 2, 1, -8, 9,
    -- filter=92 channel=85
    5, 5, 5, -3, 6, -5, 5, 2, 7,
    -- filter=92 channel=86
    -5, -5, 8, -1, -2, 1, 5, 3, 3,
    -- filter=92 channel=87
    3, 1, -2, -9, -12, 1, 0, -6, -7,
    -- filter=92 channel=88
    1, 0, -12, 4, -6, -12, -10, -15, -10,
    -- filter=92 channel=89
    -12, -1, 2, 3, -8, 4, 2, 1, 1,
    -- filter=92 channel=90
    5, -6, -3, 3, -9, 0, -10, -8, -1,
    -- filter=92 channel=91
    -8, 0, 4, 0, 0, 0, 1, 0, 3,
    -- filter=92 channel=92
    -6, -4, -3, -4, -3, -8, 4, 3, -5,
    -- filter=92 channel=93
    4, 9, 2, 8, 16, 15, 6, 9, 5,
    -- filter=92 channel=94
    5, 5, 4, 7, 7, -3, 2, 6, 0,
    -- filter=92 channel=95
    -8, 3, -1, 0, -5, -1, -4, -2, 2,
    -- filter=92 channel=96
    -2, -6, 3, 0, 3, -6, -7, 1, -5,
    -- filter=92 channel=97
    -9, 1, -4, -3, 0, 2, 2, 0, -5,
    -- filter=92 channel=98
    0, -9, 8, 2, 5, 16, -5, 0, 17,
    -- filter=92 channel=99
    -5, -9, 4, 0, -1, 2, -7, -2, 3,
    -- filter=92 channel=100
    -6, -2, 0, -5, -9, -1, 1, -5, 0,
    -- filter=92 channel=101
    -3, -4, -9, 2, 4, 3, 1, 0, 0,
    -- filter=92 channel=102
    2, -3, -6, 3, 6, 0, -7, -2, -6,
    -- filter=92 channel=103
    -10, 0, -5, 2, 5, 0, 7, 3, 8,
    -- filter=92 channel=104
    6, -8, -3, 0, -1, -7, -1, -5, -4,
    -- filter=92 channel=105
    1, 1, 2, -4, -3, -8, 1, -10, -3,
    -- filter=92 channel=106
    -1, -8, -9, -9, -5, -4, 0, -9, -9,
    -- filter=92 channel=107
    -13, -2, 6, 0, 0, 6, 1, -2, 3,
    -- filter=92 channel=108
    -7, 0, -6, -2, 0, -8, -2, 4, -6,
    -- filter=92 channel=109
    -3, 2, 3, 7, 5, 14, 5, -4, 12,
    -- filter=92 channel=110
    -6, 2, 0, -8, 2, 0, 5, -1, 1,
    -- filter=92 channel=111
    0, 4, 0, -7, -7, 2, -2, 2, 3,
    -- filter=92 channel=112
    -2, 9, 0, 5, 5, 10, 0, 0, 12,
    -- filter=92 channel=113
    -9, -5, -8, -2, -5, 4, 0, 1, 0,
    -- filter=92 channel=114
    -14, -8, 7, 1, 0, 15, 3, -1, 4,
    -- filter=92 channel=115
    5, 0, -5, -4, 1, 1, 6, -1, -5,
    -- filter=92 channel=116
    -3, -5, -5, 1, -2, 0, -5, 0, -3,
    -- filter=92 channel=117
    -6, -3, -6, 3, -7, 2, -4, -1, -7,
    -- filter=92 channel=118
    -3, -3, 0, -6, -2, -3, -7, 0, 0,
    -- filter=92 channel=119
    -1, -2, 6, 1, -5, -5, 1, -2, -1,
    -- filter=92 channel=120
    -7, 5, 9, 9, 6, 6, -8, 7, 11,
    -- filter=92 channel=121
    2, -10, -6, -3, 2, -2, 1, -7, 7,
    -- filter=92 channel=122
    -2, -2, -10, -1, -2, -9, -1, -5, 2,
    -- filter=92 channel=123
    6, -2, 0, 2, -3, -6, 3, 2, -3,
    -- filter=92 channel=124
    4, -4, 0, 3, -9, -6, -9, -4, -2,
    -- filter=92 channel=125
    3, -8, 6, 5, 4, -1, -5, -12, 5,
    -- filter=92 channel=126
    -6, -18, 2, 2, -1, 2, 0, 1, 3,
    -- filter=92 channel=127
    0, 0, 3, 6, -3, 0, -6, -8, 6,
    -- filter=93 channel=0
    5, -6, 5, 9, -13, -8, 11, 8, 3,
    -- filter=93 channel=1
    10, 2, -3, 0, -2, -15, 6, -5, -10,
    -- filter=93 channel=2
    -7, 6, 6, -4, -1, -2, 0, -2, -10,
    -- filter=93 channel=3
    3, -13, 5, -12, -13, -2, -3, 3, 2,
    -- filter=93 channel=4
    0, -5, 11, -9, -15, -5, -2, -14, -1,
    -- filter=93 channel=5
    5, 4, 4, 1, -6, -3, 13, -3, -1,
    -- filter=93 channel=6
    -6, -2, -2, -8, -10, -2, -9, 0, 5,
    -- filter=93 channel=7
    0, 2, 6, 5, -2, -6, -1, 1, -7,
    -- filter=93 channel=8
    3, 0, 0, -4, -9, -10, 0, -4, -10,
    -- filter=93 channel=9
    -3, 9, 2, 4, 1, -2, -4, 1, 2,
    -- filter=93 channel=10
    8, 0, -5, 10, 14, -4, 0, 0, 2,
    -- filter=93 channel=11
    0, -8, -2, -1, -2, 13, -2, 4, 14,
    -- filter=93 channel=12
    6, -2, -6, -1, -11, -12, 0, -10, -5,
    -- filter=93 channel=13
    9, -1, -1, 1, -2, 2, -13, -6, -8,
    -- filter=93 channel=14
    5, 0, -6, 1, 2, 4, 0, 5, 4,
    -- filter=93 channel=15
    0, -15, -4, 1, -2, 9, -11, -5, 14,
    -- filter=93 channel=16
    -2, 3, -6, -2, 0, -5, -11, -11, -17,
    -- filter=93 channel=17
    0, 2, 2, 0, -7, -1, 1, -5, 3,
    -- filter=93 channel=18
    -1, -10, 0, -5, -2, -3, -3, -5, 16,
    -- filter=93 channel=19
    7, 1, 3, 7, 1, -6, -5, -4, -3,
    -- filter=93 channel=20
    -14, -8, 10, -13, -8, 0, -15, -2, 20,
    -- filter=93 channel=21
    6, 13, -8, 1, 16, 0, -1, -7, -9,
    -- filter=93 channel=22
    -3, -2, -5, 3, -7, -5, 7, -4, 0,
    -- filter=93 channel=23
    10, -5, -2, 2, -10, -1, -3, -5, 5,
    -- filter=93 channel=24
    -4, -4, 4, 2, 6, -6, 7, 0, -2,
    -- filter=93 channel=25
    8, 9, 1, 10, 15, 1, -8, -2, -11,
    -- filter=93 channel=26
    0, 7, 5, 2, 0, -2, -4, 0, 1,
    -- filter=93 channel=27
    16, -5, -7, 6, 11, -1, 5, -8, 3,
    -- filter=93 channel=28
    0, 6, -1, 7, 0, -7, 1, -7, -4,
    -- filter=93 channel=29
    -6, -6, 2, -16, -3, -1, -7, 3, 21,
    -- filter=93 channel=30
    9, 0, 6, -1, 7, 5, 8, 4, 6,
    -- filter=93 channel=31
    11, 10, -1, 11, 19, 5, -3, 0, 4,
    -- filter=93 channel=32
    9, 0, -2, -5, -6, 6, 0, -3, 10,
    -- filter=93 channel=33
    11, 0, -6, 6, 3, 5, 8, 0, -5,
    -- filter=93 channel=34
    0, -19, -5, 0, -16, -13, -5, -21, -12,
    -- filter=93 channel=35
    4, 5, 6, 6, -2, -5, 0, 3, 3,
    -- filter=93 channel=36
    1, 0, -4, -8, -2, -10, -12, -13, -6,
    -- filter=93 channel=37
    7, -4, -5, -1, -3, -10, 4, -1, -3,
    -- filter=93 channel=38
    5, 6, -7, 10, 7, 0, -6, 7, 3,
    -- filter=93 channel=39
    -8, -5, 11, -10, -7, 0, -10, -4, 9,
    -- filter=93 channel=40
    -12, -4, 1, -9, -8, -3, 2, -3, 2,
    -- filter=93 channel=41
    3, -3, 0, -1, -18, -22, -14, -14, -13,
    -- filter=93 channel=42
    8, 7, 5, 0, 6, 1, 1, 4, 4,
    -- filter=93 channel=43
    -5, -4, 3, 0, -4, -8, 2, 5, 0,
    -- filter=93 channel=44
    9, 7, -3, 0, -2, -4, 1, 3, -1,
    -- filter=93 channel=45
    -4, 1, -2, -4, -6, 1, -4, 0, -2,
    -- filter=93 channel=46
    2, 0, -2, 0, -7, 2, 0, -10, 0,
    -- filter=93 channel=47
    0, 8, -1, 6, 3, -9, -6, 7, -5,
    -- filter=93 channel=48
    17, 8, -1, 10, 17, 0, 3, -10, -5,
    -- filter=93 channel=49
    7, 0, 0, 1, 6, 3, 0, -1, 10,
    -- filter=93 channel=50
    12, 2, -7, 2, 11, -5, 5, 10, 9,
    -- filter=93 channel=51
    6, -3, 2, 2, 1, -7, -4, -3, -5,
    -- filter=93 channel=52
    1, -4, -4, -3, -8, -8, 4, -12, -3,
    -- filter=93 channel=53
    -6, -3, 2, -4, 0, 2, 0, 7, 11,
    -- filter=93 channel=54
    -6, -3, -1, -6, 3, 6, 7, -6, -3,
    -- filter=93 channel=55
    -3, -4, -6, -8, -5, 1, -6, 2, 5,
    -- filter=93 channel=56
    2, 1, 1, -1, -1, -1, 0, -3, -9,
    -- filter=93 channel=57
    -7, 5, -1, -3, -10, -1, 0, -6, -4,
    -- filter=93 channel=58
    -5, -2, 5, 1, -6, 1, 4, 3, 5,
    -- filter=93 channel=59
    10, 11, -6, 9, 15, -2, -6, 0, -1,
    -- filter=93 channel=60
    6, 7, -5, 1, 5, 1, 3, 1, 4,
    -- filter=93 channel=61
    -2, -5, -4, -1, -6, 0, -6, -4, -7,
    -- filter=93 channel=62
    5, -6, -7, 1, -4, 3, 3, -1, -1,
    -- filter=93 channel=63
    1, 2, 9, -4, -5, -3, -3, 2, -4,
    -- filter=93 channel=64
    -1, -8, 0, -1, -9, -5, -4, 2, 6,
    -- filter=93 channel=65
    0, 7, 7, 5, 4, -5, -4, -1, -1,
    -- filter=93 channel=66
    -6, -10, -6, -10, -13, -2, -11, -2, -1,
    -- filter=93 channel=67
    0, -5, 5, 0, -6, 1, -1, -5, 5,
    -- filter=93 channel=68
    3, -1, 5, 1, -2, -6, -6, -1, -8,
    -- filter=93 channel=69
    -5, -6, 6, 3, 1, -2, -2, 5, 0,
    -- filter=93 channel=70
    6, -4, -6, 7, -3, -4, 1, -5, 3,
    -- filter=93 channel=71
    7, 0, -5, 2, -3, -6, -6, -3, -10,
    -- filter=93 channel=72
    11, 1, -9, 4, 19, -1, -8, -3, 0,
    -- filter=93 channel=73
    0, -2, -3, 2, 3, 2, -4, -7, 0,
    -- filter=93 channel=74
    2, -7, 0, 10, -10, -9, 10, -3, 4,
    -- filter=93 channel=75
    5, -1, -7, 7, -12, -11, 7, 0, 0,
    -- filter=93 channel=76
    -3, -8, 2, -14, -5, 5, -17, -5, 11,
    -- filter=93 channel=77
    1, 1, 0, -4, -4, 0, -5, 1, -6,
    -- filter=93 channel=78
    4, -3, 5, 3, 0, 2, 1, -4, 8,
    -- filter=93 channel=79
    8, -9, -10, 4, -5, 1, -1, 5, 10,
    -- filter=93 channel=80
    19, 20, 0, 7, 30, 9, -2, 1, -8,
    -- filter=93 channel=81
    -4, -4, 0, 3, 6, -5, -3, 0, 0,
    -- filter=93 channel=82
    -5, 5, 6, -2, -3, -2, 7, 1, 2,
    -- filter=93 channel=83
    4, 14, 4, 4, 13, 8, 1, 2, 6,
    -- filter=93 channel=84
    2, -9, -2, -8, -1, -2, -12, 0, -1,
    -- filter=93 channel=85
    0, 5, 1, -2, 3, 6, -6, 6, 5,
    -- filter=93 channel=86
    -6, -5, -2, -1, -9, -3, 4, -6, 1,
    -- filter=93 channel=87
    0, -18, 2, -3, -9, 4, -8, -5, 4,
    -- filter=93 channel=88
    -9, 1, 3, -4, -1, -2, -4, -13, -1,
    -- filter=93 channel=89
    17, -2, -5, 6, 15, 8, -11, -3, -2,
    -- filter=93 channel=90
    -3, -8, -7, -2, -8, -5, -5, -13, -9,
    -- filter=93 channel=91
    11, -9, 6, -4, 9, 2, 0, -3, -2,
    -- filter=93 channel=92
    -9, 1, 5, -4, -15, -1, -9, -7, -7,
    -- filter=93 channel=93
    2, 3, -1, 7, 1, -1, -6, -1, -2,
    -- filter=93 channel=94
    -2, -6, 3, -4, -2, 2, -4, -7, 0,
    -- filter=93 channel=95
    3, -7, 7, 1, 5, -2, 3, 5, -7,
    -- filter=93 channel=96
    8, 6, 5, 7, -3, 6, -1, 0, 5,
    -- filter=93 channel=97
    -4, 3, -6, 7, -3, 0, -4, 7, -2,
    -- filter=93 channel=98
    15, 12, 3, 10, 17, 5, -2, 9, 3,
    -- filter=93 channel=99
    7, 0, 5, 9, 9, 2, 0, 2, 0,
    -- filter=93 channel=100
    -6, -6, 0, -4, -4, -9, -8, 1, 2,
    -- filter=93 channel=101
    -8, -1, 8, -16, -7, 0, 2, -5, -2,
    -- filter=93 channel=102
    4, -2, 4, 6, -5, -2, -1, 2, -6,
    -- filter=93 channel=103
    2, 13, -8, 0, 16, -1, -1, 0, -16,
    -- filter=93 channel=104
    15, 9, -7, 13, 26, -3, -4, 0, 0,
    -- filter=93 channel=105
    -6, -6, -8, -1, -11, -2, 0, 4, 5,
    -- filter=93 channel=106
    -8, 3, 0, -8, 0, -8, -9, 4, 2,
    -- filter=93 channel=107
    0, -12, 1, 0, -13, 9, -8, -3, 19,
    -- filter=93 channel=108
    4, 4, -5, -2, 0, 0, -5, -6, 0,
    -- filter=93 channel=109
    13, 2, 1, 11, 11, -3, -2, -6, -7,
    -- filter=93 channel=110
    5, -5, 4, 2, 9, 2, 1, -3, -6,
    -- filter=93 channel=111
    7, 2, 4, -5, -3, -5, 4, -6, -4,
    -- filter=93 channel=112
    5, 4, -2, 12, 2, -1, 5, 6, -6,
    -- filter=93 channel=113
    11, 5, -2, 11, 0, -6, 7, 5, 2,
    -- filter=93 channel=114
    1, -10, 10, -5, -1, -4, 4, 2, 12,
    -- filter=93 channel=115
    7, 5, -3, -3, 0, 1, 7, -5, 5,
    -- filter=93 channel=116
    11, 9, -5, -2, 17, 4, -7, 1, 4,
    -- filter=93 channel=117
    0, 0, -2, 4, -3, 2, 2, -2, 4,
    -- filter=93 channel=118
    7, 4, 4, -1, 6, -4, 1, 3, -6,
    -- filter=93 channel=119
    -10, -12, 0, -3, -19, -13, -2, -9, -2,
    -- filter=93 channel=120
    5, -9, 9, 8, 0, 9, 5, 5, 10,
    -- filter=93 channel=121
    6, 4, -4, 1, -2, 2, -2, -9, -11,
    -- filter=93 channel=122
    -2, 4, -11, 1, 1, -18, -7, -12, -26,
    -- filter=93 channel=123
    -8, -2, -2, 2, -8, -12, 2, -6, -8,
    -- filter=93 channel=124
    -8, 0, -7, -9, 1, -3, -10, 5, 10,
    -- filter=93 channel=125
    13, -2, 5, 5, 13, -3, 3, -1, -2,
    -- filter=93 channel=126
    12, -5, -4, 7, 7, -3, -7, 0, 3,
    -- filter=93 channel=127
    0, 0, 6, 4, -4, -8, -8, -7, 0,
    -- filter=94 channel=0
    -4, 3, -7, 21, 27, -11, 7, 9, -3,
    -- filter=94 channel=1
    -6, 0, -7, 23, 24, -6, 7, 9, -10,
    -- filter=94 channel=2
    5, -6, 5, -5, -2, 0, -4, 0, -3,
    -- filter=94 channel=3
    -4, 7, -4, 0, -2, 9, 4, 4, 9,
    -- filter=94 channel=4
    -3, 6, 5, -4, 7, 12, -12, 4, -2,
    -- filter=94 channel=5
    0, -9, -18, 15, 13, -10, 6, 4, -5,
    -- filter=94 channel=6
    0, -1, 1, 0, 1, 1, -7, -10, 6,
    -- filter=94 channel=7
    -1, 1, -4, 7, -5, -5, -7, -4, 1,
    -- filter=94 channel=8
    -4, -8, 5, -5, 0, 8, -8, 2, 1,
    -- filter=94 channel=9
    4, -2, -1, 4, 3, -1, -2, -1, -8,
    -- filter=94 channel=10
    -5, -6, 2, -9, -8, -1, -9, -1, 11,
    -- filter=94 channel=11
    1, -4, 12, -11, -13, 3, -12, -3, -1,
    -- filter=94 channel=12
    5, -6, -3, 2, -2, 6, 0, -8, 1,
    -- filter=94 channel=13
    -3, 2, 1, 1, 0, 3, -10, -4, 9,
    -- filter=94 channel=14
    6, 2, 7, -4, 5, -7, 0, 0, -3,
    -- filter=94 channel=15
    -4, -5, 5, -2, -6, 0, -1, -9, 1,
    -- filter=94 channel=16
    -1, -6, -8, 6, 2, 0, -3, 1, 1,
    -- filter=94 channel=17
    0, 7, -6, -5, -5, 0, 2, -1, -2,
    -- filter=94 channel=18
    -5, -3, 5, 14, 1, 6, -3, -5, -1,
    -- filter=94 channel=19
    5, -3, 7, -5, -1, 3, 3, -6, 7,
    -- filter=94 channel=20
    -5, -2, 16, -7, -18, 10, -10, -3, 9,
    -- filter=94 channel=21
    0, 4, 5, -6, 2, -3, -2, 6, 1,
    -- filter=94 channel=22
    6, -6, 0, 2, 7, 0, 11, -7, 3,
    -- filter=94 channel=23
    -2, -8, 0, -7, -10, 1, -7, -5, 13,
    -- filter=94 channel=24
    -5, -7, -1, -4, -2, 6, -7, 1, -2,
    -- filter=94 channel=25
    6, 4, -1, 10, 3, -3, 2, -1, -5,
    -- filter=94 channel=26
    -3, -6, -4, 4, -6, 0, 1, 6, -2,
    -- filter=94 channel=27
    3, 0, 2, 12, -5, -7, 7, 7, -5,
    -- filter=94 channel=28
    -7, 2, 1, 1, 6, -7, 0, 4, -2,
    -- filter=94 channel=29
    -7, 3, 1, -7, -12, 3, -14, -12, 6,
    -- filter=94 channel=30
    -6, 3, -7, 12, 1, 2, 4, 2, -4,
    -- filter=94 channel=31
    -10, 3, 13, -19, -5, -1, -1, 3, 5,
    -- filter=94 channel=32
    5, 1, 1, 2, -10, -5, -2, -3, 2,
    -- filter=94 channel=33
    0, -4, 2, 1, -4, -9, 9, 7, 5,
    -- filter=94 channel=34
    5, -8, 3, 6, -4, -2, 3, -1, 8,
    -- filter=94 channel=35
    -5, -4, -3, 6, -3, 0, 4, 0, 3,
    -- filter=94 channel=36
    -8, -7, 8, -12, -13, 5, -12, -3, 11,
    -- filter=94 channel=37
    2, -2, -16, 18, 30, -5, 8, 15, -3,
    -- filter=94 channel=38
    4, 1, 2, 5, -7, -9, -3, 1, 3,
    -- filter=94 channel=39
    1, -6, 6, -1, -1, 4, 0, 2, 9,
    -- filter=94 channel=40
    1, 8, 10, -5, 0, 3, 8, 0, 6,
    -- filter=94 channel=41
    7, -12, 2, -1, -10, -2, -7, -9, -5,
    -- filter=94 channel=42
    -8, 6, -6, 3, 8, 2, 0, 4, 3,
    -- filter=94 channel=43
    4, 0, -3, -8, 6, 1, -3, -1, 9,
    -- filter=94 channel=44
    9, 0, -5, 6, 5, -4, 0, 11, -7,
    -- filter=94 channel=45
    4, 0, 0, 8, 0, 0, 1, 4, 6,
    -- filter=94 channel=46
    7, -3, -6, 0, 6, 3, 5, -1, -2,
    -- filter=94 channel=47
    -5, 1, -3, 2, -2, 0, 4, 0, 4,
    -- filter=94 channel=48
    -2, 6, -6, 2, 0, -9, 0, 7, 1,
    -- filter=94 channel=49
    7, -1, 5, 0, 1, -2, 1, 0, -5,
    -- filter=94 channel=50
    3, 6, 6, -2, 4, 0, 2, -1, -2,
    -- filter=94 channel=51
    -6, -5, 3, 7, -2, 2, 2, 5, 0,
    -- filter=94 channel=52
    3, 0, 0, -7, 0, 9, -3, -3, 0,
    -- filter=94 channel=53
    -2, 0, 3, -12, -3, 8, -9, 2, -1,
    -- filter=94 channel=54
    6, 3, 4, 4, 1, 6, -2, -2, 6,
    -- filter=94 channel=55
    -11, -6, 13, -15, -24, 4, -12, -15, 2,
    -- filter=94 channel=56
    -2, -7, 6, -6, 0, -1, 0, -2, -4,
    -- filter=94 channel=57
    -5, -3, -4, 6, -5, 0, -1, 0, 0,
    -- filter=94 channel=58
    -1, -4, -3, -2, 2, -10, -3, -3, -4,
    -- filter=94 channel=59
    -1, -6, -6, 0, -9, -3, 1, 4, 0,
    -- filter=94 channel=60
    -1, -1, 2, -4, 2, 4, -6, -7, 6,
    -- filter=94 channel=61
    -5, -3, 1, -2, 0, 5, 0, 5, 2,
    -- filter=94 channel=62
    6, -5, 7, -4, 1, -3, 3, -6, -2,
    -- filter=94 channel=63
    0, -2, -3, 2, 2, 0, -9, -2, 1,
    -- filter=94 channel=64
    -5, -4, 7, -3, -6, 0, -4, 3, 4,
    -- filter=94 channel=65
    6, 1, 2, 4, 3, -4, -1, 7, -3,
    -- filter=94 channel=66
    0, 2, 0, 0, -6, 2, -3, -8, -1,
    -- filter=94 channel=67
    4, 0, -6, -6, 5, 7, -2, 5, 4,
    -- filter=94 channel=68
    -7, 4, -2, 1, 1, 6, -5, -3, 3,
    -- filter=94 channel=69
    -4, 0, 4, 1, 2, -4, 3, 2, -3,
    -- filter=94 channel=70
    4, 12, 0, 6, -2, -2, -2, 8, 1,
    -- filter=94 channel=71
    0, 2, -4, 1, 6, 4, 5, -2, 4,
    -- filter=94 channel=72
    -10, -8, 0, -5, -10, 1, -3, -5, 10,
    -- filter=94 channel=73
    4, -1, 1, -7, 0, -2, -2, -8, 6,
    -- filter=94 channel=74
    0, 2, 0, 3, 0, -5, 4, -2, 8,
    -- filter=94 channel=75
    -1, 6, -8, 8, 14, 0, 14, 14, -2,
    -- filter=94 channel=76
    0, -5, 7, -6, -13, 12, -8, -5, 2,
    -- filter=94 channel=77
    -3, -4, -1, -4, -3, 7, -2, -5, -6,
    -- filter=94 channel=78
    -3, -2, -9, -6, -4, 0, -7, 5, -2,
    -- filter=94 channel=79
    -3, 0, 11, 13, 6, -3, 9, -7, 9,
    -- filter=94 channel=80
    -9, 4, 7, -4, -6, 4, -9, 0, 7,
    -- filter=94 channel=81
    -2, 0, 4, 2, -3, 5, 7, 0, 0,
    -- filter=94 channel=82
    7, -1, -6, 2, -3, 2, 7, 1, 1,
    -- filter=94 channel=83
    2, 0, 0, 6, -3, 4, 0, 8, 0,
    -- filter=94 channel=84
    3, 8, 9, 9, 2, 8, 1, -2, 0,
    -- filter=94 channel=85
    -2, -1, -1, 0, 2, 5, -5, -3, -1,
    -- filter=94 channel=86
    -2, -4, 6, -5, 7, 0, 1, 5, 0,
    -- filter=94 channel=87
    -3, -5, 7, -2, -3, 11, -2, 1, 0,
    -- filter=94 channel=88
    -2, 4, 14, -1, -11, 8, -2, -5, 12,
    -- filter=94 channel=89
    -5, 1, 11, -9, -3, 2, -3, -3, 0,
    -- filter=94 channel=90
    4, -8, 2, -11, -14, 3, 2, -5, 0,
    -- filter=94 channel=91
    -2, 9, 3, -3, -8, 0, 2, -7, 8,
    -- filter=94 channel=92
    -7, -3, -6, 1, 4, -6, -5, -1, 0,
    -- filter=94 channel=93
    -3, -4, -7, 4, 14, -11, 5, 14, -6,
    -- filter=94 channel=94
    1, -4, -7, -4, 3, 4, -5, -2, 0,
    -- filter=94 channel=95
    0, -7, 0, -3, -2, 1, 1, -4, 5,
    -- filter=94 channel=96
    4, -4, -7, 4, 4, -4, -1, 2, 4,
    -- filter=94 channel=97
    -8, -1, 0, -4, 5, -4, -5, 7, -2,
    -- filter=94 channel=98
    -7, -8, -6, -2, -6, -3, -3, 5, -2,
    -- filter=94 channel=99
    -7, -2, 6, -14, -17, 9, -11, -5, 3,
    -- filter=94 channel=100
    4, 2, 4, 2, 0, 4, -2, 0, -8,
    -- filter=94 channel=101
    6, -3, 9, -6, 1, 10, -8, -1, 6,
    -- filter=94 channel=102
    -3, 1, 2, 0, -1, 6, 0, 6, -5,
    -- filter=94 channel=103
    -4, -5, -3, 8, 3, -5, 8, 3, -3,
    -- filter=94 channel=104
    -5, -8, -3, -9, -5, 5, 3, 4, 1,
    -- filter=94 channel=105
    0, -5, 8, -8, -7, 8, -4, -9, 0,
    -- filter=94 channel=106
    -1, -5, 8, -6, -9, -4, -2, -6, 5,
    -- filter=94 channel=107
    -1, 3, -2, 0, 2, 8, 0, -5, 9,
    -- filter=94 channel=108
    -5, -10, -1, -5, 6, -7, -4, -9, -5,
    -- filter=94 channel=109
    6, 1, 1, 2, 0, -2, -4, 0, -3,
    -- filter=94 channel=110
    -9, 0, -2, -12, -13, 3, -4, -6, 13,
    -- filter=94 channel=111
    5, -3, -5, 6, -8, 2, 4, -2, 0,
    -- filter=94 channel=112
    5, 1, -4, 11, 0, 1, 5, 6, -1,
    -- filter=94 channel=113
    -7, -2, 2, -8, -7, 0, -4, 0, 7,
    -- filter=94 channel=114
    -3, 9, -7, 23, 3, -9, 10, 6, -6,
    -- filter=94 channel=115
    -1, 4, -2, 5, -2, 2, -5, 2, 5,
    -- filter=94 channel=116
    -3, -2, 3, 1, -13, -6, -9, -5, -3,
    -- filter=94 channel=117
    2, 6, -2, 0, -4, 7, -3, 3, 9,
    -- filter=94 channel=118
    6, -1, -5, 5, -4, -2, -4, 5, 2,
    -- filter=94 channel=119
    -2, -6, 5, 0, -3, 3, -8, -3, 6,
    -- filter=94 channel=120
    4, -3, 0, 0, -14, 6, -2, 0, 7,
    -- filter=94 channel=121
    2, -11, 6, -5, -7, 6, 0, 3, -1,
    -- filter=94 channel=122
    0, -9, -1, -4, 8, -12, 2, 9, -8,
    -- filter=94 channel=123
    4, -5, 6, 6, 1, 3, -4, 1, -6,
    -- filter=94 channel=124
    -5, 3, 3, -2, -4, 9, 5, 2, 2,
    -- filter=94 channel=125
    -2, -4, 2, -6, -7, -5, -11, 0, -2,
    -- filter=94 channel=126
    4, -6, -4, 6, -4, -6, -2, -4, 0,
    -- filter=94 channel=127
    0, -9, 3, -3, -1, -3, -4, 3, 2,
    -- filter=95 channel=0
    -11, -2, -5, 10, 14, 9, 2, -6, -5,
    -- filter=95 channel=1
    -9, -10, 6, -1, 0, 0, 11, 4, 9,
    -- filter=95 channel=2
    -1, 13, -5, -2, -4, -1, 1, 14, 15,
    -- filter=95 channel=3
    -14, -18, -16, 11, 40, 28, 5, 0, -2,
    -- filter=95 channel=4
    0, 19, 2, -6, -14, 4, 19, 40, 35,
    -- filter=95 channel=5
    -7, -14, -4, 0, 6, 9, -2, 1, -1,
    -- filter=95 channel=6
    -7, 2, -7, -1, -6, -3, 7, 4, -6,
    -- filter=95 channel=7
    2, -4, 5, -6, -6, 0, 5, 5, -3,
    -- filter=95 channel=8
    3, 8, -3, -3, -2, 2, 1, 8, 2,
    -- filter=95 channel=9
    0, 6, 6, -5, 1, 0, -1, 12, 5,
    -- filter=95 channel=10
    -8, -4, -1, 8, 11, 6, -12, -3, -5,
    -- filter=95 channel=11
    -1, 10, -3, 3, -1, -3, 0, 7, 0,
    -- filter=95 channel=12
    -2, -6, 2, -1, -1, -8, -10, -12, -5,
    -- filter=95 channel=13
    1, -3, 4, 0, 0, -17, -4, 4, 0,
    -- filter=95 channel=14
    6, 0, 1, -6, -3, -1, -1, 1, -5,
    -- filter=95 channel=15
    7, -6, -4, 0, 11, -2, -9, -5, -8,
    -- filter=95 channel=16
    -3, -6, 3, -2, -4, -7, -2, 6, -2,
    -- filter=95 channel=17
    5, 2, -2, -2, 2, -2, 6, 0, 2,
    -- filter=95 channel=18
    0, 3, 0, 4, -7, -10, 1, -7, 4,
    -- filter=95 channel=19
    -3, -1, 2, -5, -6, 0, -7, -3, -4,
    -- filter=95 channel=20
    -1, 7, 2, 0, -6, -7, 2, 7, 7,
    -- filter=95 channel=21
    2, 1, 5, -6, -10, -4, 4, 6, 2,
    -- filter=95 channel=22
    -2, 1, -5, -3, 9, 0, 3, -3, -9,
    -- filter=95 channel=23
    -9, -8, -6, 11, 7, 3, -2, 3, -11,
    -- filter=95 channel=24
    -1, 2, 0, 6, 6, 0, -4, 1, 7,
    -- filter=95 channel=25
    -2, 4, 10, -6, -24, -16, 4, 16, 22,
    -- filter=95 channel=26
    -3, 7, -3, 2, 1, -4, -1, 6, 9,
    -- filter=95 channel=27
    0, 5, 13, -8, -35, -34, -1, 12, 14,
    -- filter=95 channel=28
    0, -2, -2, 7, 0, -5, 5, 0, 2,
    -- filter=95 channel=29
    0, 0, -4, -1, -5, 2, 5, 5, -1,
    -- filter=95 channel=30
    0, 0, 0, -9, -22, -19, 0, 26, 22,
    -- filter=95 channel=31
    -3, 5, 9, -6, -11, -8, 2, 2, -5,
    -- filter=95 channel=32
    -2, 4, 10, 2, -12, -14, 6, 14, 0,
    -- filter=95 channel=33
    -2, -6, -8, 15, 13, 4, -11, -10, -7,
    -- filter=95 channel=34
    4, 7, 1, -5, -16, -14, -5, -11, -3,
    -- filter=95 channel=35
    4, 2, 4, -3, 7, -4, 3, 2, -1,
    -- filter=95 channel=36
    6, 11, 0, -7, -7, -4, -5, 10, 7,
    -- filter=95 channel=37
    -9, 0, 0, 0, -12, 0, -1, 11, 6,
    -- filter=95 channel=38
    2, -3, -5, 4, 10, -4, -4, -3, 0,
    -- filter=95 channel=39
    3, 0, 3, -4, -8, -9, -2, 10, 4,
    -- filter=95 channel=40
    -7, -4, 3, -1, -1, 7, -6, -2, -11,
    -- filter=95 channel=41
    12, -4, 1, -3, 4, -11, -2, -12, -6,
    -- filter=95 channel=42
    -8, 2, -5, 3, -6, 1, 8, 11, 9,
    -- filter=95 channel=43
    -1, -10, -6, 15, 27, 12, 0, -6, 0,
    -- filter=95 channel=44
    0, -1, 9, -2, -15, -8, 1, 6, 8,
    -- filter=95 channel=45
    -8, 5, 0, -5, -4, -3, 8, 2, 2,
    -- filter=95 channel=46
    4, 6, -3, -1, -4, 1, -7, 1, 1,
    -- filter=95 channel=47
    -12, -5, 2, 8, 3, -6, -2, 8, 6,
    -- filter=95 channel=48
    1, 20, 15, -16, -27, -31, 11, 25, 32,
    -- filter=95 channel=49
    -5, 13, -4, -8, -23, -7, 6, 22, 10,
    -- filter=95 channel=50
    -5, -6, -2, 1, -5, -7, -3, 11, 0,
    -- filter=95 channel=51
    -4, 4, -5, 2, 4, 5, 2, 5, -3,
    -- filter=95 channel=52
    -1, 0, 2, -5, -12, 5, 0, 2, -8,
    -- filter=95 channel=53
    7, -2, -2, 1, -7, 5, -4, -1, 6,
    -- filter=95 channel=54
    4, 4, 2, -5, -4, 0, -3, -5, 3,
    -- filter=95 channel=55
    1, 0, 4, 5, 3, -11, -1, -2, -1,
    -- filter=95 channel=56
    9, 1, -6, -4, -3, 3, 3, 6, -2,
    -- filter=95 channel=57
    0, -1, 2, 0, -4, -2, 5, 2, 9,
    -- filter=95 channel=58
    -7, -1, -5, -3, 7, 13, -5, 9, -2,
    -- filter=95 channel=59
    8, 2, 11, -7, -3, -23, -2, 8, 0,
    -- filter=95 channel=60
    1, -2, -1, -7, -7, 4, 6, 5, 4,
    -- filter=95 channel=61
    0, 4, 6, 1, 1, 3, 0, 7, 2,
    -- filter=95 channel=62
    -6, 2, -4, 5, 9, 4, 2, 5, 5,
    -- filter=95 channel=63
    -8, -3, -6, 4, -2, 8, 4, 3, 1,
    -- filter=95 channel=64
    3, 9, 6, -4, -2, 5, -6, 3, 5,
    -- filter=95 channel=65
    6, -3, 6, -2, -2, 0, -4, -6, 1,
    -- filter=95 channel=66
    -2, 3, 4, -6, -6, -9, -6, -15, 0,
    -- filter=95 channel=67
    -6, -5, -3, 1, 4, -4, -3, -2, 4,
    -- filter=95 channel=68
    0, -3, 4, 0, 0, -1, -5, 12, 10,
    -- filter=95 channel=69
    -1, -1, -7, 0, 2, -5, 3, -4, 1,
    -- filter=95 channel=70
    1, 3, -1, 3, -4, -12, -2, -3, -4,
    -- filter=95 channel=71
    -2, -3, -6, 8, 11, 10, -8, -11, -11,
    -- filter=95 channel=72
    0, 14, 7, 2, -6, -15, -8, 0, 5,
    -- filter=95 channel=73
    -5, 16, 11, -4, -8, -22, -6, 10, 4,
    -- filter=95 channel=74
    4, 8, 6, -2, -21, -20, -1, 8, -7,
    -- filter=95 channel=75
    -7, -16, -6, 15, 22, 20, -1, -9, 1,
    -- filter=95 channel=76
    0, -2, 5, 0, 8, -5, -8, -2, -5,
    -- filter=95 channel=77
    0, -2, -1, -2, -3, 5, -1, -5, 0,
    -- filter=95 channel=78
    3, -6, 0, 5, 6, -2, 1, -6, 5,
    -- filter=95 channel=79
    -3, -2, 4, 11, 3, -16, 2, 1, 4,
    -- filter=95 channel=80
    2, 3, 6, 0, -13, -16, -3, 6, 15,
    -- filter=95 channel=81
    -2, -5, 0, 5, 7, 1, -7, 3, 5,
    -- filter=95 channel=82
    -1, -1, -1, 6, 0, 13, -5, -5, -6,
    -- filter=95 channel=83
    9, 4, -2, -8, -17, -7, 7, 8, 0,
    -- filter=95 channel=84
    9, 16, 9, -13, -14, -22, 0, 16, 13,
    -- filter=95 channel=85
    3, -5, -3, 7, 7, 0, -2, 6, -4,
    -- filter=95 channel=86
    0, 4, -7, 0, -7, 0, -1, 2, 0,
    -- filter=95 channel=87
    -1, 9, 0, -5, -12, 1, 6, -3, 0,
    -- filter=95 channel=88
    5, 1, 2, 0, -18, -2, -1, 11, 4,
    -- filter=95 channel=89
    -4, 0, 7, 10, 5, -2, 2, -8, 1,
    -- filter=95 channel=90
    9, 2, 6, -3, 5, -1, -6, -12, -2,
    -- filter=95 channel=91
    4, 11, -1, -10, -25, -23, 11, 28, 26,
    -- filter=95 channel=92
    -2, -3, -1, 2, 2, 0, 6, -9, -6,
    -- filter=95 channel=93
    -5, 12, 6, -4, -22, -6, 10, 30, 17,
    -- filter=95 channel=94
    2, -1, -6, -4, 3, -3, 6, 4, 0,
    -- filter=95 channel=95
    -1, 0, -7, 6, 6, 4, 4, -8, -1,
    -- filter=95 channel=96
    5, -2, -5, -1, -2, 1, 3, 2, 3,
    -- filter=95 channel=97
    -2, -13, -5, 11, 25, 28, -10, -6, -1,
    -- filter=95 channel=98
    0, -5, 15, 10, 5, -19, 1, 3, 13,
    -- filter=95 channel=99
    2, 23, 8, 4, -10, -19, -2, 13, 0,
    -- filter=95 channel=100
    3, -4, -5, -5, -6, -9, 2, -1, 3,
    -- filter=95 channel=101
    1, 17, 1, -1, -8, -5, 13, 17, 23,
    -- filter=95 channel=102
    2, -5, 3, -1, 0, -6, -4, 3, 4,
    -- filter=95 channel=103
    -17, -13, 7, 1, 12, 15, -9, -8, -6,
    -- filter=95 channel=104
    4, 12, 8, -9, -5, -13, -6, 7, 4,
    -- filter=95 channel=105
    2, 4, 1, 10, 5, -2, -6, 4, -2,
    -- filter=95 channel=106
    -6, -1, -3, 5, 7, -3, 2, -4, 2,
    -- filter=95 channel=107
    -7, -6, 0, 0, -1, -1, -3, 7, -5,
    -- filter=95 channel=108
    1, 2, -3, 0, 12, -2, 5, 0, 4,
    -- filter=95 channel=109
    10, 18, 18, -3, -36, -37, -3, 9, 10,
    -- filter=95 channel=110
    -5, -5, -1, 1, 8, 0, -7, -3, 3,
    -- filter=95 channel=111
    8, 5, -7, -7, -4, 0, 0, 3, -6,
    -- filter=95 channel=112
    4, 3, 3, -9, -10, -5, -2, 7, 0,
    -- filter=95 channel=113
    -10, -16, -12, 4, 20, 8, 1, -6, -11,
    -- filter=95 channel=114
    -8, 10, 8, 8, -19, -25, 1, 21, 25,
    -- filter=95 channel=115
    -7, 7, 5, 2, -2, -2, 2, 4, -3,
    -- filter=95 channel=116
    -5, 14, 6, -15, -31, -32, 6, 14, 26,
    -- filter=95 channel=117
    1, 5, 0, -7, -5, -10, 4, 11, 6,
    -- filter=95 channel=118
    -5, 4, 2, -1, 6, 5, 2, -1, -6,
    -- filter=95 channel=119
    11, 3, 7, -8, -10, -16, 0, -7, -5,
    -- filter=95 channel=120
    -1, 25, 1, -13, -40, -25, -4, 18, 13,
    -- filter=95 channel=121
    -6, -1, 1, 6, 7, 5, -10, -8, -5,
    -- filter=95 channel=122
    -11, -1, 12, -11, 0, -11, -1, 6, 0,
    -- filter=95 channel=123
    1, -5, -6, 0, 6, 0, 6, -12, -10,
    -- filter=95 channel=124
    -1, 6, -5, -3, 5, -1, 0, -4, 5,
    -- filter=95 channel=125
    3, 22, 8, -14, -27, -31, -10, 5, 16,
    -- filter=95 channel=126
    -10, -10, -4, 16, 14, 0, -1, -5, -5,
    -- filter=95 channel=127
    8, 1, -1, -3, 1, -1, -4, 5, -5,
    -- filter=96 channel=0
    -2, 3, 3, -4, 18, -6, 0, 1, -10,
    -- filter=96 channel=1
    -8, -5, -7, 4, 16, -5, 8, 12, -5,
    -- filter=96 channel=2
    0, -2, -8, -2, -9, -2, -6, -3, 0,
    -- filter=96 channel=3
    -2, 3, -3, 3, -1, 9, 3, 0, 3,
    -- filter=96 channel=4
    -7, -1, -4, -7, -4, 2, -1, 9, 5,
    -- filter=96 channel=5
    -5, 6, 3, -1, 19, -7, -1, 7, -15,
    -- filter=96 channel=6
    -4, -4, -6, 6, -3, 3, 2, 6, 1,
    -- filter=96 channel=7
    5, 3, 5, 0, 7, 5, 5, -1, 2,
    -- filter=96 channel=8
    -3, -5, 2, -7, 7, 7, -1, 0, 10,
    -- filter=96 channel=9
    -4, -2, 3, -6, 7, 0, 3, 3, 3,
    -- filter=96 channel=10
    0, 4, 4, -2, -3, 5, 3, -8, 5,
    -- filter=96 channel=11
    -5, 3, -1, 2, 2, 6, -1, -6, -2,
    -- filter=96 channel=12
    -5, 3, -4, 6, -1, -5, -5, 7, 8,
    -- filter=96 channel=13
    1, 4, 5, 4, 0, 2, 0, -6, 3,
    -- filter=96 channel=14
    0, 4, 1, 1, 1, 0, 0, 1, 1,
    -- filter=96 channel=15
    2, 7, 5, -6, -11, 2, -4, -12, 12,
    -- filter=96 channel=16
    2, 6, 2, -2, 11, 1, 3, 10, -8,
    -- filter=96 channel=17
    -5, 0, 6, -2, -3, 3, -5, 2, 0,
    -- filter=96 channel=18
    7, 1, -4, -4, 0, -2, -5, -10, 0,
    -- filter=96 channel=19
    -4, 0, 2, 4, -6, 2, 1, -3, -5,
    -- filter=96 channel=20
    -3, 7, -4, -7, -7, 6, -2, -11, 9,
    -- filter=96 channel=21
    -2, 1, -6, 7, 6, -7, 8, -5, -13,
    -- filter=96 channel=22
    -5, 2, 1, 1, 5, 1, 4, 0, 5,
    -- filter=96 channel=23
    1, 3, 3, -10, 5, -3, 0, -6, 12,
    -- filter=96 channel=24
    -6, 7, 3, -2, -4, -1, -1, -4, -5,
    -- filter=96 channel=25
    3, 8, -6, 5, -1, 3, 2, -3, 6,
    -- filter=96 channel=26
    -3, 0, -10, 6, 3, 4, 5, 6, 0,
    -- filter=96 channel=27
    0, 0, -3, -1, 1, -1, -5, -7, 0,
    -- filter=96 channel=28
    6, -2, 1, -4, -5, -1, 0, 0, -5,
    -- filter=96 channel=29
    1, -1, 3, -5, -8, -2, 4, -9, 0,
    -- filter=96 channel=30
    -4, 0, -2, -7, 10, -4, 5, -1, 0,
    -- filter=96 channel=31
    -3, 0, 8, -9, 6, 0, 2, -10, -5,
    -- filter=96 channel=32
    -8, 9, 7, 6, -2, 0, 2, -7, 11,
    -- filter=96 channel=33
    -4, 0, 8, 2, 0, 1, 3, -3, -3,
    -- filter=96 channel=34
    0, -6, -4, -1, -2, -1, 5, 11, 6,
    -- filter=96 channel=35
    -3, -2, -7, 4, 1, -2, -1, 7, 5,
    -- filter=96 channel=36
    7, 0, -6, 1, -3, 2, 5, 2, 0,
    -- filter=96 channel=37
    -14, 4, -6, -10, 10, 2, 1, 9, -1,
    -- filter=96 channel=38
    6, 0, -5, -6, 0, -8, 1, -7, -4,
    -- filter=96 channel=39
    0, 0, -4, -7, 2, 8, -7, 2, 0,
    -- filter=96 channel=40
    2, 2, 2, -8, -10, 1, -2, -10, -4,
    -- filter=96 channel=41
    -4, 1, -6, 2, -8, 0, 4, 11, -6,
    -- filter=96 channel=42
    2, 6, -6, -1, 0, 0, -4, 0, 5,
    -- filter=96 channel=43
    0, 7, 3, -3, 0, 0, -4, -5, 5,
    -- filter=96 channel=44
    -4, 1, 0, 1, 12, -9, -6, -5, 3,
    -- filter=96 channel=45
    0, 4, 3, 2, 2, -5, 0, 6, 2,
    -- filter=96 channel=46
    -2, 2, 4, -1, 7, -5, -4, 1, -4,
    -- filter=96 channel=47
    -4, 0, 0, -4, 17, -4, 4, 5, -12,
    -- filter=96 channel=48
    -1, -1, 0, -2, -6, 2, 6, 0, 1,
    -- filter=96 channel=49
    -6, -9, -1, -1, 0, 8, -8, -5, 13,
    -- filter=96 channel=50
    -1, 2, -2, -5, 0, -2, 4, -5, 2,
    -- filter=96 channel=51
    -5, 0, 0, -3, -4, 4, 0, 2, 5,
    -- filter=96 channel=52
    7, 0, 5, 0, 4, -1, 5, 6, 8,
    -- filter=96 channel=53
    -1, 8, -4, -4, -4, 7, -4, 1, 6,
    -- filter=96 channel=54
    5, 0, -5, -6, 0, 0, 4, -3, 6,
    -- filter=96 channel=55
    6, 6, 5, 5, 0, -2, -5, -14, 12,
    -- filter=96 channel=56
    1, 6, -3, 0, 2, 6, 2, 0, -1,
    -- filter=96 channel=57
    -7, 4, -4, 5, 2, -2, 4, -2, 5,
    -- filter=96 channel=58
    -6, 5, 3, 3, 3, 1, 2, 4, -4,
    -- filter=96 channel=59
    -5, 6, 6, 6, -5, -4, -1, -8, 0,
    -- filter=96 channel=60
    4, 6, -2, 4, 0, -2, -5, 7, -2,
    -- filter=96 channel=61
    -2, 1, 7, -6, 2, -7, 8, 4, 4,
    -- filter=96 channel=62
    -1, -4, 5, 1, -7, -4, 5, 4, 3,
    -- filter=96 channel=63
    4, 4, -4, 8, 3, 0, 1, 0, -2,
    -- filter=96 channel=64
    2, 2, 0, -4, -9, 1, -4, -8, -1,
    -- filter=96 channel=65
    -1, 0, -6, 3, -2, 5, -5, 0, 5,
    -- filter=96 channel=66
    -7, -1, 0, 1, 8, 2, 9, 3, 2,
    -- filter=96 channel=67
    -2, -3, 6, -3, -6, -2, 5, -6, -6,
    -- filter=96 channel=68
    0, -9, -8, 0, 1, 0, 6, -3, 3,
    -- filter=96 channel=69
    0, 3, 0, -3, 7, -7, -4, 0, 0,
    -- filter=96 channel=70
    -6, -5, -1, 0, -8, -1, 1, -6, 10,
    -- filter=96 channel=71
    -2, 0, 6, 3, 3, -1, 2, 3, 1,
    -- filter=96 channel=72
    4, 1, 7, -1, -2, -1, 5, -4, 2,
    -- filter=96 channel=73
    -1, -2, -6, 3, -3, -5, 1, 5, 10,
    -- filter=96 channel=74
    1, 1, 4, 0, 1, 0, 3, 4, 5,
    -- filter=96 channel=75
    -5, 0, -5, -1, 20, -6, 4, 6, -15,
    -- filter=96 channel=76
    2, -3, -4, -3, -7, -4, -3, -1, -1,
    -- filter=96 channel=77
    -7, -6, -2, 6, 0, -6, -2, -3, -4,
    -- filter=96 channel=78
    -2, -2, 1, 2, 11, -6, 3, -4, -4,
    -- filter=96 channel=79
    4, -4, 8, -4, -5, -3, 7, -8, 15,
    -- filter=96 channel=80
    -9, -2, 5, 1, 0, -5, -2, 0, -6,
    -- filter=96 channel=81
    0, -5, -3, 3, 2, 3, -3, 2, 1,
    -- filter=96 channel=82
    3, 6, 1, 0, 4, -4, 3, 2, -6,
    -- filter=96 channel=83
    -2, 2, 5, 1, -6, 2, 5, 3, -2,
    -- filter=96 channel=84
    4, -2, 0, 6, -4, -2, -3, 2, 8,
    -- filter=96 channel=85
    -3, 6, 7, 2, 1, -1, -3, -6, -1,
    -- filter=96 channel=86
    -3, 0, 2, -2, 6, 2, -7, 0, 8,
    -- filter=96 channel=87
    0, -3, 4, -5, -3, 4, 2, -4, 4,
    -- filter=96 channel=88
    -3, -5, -4, 0, -4, -7, -4, -1, -2,
    -- filter=96 channel=89
    -2, 0, 5, 7, -3, 0, -2, -14, 0,
    -- filter=96 channel=90
    1, 7, 7, -8, 3, 1, 1, -2, -6,
    -- filter=96 channel=91
    4, -6, 1, -10, 0, -5, 0, 4, 11,
    -- filter=96 channel=92
    -5, -4, -5, 3, -1, 1, -2, 6, -7,
    -- filter=96 channel=93
    -11, 1, -7, -7, 8, -5, 1, 11, -2,
    -- filter=96 channel=94
    -1, 0, 0, 7, -3, 4, 1, 2, 1,
    -- filter=96 channel=95
    -8, 0, -5, 2, 3, 4, 3, 6, 4,
    -- filter=96 channel=96
    0, 0, -2, -7, 0, 0, 0, -6, 1,
    -- filter=96 channel=97
    -6, 4, -5, 0, 0, 5, -8, -1, 0,
    -- filter=96 channel=98
    4, 7, -3, -2, -2, 0, 0, -9, 9,
    -- filter=96 channel=99
    6, 2, 0, 1, 5, -2, 6, -9, -2,
    -- filter=96 channel=100
    -2, -4, 0, 6, -1, 8, -5, 6, 8,
    -- filter=96 channel=101
    -8, -3, -1, -5, 0, 2, 4, 6, 0,
    -- filter=96 channel=102
    7, 2, 5, 7, 3, -3, 4, -2, 2,
    -- filter=96 channel=103
    0, 0, 2, 5, 19, -9, 4, -5, -5,
    -- filter=96 channel=104
    4, -5, -4, 5, 0, -9, 3, 1, -2,
    -- filter=96 channel=105
    0, -8, -1, 6, 3, -1, -8, -7, 6,
    -- filter=96 channel=106
    4, 5, 1, 2, -9, 7, -2, 0, 0,
    -- filter=96 channel=107
    7, -2, -5, 4, -6, -2, 3, -4, 8,
    -- filter=96 channel=108
    2, -6, -8, 0, 2, 0, 5, 7, -1,
    -- filter=96 channel=109
    -1, 3, 1, -3, -1, -9, 5, -8, 2,
    -- filter=96 channel=110
    -6, 5, 2, 2, 7, -2, -2, 3, -4,
    -- filter=96 channel=111
    5, -4, -8, 0, 2, -8, 0, -1, -2,
    -- filter=96 channel=112
    -1, 7, -3, 3, 4, -8, 0, -6, -1,
    -- filter=96 channel=113
    1, 4, 8, -4, -2, 0, 6, -10, 5,
    -- filter=96 channel=114
    -2, -4, -5, 0, 1, -4, 3, 4, 10,
    -- filter=96 channel=115
    -6, -1, -6, 7, 7, 0, -6, -4, -6,
    -- filter=96 channel=116
    4, -4, 7, 4, 1, -5, 2, 0, 10,
    -- filter=96 channel=117
    -6, -2, 5, 4, 2, -3, 5, 5, -3,
    -- filter=96 channel=118
    3, 5, 3, -1, -6, -5, 6, 1, 6,
    -- filter=96 channel=119
    3, -1, 4, 7, 0, 3, -4, 5, -7,
    -- filter=96 channel=120
    2, 4, -1, -10, -2, -6, -5, -7, 9,
    -- filter=96 channel=121
    5, 4, 1, -4, 0, -3, 1, 5, 0,
    -- filter=96 channel=122
    -12, 9, -4, 0, 12, -3, 4, 7, -16,
    -- filter=96 channel=123
    2, -3, 6, -4, 2, 4, -4, 2, 5,
    -- filter=96 channel=124
    0, 4, 4, -3, -7, -5, 3, -7, 7,
    -- filter=96 channel=125
    -4, 1, 0, 0, 0, -2, 8, -5, -3,
    -- filter=96 channel=126
    0, 4, 0, 1, 1, 3, -3, 3, 2,
    -- filter=96 channel=127
    1, -1, 0, 1, 1, -1, 0, 5, -7,
    -- filter=97 channel=0
    -16, 8, 2, -30, 13, -10, -7, 18, 0,
    -- filter=97 channel=1
    -8, 7, -3, -29, 21, -5, -13, 13, 2,
    -- filter=97 channel=2
    -5, 3, 5, 8, 1, 0, 1, -2, -5,
    -- filter=97 channel=3
    0, -11, 3, -5, -13, 2, 0, 0, 0,
    -- filter=97 channel=4
    0, 0, 6, 0, -9, -2, 1, 0, -4,
    -- filter=97 channel=5
    -9, 9, 6, -15, 14, 3, -1, 8, -4,
    -- filter=97 channel=6
    2, 10, -6, 1, 0, 1, -7, 4, -8,
    -- filter=97 channel=7
    0, -1, -3, 7, -4, -1, 6, 5, 6,
    -- filter=97 channel=8
    0, -7, 0, 5, -3, 15, 2, -2, 13,
    -- filter=97 channel=9
    0, 4, -2, 4, 6, -9, -6, -1, -2,
    -- filter=97 channel=10
    -2, 8, -5, -3, 13, -8, -3, -1, 2,
    -- filter=97 channel=11
    10, 9, -8, 13, 12, -11, -2, -9, -7,
    -- filter=97 channel=12
    -2, 3, 10, -4, 12, 9, 0, 12, 0,
    -- filter=97 channel=13
    0, 0, -4, -6, 21, -5, -7, 9, -2,
    -- filter=97 channel=14
    -1, -4, -4, 7, -7, 1, 6, -3, -2,
    -- filter=97 channel=15
    5, -3, -3, 6, 8, -1, -12, 2, -7,
    -- filter=97 channel=16
    4, 6, -4, -12, 10, -5, 2, -1, -6,
    -- filter=97 channel=17
    4, 3, 3, -3, -4, 4, 6, -1, 3,
    -- filter=97 channel=18
    -1, 18, -15, 2, 30, -9, -10, 11, -15,
    -- filter=97 channel=19
    0, -7, -2, 1, -4, -3, -3, -6, -2,
    -- filter=97 channel=20
    11, 6, -8, 12, 10, -13, -8, 0, -17,
    -- filter=97 channel=21
    -6, -7, 0, -9, -5, -1, 0, 0, -1,
    -- filter=97 channel=22
    -1, 3, -2, -6, -1, 0, 0, 2, 0,
    -- filter=97 channel=23
    0, -10, 1, 6, -8, -9, 0, -5, 3,
    -- filter=97 channel=24
    -5, -5, -3, 5, 0, -3, 0, -1, 2,
    -- filter=97 channel=25
    -2, 6, -8, -9, 19, -6, -7, 12, 0,
    -- filter=97 channel=26
    -9, 5, 0, -9, 0, -3, 4, 0, 9,
    -- filter=97 channel=27
    -2, -8, -8, -9, 14, -9, -12, -2, -5,
    -- filter=97 channel=28
    1, -4, -2, 3, 0, 0, 6, 7, 3,
    -- filter=97 channel=29
    7, 12, 0, 6, 15, -10, -16, -1, -17,
    -- filter=97 channel=30
    -10, 2, 6, -6, 11, 6, -8, 6, 1,
    -- filter=97 channel=31
    -7, -12, -4, -7, -1, 2, -7, -5, 14,
    -- filter=97 channel=32
    0, 11, -7, 1, 29, -1, -5, 9, -15,
    -- filter=97 channel=33
    -4, 4, -7, -11, 2, -3, -10, 13, -9,
    -- filter=97 channel=34
    11, 7, 11, 8, 9, 24, -2, 5, 24,
    -- filter=97 channel=35
    -4, 4, -2, 2, 1, 3, -5, 1, -4,
    -- filter=97 channel=36
    -4, 6, 0, 5, 1, 2, 4, -6, 7,
    -- filter=97 channel=37
    -15, 6, -1, -17, 8, -8, -15, 0, 5,
    -- filter=97 channel=38
    -6, -4, -8, -7, 8, -2, 0, 7, -7,
    -- filter=97 channel=39
    -1, -4, 2, 4, 8, -8, -10, -8, -11,
    -- filter=97 channel=40
    -5, -1, -7, 3, -2, -10, 0, 3, -7,
    -- filter=97 channel=41
    10, 25, -1, 10, 34, 6, 15, 32, -3,
    -- filter=97 channel=42
    -6, 0, 1, -8, -9, -1, 1, 3, 5,
    -- filter=97 channel=43
    -4, -6, 6, -6, 4, 0, 4, 3, -9,
    -- filter=97 channel=44
    -7, -6, -5, -6, 0, 4, 2, 3, -3,
    -- filter=97 channel=45
    -3, -5, -3, -4, 5, 2, -10, 4, -10,
    -- filter=97 channel=46
    3, 5, 4, -2, 6, 0, 0, 1, 3,
    -- filter=97 channel=47
    -11, -2, -9, -12, 3, -11, 5, 7, -3,
    -- filter=97 channel=48
    -14, -1, -7, -8, -1, -8, 6, -9, -4,
    -- filter=97 channel=49
    -7, 2, 0, 4, 0, -7, 0, -1, -3,
    -- filter=97 channel=50
    2, -13, -5, -5, -5, 0, 1, -6, 2,
    -- filter=97 channel=51
    -2, -6, -2, -6, -3, -6, -4, -2, 1,
    -- filter=97 channel=52
    1, 6, 0, 7, 6, 7, -6, -4, 12,
    -- filter=97 channel=53
    2, 10, -5, 7, 6, 2, -2, -8, 3,
    -- filter=97 channel=54
    0, 0, -1, -5, -3, -3, 1, 0, -5,
    -- filter=97 channel=55
    7, 14, -7, 8, 21, -11, -9, 1, -7,
    -- filter=97 channel=56
    0, 9, 6, 13, 2, 11, 5, 4, 9,
    -- filter=97 channel=57
    5, 3, -4, -5, 11, -1, -3, 2, 0,
    -- filter=97 channel=58
    -7, 9, 10, 0, 9, 9, 6, 9, 4,
    -- filter=97 channel=59
    -3, 1, -11, -11, 8, -4, 0, 10, -7,
    -- filter=97 channel=60
    -5, -4, -4, -3, 0, -1, 0, -4, 1,
    -- filter=97 channel=61
    1, 5, 2, 4, 5, 5, 6, 8, 2,
    -- filter=97 channel=62
    5, 1, -7, -1, 5, 3, 4, -4, 2,
    -- filter=97 channel=63
    3, 12, 4, -4, 11, 2, 5, 1, -2,
    -- filter=97 channel=64
    -3, -6, -3, 2, 7, -2, -6, 0, 1,
    -- filter=97 channel=65
    -2, -2, 5, -1, -4, 0, -3, 1, 7,
    -- filter=97 channel=66
    0, 18, 10, 0, 27, 8, 8, 15, 0,
    -- filter=97 channel=67
    3, 3, 3, 1, 4, 5, 1, -3, -6,
    -- filter=97 channel=68
    -7, 8, 4, 0, 0, -10, 4, 3, -1,
    -- filter=97 channel=69
    3, 6, -4, 3, 11, 0, -1, 3, 6,
    -- filter=97 channel=70
    -9, -13, 4, -2, -5, -1, -5, -9, 9,
    -- filter=97 channel=71
    -5, -9, 3, -5, -1, -6, -3, 3, 2,
    -- filter=97 channel=72
    7, -5, 4, 3, 1, -7, 0, 0, -1,
    -- filter=97 channel=73
    3, 1, 0, 5, 10, 1, -1, -7, -8,
    -- filter=97 channel=74
    -1, -1, -3, 7, -1, 17, 5, -7, 17,
    -- filter=97 channel=75
    -16, 10, 0, -14, 20, -9, -5, 24, -11,
    -- filter=97 channel=76
    -1, 11, -7, 1, 16, -8, -2, 3, -16,
    -- filter=97 channel=77
    -6, -5, 3, -4, 1, 5, 4, -4, 3,
    -- filter=97 channel=78
    2, -3, 0, 4, 4, -2, 7, 2, 0,
    -- filter=97 channel=79
    0, 8, -1, -13, 21, -10, -5, 18, -14,
    -- filter=97 channel=80
    -11, -4, -7, -10, 4, -2, -2, -4, 0,
    -- filter=97 channel=81
    -6, -6, -3, 0, 4, -1, 7, 4, 0,
    -- filter=97 channel=82
    2, -3, 0, -1, 0, -7, -3, 0, -9,
    -- filter=97 channel=83
    2, 3, -3, -2, -2, 0, -1, -6, -5,
    -- filter=97 channel=84
    5, 1, 1, 7, 14, 3, -6, 11, -3,
    -- filter=97 channel=85
    0, -5, -2, -4, 3, -4, -5, -2, -6,
    -- filter=97 channel=86
    -4, 12, 6, -4, 5, 12, 0, 15, 13,
    -- filter=97 channel=87
    0, 4, 0, 1, 6, 6, 1, 6, 4,
    -- filter=97 channel=88
    2, -7, -2, 6, -3, 8, 1, -1, 4,
    -- filter=97 channel=89
    5, 10, -10, -12, 18, -13, -1, 11, -3,
    -- filter=97 channel=90
    4, -1, 4, 0, -6, 2, 5, -6, 14,
    -- filter=97 channel=91
    2, -1, -2, 6, 0, -5, -12, -5, 2,
    -- filter=97 channel=92
    1, -4, 8, 7, -7, -1, 6, 4, 3,
    -- filter=97 channel=93
    -7, 10, -1, -16, 5, 0, 4, 4, 8,
    -- filter=97 channel=94
    0, -5, 1, 5, -3, 0, 3, 4, -4,
    -- filter=97 channel=95
    -4, 0, -2, 5, -3, -2, -3, -3, -3,
    -- filter=97 channel=96
    -8, -8, -6, -10, -1, -5, 4, -4, -2,
    -- filter=97 channel=97
    -4, -3, 0, -6, -3, -4, -3, -3, 3,
    -- filter=97 channel=98
    -8, -6, 0, -8, 5, -6, 0, -1, -2,
    -- filter=97 channel=99
    -3, 1, 8, 6, 11, 4, 0, -8, 11,
    -- filter=97 channel=100
    9, 3, 8, 5, -3, 10, 10, 6, 1,
    -- filter=97 channel=101
    5, -3, -4, 3, -7, -3, -6, -10, -7,
    -- filter=97 channel=102
    5, 0, 5, 5, 0, -5, -2, -5, 0,
    -- filter=97 channel=103
    -9, 6, -5, -6, -5, -7, 0, -5, -6,
    -- filter=97 channel=104
    -6, 2, 0, -8, 1, -4, -5, -5, -7,
    -- filter=97 channel=105
    6, 7, -9, 9, 7, -5, -1, -6, -13,
    -- filter=97 channel=106
    2, 0, -9, 5, 0, -8, -3, -2, -1,
    -- filter=97 channel=107
    -3, 0, 3, 11, 0, 2, -3, -9, -9,
    -- filter=97 channel=108
    6, 0, 4, 0, 9, 5, 5, 14, -2,
    -- filter=97 channel=109
    -1, 0, 0, 0, 22, -8, -5, -4, -1,
    -- filter=97 channel=110
    -1, -2, 5, 2, -3, -1, 1, 3, 0,
    -- filter=97 channel=111
    -6, 10, -3, 0, 11, -4, 3, 1, -4,
    -- filter=97 channel=112
    -4, 0, -6, -5, -2, 1, -8, -3, 2,
    -- filter=97 channel=113
    1, 0, -6, -6, -2, 0, 1, 6, 4,
    -- filter=97 channel=114
    -11, 22, 1, -13, 27, -14, -11, 16, -10,
    -- filter=97 channel=115
    -3, 0, -6, 0, 7, 7, 4, 4, 3,
    -- filter=97 channel=116
    -6, 0, -7, -2, 5, -11, -5, -8, 2,
    -- filter=97 channel=117
    -4, 0, 2, -5, -3, -7, -5, -5, -7,
    -- filter=97 channel=118
    1, 5, -1, -1, 1, 1, 1, 1, -1,
    -- filter=97 channel=119
    6, 7, 4, 21, 2, 15, 15, 4, 11,
    -- filter=97 channel=120
    1, -11, 3, 1, -3, -1, 0, -12, 0,
    -- filter=97 channel=121
    2, 3, 4, -7, 16, -2, 1, 12, -5,
    -- filter=97 channel=122
    -1, -1, -2, -15, -11, -9, -5, 0, 0,
    -- filter=97 channel=123
    1, 1, 8, 10, 0, 12, 2, 0, 11,
    -- filter=97 channel=124
    -3, 5, -8, 0, 0, -13, -11, 1, -15,
    -- filter=97 channel=125
    -2, 2, 3, 1, 4, -1, 3, 7, 7,
    -- filter=97 channel=126
    -3, 6, -2, -6, 7, -5, 1, 9, -13,
    -- filter=97 channel=127
    -1, 11, 5, 6, 10, -7, 5, 3, 2,
    -- filter=98 channel=0
    13, 11, 1, 15, 5, -4, -2, -11, -16,
    -- filter=98 channel=1
    11, 10, -3, 9, 3, -10, -13, -16, -10,
    -- filter=98 channel=2
    4, 0, 2, -4, -5, -4, -6, -1, 0,
    -- filter=98 channel=3
    9, 19, 15, 2, 1, 10, 1, 7, -3,
    -- filter=98 channel=4
    3, 3, 8, -5, 8, 6, -5, 6, 7,
    -- filter=98 channel=5
    7, 11, 6, -2, 4, 1, -13, -12, 1,
    -- filter=98 channel=6
    11, 7, 0, -7, 0, 2, 6, -7, -2,
    -- filter=98 channel=7
    0, 0, 3, -4, -6, 0, 6, -4, -2,
    -- filter=98 channel=8
    2, -3, -2, 1, -9, -4, -10, 1, 2,
    -- filter=98 channel=9
    2, 7, 4, 2, 2, -1, 7, 10, 3,
    -- filter=98 channel=10
    0, 7, 9, -11, -13, -5, -3, -7, 3,
    -- filter=98 channel=11
    2, 10, 3, 0, -5, 0, 1, 7, 4,
    -- filter=98 channel=12
    -1, -4, -6, -10, -7, 0, -1, -5, -7,
    -- filter=98 channel=13
    6, 1, 12, -12, -7, -14, -1, 0, -5,
    -- filter=98 channel=14
    5, 0, 5, 6, 7, -3, 3, 3, -7,
    -- filter=98 channel=15
    9, 11, 12, -5, -14, -14, 0, 2, -5,
    -- filter=98 channel=16
    -2, -2, -6, -3, -3, -4, -8, -5, -1,
    -- filter=98 channel=17
    -5, 5, 4, -3, 1, 0, 2, 4, 7,
    -- filter=98 channel=18
    24, 20, 12, 2, -10, -25, 5, -1, -5,
    -- filter=98 channel=19
    -2, 1, 7, 2, -1, -4, 1, 0, 7,
    -- filter=98 channel=20
    -3, 18, 15, -10, -3, -10, 7, 8, 11,
    -- filter=98 channel=21
    -3, -8, 4, 3, -7, 9, 8, -2, 15,
    -- filter=98 channel=22
    -1, 5, 4, -9, -12, -10, -7, -2, -10,
    -- filter=98 channel=23
    8, 29, 15, -13, -26, -20, 0, 14, 0,
    -- filter=98 channel=24
    -6, 2, -6, -2, 5, 2, -6, -4, -6,
    -- filter=98 channel=25
    1, 1, 10, -2, -12, -17, -3, 2, 7,
    -- filter=98 channel=26
    -8, 0, 0, 3, 3, 12, 2, 0, -4,
    -- filter=98 channel=27
    16, 15, 7, -15, -13, -30, 0, 5, 4,
    -- filter=98 channel=28
    -7, 0, 0, -2, 2, -1, 0, 5, 3,
    -- filter=98 channel=29
    11, 13, 0, -7, 0, -3, -4, 9, 7,
    -- filter=98 channel=30
    8, 12, 0, 3, -7, -7, -9, 2, 2,
    -- filter=98 channel=31
    -1, 4, 12, -11, -14, -4, 6, 11, 5,
    -- filter=98 channel=32
    10, 15, 15, -6, -17, -25, -3, 0, -7,
    -- filter=98 channel=33
    18, 13, 10, 0, -17, -20, 0, -5, -5,
    -- filter=98 channel=34
    -5, -6, -7, -17, -12, -13, -16, 3, -7,
    -- filter=98 channel=35
    5, 3, -5, -5, -6, 4, -5, 6, 6,
    -- filter=98 channel=36
    -9, -13, 6, -11, 0, 9, -4, -3, 0,
    -- filter=98 channel=37
    1, 13, 0, 8, 0, -6, -8, -4, -8,
    -- filter=98 channel=38
    0, 15, 5, -8, -6, -7, -2, 0, 0,
    -- filter=98 channel=39
    3, -2, 8, -9, -3, -1, 2, 0, 2,
    -- filter=98 channel=40
    -4, 6, 10, -10, 0, -7, 0, 5, -7,
    -- filter=98 channel=41
    -4, -1, 3, 1, -1, -9, -5, -13, 0,
    -- filter=98 channel=42
    3, 7, 6, 10, -2, -3, 2, 0, -2,
    -- filter=98 channel=43
    6, 19, 1, -1, -11, -4, 0, -3, -6,
    -- filter=98 channel=44
    6, -2, -8, -6, 2, -8, -6, 0, -4,
    -- filter=98 channel=45
    0, 10, -3, -5, 3, -2, 0, 5, -5,
    -- filter=98 channel=46
    5, 4, 2, 6, 5, 1, 4, -7, -2,
    -- filter=98 channel=47
    10, 1, 0, -3, 5, 5, -7, 3, 9,
    -- filter=98 channel=48
    0, -5, 0, -5, 0, -7, 4, 8, 7,
    -- filter=98 channel=49
    4, 7, 3, -1, -5, -7, 4, 12, 9,
    -- filter=98 channel=50
    2, 13, 6, -3, 1, -9, 4, 13, 9,
    -- filter=98 channel=51
    -6, -1, 6, 2, -5, 7, 1, 0, 2,
    -- filter=98 channel=52
    -1, 0, -4, -6, -10, -12, -12, -8, -10,
    -- filter=98 channel=53
    1, 11, 1, -1, 5, -5, 1, 1, -2,
    -- filter=98 channel=54
    2, 3, 1, -3, 0, 4, 5, 2, 0,
    -- filter=98 channel=55
    4, 15, 4, -14, -16, -10, 7, 13, 8,
    -- filter=98 channel=56
    -5, -5, -6, 0, 0, -13, 0, 0, -2,
    -- filter=98 channel=57
    -2, 3, -7, 6, -5, -6, 2, 0, 2,
    -- filter=98 channel=58
    0, 0, 0, -2, -1, -1, -6, -9, -1,
    -- filter=98 channel=59
    8, 2, 9, -5, -8, -14, 1, 1, 11,
    -- filter=98 channel=60
    -4, 2, 0, 6, -4, -6, -5, 0, 0,
    -- filter=98 channel=61
    -3, -6, -6, -11, 1, -1, -6, -3, -5,
    -- filter=98 channel=62
    4, 2, 9, 0, -7, 7, 5, -4, -8,
    -- filter=98 channel=63
    -2, 10, -4, 0, -3, 9, -5, 2, -3,
    -- filter=98 channel=64
    -5, 0, -3, -6, -2, -1, 0, 0, 9,
    -- filter=98 channel=65
    0, -3, -5, -1, -1, 4, 4, 2, -3,
    -- filter=98 channel=66
    -2, -8, -9, -15, -9, -12, -1, -11, -8,
    -- filter=98 channel=67
    -6, -7, 0, -4, 4, -5, -3, 6, 0,
    -- filter=98 channel=68
    -1, 5, 4, -4, -2, 3, -6, -1, 0,
    -- filter=98 channel=69
    -3, 0, -5, -1, 7, -4, -2, -3, -6,
    -- filter=98 channel=70
    14, 3, 6, -9, -13, -20, 5, 6, -11,
    -- filter=98 channel=71
    0, 8, 2, 2, -3, -1, 2, 0, -1,
    -- filter=98 channel=72
    -5, 7, 3, -10, -2, -1, 10, 12, 15,
    -- filter=98 channel=73
    11, -1, -5, -6, -9, -4, 3, 7, 4,
    -- filter=98 channel=74
    -9, -6, -12, -12, -14, -9, 0, 4, -9,
    -- filter=98 channel=75
    14, 16, 8, 12, 1, -2, -9, -19, -6,
    -- filter=98 channel=76
    -3, 13, 17, -14, -1, -2, 0, 4, 0,
    -- filter=98 channel=77
    -7, 4, 6, 1, -3, 7, 1, 3, 3,
    -- filter=98 channel=78
    1, 10, 1, -8, -5, -2, 0, -8, 2,
    -- filter=98 channel=79
    16, 19, 4, 0, -21, -31, 6, -4, -1,
    -- filter=98 channel=80
    11, 0, 8, 6, -7, 0, 9, 7, 14,
    -- filter=98 channel=81
    3, 2, -2, -2, -6, -6, 5, -6, 7,
    -- filter=98 channel=82
    -1, 6, -3, 4, 4, 0, -1, -4, -4,
    -- filter=98 channel=83
    -3, 1, -10, -1, 4, 5, 8, 1, 7,
    -- filter=98 channel=84
    5, 8, 5, -11, -6, -12, -6, 3, -6,
    -- filter=98 channel=85
    1, 4, -5, 5, -1, 0, -3, 0, 4,
    -- filter=98 channel=86
    -5, -4, 0, -8, -13, 2, -1, -12, -5,
    -- filter=98 channel=87
    -3, -4, 6, -2, -12, -13, -6, -4, -3,
    -- filter=98 channel=88
    -12, -12, -7, -9, -3, -2, -4, -4, 5,
    -- filter=98 channel=89
    11, 14, 21, -14, -17, -5, 1, 0, 7,
    -- filter=98 channel=90
    0, -5, -2, -15, 0, 5, -8, 0, 4,
    -- filter=98 channel=91
    0, 10, 1, -12, -12, -19, 2, 13, 4,
    -- filter=98 channel=92
    -6, 4, -4, -6, -5, 0, 4, -6, -9,
    -- filter=98 channel=93
    9, 0, 2, 4, 2, -7, -8, -6, 6,
    -- filter=98 channel=94
    6, 5, 5, 5, -2, 2, -1, 5, -4,
    -- filter=98 channel=95
    1, -1, -2, -1, 1, -6, 3, 4, 4,
    -- filter=98 channel=96
    3, 0, -5, -2, 2, -4, 5, 5, -5,
    -- filter=98 channel=97
    0, 13, 6, 0, 1, 4, -2, 0, -7,
    -- filter=98 channel=98
    11, 21, 10, 0, -17, -12, 5, 11, 5,
    -- filter=98 channel=99
    4, 15, 7, -21, -17, -16, -4, 9, 12,
    -- filter=98 channel=100
    -4, 0, 4, 5, 0, -6, -8, 1, -8,
    -- filter=98 channel=101
    8, 3, 10, 1, 9, 7, -5, 1, 6,
    -- filter=98 channel=102
    -1, -1, 6, 6, 7, -5, -4, 0, -2,
    -- filter=98 channel=103
    13, 18, -1, 6, 7, 9, 0, -8, 0,
    -- filter=98 channel=104
    4, -9, -3, 2, -5, -4, 4, 7, 18,
    -- filter=98 channel=105
    0, 2, 10, 1, -6, -10, -2, 1, 4,
    -- filter=98 channel=106
    7, 3, 0, 2, 1, -2, 0, 0, -1,
    -- filter=98 channel=107
    -1, 5, -1, -8, -4, -15, -1, 1, -5,
    -- filter=98 channel=108
    -2, 6, 2, 3, -5, 2, 4, -10, 2,
    -- filter=98 channel=109
    4, 13, -5, -4, -10, -22, -1, 5, -3,
    -- filter=98 channel=110
    4, 8, 4, -12, -7, 5, 1, 2, -3,
    -- filter=98 channel=111
    3, -4, -5, -3, 5, 2, -5, -3, 4,
    -- filter=98 channel=112
    2, 8, -7, -8, 3, -4, -6, 9, -2,
    -- filter=98 channel=113
    3, 12, 4, -3, -5, -5, 1, 1, 0,
    -- filter=98 channel=114
    16, 22, 9, 8, -3, -24, -2, 6, -6,
    -- filter=98 channel=115
    -1, -3, -5, -5, 2, -1, 0, -6, -6,
    -- filter=98 channel=116
    -1, 7, 0, -2, -10, -10, 1, 9, 12,
    -- filter=98 channel=117
    4, -1, 6, -1, -7, 1, 6, 6, 8,
    -- filter=98 channel=118
    1, 1, -3, 5, -4, -5, -5, 6, -2,
    -- filter=98 channel=119
    -8, 0, -9, -10, -12, -17, -7, -4, -9,
    -- filter=98 channel=120
    3, 3, -7, -15, -14, -19, -1, 10, -1,
    -- filter=98 channel=121
    3, 0, 11, -1, -8, -11, 4, -1, 0,
    -- filter=98 channel=122
    -6, 1, 0, 7, 6, 0, -7, 2, 10,
    -- filter=98 channel=123
    -1, 0, -8, -1, -1, -8, -5, -5, -10,
    -- filter=98 channel=124
    2, 1, -2, -9, -4, -1, -2, 7, -7,
    -- filter=98 channel=125
    2, 2, 7, -10, -1, -8, -6, 4, 17,
    -- filter=98 channel=126
    8, 17, 11, 3, 0, -5, 8, 0, 0,
    -- filter=98 channel=127
    -2, 0, 4, -7, 5, -6, -7, 2, 6,
    -- filter=99 channel=0
    5, 4, -1, -6, -11, 4, 3, 3, 10,
    -- filter=99 channel=1
    3, -10, 9, 2, -14, 2, -6, -5, 9,
    -- filter=99 channel=2
    2, 2, -3, -2, -1, 0, 2, 2, -7,
    -- filter=99 channel=3
    -6, 6, 4, -7, -8, 3, -1, 0, 2,
    -- filter=99 channel=4
    -8, -7, -5, -5, -12, -4, 0, -8, 0,
    -- filter=99 channel=5
    -1, 0, 1, 1, 1, 2, 6, -2, 4,
    -- filter=99 channel=6
    -5, 0, -4, 6, 1, 6, 1, 4, -2,
    -- filter=99 channel=7
    0, 1, 2, 2, 5, -5, 0, 5, -1,
    -- filter=99 channel=8
    -5, 4, -2, -9, -1, 2, 3, -7, 6,
    -- filter=99 channel=9
    -5, 3, -5, 0, 0, 3, -4, -4, 1,
    -- filter=99 channel=10
    8, -3, -2, 0, -5, -7, -8, -10, 2,
    -- filter=99 channel=11
    -5, 8, 3, 1, 14, 7, -1, 0, 3,
    -- filter=99 channel=12
    -8, 0, 4, -7, -8, 0, -1, 4, -2,
    -- filter=99 channel=13
    -3, -2, 3, 0, -3, -4, -3, -4, 0,
    -- filter=99 channel=14
    0, -2, -3, -6, 4, -2, 4, -3, 3,
    -- filter=99 channel=15
    -9, 9, 7, 1, 11, 8, 2, -4, -7,
    -- filter=99 channel=16
    -1, 2, 4, -4, -3, 3, 4, -5, -9,
    -- filter=99 channel=17
    -1, 7, 6, 6, -6, -2, 3, 1, -4,
    -- filter=99 channel=18
    -8, 4, 15, -5, 6, 10, -12, 0, 0,
    -- filter=99 channel=19
    3, -1, -6, -3, -4, 6, -2, 7, -6,
    -- filter=99 channel=20
    -11, 10, -1, -5, 15, 9, 1, 3, 3,
    -- filter=99 channel=21
    1, -2, -1, 0, -7, -7, -4, 0, -3,
    -- filter=99 channel=22
    1, -1, 0, -3, 0, 5, 0, -4, 5,
    -- filter=99 channel=23
    4, 1, 16, -1, 6, 16, -4, -8, -5,
    -- filter=99 channel=24
    5, 0, 4, -2, 2, 2, 7, 4, -3,
    -- filter=99 channel=25
    5, 1, 0, -1, -6, 0, -2, -7, 2,
    -- filter=99 channel=26
    2, 4, -6, 0, 6, 3, 7, 4, 4,
    -- filter=99 channel=27
    -5, 6, 8, 2, -7, 10, 2, -12, -8,
    -- filter=99 channel=28
    0, 5, 0, -2, 3, 0, 0, -1, 2,
    -- filter=99 channel=29
    -7, 6, 6, -1, 11, 3, -7, 6, -6,
    -- filter=99 channel=30
    3, 6, -1, -6, -5, 1, -4, 1, 1,
    -- filter=99 channel=31
    7, -4, -2, -4, -16, -3, -4, -3, -4,
    -- filter=99 channel=32
    -2, -6, 17, -2, 4, 9, -9, 0, -3,
    -- filter=99 channel=33
    0, -3, 4, -2, 0, 4, -1, -6, 2,
    -- filter=99 channel=34
    -8, 0, 0, -1, -10, 10, -7, -1, 0,
    -- filter=99 channel=35
    6, -3, 5, -5, 2, -1, 6, 4, -6,
    -- filter=99 channel=36
    0, -6, -5, -2, 0, 4, -7, 3, -6,
    -- filter=99 channel=37
    2, -4, -1, 1, -12, -2, -8, 0, 5,
    -- filter=99 channel=38
    4, 7, 9, 7, -2, -2, 0, 1, -7,
    -- filter=99 channel=39
    -2, 4, 3, 5, 6, 6, 5, -3, -5,
    -- filter=99 channel=40
    -3, 6, 6, 4, -4, 0, 3, 3, -7,
    -- filter=99 channel=41
    -3, -3, 9, -15, -4, 3, -7, -2, -3,
    -- filter=99 channel=42
    2, 1, 1, 3, 3, -2, 4, 0, -1,
    -- filter=99 channel=43
    -8, 10, 1, 5, 0, 0, 0, 4, 8,
    -- filter=99 channel=44
    -5, -9, -7, -6, -6, 3, -8, -11, 5,
    -- filter=99 channel=45
    -4, -6, -2, 0, -4, 1, 5, -4, -1,
    -- filter=99 channel=46
    0, 0, 0, -4, -1, -4, -6, -4, 1,
    -- filter=99 channel=47
    2, -7, -6, -4, -15, -3, 4, -13, -9,
    -- filter=99 channel=48
    6, 0, -1, -8, -15, -4, 3, -8, -4,
    -- filter=99 channel=49
    -3, 1, 2, -3, 8, 2, -5, 1, 1,
    -- filter=99 channel=50
    -3, -6, 9, 0, -10, -2, 5, -4, -1,
    -- filter=99 channel=51
    1, 4, 5, -4, -6, -1, -2, 2, 6,
    -- filter=99 channel=52
    3, -3, 9, 3, -7, 7, -5, -7, 3,
    -- filter=99 channel=53
    6, 4, 3, 2, 0, 2, 1, -6, -5,
    -- filter=99 channel=54
    4, 1, -3, 2, -4, 4, -4, -4, 3,
    -- filter=99 channel=55
    0, 5, 4, 1, -1, 0, -1, -7, -6,
    -- filter=99 channel=56
    -6, -3, -1, 1, -5, 7, -6, 2, -6,
    -- filter=99 channel=57
    -1, 0, 0, -5, 0, -5, -7, 2, -6,
    -- filter=99 channel=58
    7, 5, 3, -4, 2, -3, -4, 0, 5,
    -- filter=99 channel=59
    0, -2, 5, 0, -6, 0, -9, -3, -3,
    -- filter=99 channel=60
    5, 2, -5, 0, 1, 7, 4, 6, -4,
    -- filter=99 channel=61
    6, 5, 2, 0, -6, 0, 3, -1, -4,
    -- filter=99 channel=62
    2, 4, -6, 3, -3, 6, -5, 7, 2,
    -- filter=99 channel=63
    -3, 0, -1, 1, 3, 1, 4, -3, -3,
    -- filter=99 channel=64
    -2, 1, 1, -5, 0, -4, 6, -7, -4,
    -- filter=99 channel=65
    -4, 0, 5, 3, 3, -6, -7, 0, 4,
    -- filter=99 channel=66
    0, 3, 9, -7, -6, 4, -1, -5, 6,
    -- filter=99 channel=67
    3, -3, -1, 3, 5, -4, -2, -6, 7,
    -- filter=99 channel=68
    2, -4, 3, -5, 5, -6, -1, -4, 3,
    -- filter=99 channel=69
    7, -6, 3, 1, -1, 8, 5, -2, -4,
    -- filter=99 channel=70
    1, 1, 12, -6, -2, -1, 1, -7, 0,
    -- filter=99 channel=71
    5, 4, -5, -6, 3, 4, 1, 5, 4,
    -- filter=99 channel=72
    8, -5, -1, 5, -6, -2, -4, -2, 0,
    -- filter=99 channel=73
    1, -5, 10, -3, 3, 1, -4, -5, 3,
    -- filter=99 channel=74
    0, -5, 7, -1, -5, 2, -5, -8, -5,
    -- filter=99 channel=75
    -4, -3, 7, -6, -1, -7, -3, 0, 0,
    -- filter=99 channel=76
    -8, 7, 8, -6, 12, 1, -3, 3, 2,
    -- filter=99 channel=77
    -3, 0, 7, 1, -2, -5, 0, 5, 5,
    -- filter=99 channel=78
    4, -3, 3, -6, -5, -2, -6, 1, 0,
    -- filter=99 channel=79
    -3, 6, 11, -9, -5, 14, -7, -8, 0,
    -- filter=99 channel=80
    -4, 1, 5, -8, -2, -8, 1, -6, -13,
    -- filter=99 channel=81
    -1, 0, 5, 6, 5, 2, -5, 0, -5,
    -- filter=99 channel=82
    0, -5, 5, -6, 1, 2, -6, -3, -3,
    -- filter=99 channel=83
    1, -6, -2, 5, -9, -1, -2, 2, 3,
    -- filter=99 channel=84
    4, 2, -2, -6, -7, -3, 0, -10, 0,
    -- filter=99 channel=85
    5, -4, -5, -6, -6, -6, 7, 7, -6,
    -- filter=99 channel=86
    -2, -7, -3, -1, 1, -4, -4, -5, -4,
    -- filter=99 channel=87
    -2, -5, -5, -7, -4, 11, 0, 6, 4,
    -- filter=99 channel=88
    -2, -1, 5, 6, -7, 0, 7, 3, 0,
    -- filter=99 channel=89
    4, -1, 10, -7, -7, 6, -2, -6, -11,
    -- filter=99 channel=90
    -6, -8, -4, -6, -5, -1, -3, 2, 6,
    -- filter=99 channel=91
    5, -6, 11, 3, 3, 9, 0, -11, -7,
    -- filter=99 channel=92
    0, -3, 5, -6, -2, 0, -1, 0, 3,
    -- filter=99 channel=93
    -2, -6, 3, -9, -6, -5, -4, -2, -6,
    -- filter=99 channel=94
    0, 3, -1, 0, 2, -1, 3, -6, -5,
    -- filter=99 channel=95
    4, 7, 6, 4, -7, -6, 4, 2, 3,
    -- filter=99 channel=96
    7, 0, 4, -3, 6, -2, 4, -4, -3,
    -- filter=99 channel=97
    3, 0, 4, 1, 3, -1, 0, 0, -3,
    -- filter=99 channel=98
    1, 0, 11, -3, -12, 0, 2, -10, -11,
    -- filter=99 channel=99
    -6, -4, 1, -2, -8, 6, -2, -11, -4,
    -- filter=99 channel=100
    -3, -6, -2, -1, -5, 1, -7, 5, 2,
    -- filter=99 channel=101
    -1, 3, -2, 5, -7, -3, -1, 0, 0,
    -- filter=99 channel=102
    -3, -1, 4, 6, -4, -6, -1, -3, -2,
    -- filter=99 channel=103
    -1, -10, 3, -2, -9, -7, -6, -9, -5,
    -- filter=99 channel=104
    -5, -9, -5, -5, -5, -1, 0, -5, -2,
    -- filter=99 channel=105
    -4, 7, 5, 4, 14, 0, -3, 4, 0,
    -- filter=99 channel=106
    -5, 5, -7, -5, 8, 2, -6, -4, 2,
    -- filter=99 channel=107
    -1, 9, 3, -1, 3, 5, 2, -3, 2,
    -- filter=99 channel=108
    -1, -6, -3, 1, -5, -3, -8, 1, -6,
    -- filter=99 channel=109
    -2, -3, 11, -4, -11, 7, -6, 0, -6,
    -- filter=99 channel=110
    0, 0, 1, 4, 1, -8, 2, -8, -4,
    -- filter=99 channel=111
    -7, 0, 0, -8, -1, -2, -5, 6, 1,
    -- filter=99 channel=112
    3, -6, 3, 6, -11, 5, 5, 4, 1,
    -- filter=99 channel=113
    7, -4, -2, 1, -7, 4, 0, -8, -6,
    -- filter=99 channel=114
    -7, 3, 20, -6, 4, 18, -4, 0, 4,
    -- filter=99 channel=115
    -7, -1, 0, -7, -3, 0, 0, 0, -4,
    -- filter=99 channel=116
    8, 5, -1, 4, 0, 0, -7, -8, -5,
    -- filter=99 channel=117
    3, -2, -5, -2, -3, -8, 3, -7, -4,
    -- filter=99 channel=118
    4, -6, -4, -4, 0, -3, -6, 4, 5,
    -- filter=99 channel=119
    -9, 0, 5, 0, -7, 0, -2, -2, 4,
    -- filter=99 channel=120
    4, 0, 14, 2, 2, 5, 3, -3, -4,
    -- filter=99 channel=121
    4, -5, 5, 0, 0, 0, 1, -9, 5,
    -- filter=99 channel=122
    -10, -6, 0, 2, -17, -7, 0, -10, -4,
    -- filter=99 channel=123
    -5, -4, 0, -6, -4, 6, -5, -3, -2,
    -- filter=99 channel=124
    -2, 1, -3, 0, -1, 3, 4, -1, 3,
    -- filter=99 channel=125
    0, 0, 2, 3, -5, 3, -6, -1, 2,
    -- filter=99 channel=126
    7, 0, 6, 2, -3, -3, 0, 3, 5,
    -- filter=99 channel=127
    1, -6, -4, 5, -3, -2, -1, 0, -5,
    -- filter=100 channel=0
    7, 4, -13, 14, 7, -14, 19, 11, -5,
    -- filter=100 channel=1
    0, -4, -8, 0, 0, -10, 12, 7, -2,
    -- filter=100 channel=2
    -5, -7, 2, -1, -7, -2, -1, -2, 1,
    -- filter=100 channel=3
    0, -4, 8, -1, -5, -8, -5, 5, -9,
    -- filter=100 channel=4
    -3, -6, -13, 0, -2, -7, 6, 1, 4,
    -- filter=100 channel=5
    3, 2, -7, 5, 3, -15, 5, 1, -6,
    -- filter=100 channel=6
    -8, 3, 1, -1, -4, 0, -6, -3, 2,
    -- filter=100 channel=7
    1, 6, -6, -5, -4, -5, 2, 0, 5,
    -- filter=100 channel=8
    -2, -2, -4, 4, 5, -2, -6, -2, 0,
    -- filter=100 channel=9
    0, 5, 0, 6, 3, -6, 5, 0, -1,
    -- filter=100 channel=10
    1, -2, 1, 4, 6, 4, 0, 5, 1,
    -- filter=100 channel=11
    1, 3, -8, 2, 11, 0, -3, 5, -5,
    -- filter=100 channel=12
    1, 3, 1, -11, 8, 6, -1, 11, -4,
    -- filter=100 channel=13
    -1, 11, 1, -9, 6, 0, -6, 4, -6,
    -- filter=100 channel=14
    -4, -5, 0, -1, 7, 0, -3, 2, -1,
    -- filter=100 channel=15
    8, 1, -3, -1, 2, -12, 6, 0, -12,
    -- filter=100 channel=16
    2, -1, -8, 0, 5, 0, 2, 1, -1,
    -- filter=100 channel=17
    1, 5, -7, -2, 2, -2, 5, -5, -3,
    -- filter=100 channel=18
    5, 8, 4, -3, 5, -13, 11, 2, -2,
    -- filter=100 channel=19
    -4, 2, -2, -7, -2, -5, -3, 4, 4,
    -- filter=100 channel=20
    -4, 10, -3, -10, 12, -11, -7, 7, 1,
    -- filter=100 channel=21
    5, -10, -6, -3, 4, -6, -10, -5, -2,
    -- filter=100 channel=22
    2, 0, -5, -3, 4, 1, -3, 1, -7,
    -- filter=100 channel=23
    0, 12, 0, -7, 0, -23, -6, 2, -10,
    -- filter=100 channel=24
    -3, 7, 6, 5, -6, 6, -5, -5, 2,
    -- filter=100 channel=25
    6, 0, -4, 4, 2, -19, 5, 9, -14,
    -- filter=100 channel=26
    -5, -6, 0, -2, 1, -4, 2, 4, 5,
    -- filter=100 channel=27
    1, 2, -9, 4, 4, -29, 3, -2, -21,
    -- filter=100 channel=28
    -6, -3, 7, -6, 1, -6, -6, -7, -1,
    -- filter=100 channel=29
    1, -3, 2, -3, 3, -1, 0, 5, -9,
    -- filter=100 channel=30
    5, -4, 2, 4, 1, -5, 9, 4, -12,
    -- filter=100 channel=31
    11, 6, -9, 2, 0, -9, -1, 5, -20,
    -- filter=100 channel=32
    13, 4, -7, -6, 2, -18, 4, -2, -3,
    -- filter=100 channel=33
    15, 0, 1, 0, 6, -8, -5, -1, -19,
    -- filter=100 channel=34
    0, 10, 11, -7, 8, 8, -6, 4, 1,
    -- filter=100 channel=35
    4, 4, 6, 2, -1, 2, 5, 5, 0,
    -- filter=100 channel=36
    -8, 5, 1, -2, 6, 0, 4, -4, 9,
    -- filter=100 channel=37
    -8, -7, -14, -3, 5, -12, 10, 12, -12,
    -- filter=100 channel=38
    -1, 8, 0, 0, 3, -13, -5, 3, -7,
    -- filter=100 channel=39
    -5, 0, 0, -4, 0, -9, 4, 5, -1,
    -- filter=100 channel=40
    -3, 2, 9, -4, 4, 4, -5, 6, -1,
    -- filter=100 channel=41
    -13, 14, 11, -14, 14, 39, -5, 3, 40,
    -- filter=100 channel=42
    -1, -1, -2, 10, 4, 2, 3, 6, 1,
    -- filter=100 channel=43
    3, 3, 15, 6, 5, 0, -2, 5, 6,
    -- filter=100 channel=44
    1, 2, -10, -4, -1, -4, -3, -1, -12,
    -- filter=100 channel=45
    0, -3, -1, 1, 1, -7, 2, -1, -8,
    -- filter=100 channel=46
    4, 0, 9, -6, -2, 0, 0, -8, 10,
    -- filter=100 channel=47
    0, -1, -4, 3, -4, -9, -4, -5, -17,
    -- filter=100 channel=48
    0, 5, -9, 8, 0, -13, 8, 7, -13,
    -- filter=100 channel=49
    3, 3, -6, -4, -2, -11, -1, -3, 0,
    -- filter=100 channel=50
    10, 4, 0, 7, 0, -15, -4, -3, -14,
    -- filter=100 channel=51
    6, -6, 5, -3, -6, 0, 3, 1, -2,
    -- filter=100 channel=52
    -11, 10, -3, -6, 10, 7, -9, -3, 1,
    -- filter=100 channel=53
    6, 0, -4, -4, 11, 1, -5, 0, 0,
    -- filter=100 channel=54
    2, -5, 7, -2, -7, 1, -4, -4, -6,
    -- filter=100 channel=55
    8, 6, 5, 4, 2, -3, -3, 5, -6,
    -- filter=100 channel=56
    -8, 4, -3, -9, -1, 0, 2, -3, 0,
    -- filter=100 channel=57
    1, -4, 8, 0, 0, 9, 2, -6, 9,
    -- filter=100 channel=58
    6, 4, -5, 6, 4, 3, 8, 3, 3,
    -- filter=100 channel=59
    8, 5, -5, -4, 5, -5, -2, -1, -9,
    -- filter=100 channel=60
    5, 4, -3, 0, 4, -3, 1, 0, 8,
    -- filter=100 channel=61
    -2, 3, -1, -8, 1, -6, -6, -2, -1,
    -- filter=100 channel=62
    -2, 6, 2, 2, -5, 0, 4, -1, -5,
    -- filter=100 channel=63
    9, 6, -6, 4, 8, -6, 9, 10, 2,
    -- filter=100 channel=64
    -6, 5, -3, 4, -1, -3, -5, 3, 5,
    -- filter=100 channel=65
    -2, -5, -6, -2, 0, -5, 5, 4, 5,
    -- filter=100 channel=66
    -5, 14, 5, -11, 8, 3, 1, 4, 15,
    -- filter=100 channel=67
    4, 4, 5, 5, -4, -1, 0, -5, -2,
    -- filter=100 channel=68
    -4, 1, -9, 1, -7, 0, -2, 1, -5,
    -- filter=100 channel=69
    1, 5, 4, -2, 8, 3, 7, 4, 7,
    -- filter=100 channel=70
    0, 3, 5, -6, 4, -7, -2, 7, -18,
    -- filter=100 channel=71
    1, 5, 3, 5, 4, -5, 0, 1, 0,
    -- filter=100 channel=72
    8, 7, -7, 3, -1, -11, -4, 3, -7,
    -- filter=100 channel=73
    -7, 0, 3, -9, 10, -9, 2, -4, -11,
    -- filter=100 channel=74
    -11, 0, 6, 0, 10, 0, -3, 11, -10,
    -- filter=100 channel=75
    3, 0, -7, 0, -3, -4, 8, 7, -11,
    -- filter=100 channel=76
    3, 6, 4, 3, 2, -4, 4, 0, 9,
    -- filter=100 channel=77
    0, 6, 0, -2, 3, 8, 0, 1, -1,
    -- filter=100 channel=78
    -5, 8, -3, 7, 5, 2, 1, 9, 6,
    -- filter=100 channel=79
    10, 7, -1, 8, 17, -23, 1, 9, -10,
    -- filter=100 channel=80
    12, 5, -4, 1, 6, -18, -3, -2, -21,
    -- filter=100 channel=81
    5, -4, -1, -5, 0, 1, 0, -5, 0,
    -- filter=100 channel=82
    3, 0, 0, 6, 2, 1, -6, -1, 6,
    -- filter=100 channel=83
    -2, -7, 1, 4, -2, -7, 10, -7, -4,
    -- filter=100 channel=84
    -9, 2, -1, 1, 9, -10, 2, 10, -2,
    -- filter=100 channel=85
    4, 0, -1, 4, 4, 0, -4, 6, 2,
    -- filter=100 channel=86
    1, 9, -4, -3, 0, -7, 6, 5, -5,
    -- filter=100 channel=87
    0, 9, 9, 2, 10, 4, -4, 4, 4,
    -- filter=100 channel=88
    0, 2, 4, -1, 2, 8, 1, -1, -5,
    -- filter=100 channel=89
    4, 0, 5, 0, 10, -10, -2, 0, -14,
    -- filter=100 channel=90
    -10, 5, 2, -10, 3, 4, -6, 1, 0,
    -- filter=100 channel=91
    2, 4, -4, -9, 3, -20, -3, 5, -13,
    -- filter=100 channel=92
    1, 1, 11, 1, 3, 10, -8, 5, 7,
    -- filter=100 channel=93
    -7, -2, -12, 3, -3, -15, 3, -2, -17,
    -- filter=100 channel=94
    -3, -7, -6, 5, -6, 0, -3, 0, 7,
    -- filter=100 channel=95
    7, 0, 5, 0, -3, 4, 5, 2, 0,
    -- filter=100 channel=96
    0, 0, -5, -6, 0, -2, 5, 1, 2,
    -- filter=100 channel=97
    5, -2, 2, 0, 4, 1, -4, 2, -4,
    -- filter=100 channel=98
    17, 5, -1, 1, 13, -13, 5, 3, -15,
    -- filter=100 channel=99
    0, 3, -4, -8, 1, -13, -2, 1, -10,
    -- filter=100 channel=100
    5, 5, 12, 3, -4, 14, -9, 7, 9,
    -- filter=100 channel=101
    -1, -6, -7, -10, -2, -5, 7, 7, 0,
    -- filter=100 channel=102
    -1, 6, 2, -5, 7, 4, -4, -3, -4,
    -- filter=100 channel=103
    0, -8, -3, -5, -9, -9, -4, -3, -22,
    -- filter=100 channel=104
    9, 3, -6, -1, 2, -13, 2, 6, -12,
    -- filter=100 channel=105
    0, 6, 0, 3, 4, 6, -5, 3, 5,
    -- filter=100 channel=106
    -4, 6, 0, -5, 6, 6, -8, 2, 14,
    -- filter=100 channel=107
    1, 4, 0, 2, 1, -10, -3, 9, 2,
    -- filter=100 channel=108
    -5, 0, 8, -3, 0, 7, 1, -2, 14,
    -- filter=100 channel=109
    8, 5, 0, 4, 10, -16, 7, 8, -19,
    -- filter=100 channel=110
    -2, 3, -1, -3, 8, -1, -3, -3, 0,
    -- filter=100 channel=111
    5, 0, 6, 2, -2, 8, -2, -5, 5,
    -- filter=100 channel=112
    9, 0, -6, 7, 2, -6, -6, 1, -9,
    -- filter=100 channel=113
    11, -1, 5, -1, -3, -7, 0, -5, -6,
    -- filter=100 channel=114
    0, 9, -14, 6, 13, -26, 17, 17, -18,
    -- filter=100 channel=115
    -2, -1, 0, 3, -1, 3, -5, -3, -7,
    -- filter=100 channel=116
    8, 4, 0, -4, 8, -14, 1, 1, 0,
    -- filter=100 channel=117
    1, -5, -7, -5, 0, -3, 0, -1, -1,
    -- filter=100 channel=118
    -2, -6, 1, -1, -7, -3, 3, 1, 6,
    -- filter=100 channel=119
    -13, 11, 10, -8, 12, 9, -8, 8, 6,
    -- filter=100 channel=120
    -9, 0, 0, -8, 13, -21, -5, -1, -27,
    -- filter=100 channel=121
    7, 0, 11, -3, 10, 9, -7, 1, 0,
    -- filter=100 channel=122
    -13, -12, -10, -10, -10, -11, -7, -8, -13,
    -- filter=100 channel=123
    -9, 0, 10, 0, 2, -2, -4, -3, 9,
    -- filter=100 channel=124
    -5, 2, 4, -9, -3, -10, 4, 6, -8,
    -- filter=100 channel=125
    9, -2, -2, 6, 4, -15, -1, 0, -8,
    -- filter=100 channel=126
    7, 3, 3, -3, 0, 1, 1, -3, 8,
    -- filter=100 channel=127
    -3, 4, 5, -3, -2, 11, 4, -5, 10,
    -- filter=101 channel=0
    -2, -9, 0, -9, -9, 1, 4, -6, 5,
    -- filter=101 channel=1
    -4, -2, 0, -2, 0, -4, 4, -4, -4,
    -- filter=101 channel=2
    1, -1, -1, -5, 3, 0, -1, 6, 7,
    -- filter=101 channel=3
    3, -4, 3, 0, 1, 3, -4, 0, 5,
    -- filter=101 channel=4
    -4, 1, 3, -9, -1, 7, -2, 3, -1,
    -- filter=101 channel=5
    -5, 6, -1, 2, -3, -3, 2, 4, -2,
    -- filter=101 channel=6
    0, 2, 4, 0, 11, 7, 6, 12, -4,
    -- filter=101 channel=7
    -6, -2, -3, -4, 6, 6, 0, 0, -5,
    -- filter=101 channel=8
    5, 3, 4, 4, -3, -2, 2, 3, 5,
    -- filter=101 channel=9
    -8, 1, 0, 0, -2, -4, -2, 4, 0,
    -- filter=101 channel=10
    -8, -6, 2, 0, -12, -4, 0, -2, -1,
    -- filter=101 channel=11
    2, 13, 1, 11, 16, 4, 0, 7, 3,
    -- filter=101 channel=12
    6, -10, 2, 6, 0, 4, 5, 1, -3,
    -- filter=101 channel=13
    -10, -11, -4, -1, -12, 2, 2, -11, -6,
    -- filter=101 channel=14
    6, -1, -3, -5, -6, -5, 1, 0, 0,
    -- filter=101 channel=15
    -10, -1, -4, 4, 4, 11, 2, 0, 5,
    -- filter=101 channel=16
    -4, -8, 5, 1, -9, 6, -5, -1, 2,
    -- filter=101 channel=17
    6, 5, -5, 1, 0, 3, -4, -1, 6,
    -- filter=101 channel=18
    -7, -3, -8, 0, 6, -2, 3, 5, -6,
    -- filter=101 channel=19
    -5, 0, 5, 6, 5, 2, 0, -5, -5,
    -- filter=101 channel=20
    8, 19, 5, 10, 21, 10, 11, 25, 14,
    -- filter=101 channel=21
    1, 0, 5, -10, -2, -8, 0, -5, -7,
    -- filter=101 channel=22
    2, 1, -7, 0, 5, -3, -4, 0, 0,
    -- filter=101 channel=23
    -4, 0, 1, -4, 1, 6, -3, 7, 6,
    -- filter=101 channel=24
    3, 0, 5, 0, 0, 4, 2, 4, 0,
    -- filter=101 channel=25
    -12, -8, -4, -8, -21, 0, -8, -12, -6,
    -- filter=101 channel=26
    7, 7, 6, 4, -5, 5, -6, -3, 3,
    -- filter=101 channel=27
    -16, -8, -4, -12, -25, 7, -7, -16, -4,
    -- filter=101 channel=28
    4, -2, -1, 3, -3, -4, 5, 0, 1,
    -- filter=101 channel=29
    7, 7, 0, 7, 30, 14, 4, 15, 2,
    -- filter=101 channel=30
    -1, 3, 0, -5, -12, 5, 3, -7, 7,
    -- filter=101 channel=31
    -13, -12, -10, -10, -16, 1, -14, -5, 3,
    -- filter=101 channel=32
    -15, -12, -2, -5, -9, 0, -2, 3, 7,
    -- filter=101 channel=33
    -14, -3, 0, -5, -20, -7, -1, -11, -7,
    -- filter=101 channel=34
    -4, 2, 4, 2, -4, 2, 3, -4, -4,
    -- filter=101 channel=35
    0, 6, 3, -3, -4, -3, -5, -3, -6,
    -- filter=101 channel=36
    5, 2, 1, 2, 1, 0, -2, 0, 4,
    -- filter=101 channel=37
    -7, -2, 3, -7, -11, -1, 5, -7, 4,
    -- filter=101 channel=38
    -2, -3, -1, -7, -7, 5, 3, -2, 0,
    -- filter=101 channel=39
    5, 2, -2, 11, 18, 8, -4, 6, 5,
    -- filter=101 channel=40
    5, -6, -6, 3, 11, 5, 6, 3, 5,
    -- filter=101 channel=41
    -9, -7, 4, -9, -13, -10, -1, -14, -9,
    -- filter=101 channel=42
    -4, 3, 6, -8, 1, -3, -6, -7, -3,
    -- filter=101 channel=43
    -2, 9, 7, 9, 7, 1, -2, 3, 9,
    -- filter=101 channel=44
    -10, -11, -1, -4, -4, 7, 0, -1, 0,
    -- filter=101 channel=45
    0, 0, 2, 0, 2, -1, -4, 10, 8,
    -- filter=101 channel=46
    0, 5, -2, -3, -7, 2, 1, -4, 0,
    -- filter=101 channel=47
    -1, -9, -1, -2, -11, -4, -6, -3, -5,
    -- filter=101 channel=48
    -11, -10, -9, -5, -18, -8, 2, -5, -4,
    -- filter=101 channel=49
    2, -2, 0, -2, -1, 10, 8, 1, 2,
    -- filter=101 channel=50
    -6, -4, 0, -1, -4, -3, -12, -1, 3,
    -- filter=101 channel=51
    0, -2, -6, -5, 0, 0, -4, -1, 3,
    -- filter=101 channel=52
    -5, 2, 0, 3, 7, 7, -4, -3, -2,
    -- filter=101 channel=53
    -1, 2, 0, 0, 9, 11, 6, 7, -1,
    -- filter=101 channel=54
    4, 6, 4, -3, 6, -5, 6, -6, -4,
    -- filter=101 channel=55
    -13, -2, 3, -7, 0, 0, -7, 1, 0,
    -- filter=101 channel=56
    0, 0, -6, 0, -2, 3, 0, 5, -1,
    -- filter=101 channel=57
    1, 0, 3, 6, -5, 3, 0, -2, 3,
    -- filter=101 channel=58
    -2, -1, -3, 5, -3, 7, 0, -4, 0,
    -- filter=101 channel=59
    -10, -11, 3, -6, -16, -8, -9, -7, -7,
    -- filter=101 channel=60
    0, -4, 7, 6, 5, 3, 1, -1, 1,
    -- filter=101 channel=61
    8, 0, 7, 4, -6, 3, 4, -5, -3,
    -- filter=101 channel=62
    -5, -5, 5, -6, -4, 4, 1, -1, 1,
    -- filter=101 channel=63
    7, 5, -4, 0, 6, -2, 3, 5, 6,
    -- filter=101 channel=64
    5, -1, 7, 3, 3, 0, 6, 1, -2,
    -- filter=101 channel=65
    1, 3, 1, 2, 3, 3, 4, -7, 6,
    -- filter=101 channel=66
    0, -5, 6, -1, -14, -6, 0, 0, -4,
    -- filter=101 channel=67
    2, 8, 0, 5, -3, 7, 0, 4, 5,
    -- filter=101 channel=68
    3, 1, -4, -4, 0, -2, -5, 6, 0,
    -- filter=101 channel=69
    -5, -6, 7, 1, -8, 6, -5, 5, -4,
    -- filter=101 channel=70
    -9, -1, -5, -3, -12, -4, -8, -11, 0,
    -- filter=101 channel=71
    0, 0, -6, -3, 5, -1, -2, -8, -2,
    -- filter=101 channel=72
    -12, -14, -7, -14, -8, -1, -3, -7, -4,
    -- filter=101 channel=73
    -12, 0, -7, 0, 6, 10, -3, 4, 6,
    -- filter=101 channel=74
    -9, -4, -2, -6, -7, 9, -9, 0, -4,
    -- filter=101 channel=75
    -4, -6, -4, -11, 0, -5, 5, -6, -5,
    -- filter=101 channel=76
    0, 7, 0, 9, 17, 17, 2, 12, 5,
    -- filter=101 channel=77
    2, -5, 1, 0, -3, -7, -4, 4, 4,
    -- filter=101 channel=78
    2, 2, -5, 4, -5, 1, 0, -3, 6,
    -- filter=101 channel=79
    -11, -9, 2, -9, -7, 0, 0, -3, -4,
    -- filter=101 channel=80
    -15, -10, 5, -12, -23, 1, -12, -7, -5,
    -- filter=101 channel=81
    -5, -5, 7, -3, -4, -7, 4, 1, 4,
    -- filter=101 channel=82
    4, 7, 0, -3, 2, -2, 6, -4, -5,
    -- filter=101 channel=83
    -6, -6, -2, 0, -9, 6, -5, -7, 0,
    -- filter=101 channel=84
    -2, -8, 0, -1, 8, 3, -1, 6, 7,
    -- filter=101 channel=85
    -4, -1, 7, -5, 6, 5, 4, 4, 7,
    -- filter=101 channel=86
    6, 1, 2, 4, -1, 9, 5, -9, 0,
    -- filter=101 channel=87
    8, -2, -2, 0, 9, 12, 8, 13, 0,
    -- filter=101 channel=88
    3, 3, 1, 2, 5, 10, -5, -3, 8,
    -- filter=101 channel=89
    -11, -10, -11, -12, -12, -1, 0, -9, -2,
    -- filter=101 channel=90
    -6, -6, -8, -6, 2, 6, -9, 4, -5,
    -- filter=101 channel=91
    -8, -12, 3, -10, -4, 8, -3, -4, -1,
    -- filter=101 channel=92
    5, 1, -4, 3, 6, 6, 6, 4, 3,
    -- filter=101 channel=93
    -8, -3, 3, 2, -12, -2, -1, -5, -6,
    -- filter=101 channel=94
    -2, -3, 4, -5, 5, -1, 0, -6, 1,
    -- filter=101 channel=95
    3, 2, 5, -5, -3, -6, 0, -8, 2,
    -- filter=101 channel=96
    -5, 0, -5, -2, 0, -2, 1, 2, 0,
    -- filter=101 channel=97
    -5, 0, 5, 2, -2, -8, 1, 0, -4,
    -- filter=101 channel=98
    -10, -2, -3, -14, -16, -10, 0, -1, -2,
    -- filter=101 channel=99
    -5, -10, -4, 1, -1, 0, -8, 4, 9,
    -- filter=101 channel=100
    1, -6, 1, -4, -2, -9, -1, 3, -2,
    -- filter=101 channel=101
    6, -7, 4, -7, 9, 11, -6, 7, 1,
    -- filter=101 channel=102
    -3, 5, -3, -2, -6, -7, 3, 0, -7,
    -- filter=101 channel=103
    -6, -6, -6, -8, -10, -6, 0, -7, -5,
    -- filter=101 channel=104
    0, -2, 0, -13, -10, -6, -3, -14, 0,
    -- filter=101 channel=105
    2, 15, 0, 12, 25, 7, 5, 7, 3,
    -- filter=101 channel=106
    7, 0, -2, 6, 2, 3, -1, 5, -1,
    -- filter=101 channel=107
    3, 3, 1, 12, 11, 14, 7, 10, 2,
    -- filter=101 channel=108
    3, 0, -3, 0, 3, 6, 8, 1, 5,
    -- filter=101 channel=109
    -4, -11, 3, -9, -9, 2, -8, -6, -7,
    -- filter=101 channel=110
    -10, -5, -7, -4, 0, 1, -5, 1, 6,
    -- filter=101 channel=111
    -7, -2, 6, 6, 0, 0, 0, -7, -1,
    -- filter=101 channel=112
    -7, 3, 3, -2, -13, -1, -7, -5, -2,
    -- filter=101 channel=113
    -2, -11, 2, -2, -9, 4, -2, -9, -1,
    -- filter=101 channel=114
    -14, -4, -3, -2, -2, 11, 1, 7, 9,
    -- filter=101 channel=115
    5, 0, 5, 3, -6, 7, 0, 4, 5,
    -- filter=101 channel=116
    -12, -8, -7, -1, -5, 2, 0, -7, 3,
    -- filter=101 channel=117
    -5, -5, 5, -4, -2, 4, -2, -8, 3,
    -- filter=101 channel=118
    -6, -3, 6, -5, 2, -5, 2, 2, 0,
    -- filter=101 channel=119
    0, 4, -2, -1, 4, 3, 0, -5, 7,
    -- filter=101 channel=120
    -1, -2, 4, 2, 2, 5, -7, 1, 7,
    -- filter=101 channel=121
    -8, -3, -5, -10, -15, 0, -2, -12, -3,
    -- filter=101 channel=122
    -2, -9, -5, -12, -14, -1, -8, -5, -8,
    -- filter=101 channel=123
    4, -6, -7, 2, -6, 0, -7, -7, -5,
    -- filter=101 channel=124
    6, 14, 2, 12, 18, 9, 8, 14, 3,
    -- filter=101 channel=125
    -12, -4, -9, -11, -5, -5, -8, -14, 1,
    -- filter=101 channel=126
    -6, -1, 4, -3, -6, 0, 0, -9, 0,
    -- filter=101 channel=127
    -3, 0, -5, -2, -4, 5, 0, -5, -4,
    -- filter=102 channel=0
    14, -1, -7, 14, 8, 2, -4, 4, 4,
    -- filter=102 channel=1
    0, 0, -2, 3, -2, -14, -13, 0, -7,
    -- filter=102 channel=2
    -6, -9, -4, -6, -3, -11, -4, -7, -2,
    -- filter=102 channel=3
    11, 5, 10, 5, 4, 4, 5, 5, 0,
    -- filter=102 channel=4
    0, -7, -5, -13, -20, -16, -16, -17, -27,
    -- filter=102 channel=5
    4, -2, 4, 4, 12, 12, 6, 16, 10,
    -- filter=102 channel=6
    -3, 3, 5, -8, 1, 5, 0, 0, 10,
    -- filter=102 channel=7
    -7, -4, 2, 4, 1, -2, -2, 0, 4,
    -- filter=102 channel=8
    -4, -1, 1, -9, -5, 0, -5, -11, -1,
    -- filter=102 channel=9
    8, 5, -5, 3, 0, 9, -4, 3, -4,
    -- filter=102 channel=10
    9, 13, -1, 5, 4, 7, -1, -5, -9,
    -- filter=102 channel=11
    0, -3, 11, 0, 0, 19, 11, 4, 11,
    -- filter=102 channel=12
    -13, 3, -7, -10, -6, -1, 2, -6, -1,
    -- filter=102 channel=13
    4, 11, 1, -4, -4, -4, 1, -9, -10,
    -- filter=102 channel=14
    0, 0, -6, 0, 0, -3, -5, -2, -5,
    -- filter=102 channel=15
    13, 12, 12, -11, -7, 15, -7, -12, -7,
    -- filter=102 channel=16
    -8, -2, -8, -1, 0, 0, 4, 11, -3,
    -- filter=102 channel=17
    -1, -4, 4, 1, 1, -5, -5, 1, -3,
    -- filter=102 channel=18
    20, 17, 5, -2, 2, 14, -6, -12, -12,
    -- filter=102 channel=19
    -4, 3, 5, -2, 0, -1, 3, 3, 4,
    -- filter=102 channel=20
    -2, 2, 11, -11, -3, 24, 10, 4, 15,
    -- filter=102 channel=21
    -3, -4, -4, -1, -1, -1, -3, 9, 0,
    -- filter=102 channel=22
    5, 2, -1, 0, -7, 6, 0, -4, 2,
    -- filter=102 channel=23
    15, 10, 7, -14, -6, 17, -3, -14, 0,
    -- filter=102 channel=24
    0, -3, 2, -4, -2, -4, -2, 1, -4,
    -- filter=102 channel=25
    5, 0, 0, 5, 0, -10, -3, -11, -11,
    -- filter=102 channel=26
    -7, -4, -5, 8, 0, -7, 8, 4, 5,
    -- filter=102 channel=27
    9, 9, 5, -8, 0, 11, -9, -20, -20,
    -- filter=102 channel=28
    -2, 2, -1, -5, -5, -4, -3, -1, -5,
    -- filter=102 channel=29
    9, 2, 14, -7, 3, 24, 10, 1, 11,
    -- filter=102 channel=30
    0, 1, 0, -5, 6, -2, -11, -5, -9,
    -- filter=102 channel=31
    3, 7, 7, -7, 8, -2, -4, 1, -12,
    -- filter=102 channel=32
    0, 17, 12, -3, -4, 11, -12, -21, -8,
    -- filter=102 channel=33
    24, 11, 13, 1, 1, 3, 2, -10, -10,
    -- filter=102 channel=34
    -14, -3, -6, -3, 0, 6, -11, -5, -3,
    -- filter=102 channel=35
    0, 1, -3, 1, 6, 5, 0, 5, 3,
    -- filter=102 channel=36
    -4, -4, -5, -8, -12, -6, 6, -3, -3,
    -- filter=102 channel=37
    4, -8, -16, 7, 9, -15, -14, -2, -5,
    -- filter=102 channel=38
    11, 14, -1, 5, 0, 0, 7, -8, -5,
    -- filter=102 channel=39
    -7, -1, 0, -3, -7, 3, 0, -2, 6,
    -- filter=102 channel=40
    6, 8, 2, -10, -8, 8, -1, -7, -2,
    -- filter=102 channel=41
    -10, -2, 1, 4, -4, -9, -5, 7, -14,
    -- filter=102 channel=42
    6, 5, 7, 7, 3, 0, 0, 1, -6,
    -- filter=102 channel=43
    9, 5, 2, 3, -6, 6, 6, 2, 11,
    -- filter=102 channel=44
    -2, -2, 0, 0, 5, -5, -9, -3, -13,
    -- filter=102 channel=45
    5, -1, 7, 6, 8, -2, 6, 0, 0,
    -- filter=102 channel=46
    6, 4, -2, 0, -2, -8, 2, 6, -5,
    -- filter=102 channel=47
    0, 1, -7, 14, 2, -4, 5, 4, 3,
    -- filter=102 channel=48
    1, -3, -8, 10, -3, -10, -4, -6, -21,
    -- filter=102 channel=49
    4, -6, 1, -4, -3, -5, -11, -12, -7,
    -- filter=102 channel=50
    1, 2, 1, -3, 3, 1, 3, -9, -15,
    -- filter=102 channel=51
    3, -1, 4, 5, 7, -5, 0, 5, -6,
    -- filter=102 channel=52
    2, -2, -7, -5, -5, 5, -1, -12, 4,
    -- filter=102 channel=53
    2, -1, 7, -9, -2, 12, 1, 4, 3,
    -- filter=102 channel=54
    6, 4, -3, 1, 4, 0, 1, -5, -5,
    -- filter=102 channel=55
    14, 6, 16, -11, -4, 17, 0, -13, -8,
    -- filter=102 channel=56
    -5, -8, 0, -7, -10, -3, -6, -2, -1,
    -- filter=102 channel=57
    -6, 1, 4, -1, -4, -10, -1, -3, -4,
    -- filter=102 channel=58
    2, 0, -3, 0, 4, 4, 2, 3, 3,
    -- filter=102 channel=59
    3, 5, 4, 2, -2, -1, 2, -12, -11,
    -- filter=102 channel=60
    6, 5, 7, 2, 7, 5, -1, -1, 6,
    -- filter=102 channel=61
    -4, -10, -6, -3, -3, -2, 3, -6, 6,
    -- filter=102 channel=62
    3, 4, 0, 0, 6, -4, -1, 3, -6,
    -- filter=102 channel=63
    1, 5, 6, 6, 11, 10, 7, 4, 10,
    -- filter=102 channel=64
    -6, -1, 0, 5, 0, 4, 8, 0, -5,
    -- filter=102 channel=65
    7, -6, -4, 3, 1, 6, 1, -4, -1,
    -- filter=102 channel=66
    -13, 2, 0, -8, 0, -1, -5, -1, -4,
    -- filter=102 channel=67
    0, 3, 7, 4, 2, 5, 1, 7, -2,
    -- filter=102 channel=68
    -4, 0, -7, -7, -6, 0, 7, -6, -1,
    -- filter=102 channel=69
    -3, 6, 4, 4, 1, 4, 5, 4, -3,
    -- filter=102 channel=70
    7, 12, -1, -12, -3, -4, -12, -16, -12,
    -- filter=102 channel=71
    9, 3, 3, 6, 0, 5, -4, 5, 5,
    -- filter=102 channel=72
    0, 1, 0, -2, -4, 3, -4, -1, -6,
    -- filter=102 channel=73
    -6, 6, 1, -7, -5, 3, -5, -11, -12,
    -- filter=102 channel=74
    0, 2, -2, -10, 3, 3, -10, -2, -5,
    -- filter=102 channel=75
    14, 11, 0, 15, 9, 6, -6, -2, 0,
    -- filter=102 channel=76
    7, -3, 15, 0, -4, 14, 15, 8, 6,
    -- filter=102 channel=77
    -4, 4, -2, 0, -2, -2, 6, -4, 2,
    -- filter=102 channel=78
    1, 3, 4, 6, 7, 12, 1, 0, 7,
    -- filter=102 channel=79
    25, 13, 16, -1, 3, 15, -6, -27, -13,
    -- filter=102 channel=80
    4, 9, 2, 12, 11, 6, -3, 2, -5,
    -- filter=102 channel=81
    -5, -1, 0, 2, 0, -6, 5, -5, 1,
    -- filter=102 channel=82
    7, 5, 1, -5, 1, 4, -1, 8, 6,
    -- filter=102 channel=83
    0, 0, 9, 0, 0, -1, -5, -11, -3,
    -- filter=102 channel=84
    -3, 6, 7, -6, -6, 0, -13, -15, -16,
    -- filter=102 channel=85
    -2, -2, -3, -6, -5, -6, 7, 7, -3,
    -- filter=102 channel=86
    -2, -4, -7, 0, 1, -1, 0, -2, 7,
    -- filter=102 channel=87
    -3, -11, -2, -12, 0, 2, 2, -6, -1,
    -- filter=102 channel=88
    -6, -1, 0, -11, -3, -11, -3, -4, 2,
    -- filter=102 channel=89
    13, 16, 3, -1, -3, -1, 0, -9, -7,
    -- filter=102 channel=90
    -7, -10, -1, -12, -9, -5, 1, -2, 2,
    -- filter=102 channel=91
    -4, 0, 3, -8, -4, 1, -19, -24, -22,
    -- filter=102 channel=92
    6, -1, 8, -4, 3, 1, -7, -7, 2,
    -- filter=102 channel=93
    -10, -6, -3, 11, -3, -12, -7, -3, -11,
    -- filter=102 channel=94
    0, -7, -3, -3, 3, -6, -6, 1, 0,
    -- filter=102 channel=95
    -3, 4, 0, 4, -4, 0, 6, -2, 2,
    -- filter=102 channel=96
    -3, 4, -4, 8, 2, -2, 7, -4, 2,
    -- filter=102 channel=97
    18, 4, 7, 4, 0, -4, 4, 10, -2,
    -- filter=102 channel=98
    14, 12, 6, 1, 0, 6, 5, -12, -11,
    -- filter=102 channel=99
    3, 4, 9, -10, -5, 15, -6, -16, 0,
    -- filter=102 channel=100
    -1, -6, 5, 3, -5, 6, -6, -4, -8,
    -- filter=102 channel=101
    2, -6, 0, -12, -15, -10, 0, -3, -5,
    -- filter=102 channel=102
    0, 1, -1, -7, 3, -1, 2, -4, 0,
    -- filter=102 channel=103
    10, 0, -7, 10, 14, 4, -3, 5, -1,
    -- filter=102 channel=104
    -1, 10, 2, -4, 0, 2, -2, -6, -14,
    -- filter=102 channel=105
    9, 0, 2, -5, 1, 15, 2, 8, 11,
    -- filter=102 channel=106
    -2, 0, 2, 1, -8, 5, 11, 7, -2,
    -- filter=102 channel=107
    2, 5, 10, -16, -11, 6, -11, -14, 11,
    -- filter=102 channel=108
    -2, 3, -4, -2, 1, 7, 1, 3, 2,
    -- filter=102 channel=109
    4, 14, 3, 3, -4, 7, -7, -19, -11,
    -- filter=102 channel=110
    4, 5, 6, 4, 3, 1, -2, 1, 2,
    -- filter=102 channel=111
    -4, 5, 3, -1, -3, 0, 1, -5, 0,
    -- filter=102 channel=112
    8, 0, 0, -9, 8, 6, 1, -9, -7,
    -- filter=102 channel=113
    15, 11, 9, -3, 0, 3, 2, -1, -7,
    -- filter=102 channel=114
    8, 4, 6, 0, -7, 12, -5, -23, -13,
    -- filter=102 channel=115
    0, -5, -3, -6, 2, 0, 1, 0, -4,
    -- filter=102 channel=116
    0, 2, 1, -7, 1, -6, -6, -5, -11,
    -- filter=102 channel=117
    -5, 0, -7, 1, 0, -3, -8, 0, -7,
    -- filter=102 channel=118
    5, 0, -3, 1, -5, 1, -6, 0, -1,
    -- filter=102 channel=119
    -12, -8, -3, -1, -10, -6, -10, -12, -7,
    -- filter=102 channel=120
    -1, 0, 14, -14, -7, 11, -9, -19, -24,
    -- filter=102 channel=121
    -1, 7, 4, -1, -1, -1, 0, 0, 0,
    -- filter=102 channel=122
    -19, -8, -13, 7, 4, -15, -7, 2, -5,
    -- filter=102 channel=123
    -2, -4, 5, -7, -3, 1, -10, -8, -1,
    -- filter=102 channel=124
    3, 4, 8, -4, 4, 11, 9, 5, 8,
    -- filter=102 channel=125
    0, 3, 0, -5, -7, 8, -5, -11, -8,
    -- filter=102 channel=126
    21, 7, 7, 7, -3, 6, 6, 0, 1,
    -- filter=102 channel=127
    -4, 1, -4, 1, 7, -9, 6, -2, -1,
    -- filter=103 channel=0
    -22, -2, 7, -31, 7, 21, -25, 3, 20,
    -- filter=103 channel=1
    -31, -4, 8, -24, 10, 25, -11, 4, 7,
    -- filter=103 channel=2
    5, 0, 0, 1, 7, -5, 7, 0, -6,
    -- filter=103 channel=3
    -5, -4, -3, -7, -6, -5, -3, -7, 3,
    -- filter=103 channel=4
    0, -7, 3, -7, 5, 8, 9, 5, 5,
    -- filter=103 channel=5
    -24, -9, 11, -20, 5, 25, -5, 10, 17,
    -- filter=103 channel=6
    9, 4, 1, 2, 8, 4, 2, -4, 1,
    -- filter=103 channel=7
    0, 1, 4, 7, -6, -2, 0, 1, 2,
    -- filter=103 channel=8
    2, 3, 0, -4, 2, 5, 7, -8, 0,
    -- filter=103 channel=9
    3, 0, 10, -10, -2, 8, 1, 8, 8,
    -- filter=103 channel=10
    9, -3, -4, -7, -2, -10, 2, -5, 0,
    -- filter=103 channel=11
    18, 4, -5, 9, 0, -8, 7, -7, -9,
    -- filter=103 channel=12
    0, -3, -6, 1, 2, -7, 6, 1, 2,
    -- filter=103 channel=13
    -1, -5, -10, 6, -5, -7, -6, 0, -2,
    -- filter=103 channel=14
    4, -4, -4, 4, 5, -6, -5, 7, -7,
    -- filter=103 channel=15
    2, 16, -2, 2, 9, -8, -12, -9, -8,
    -- filter=103 channel=16
    -11, -16, 5, -5, -1, 11, -2, 10, 3,
    -- filter=103 channel=17
    0, -6, -3, -2, -2, -4, 2, 0, -4,
    -- filter=103 channel=18
    -2, 16, -5, -4, 2, -3, -19, 0, -14,
    -- filter=103 channel=19
    -2, -2, 0, 1, 0, 7, 7, 3, 4,
    -- filter=103 channel=20
    10, 28, 0, 14, -3, -15, -4, -11, -18,
    -- filter=103 channel=21
    3, -12, -2, -11, -11, 8, 12, 5, 6,
    -- filter=103 channel=22
    -8, 8, 3, -2, 9, 5, 1, 4, 3,
    -- filter=103 channel=23
    12, 3, -7, 6, -5, -16, -4, 0, -16,
    -- filter=103 channel=24
    -1, 0, 2, 3, -1, 7, 6, -5, 3,
    -- filter=103 channel=25
    -14, 4, 2, -9, 1, 8, -2, 3, 11,
    -- filter=103 channel=26
    -11, -7, 7, -1, 0, 7, 0, 7, 3,
    -- filter=103 channel=27
    -18, 12, 2, -16, 5, 4, -9, 17, 10,
    -- filter=103 channel=28
    -1, -4, -5, 7, -2, -7, 5, -5, 4,
    -- filter=103 channel=29
    20, 28, 5, 17, -2, -22, 2, -17, -18,
    -- filter=103 channel=30
    -17, 1, 11, -20, -5, 19, -1, 3, 1,
    -- filter=103 channel=31
    4, -16, -9, -4, -19, 6, 11, -2, 12,
    -- filter=103 channel=32
    -2, 4, -4, -1, 4, 3, -1, 5, -1,
    -- filter=103 channel=33
    -5, -8, -1, -10, 6, -2, -6, 5, 8,
    -- filter=103 channel=34
    -1, -2, 3, -1, 0, 12, 0, 5, 9,
    -- filter=103 channel=35
    -4, 0, 7, -6, 0, 6, 2, -6, 1,
    -- filter=103 channel=36
    0, -7, -1, 12, -6, -12, -1, -2, -2,
    -- filter=103 channel=37
    -27, -7, 15, -35, 0, 32, -16, 12, 23,
    -- filter=103 channel=38
    4, -2, 3, -5, -3, 4, -7, 1, -2,
    -- filter=103 channel=39
    9, 4, -8, 9, 6, -8, -6, 1, -15,
    -- filter=103 channel=40
    6, 2, -5, 10, 4, -3, -3, 0, -11,
    -- filter=103 channel=41
    -10, -3, -5, -18, -10, -4, -9, -7, -7,
    -- filter=103 channel=42
    -11, -9, 9, -1, 0, 9, -1, 2, 9,
    -- filter=103 channel=43
    -7, 9, -2, 0, 1, -7, -6, 2, -1,
    -- filter=103 channel=44
    -8, -18, 9, -10, -7, 22, 0, 10, 13,
    -- filter=103 channel=45
    4, -4, 4, 3, 4, 5, 0, 2, 7,
    -- filter=103 channel=46
    -4, 0, -1, 2, 7, -1, -5, 5, -4,
    -- filter=103 channel=47
    -14, -13, 1, -13, -2, 22, -5, 7, 18,
    -- filter=103 channel=48
    -15, -13, 2, -5, 2, 15, -1, 18, 7,
    -- filter=103 channel=49
    4, 5, -3, 1, 5, -13, -6, -6, -11,
    -- filter=103 channel=50
    -5, -7, 7, -7, -7, 6, -6, 7, 2,
    -- filter=103 channel=51
    5, 7, -5, 0, -6, 6, -1, 7, 5,
    -- filter=103 channel=52
    -5, 1, 0, -1, 5, -3, 6, -8, -2,
    -- filter=103 channel=53
    0, 11, 5, 0, 4, -4, 7, -6, -4,
    -- filter=103 channel=54
    0, 0, 7, -4, 5, -5, -1, 1, 1,
    -- filter=103 channel=55
    4, 15, -3, 8, 9, -25, -2, -7, -15,
    -- filter=103 channel=56
    -1, 0, -4, -1, 5, -5, 7, -4, 3,
    -- filter=103 channel=57
    -3, -8, 4, -1, -3, -3, -7, 0, -5,
    -- filter=103 channel=58
    -7, -5, 4, -13, 3, 16, -8, -1, 6,
    -- filter=103 channel=59
    -8, -9, 2, -8, -4, 9, 1, 6, 12,
    -- filter=103 channel=60
    6, -5, 3, 6, -2, -4, -2, 3, 6,
    -- filter=103 channel=61
    8, 0, 4, 9, -6, -1, 4, 4, 1,
    -- filter=103 channel=62
    2, -6, -2, 0, 6, -5, 4, 3, -8,
    -- filter=103 channel=63
    -4, -7, 11, -10, -5, 11, 3, 7, 11,
    -- filter=103 channel=64
    10, 6, 0, -3, -6, -2, -1, -10, 0,
    -- filter=103 channel=65
    7, 0, 2, -2, -7, -3, -2, -6, -3,
    -- filter=103 channel=66
    -1, -4, 5, 4, -5, 0, 3, -8, -3,
    -- filter=103 channel=67
    4, 5, 5, -2, 1, -1, 6, -2, -3,
    -- filter=103 channel=68
    2, -4, -3, 0, 0, -4, -4, -1, 0,
    -- filter=103 channel=69
    -5, -7, 5, -5, 0, 5, 1, -6, 0,
    -- filter=103 channel=70
    -3, -5, -3, -10, 8, -2, -3, 6, -6,
    -- filter=103 channel=71
    5, -4, -10, -4, 1, -10, -4, -9, -3,
    -- filter=103 channel=72
    5, -10, 4, 0, -12, 0, 7, -1, 1,
    -- filter=103 channel=73
    3, 0, -4, 5, 2, 0, 4, -3, -10,
    -- filter=103 channel=74
    -10, -4, 7, -8, 7, 4, -2, -3, 0,
    -- filter=103 channel=75
    -16, -11, 14, -26, -6, 34, -12, 13, 20,
    -- filter=103 channel=76
    19, 15, -9, 20, 5, -27, 0, -7, -26,
    -- filter=103 channel=77
    -6, -1, 2, -4, 1, 5, -7, -7, 3,
    -- filter=103 channel=78
    -6, 1, 1, -2, -2, 11, -4, 6, 8,
    -- filter=103 channel=79
    -12, 6, -9, -13, 11, -7, -18, -2, -8,
    -- filter=103 channel=80
    3, -10, 5, -10, -18, 5, 9, 6, 8,
    -- filter=103 channel=81
    5, -4, -4, 0, 6, -7, 2, 5, 0,
    -- filter=103 channel=82
    5, 6, 0, -2, 3, -1, -5, -6, 6,
    -- filter=103 channel=83
    -6, -1, 0, 0, 6, 1, 0, 8, 0,
    -- filter=103 channel=84
    1, 0, 6, -2, 11, 3, -9, 4, 1,
    -- filter=103 channel=85
    1, -6, 2, 6, 5, 1, 0, 4, 6,
    -- filter=103 channel=86
    2, -4, 6, -5, -6, 11, 0, 4, 0,
    -- filter=103 channel=87
    9, 9, -5, 13, 4, -7, 3, 3, -12,
    -- filter=103 channel=88
    11, 2, 0, 0, -4, -14, -2, 3, 0,
    -- filter=103 channel=89
    -1, 1, -10, 0, -6, -18, 4, 1, -7,
    -- filter=103 channel=90
    4, -6, -6, 7, -12, -13, 10, 1, -8,
    -- filter=103 channel=91
    5, 12, -5, 6, -2, 2, 7, -2, -5,
    -- filter=103 channel=92
    -2, 2, 2, 5, 0, -1, -1, 4, 0,
    -- filter=103 channel=93
    -9, -12, 3, -12, 4, 16, -6, 14, 18,
    -- filter=103 channel=94
    -4, -1, -6, 1, -2, 4, 4, 1, 4,
    -- filter=103 channel=95
    -3, -8, -2, 4, 0, 6, 4, -8, 0,
    -- filter=103 channel=96
    2, 4, 3, -9, -2, 5, -5, -5, 0,
    -- filter=103 channel=97
    -1, 1, -5, -10, -1, 5, -1, 0, 0,
    -- filter=103 channel=98
    -10, -6, -6, -3, -9, 10, -5, 3, 4,
    -- filter=103 channel=99
    10, 5, -7, 5, 2, -11, 14, -3, -11,
    -- filter=103 channel=100
    0, -3, 0, -6, 6, -7, 0, -7, -2,
    -- filter=103 channel=101
    5, 0, 3, 7, -3, -5, -4, 0, 6,
    -- filter=103 channel=102
    3, -4, 0, 7, 1, 3, 3, -7, 3,
    -- filter=103 channel=103
    -8, -4, -2, -21, -9, 23, 2, 3, 11,
    -- filter=103 channel=104
    6, -7, 2, -2, -6, 4, 6, 9, 1,
    -- filter=103 channel=105
    12, 19, -6, 14, 0, -8, -4, -11, -17,
    -- filter=103 channel=106
    9, 1, 0, 2, 5, -1, -5, -5, -4,
    -- filter=103 channel=107
    0, 19, -6, 8, 14, 1, -2, 0, -11,
    -- filter=103 channel=108
    -5, 2, 7, -12, -3, 1, 0, 0, -5,
    -- filter=103 channel=109
    -15, 14, 3, -6, 11, 1, 2, 12, 3,
    -- filter=103 channel=110
    0, 0, -4, 7, -13, 2, -1, 0, 5,
    -- filter=103 channel=111
    -4, 0, 5, 3, -4, -5, 0, -7, -6,
    -- filter=103 channel=112
    -10, -4, 1, -9, 0, 4, 2, 5, 8,
    -- filter=103 channel=113
    -3, -9, -10, -9, -5, 0, -8, -3, 7,
    -- filter=103 channel=114
    -24, 6, 16, -11, 21, 15, -19, 4, 3,
    -- filter=103 channel=115
    -4, 3, 6, 2, 1, 5, 0, -1, -1,
    -- filter=103 channel=116
    3, 0, -5, 4, 0, -9, 0, 6, -3,
    -- filter=103 channel=117
    -1, 0, -6, 7, -4, 0, 8, -7, 0,
    -- filter=103 channel=118
    1, -1, 3, 6, -5, -7, -6, 4, -6,
    -- filter=103 channel=119
    -4, 2, 0, 2, 3, -2, -4, -2, 11,
    -- filter=103 channel=120
    4, 8, 4, 8, 8, -5, -4, 3, 2,
    -- filter=103 channel=121
    0, -10, -5, -3, -8, -1, 1, 0, 5,
    -- filter=103 channel=122
    -15, -26, 6, -11, -4, 20, 2, 8, 15,
    -- filter=103 channel=123
    -5, 1, -6, 4, -2, 3, -8, 3, 7,
    -- filter=103 channel=124
    1, 15, -5, 7, 5, -1, -2, -9, -13,
    -- filter=103 channel=125
    2, -2, 6, 0, -5, -5, 6, 3, 9,
    -- filter=103 channel=126
    0, -5, 0, -6, -2, 3, -10, -12, -2,
    -- filter=103 channel=127
    0, 0, 4, 0, 3, 7, 1, 0, 5,
    -- filter=104 channel=0
    -3, -3, 5, 6, 0, 4, 1, 14, 0,
    -- filter=104 channel=1
    -2, -5, 5, 5, -5, 5, 0, 2, 2,
    -- filter=104 channel=2
    -2, -3, 0, -2, -7, -6, -5, -3, 3,
    -- filter=104 channel=3
    3, 4, 5, 0, 9, 6, 7, 4, -3,
    -- filter=104 channel=4
    6, 8, -3, -3, -4, 2, 0, -7, -4,
    -- filter=104 channel=5
    -5, 4, 0, -3, 7, 2, 6, 1, 6,
    -- filter=104 channel=6
    4, -5, 3, -1, -4, 3, 6, 7, 1,
    -- filter=104 channel=7
    2, -6, 0, -6, -4, -5, -1, -3, 2,
    -- filter=104 channel=8
    5, -2, 0, 4, -3, 6, 5, -8, 0,
    -- filter=104 channel=9
    -4, 0, 0, 3, -3, 5, -2, -7, 0,
    -- filter=104 channel=10
    12, 8, -3, 0, -4, -10, 1, -9, -4,
    -- filter=104 channel=11
    0, 1, 4, 2, 1, 6, -1, -4, 6,
    -- filter=104 channel=12
    0, -4, -2, -1, -4, -4, -4, 5, -4,
    -- filter=104 channel=13
    8, 0, 3, 1, 0, -1, 4, 0, -6,
    -- filter=104 channel=14
    0, 4, 5, -6, 7, 0, -5, 4, 0,
    -- filter=104 channel=15
    -1, -2, 3, 0, 2, -7, 4, 0, 0,
    -- filter=104 channel=16
    -5, -1, -1, -7, -2, 6, 0, -4, -1,
    -- filter=104 channel=17
    1, 1, 3, 3, 5, -6, 1, -4, -5,
    -- filter=104 channel=18
    11, 9, -6, 8, -1, -9, 5, -7, -15,
    -- filter=104 channel=19
    3, -2, -5, -2, 0, 5, -6, 0, 6,
    -- filter=104 channel=20
    -6, 5, 3, 13, 2, -4, 2, 6, 9,
    -- filter=104 channel=21
    -4, -4, 6, -8, -12, -2, -9, -7, -10,
    -- filter=104 channel=22
    4, -8, 8, 0, -3, 9, 4, 5, 2,
    -- filter=104 channel=23
    12, 6, -1, 2, -13, -1, -3, -14, -7,
    -- filter=104 channel=24
    -6, -2, -1, 5, -1, 5, 3, -3, 1,
    -- filter=104 channel=25
    1, -5, -3, 3, -4, -7, 0, -12, -12,
    -- filter=104 channel=26
    -1, -1, 1, -1, -2, 1, -2, -6, 1,
    -- filter=104 channel=27
    1, -9, -6, 9, -9, -3, -5, -28, -15,
    -- filter=104 channel=28
    -6, -7, 3, 2, -6, -4, 0, 2, -6,
    -- filter=104 channel=29
    -4, -2, 0, 1, 0, -8, 7, -2, -3,
    -- filter=104 channel=30
    5, 4, 1, -7, -4, 8, -3, 1, -7,
    -- filter=104 channel=31
    1, -1, 7, 6, -9, 4, 0, -12, -2,
    -- filter=104 channel=32
    4, 8, -9, 14, -5, -10, 3, -8, -13,
    -- filter=104 channel=33
    10, 0, -2, 0, 4, -4, 2, 0, -10,
    -- filter=104 channel=34
    -3, 0, -2, -5, -4, 5, -1, -5, 0,
    -- filter=104 channel=35
    -6, 7, -7, 0, 2, 4, -3, -6, -4,
    -- filter=104 channel=36
    -3, 4, 6, 1, -3, 0, 0, -8, -1,
    -- filter=104 channel=37
    1, -9, 9, 0, -5, 6, -2, 2, 8,
    -- filter=104 channel=38
    7, 3, 5, 8, -9, -5, -4, -11, -2,
    -- filter=104 channel=39
    4, -3, 1, 3, -6, -4, 6, 0, 2,
    -- filter=104 channel=40
    4, -1, 6, -3, 1, 6, 0, 6, 0,
    -- filter=104 channel=41
    3, 4, -5, 16, 9, -2, 13, 5, -15,
    -- filter=104 channel=42
    1, -7, 0, -5, 4, -5, 3, -6, -5,
    -- filter=104 channel=43
    -4, 7, 0, 5, 0, 1, 0, 7, 8,
    -- filter=104 channel=44
    -2, 0, 3, -10, 0, 3, -2, -13, 1,
    -- filter=104 channel=45
    -6, -2, 5, -2, -1, -5, -4, 6, -2,
    -- filter=104 channel=46
    4, 5, 1, 4, 6, -6, -2, 0, 6,
    -- filter=104 channel=47
    0, -5, -3, -13, -1, 0, -6, -17, -9,
    -- filter=104 channel=48
    -3, 1, -5, -2, -1, -2, -12, -14, -7,
    -- filter=104 channel=49
    -5, 3, 2, 0, -1, -12, -5, -3, -9,
    -- filter=104 channel=50
    3, -6, 3, -2, -13, -7, 1, -16, -4,
    -- filter=104 channel=51
    -2, -1, -2, -5, -1, -7, 3, -4, -6,
    -- filter=104 channel=52
    0, -7, -6, 7, -2, 4, 4, 0, 7,
    -- filter=104 channel=53
    2, 0, -5, 5, 7, 1, 5, 4, 3,
    -- filter=104 channel=54
    6, -6, 6, 1, 2, 6, 1, 0, 7,
    -- filter=104 channel=55
    0, 7, 0, 14, -2, -2, 0, -9, -5,
    -- filter=104 channel=56
    0, 2, 6, -6, -2, -4, 7, 0, -5,
    -- filter=104 channel=57
    0, -1, -5, 1, -1, 5, 0, 1, 0,
    -- filter=104 channel=58
    1, 0, 5, 1, 6, 11, 3, 3, 5,
    -- filter=104 channel=59
    -1, -6, 0, -1, -2, -9, -4, -13, -4,
    -- filter=104 channel=60
    1, -1, 2, -1, -5, -2, -5, -5, 1,
    -- filter=104 channel=61
    -1, 1, -1, -4, 0, 7, -3, 0, -4,
    -- filter=104 channel=62
    -3, 3, -5, -2, -3, 3, 2, 4, 0,
    -- filter=104 channel=63
    -2, -4, 2, -2, 1, 11, 8, 2, -1,
    -- filter=104 channel=64
    6, -5, 2, -3, -4, -7, 0, 5, -3,
    -- filter=104 channel=65
    -4, -6, -3, -1, 1, -5, -3, 2, 7,
    -- filter=104 channel=66
    -1, -2, -8, -1, 6, -9, 9, -1, -4,
    -- filter=104 channel=67
    1, 0, -4, -4, 0, -5, 4, -5, -2,
    -- filter=104 channel=68
    7, -2, -6, -7, 6, -3, 0, -5, 4,
    -- filter=104 channel=69
    6, 7, 0, -1, -5, 6, 1, -1, 6,
    -- filter=104 channel=70
    0, 5, 6, 4, -6, 2, -5, -11, -2,
    -- filter=104 channel=71
    -3, 4, 3, 5, -1, -1, 6, -4, 1,
    -- filter=104 channel=72
    4, -2, -2, 4, -1, 0, -9, -14, -13,
    -- filter=104 channel=73
    3, -5, -3, 4, 1, -8, 0, -10, -6,
    -- filter=104 channel=74
    6, 3, 1, 0, -4, 10, -9, -14, 0,
    -- filter=104 channel=75
    7, -6, 6, 7, 9, 0, 9, -1, 6,
    -- filter=104 channel=76
    6, 11, -9, 14, 8, -10, 4, -1, 0,
    -- filter=104 channel=77
    6, 3, 1, -1, 0, 7, 3, -2, -1,
    -- filter=104 channel=78
    0, 6, 7, 1, 3, 10, -5, -4, 0,
    -- filter=104 channel=79
    14, 6, -5, 17, -3, -10, 0, -5, -7,
    -- filter=104 channel=80
    3, 0, 6, 7, -8, -5, -4, -15, -15,
    -- filter=104 channel=81
    5, 2, -6, 6, 6, 6, -3, 6, 0,
    -- filter=104 channel=82
    -6, -3, 0, 2, 1, -4, 3, -1, 8,
    -- filter=104 channel=83
    2, 1, 2, 4, -1, 2, 1, -4, -8,
    -- filter=104 channel=84
    2, -2, -9, 9, 1, -6, -5, -10, -5,
    -- filter=104 channel=85
    0, 0, -7, -3, -7, 0, -2, -1, 0,
    -- filter=104 channel=86
    -1, 3, 7, 8, 0, -1, 9, 6, 5,
    -- filter=104 channel=87
    -6, 0, 3, 1, -2, -1, 9, -7, 9,
    -- filter=104 channel=88
    -1, 5, 3, 5, 2, 6, 1, 3, -1,
    -- filter=104 channel=89
    13, 5, 3, 11, 3, -7, 0, -13, -13,
    -- filter=104 channel=90
    5, -3, 2, 1, -5, 8, -1, -4, 10,
    -- filter=104 channel=91
    4, 5, -6, 9, -14, 2, -3, -11, -12,
    -- filter=104 channel=92
    0, 0, 8, 3, 0, 4, 2, 0, 0,
    -- filter=104 channel=93
    -8, 0, -2, -3, -7, 1, -6, -3, -4,
    -- filter=104 channel=94
    -1, 1, -2, -7, 2, 1, 0, -1, -5,
    -- filter=104 channel=95
    2, 6, 1, 3, -6, 6, 3, -5, -1,
    -- filter=104 channel=96
    2, 7, 5, 8, -3, 3, 6, 0, 3,
    -- filter=104 channel=97
    0, -6, 1, 0, 2, 5, 6, -2, 1,
    -- filter=104 channel=98
    8, -2, 5, 3, -8, 1, -9, -4, -4,
    -- filter=104 channel=99
    13, 4, -5, 7, -8, 8, -5, -12, 0,
    -- filter=104 channel=100
    -2, -4, 3, -2, 1, -4, 4, -5, -1,
    -- filter=104 channel=101
    0, 1, 5, -5, -7, -4, -5, -7, 1,
    -- filter=104 channel=102
    0, -3, 0, -6, 3, -6, 7, -1, -7,
    -- filter=104 channel=103
    1, -2, 2, -4, -10, 6, -2, -6, -5,
    -- filter=104 channel=104
    0, 2, 0, 0, -4, -4, -10, -15, 0,
    -- filter=104 channel=105
    -7, 7, -9, 2, 6, -7, 7, 7, -3,
    -- filter=104 channel=106
    0, 0, 3, 8, 0, -2, 4, 4, 6,
    -- filter=104 channel=107
    -2, 6, 0, -2, -1, 9, 4, -3, 6,
    -- filter=104 channel=108
    5, 1, 1, 9, 1, 2, 12, 6, 3,
    -- filter=104 channel=109
    4, 1, 0, 4, -4, 0, -3, -22, -13,
    -- filter=104 channel=110
    3, -7, 4, 11, 2, -2, -5, -4, 5,
    -- filter=104 channel=111
    7, -3, -5, 0, 4, 6, 3, 5, 1,
    -- filter=104 channel=112
    1, -7, 2, 0, -12, 6, 1, -12, -4,
    -- filter=104 channel=113
    7, -5, -1, 0, -2, 6, -1, -5, -9,
    -- filter=104 channel=114
    -6, -3, 1, 10, 0, 4, 0, -5, 3,
    -- filter=104 channel=115
    8, 2, -1, 7, -2, 6, 0, -4, 3,
    -- filter=104 channel=116
    4, 3, 2, 0, -8, -11, -7, -16, -17,
    -- filter=104 channel=117
    3, -4, 0, -5, 5, -1, -4, -9, -10,
    -- filter=104 channel=118
    -4, 6, -1, -5, 2, 7, -6, 6, -5,
    -- filter=104 channel=119
    0, 1, -2, 3, -6, 9, 6, -8, 4,
    -- filter=104 channel=120
    0, 0, -1, 0, -17, 2, -11, -18, -8,
    -- filter=104 channel=121
    6, 1, -7, 2, -6, -1, 6, -7, -9,
    -- filter=104 channel=122
    0, -12, -2, -11, -20, 1, -23, -10, -12,
    -- filter=104 channel=123
    3, 5, 0, -2, 4, 5, 4, 1, 4,
    -- filter=104 channel=124
    -6, 0, -6, -4, -6, -3, 5, -3, 6,
    -- filter=104 channel=125
    14, 7, -4, 9, 0, -4, -5, -15, -13,
    -- filter=104 channel=126
    9, 9, 3, 5, 11, 0, 12, 8, -4,
    -- filter=104 channel=127
    2, -4, -3, -4, -3, 1, 3, -3, 2,
    -- filter=105 channel=0
    -2, 6, -2, 6, 2, 5, -4, -6, 3,
    -- filter=105 channel=1
    8, 15, -2, -11, 6, 5, -7, -11, 5,
    -- filter=105 channel=2
    0, 4, 3, 0, -5, -4, 0, -8, 4,
    -- filter=105 channel=3
    3, -6, 5, 13, -2, -15, -5, 9, -4,
    -- filter=105 channel=4
    8, 5, 0, 1, 8, 0, 11, -1, -5,
    -- filter=105 channel=5
    2, -6, -6, 6, -6, -6, -8, -3, -2,
    -- filter=105 channel=6
    2, 4, 0, -3, 5, -8, -2, 0, 5,
    -- filter=105 channel=7
    -5, -1, 3, -5, 4, 0, 0, 6, -4,
    -- filter=105 channel=8
    -3, -2, 2, -2, 0, -9, 2, -4, 1,
    -- filter=105 channel=9
    3, 4, -3, 3, 5, 0, 0, -9, 4,
    -- filter=105 channel=10
    3, -2, -4, 5, 1, -4, -1, 3, -1,
    -- filter=105 channel=11
    -7, -10, -5, -3, 10, -2, 0, 10, 5,
    -- filter=105 channel=12
    7, -1, 5, 5, 10, 5, 1, 0, -3,
    -- filter=105 channel=13
    9, 1, -2, 6, 23, -5, -5, -1, 2,
    -- filter=105 channel=14
    6, 7, -3, 4, 2, 4, -6, 3, 0,
    -- filter=105 channel=15
    2, 1, -1, 8, 14, -6, -13, 3, -3,
    -- filter=105 channel=16
    4, 3, 10, 0, 3, 7, -6, -2, 8,
    -- filter=105 channel=17
    -2, 3, -4, -6, 3, 4, -5, 6, -1,
    -- filter=105 channel=18
    0, -4, -11, 2, 20, -1, -11, 0, 5,
    -- filter=105 channel=19
    1, -3, 0, -3, 3, 6, -2, -6, 5,
    -- filter=105 channel=20
    -11, -12, -13, 5, 15, -12, -8, 7, 3,
    -- filter=105 channel=21
    11, 1, 11, -6, -2, 6, -1, -18, 3,
    -- filter=105 channel=22
    -2, 3, 4, 9, 11, -5, -3, 11, -4,
    -- filter=105 channel=23
    0, -22, 4, 18, 20, -11, -13, 23, -4,
    -- filter=105 channel=24
    2, 6, 2, -2, 6, -2, -2, -2, 4,
    -- filter=105 channel=25
    3, 3, -5, -6, 15, 8, -14, -16, 16,
    -- filter=105 channel=26
    4, 10, -6, -8, -11, -2, 4, -4, -2,
    -- filter=105 channel=27
    5, -1, 0, -3, 24, 0, -24, -1, 4,
    -- filter=105 channel=28
    3, 2, 0, -2, -4, -5, -7, 6, 3,
    -- filter=105 channel=29
    -12, -2, -13, 1, 12, 0, -1, 9, 0,
    -- filter=105 channel=30
    5, 8, 5, 0, 1, -6, -10, -8, 4,
    -- filter=105 channel=31
    0, -5, 1, 0, 7, -13, -15, 0, 10,
    -- filter=105 channel=32
    -1, 0, -10, 0, 22, -4, -7, 0, 0,
    -- filter=105 channel=33
    13, -9, 0, 3, 7, -9, -9, -2, 11,
    -- filter=105 channel=34
    0, 0, 0, 8, 0, 5, -7, 19, -3,
    -- filter=105 channel=35
    0, 1, 0, 2, -7, 6, -4, 2, 7,
    -- filter=105 channel=36
    0, -6, 1, 2, -2, 3, 7, -1, 0,
    -- filter=105 channel=37
    9, 0, 7, 4, -8, 9, -1, -15, 9,
    -- filter=105 channel=38
    8, 2, -1, -1, 8, -2, 0, 3, 4,
    -- filter=105 channel=39
    -5, -9, -5, 4, -1, -10, -5, 5, 4,
    -- filter=105 channel=40
    0, 1, -8, 0, 11, -5, 5, 7, -8,
    -- filter=105 channel=41
    -6, 7, 0, -19, 6, 17, 19, -4, -7,
    -- filter=105 channel=42
    11, 8, -1, 0, -9, -2, 0, -7, 6,
    -- filter=105 channel=43
    -1, -3, 6, 17, 10, -8, 0, 21, 2,
    -- filter=105 channel=44
    10, 6, -3, -3, -7, -3, -11, -4, 7,
    -- filter=105 channel=45
    1, 4, -1, 1, -8, -3, -8, 0, 5,
    -- filter=105 channel=46
    -3, 4, -1, -2, -3, -4, 6, 0, -5,
    -- filter=105 channel=47
    7, 10, 0, -10, 0, 3, -6, -17, 5,
    -- filter=105 channel=48
    2, 6, 5, -1, 4, 8, -13, -10, 12,
    -- filter=105 channel=49
    7, -4, -10, -11, 11, -12, -4, -14, -1,
    -- filter=105 channel=50
    1, -7, 2, -4, 0, -8, -14, -1, 7,
    -- filter=105 channel=51
    0, -5, -2, -2, 2, 3, -3, -7, -5,
    -- filter=105 channel=52
    -4, -8, 1, 10, 2, -4, -2, 8, 4,
    -- filter=105 channel=53
    1, -4, -7, 4, 4, 1, -8, 7, -6,
    -- filter=105 channel=54
    -1, -4, -2, 3, 6, -2, 4, -5, 6,
    -- filter=105 channel=55
    4, 0, -8, 2, 27, -2, -9, 2, -1,
    -- filter=105 channel=56
    -4, 2, 1, 0, 7, 5, 4, 6, 5,
    -- filter=105 channel=57
    5, 3, 8, 3, 6, 5, 8, -1, -8,
    -- filter=105 channel=58
    3, -3, -5, 4, -8, 0, -3, -6, 3,
    -- filter=105 channel=59
    11, 4, -6, -4, -1, 0, -10, -17, 13,
    -- filter=105 channel=60
    0, 5, -4, -3, 6, -3, 1, -1, -3,
    -- filter=105 channel=61
    0, 4, 2, -6, -1, 4, 9, -4, 2,
    -- filter=105 channel=62
    1, 5, -4, 7, 3, 0, -2, 1, -2,
    -- filter=105 channel=63
    7, -8, -2, -1, -1, -6, 1, -8, 4,
    -- filter=105 channel=64
    5, -2, -5, -1, 2, 1, -4, 5, -4,
    -- filter=105 channel=65
    0, -3, 0, -1, -2, 4, 4, -1, -1,
    -- filter=105 channel=66
    1, 8, -3, 2, 11, 0, 11, -4, -5,
    -- filter=105 channel=67
    -2, 0, -7, 1, 1, 6, 4, 0, 5,
    -- filter=105 channel=68
    -1, 8, 6, -8, 6, -4, 3, 0, 0,
    -- filter=105 channel=69
    5, -1, -2, 3, 0, 5, -5, -1, -4,
    -- filter=105 channel=70
    4, -5, 7, 3, 11, 1, -9, 11, -1,
    -- filter=105 channel=71
    0, -4, 0, 10, 1, 2, -3, -4, -5,
    -- filter=105 channel=72
    7, -3, -3, 0, 3, -9, -12, -2, 6,
    -- filter=105 channel=73
    -7, -1, -7, 4, 8, 1, -1, -10, 0,
    -- filter=105 channel=74
    1, -5, 0, -3, 4, -12, -2, 13, 2,
    -- filter=105 channel=75
    4, -8, -2, 0, 2, 1, -6, -13, 5,
    -- filter=105 channel=76
    -6, 0, -11, 3, 12, -11, -7, 5, 1,
    -- filter=105 channel=77
    -3, -6, 1, 1, -4, 5, 1, -1, -2,
    -- filter=105 channel=78
    -1, -4, 4, 7, 0, 0, 0, -3, 6,
    -- filter=105 channel=79
    5, -2, 0, 3, 27, -7, -19, 1, 6,
    -- filter=105 channel=80
    14, 9, 7, -11, 2, 0, -11, -26, 16,
    -- filter=105 channel=81
    -6, 7, 6, -1, 4, 0, 6, 1, -1,
    -- filter=105 channel=82
    -3, -3, -2, -2, 5, -6, 5, 0, -7,
    -- filter=105 channel=83
    5, 1, 2, 0, -1, 7, -11, -9, 0,
    -- filter=105 channel=84
    0, 0, -9, 0, 14, -4, -4, -9, 1,
    -- filter=105 channel=85
    5, 4, -1, -1, 0, -1, 7, 7, 3,
    -- filter=105 channel=86
    -4, -3, -5, 3, 10, 3, 5, -3, 6,
    -- filter=105 channel=87
    -7, -6, 3, 0, 6, -6, 5, 16, 5,
    -- filter=105 channel=88
    0, -3, -1, -2, -4, -8, -1, 5, 1,
    -- filter=105 channel=89
    10, -1, 0, -7, 11, 0, -13, -12, -5,
    -- filter=105 channel=90
    -8, 0, 0, 5, 2, 2, 7, 5, 4,
    -- filter=105 channel=91
    0, -1, -2, 2, 11, -6, -12, -12, 6,
    -- filter=105 channel=92
    4, -3, 2, 3, -1, -2, 8, 14, -4,
    -- filter=105 channel=93
    16, 16, 7, -11, -5, 2, -7, -19, 1,
    -- filter=105 channel=94
    0, -4, 0, -2, 3, 4, 0, 4, -1,
    -- filter=105 channel=95
    0, -7, 4, 2, 7, -7, 0, 1, -3,
    -- filter=105 channel=96
    -2, 7, 0, -8, 4, 6, -2, -3, 3,
    -- filter=105 channel=97
    4, 2, 2, 5, -7, -2, -5, 3, -4,
    -- filter=105 channel=98
    6, -2, -1, 4, 4, -3, -18, -17, 2,
    -- filter=105 channel=99
    1, -9, 0, -2, 2, -6, -8, 6, 1,
    -- filter=105 channel=100
    -8, 5, 7, 3, 3, 7, -3, -2, -1,
    -- filter=105 channel=101
    1, 1, -5, 5, 5, 2, 7, -7, -2,
    -- filter=105 channel=102
    7, 6, -1, 2, 4, -5, -2, 6, -3,
    -- filter=105 channel=103
    5, -6, -5, 5, -10, 1, -16, -12, 10,
    -- filter=105 channel=104
    8, -2, -6, -5, -4, -3, -3, -9, 11,
    -- filter=105 channel=105
    -10, -7, -7, 2, 3, 3, 6, 11, -2,
    -- filter=105 channel=106
    1, 4, -6, 0, 1, 0, 6, 5, -3,
    -- filter=105 channel=107
    -5, -5, -11, 12, 14, -1, -3, 6, -6,
    -- filter=105 channel=108
    2, -6, -8, 1, -4, 7, 5, 1, 0,
    -- filter=105 channel=109
    6, 5, -9, -11, 19, -5, -19, -2, 6,
    -- filter=105 channel=110
    -2, -9, 1, 7, 0, 1, -3, 7, 1,
    -- filter=105 channel=111
    -1, 1, -2, -7, 5, 2, 0, 0, 6,
    -- filter=105 channel=112
    0, -5, 0, -3, 8, 0, -5, 0, 5,
    -- filter=105 channel=113
    5, 1, 0, 3, 11, -1, -8, 5, -3,
    -- filter=105 channel=114
    4, 5, -8, -12, 14, -2, -17, 0, -4,
    -- filter=105 channel=115
    -5, 6, -1, 5, -6, 6, 7, 0, -2,
    -- filter=105 channel=116
    3, 7, 1, -8, 12, -4, -7, -8, 9,
    -- filter=105 channel=117
    -5, 4, -4, 0, 0, 4, -5, -1, 5,
    -- filter=105 channel=118
    0, 1, -1, -7, -3, 4, 1, 4, -7,
    -- filter=105 channel=119
    -2, -3, 9, 9, -4, 6, -7, 9, -1,
    -- filter=105 channel=120
    -3, -3, -15, 3, 17, -15, -21, 3, -4,
    -- filter=105 channel=121
    6, 8, -2, -3, 3, 5, -4, -5, 1,
    -- filter=105 channel=122
    19, 11, 10, -10, -5, 3, -10, -30, 4,
    -- filter=105 channel=123
    5, -7, 3, 4, 10, 8, -5, 12, -4,
    -- filter=105 channel=124
    2, 3, -6, 7, 7, -8, 2, 9, 0,
    -- filter=105 channel=125
    2, 0, -8, -5, 14, 2, -11, -14, 1,
    -- filter=105 channel=126
    -8, 1, -7, -6, 1, 0, 0, -9, -7,
    -- filter=105 channel=127
    2, 2, 0, -2, -3, -4, 9, 2, -8,
    -- filter=106 channel=0
    -1, -2, -6, 6, -10, -5, 11, 8, -11,
    -- filter=106 channel=1
    7, 9, 4, 3, -4, -3, 13, -2, -6,
    -- filter=106 channel=2
    3, 6, -2, -2, 2, 8, -5, 4, 7,
    -- filter=106 channel=3
    9, 5, 2, 11, 4, -5, -5, -1, 2,
    -- filter=106 channel=4
    7, -2, 10, -8, 0, 1, 6, 14, 4,
    -- filter=106 channel=5
    -3, 0, -5, 7, 0, -7, 0, -2, 0,
    -- filter=106 channel=6
    0, 1, -9, -5, 3, 0, -3, 3, 0,
    -- filter=106 channel=7
    1, 3, 4, 1, 4, -7, 3, 4, -4,
    -- filter=106 channel=8
    7, -6, 4, 3, 0, -5, 9, 10, 5,
    -- filter=106 channel=9
    2, -6, 2, -6, 2, -7, 0, 5, 0,
    -- filter=106 channel=10
    -6, 0, -8, -10, -8, -4, -2, 3, 7,
    -- filter=106 channel=11
    -2, -5, -3, 0, -3, -5, 5, 1, 8,
    -- filter=106 channel=12
    5, -5, 8, -5, 0, 7, 8, 6, -4,
    -- filter=106 channel=13
    -1, -4, 5, -7, 1, 8, 4, 2, 12,
    -- filter=106 channel=14
    0, -6, 2, -2, 3, -6, 0, -5, 0,
    -- filter=106 channel=15
    -5, -10, -7, -6, -6, -8, -1, -4, 0,
    -- filter=106 channel=16
    7, -1, 4, -1, 13, 2, 6, -5, -4,
    -- filter=106 channel=17
    -2, 4, 6, 3, -2, 0, 5, -2, 7,
    -- filter=106 channel=18
    -8, 0, -4, -15, -9, -12, -10, 0, 1,
    -- filter=106 channel=19
    2, 6, 1, 3, -3, -4, 0, 3, -4,
    -- filter=106 channel=20
    2, -4, 0, 3, -6, 0, -3, 3, 9,
    -- filter=106 channel=21
    7, 9, -1, -2, 6, 2, 2, 7, -5,
    -- filter=106 channel=22
    -1, 0, -7, 3, -8, -5, 6, 0, 4,
    -- filter=106 channel=23
    -6, -5, -11, -9, -7, 0, 0, 9, 6,
    -- filter=106 channel=24
    0, -3, -2, 2, -6, 2, 0, 5, 6,
    -- filter=106 channel=25
    -6, -1, -5, -10, -9, -4, 3, 0, 5,
    -- filter=106 channel=26
    -1, -1, 1, 4, 9, 0, 8, 1, -8,
    -- filter=106 channel=27
    -7, 4, -2, -19, -10, -10, -8, 10, -1,
    -- filter=106 channel=28
    3, -5, 5, -2, 3, -3, 5, -6, -7,
    -- filter=106 channel=29
    3, -8, -2, -7, -7, 0, -4, 6, 5,
    -- filter=106 channel=30
    -6, 0, -3, 4, -3, -2, -1, 9, 1,
    -- filter=106 channel=31
    -2, 3, -11, -8, 6, 9, 0, 0, 7,
    -- filter=106 channel=32
    0, -9, 0, -17, -18, -2, 0, -2, 3,
    -- filter=106 channel=33
    -1, -7, -6, 1, -8, -7, -10, 7, 2,
    -- filter=106 channel=34
    0, 2, 6, 6, 0, 1, 9, 3, 0,
    -- filter=106 channel=35
    6, -4, 0, 1, 4, -2, 1, -3, 0,
    -- filter=106 channel=36
    -4, 10, 10, -1, 7, 15, 3, 11, 11,
    -- filter=106 channel=37
    -2, -1, 3, 9, 7, -8, 9, 5, -11,
    -- filter=106 channel=38
    3, 0, -10, 2, -1, 0, -8, -1, 5,
    -- filter=106 channel=39
    1, -7, -5, -5, 0, 0, 3, 0, 0,
    -- filter=106 channel=40
    4, 0, 3, 0, 6, 7, 3, -3, 0,
    -- filter=106 channel=41
    2, -2, 2, 1, -4, -4, 2, -10, 6,
    -- filter=106 channel=42
    -3, 2, -4, 5, 0, -8, -3, 4, 0,
    -- filter=106 channel=43
    -3, -7, 0, -3, -9, -8, 0, -3, 7,
    -- filter=106 channel=44
    -2, -1, 1, 0, 0, 0, 6, -1, 1,
    -- filter=106 channel=45
    9, 4, 0, -5, 0, 5, 1, 1, -6,
    -- filter=106 channel=46
    0, -4, -6, 4, 3, 2, 2, -6, 5,
    -- filter=106 channel=47
    0, -3, -3, 6, -1, 3, 2, 9, -1,
    -- filter=106 channel=48
    -2, -3, -10, -1, -5, 8, 6, 13, -5,
    -- filter=106 channel=49
    -1, -3, -8, 0, 0, 0, 2, -5, -6,
    -- filter=106 channel=50
    -5, -7, -4, -8, -8, 0, -8, 8, -2,
    -- filter=106 channel=51
    0, 3, 1, -5, -3, -2, 0, -1, 6,
    -- filter=106 channel=52
    8, 3, 6, 3, 4, -6, 9, 0, 6,
    -- filter=106 channel=53
    -1, -7, -9, -8, 2, -2, -7, 3, -4,
    -- filter=106 channel=54
    1, 3, 7, -7, 0, -1, 0, 5, 5,
    -- filter=106 channel=55
    1, -3, -1, -14, -4, -5, -4, -1, 8,
    -- filter=106 channel=56
    4, -5, 0, -3, 6, 1, 7, 7, -6,
    -- filter=106 channel=57
    2, -2, 1, 0, -6, -2, -2, -2, 0,
    -- filter=106 channel=58
    -5, -5, 2, 2, 8, 3, -4, -1, 3,
    -- filter=106 channel=59
    -5, 4, 0, -8, -7, 2, -8, 6, -3,
    -- filter=106 channel=60
    -4, 2, 0, 2, -6, 2, 6, 0, -7,
    -- filter=106 channel=61
    3, -2, -3, 1, 6, 0, 3, 3, -7,
    -- filter=106 channel=62
    6, -4, 0, -5, 0, -3, 0, 0, 4,
    -- filter=106 channel=63
    1, -3, -8, 2, 0, 3, 1, -8, -1,
    -- filter=106 channel=64
    2, 1, 3, -1, 5, -1, -1, 8, 2,
    -- filter=106 channel=65
    6, -5, -4, -5, -3, -5, 5, 6, 0,
    -- filter=106 channel=66
    -5, 2, 0, 6, 0, 0, 2, 2, 0,
    -- filter=106 channel=67
    -2, -7, -3, -1, 8, -6, 0, 5, -2,
    -- filter=106 channel=68
    5, 6, 8, -4, -5, 6, 7, 5, 8,
    -- filter=106 channel=69
    -5, -1, -4, -2, 0, 1, -2, -2, -4,
    -- filter=106 channel=70
    7, 4, -2, -9, 2, -2, 5, 11, 4,
    -- filter=106 channel=71
    8, 3, 5, 7, -2, 7, -6, -6, 2,
    -- filter=106 channel=72
    -6, 3, -10, -6, 2, 0, -3, 6, 1,
    -- filter=106 channel=73
    -7, -5, -8, -5, -10, 0, 2, 7, -4,
    -- filter=106 channel=74
    5, -3, -4, -3, 0, 0, 6, 9, -9,
    -- filter=106 channel=75
    0, -5, -8, 12, -8, -19, -7, -10, 3,
    -- filter=106 channel=76
    -3, 0, -7, 0, -7, -1, -6, -5, 9,
    -- filter=106 channel=77
    2, -1, 0, 1, -6, 0, 7, -4, 5,
    -- filter=106 channel=78
    -1, 0, -4, 1, 1, -9, 5, -3, -1,
    -- filter=106 channel=79
    4, 4, 0, -11, -16, -10, -3, 6, 0,
    -- filter=106 channel=80
    -4, 8, -2, 0, -2, -4, -10, 8, -4,
    -- filter=106 channel=81
    4, -6, -3, 2, -1, 7, 5, -3, 6,
    -- filter=106 channel=82
    0, -2, 0, 0, 7, -3, -4, -4, 7,
    -- filter=106 channel=83
    2, -4, -5, 2, 1, 4, 7, -1, 4,
    -- filter=106 channel=84
    -4, -5, 0, -7, -2, 5, 9, 4, -1,
    -- filter=106 channel=85
    0, -4, -1, -3, 1, 4, -2, 0, 5,
    -- filter=106 channel=86
    5, -5, 6, 0, -8, -5, 8, 6, 4,
    -- filter=106 channel=87
    3, -7, -6, -5, 1, 2, -2, 2, 1,
    -- filter=106 channel=88
    -4, 1, 0, -3, 3, 13, 0, 6, 9,
    -- filter=106 channel=89
    0, 2, -4, -2, -11, -2, -11, 6, 4,
    -- filter=106 channel=90
    -4, 8, 0, 3, 14, 10, 0, 8, 8,
    -- filter=106 channel=91
    -5, 0, -9, -11, -3, 5, -2, 6, -5,
    -- filter=106 channel=92
    6, -7, 0, -1, 2, 0, 1, 6, 2,
    -- filter=106 channel=93
    5, 4, -1, 7, 8, 4, 1, 8, -1,
    -- filter=106 channel=94
    -6, 1, 4, -5, -6, -2, -3, -6, 6,
    -- filter=106 channel=95
    -1, 4, -2, -5, 5, 4, 0, -5, 6,
    -- filter=106 channel=96
    -2, 4, 5, 1, 6, -6, -4, -3, 7,
    -- filter=106 channel=97
    4, 2, -2, 11, 10, -3, -9, 5, 5,
    -- filter=106 channel=98
    -5, 1, -18, -10, -15, -6, -7, 5, -3,
    -- filter=106 channel=99
    -1, -3, 0, -13, -7, 5, 3, 14, 0,
    -- filter=106 channel=100
    -1, 1, -6, 2, 4, -6, 0, 4, 5,
    -- filter=106 channel=101
    0, -2, 9, -3, -4, -1, 4, 6, 7,
    -- filter=106 channel=102
    1, -3, 7, 6, 0, -7, 1, 7, 3,
    -- filter=106 channel=103
    1, -1, 1, 3, 8, -1, 4, -5, 2,
    -- filter=106 channel=104
    2, -3, 1, 2, 2, 11, -8, -3, 6,
    -- filter=106 channel=105
    0, -8, -8, -5, -6, -3, -6, 1, 2,
    -- filter=106 channel=106
    -2, 3, 3, 0, 3, 5, 4, -5, 10,
    -- filter=106 channel=107
    6, -8, 0, -8, -8, -9, 2, 5, -2,
    -- filter=106 channel=108
    0, 5, 0, -2, 3, -4, 3, 3, 6,
    -- filter=106 channel=109
    -5, 4, -11, -8, -12, 1, -6, 3, -6,
    -- filter=106 channel=110
    -8, -2, -7, 3, 7, -6, -7, 0, 8,
    -- filter=106 channel=111
    4, -4, 4, 0, 4, 4, 5, -2, -3,
    -- filter=106 channel=112
    -5, -5, 1, -3, -4, -2, 2, 0, -3,
    -- filter=106 channel=113
    4, 6, 1, -9, 4, 0, -5, 3, 3,
    -- filter=106 channel=114
    0, -2, -3, -16, -19, -3, -5, -3, -10,
    -- filter=106 channel=115
    -3, -6, -5, 2, 5, 4, 2, 2, 0,
    -- filter=106 channel=116
    0, -3, -2, -10, -8, 2, 0, 2, -1,
    -- filter=106 channel=117
    7, 4, 7, -8, 1, 3, 0, 0, 6,
    -- filter=106 channel=118
    0, 0, 6, -1, 7, -5, 4, -7, -4,
    -- filter=106 channel=119
    -2, -3, -5, 0, -4, 0, 5, -1, 1,
    -- filter=106 channel=120
    -2, 0, -4, -14, -8, 9, -3, 19, 5,
    -- filter=106 channel=121
    6, -4, 7, -6, -2, -6, 2, -4, 4,
    -- filter=106 channel=122
    0, 14, -4, 4, 13, 0, 2, 7, 0,
    -- filter=106 channel=123
    5, 0, 2, 2, 2, -6, 0, -5, -1,
    -- filter=106 channel=124
    -7, -1, 1, -7, -7, 3, -4, -4, 2,
    -- filter=106 channel=125
    2, 4, -6, -4, 3, 6, 2, 2, 4,
    -- filter=106 channel=126
    -2, -1, -2, 1, -8, -6, 0, 1, 6,
    -- filter=106 channel=127
    1, 0, 5, -6, -4, 4, 6, -5, -1,
    -- filter=107 channel=0
    4, -1, 6, -1, -2, 12, 0, 3, 5,
    -- filter=107 channel=1
    1, -9, 8, 0, -7, 0, -4, -4, 9,
    -- filter=107 channel=2
    -1, 4, 0, -4, -5, 3, -7, 5, 0,
    -- filter=107 channel=3
    -3, 8, 2, -13, 1, 5, -4, -1, 1,
    -- filter=107 channel=4
    -6, 3, 2, 4, -2, 4, -8, -4, -10,
    -- filter=107 channel=5
    -6, -6, 11, -12, -4, 8, -2, 3, -2,
    -- filter=107 channel=6
    -3, 0, 2, 7, 2, -5, -1, -7, -6,
    -- filter=107 channel=7
    -1, 5, -2, 0, 2, -3, -3, -4, -4,
    -- filter=107 channel=8
    0, 1, 0, 2, -6, -4, 6, -4, -5,
    -- filter=107 channel=9
    -5, 2, 10, -3, 1, 8, 5, 5, 2,
    -- filter=107 channel=10
    0, -8, 0, -2, 2, -8, 8, -2, -4,
    -- filter=107 channel=11
    -3, 11, 3, -2, 2, 2, -7, -6, -7,
    -- filter=107 channel=12
    1, -2, -2, 6, 0, -4, 1, -7, -7,
    -- filter=107 channel=13
    2, -9, -1, -5, -10, -5, -3, 5, -4,
    -- filter=107 channel=14
    6, 0, 2, -2, 0, -4, -7, 1, 3,
    -- filter=107 channel=15
    -1, 7, 11, 4, 3, -5, -7, 2, -1,
    -- filter=107 channel=16
    -11, -3, -4, -2, -12, -5, -9, -7, 5,
    -- filter=107 channel=17
    2, -6, -6, 3, 5, -1, -5, 4, -4,
    -- filter=107 channel=18
    2, 5, 0, 2, 10, 7, -2, 2, -13,
    -- filter=107 channel=19
    2, 2, 2, 4, -5, -5, 2, 2, -6,
    -- filter=107 channel=20
    5, 12, -5, 4, -7, -10, -14, -5, -9,
    -- filter=107 channel=21
    -5, -7, -12, -12, -12, 3, -5, -5, 6,
    -- filter=107 channel=22
    -4, -4, 7, 0, -1, 4, 2, 3, -8,
    -- filter=107 channel=23
    -6, 5, 13, -2, -5, 6, 6, -3, -15,
    -- filter=107 channel=24
    6, -6, 2, -2, 6, -2, 3, -4, 1,
    -- filter=107 channel=25
    8, -6, 4, -3, 0, 7, 5, -1, -3,
    -- filter=107 channel=26
    2, -5, 0, -5, -3, -6, -7, -9, 3,
    -- filter=107 channel=27
    -3, 3, 19, 0, 4, 18, 4, 12, -7,
    -- filter=107 channel=28
    0, 5, -1, 5, 3, -6, -2, -5, 7,
    -- filter=107 channel=29
    -3, 11, -1, 1, 2, -2, -10, 0, -18,
    -- filter=107 channel=30
    2, -7, 10, -7, -4, 13, 1, 5, 5,
    -- filter=107 channel=31
    -3, -19, 5, -7, -5, 14, 3, 0, 5,
    -- filter=107 channel=32
    1, 0, 3, 1, -2, 5, 4, -2, -3,
    -- filter=107 channel=33
    -2, -1, 7, 2, -7, 8, 2, 9, 1,
    -- filter=107 channel=34
    7, -7, 0, 1, -4, 0, 3, -14, -9,
    -- filter=107 channel=35
    -4, 0, -3, 4, 4, 2, -4, 0, 2,
    -- filter=107 channel=36
    -8, -3, -9, 0, 0, 0, -6, -10, -9,
    -- filter=107 channel=37
    -6, -8, 0, -7, -5, 3, -10, -2, 1,
    -- filter=107 channel=38
    0, -4, -3, 0, -6, 7, 0, 7, 4,
    -- filter=107 channel=39
    0, -2, 4, 0, 5, -8, -8, 2, -12,
    -- filter=107 channel=40
    4, 1, 1, -10, -6, -7, -5, -2, -1,
    -- filter=107 channel=41
    -1, -7, -18, 8, -5, -22, -10, -13, -13,
    -- filter=107 channel=42
    -3, 4, 4, -9, 5, 2, -6, 0, 2,
    -- filter=107 channel=43
    0, 4, -1, -1, -7, -3, -4, 0, -4,
    -- filter=107 channel=44
    -10, -13, 2, -4, 1, 3, -6, 4, 11,
    -- filter=107 channel=45
    -5, 1, 2, 2, 5, 4, 2, -4, 0,
    -- filter=107 channel=46
    0, 3, -8, -5, -1, -7, -6, 4, 0,
    -- filter=107 channel=47
    -12, -18, 0, -17, -8, 9, -2, 4, 0,
    -- filter=107 channel=48
    -11, -12, 5, -2, -3, 14, 3, 1, 12,
    -- filter=107 channel=49
    10, 4, 0, 12, 8, 1, -1, 10, -10,
    -- filter=107 channel=50
    -8, 5, 1, -3, -3, 3, 2, 0, 7,
    -- filter=107 channel=51
    5, -6, -3, 0, 4, -5, 5, 3, 0,
    -- filter=107 channel=52
    5, 0, -2, 6, -10, -9, -1, -14, -8,
    -- filter=107 channel=53
    1, -5, 0, 6, 6, 5, 0, -9, -6,
    -- filter=107 channel=54
    3, 2, -2, 4, -1, -1, -3, -6, -6,
    -- filter=107 channel=55
    4, 1, -1, -5, 0, -4, 4, 3, -13,
    -- filter=107 channel=56
    0, 1, -1, 3, 4, 5, 5, -1, -7,
    -- filter=107 channel=57
    2, -5, 0, -6, 8, -1, 3, -1, -4,
    -- filter=107 channel=58
    -2, 0, 7, -6, -5, 2, -9, 1, 7,
    -- filter=107 channel=59
    3, -9, -5, 8, -8, -3, 12, 9, 7,
    -- filter=107 channel=60
    0, -2, -1, 0, -2, -6, -6, -2, 5,
    -- filter=107 channel=61
    2, -8, -2, -4, -4, -8, -5, -10, -7,
    -- filter=107 channel=62
    -7, 2, -5, -1, -6, 1, -5, 0, -5,
    -- filter=107 channel=63
    -7, -8, 0, -5, -6, 5, 0, 2, 1,
    -- filter=107 channel=64
    -8, -8, 2, -10, -2, -9, -9, -8, -7,
    -- filter=107 channel=65
    1, -6, 3, 3, -4, 1, 7, -3, 5,
    -- filter=107 channel=66
    4, -12, -8, 6, -11, -10, -1, -6, -10,
    -- filter=107 channel=67
    -3, 1, -5, -5, 4, -6, -4, -3, -7,
    -- filter=107 channel=68
    3, 2, 1, 5, -2, -6, -5, -1, -3,
    -- filter=107 channel=69
    -1, -5, -7, 5, -5, 3, 0, 4, 1,
    -- filter=107 channel=70
    3, 3, 14, 1, -2, 5, 2, 0, -4,
    -- filter=107 channel=71
    1, 0, 7, -1, -5, 4, -1, -2, 0,
    -- filter=107 channel=72
    1, -12, -10, 3, -3, 2, 3, 10, -1,
    -- filter=107 channel=73
    6, 9, 8, 1, 4, 4, 3, 0, -4,
    -- filter=107 channel=74
    0, -5, 8, -5, -8, -1, 4, -6, -6,
    -- filter=107 channel=75
    -1, -3, 6, -5, -8, 7, 1, -11, 5,
    -- filter=107 channel=76
    2, -1, 1, 2, -6, -4, -11, -7, -13,
    -- filter=107 channel=77
    -3, 6, 0, 1, 5, -1, -3, 5, 2,
    -- filter=107 channel=78
    -5, 6, -3, -6, 1, 6, 5, 6, 4,
    -- filter=107 channel=79
    0, 2, 11, 6, -2, 4, 9, 2, -12,
    -- filter=107 channel=80
    -5, -21, -10, 3, -7, -1, 2, 1, 0,
    -- filter=107 channel=81
    -1, 7, 1, 1, -6, -1, 4, 3, 7,
    -- filter=107 channel=82
    4, -3, -1, -4, -4, -7, 2, 5, -4,
    -- filter=107 channel=83
    -9, 0, 9, 0, -5, -2, 0, 0, 6,
    -- filter=107 channel=84
    5, -6, 9, 6, 5, -1, -5, -4, -8,
    -- filter=107 channel=85
    -4, -3, -5, 5, -1, -6, -3, 5, -3,
    -- filter=107 channel=86
    4, -5, 4, 5, -8, -6, -6, 0, -2,
    -- filter=107 channel=87
    1, -2, 2, -8, -4, -2, -3, -6, -11,
    -- filter=107 channel=88
    -2, -13, -11, -2, -2, 0, 0, 1, -9,
    -- filter=107 channel=89
    4, -7, -10, 8, -9, 0, 9, 5, -8,
    -- filter=107 channel=90
    -11, -14, 0, 0, -13, -12, -11, -8, -9,
    -- filter=107 channel=91
    -4, 5, 0, 6, 0, 8, 4, 11, -8,
    -- filter=107 channel=92
    -6, 0, 2, 5, -2, 4, 5, -2, -3,
    -- filter=107 channel=93
    -12, -10, 0, -8, 2, 7, -7, -5, 9,
    -- filter=107 channel=94
    4, 4, 2, -4, -3, 1, 7, -1, 5,
    -- filter=107 channel=95
    0, 5, 4, -1, 5, 0, 4, -5, -1,
    -- filter=107 channel=96
    0, -2, -6, -3, -4, -2, -1, 2, -3,
    -- filter=107 channel=97
    -8, -1, 8, 0, -7, -4, 2, 0, 2,
    -- filter=107 channel=98
    1, -6, -1, 6, -9, 4, 14, 11, 3,
    -- filter=107 channel=99
    -2, -14, -1, 0, 2, 3, 8, -7, -7,
    -- filter=107 channel=100
    1, 1, -4, -3, 6, -5, -3, 1, -9,
    -- filter=107 channel=101
    0, -6, 7, 6, 9, -1, -10, 0, 4,
    -- filter=107 channel=102
    -3, -3, 3, -5, 0, -2, -5, 6, -5,
    -- filter=107 channel=103
    -11, 0, 1, -7, -1, 12, -9, -6, 5,
    -- filter=107 channel=104
    -8, -14, -9, 0, -4, -1, 3, 6, 7,
    -- filter=107 channel=105
    -4, 12, 0, 3, -2, -9, -3, 0, -4,
    -- filter=107 channel=106
    -7, 4, -6, 0, 4, -9, -10, 4, -11,
    -- filter=107 channel=107
    0, 5, 10, -6, 6, -3, -3, -5, -12,
    -- filter=107 channel=108
    -3, 3, -4, 4, -7, 0, -6, -8, -5,
    -- filter=107 channel=109
    1, -8, 12, 9, 8, 12, 4, 7, -5,
    -- filter=107 channel=110
    4, 1, -11, -7, 0, -6, 0, 0, -6,
    -- filter=107 channel=111
    7, -5, -6, -5, -7, -1, 6, -8, 4,
    -- filter=107 channel=112
    -6, 4, 2, 6, 2, 0, 11, -2, -1,
    -- filter=107 channel=113
    5, -8, -3, -7, -8, 8, 2, -4, -3,
    -- filter=107 channel=114
    7, 9, 16, 1, 0, 2, 6, -2, -1,
    -- filter=107 channel=115
    2, 2, 5, 1, 1, -2, 0, 5, -4,
    -- filter=107 channel=116
    8, -2, 1, 11, 0, 0, 6, 5, -7,
    -- filter=107 channel=117
    -2, 0, -11, 2, 1, 1, 7, 0, 0,
    -- filter=107 channel=118
    2, 0, 0, 5, 1, 0, -6, 1, -3,
    -- filter=107 channel=119
    -6, -8, 5, 4, -9, 1, 3, 0, 2,
    -- filter=107 channel=120
    6, 8, 15, 12, 11, 10, 7, -4, 0,
    -- filter=107 channel=121
    2, -11, -9, 0, -11, -3, 0, -6, -5,
    -- filter=107 channel=122
    -18, -13, -16, -23, -17, -4, -14, 2, 0,
    -- filter=107 channel=123
    -1, -2, 4, 2, 1, -7, -4, 3, 3,
    -- filter=107 channel=124
    1, 3, -4, 2, 6, -1, 2, -3, -5,
    -- filter=107 channel=125
    -2, -10, -2, 0, -9, -6, 9, 8, -3,
    -- filter=107 channel=126
    7, -1, -3, 0, -9, -7, 4, 6, 0,
    -- filter=107 channel=127
    -5, 4, -10, -1, -4, -10, 2, 2, 0,
    -- filter=108 channel=0
    -2, 6, 0, -2, -3, -7, -7, -8, -2,
    -- filter=108 channel=1
    -4, 8, 0, -2, -6, -4, 4, -6, -5,
    -- filter=108 channel=2
    -3, 4, 0, -2, 6, 7, 0, 2, 4,
    -- filter=108 channel=3
    -1, 0, -4, -6, 0, 5, 2, -6, 0,
    -- filter=108 channel=4
    -3, 3, 6, 5, 6, -6, 0, 5, -4,
    -- filter=108 channel=5
    7, 3, 2, -1, -6, 5, -5, 3, -5,
    -- filter=108 channel=6
    7, -6, 5, -1, 0, 0, 5, 2, 1,
    -- filter=108 channel=7
    5, 5, 0, 2, 0, 6, -5, 2, 7,
    -- filter=108 channel=8
    -4, -2, 3, -6, 0, -5, -1, 1, -5,
    -- filter=108 channel=9
    1, -2, 0, -5, 3, -2, 1, -3, 6,
    -- filter=108 channel=10
    -5, -1, 0, 1, 1, 6, -2, 4, 5,
    -- filter=108 channel=11
    -3, -5, 3, -4, 3, 5, 7, -6, 5,
    -- filter=108 channel=12
    -7, 2, 1, 2, 3, -7, 1, -5, 7,
    -- filter=108 channel=13
    -2, 0, -2, 4, 1, 3, -5, -5, 0,
    -- filter=108 channel=14
    -2, -3, 7, -4, 3, -5, -2, 2, -6,
    -- filter=108 channel=15
    -3, 0, 6, -6, 1, 4, 2, 4, -6,
    -- filter=108 channel=16
    -6, 6, 4, -5, -6, 0, 1, -6, 2,
    -- filter=108 channel=17
    3, 0, 0, 0, 0, -1, 0, -7, 6,
    -- filter=108 channel=18
    -4, 6, 4, 0, -7, -8, -6, 1, -1,
    -- filter=108 channel=19
    1, 7, 4, 2, -3, -4, -3, -6, 2,
    -- filter=108 channel=20
    1, -2, -3, -6, -5, -6, -5, 0, -1,
    -- filter=108 channel=21
    -2, -6, 5, 3, -6, 0, 5, 1, 0,
    -- filter=108 channel=22
    -5, 0, 3, 1, -1, 1, -2, 7, -4,
    -- filter=108 channel=23
    4, 3, -1, -4, 0, 6, 3, -3, 3,
    -- filter=108 channel=24
    5, 1, 0, -5, -1, 3, 0, 5, -5,
    -- filter=108 channel=25
    1, -7, -1, 5, -3, -1, 2, 0, -2,
    -- filter=108 channel=26
    4, 3, -4, 0, 5, 1, 3, -5, 0,
    -- filter=108 channel=27
    5, 5, 3, 0, 4, -3, 2, -2, 0,
    -- filter=108 channel=28
    5, -6, 7, -4, -4, 6, 4, 4, 1,
    -- filter=108 channel=29
    -1, -2, 3, 2, -5, 1, -5, 5, -2,
    -- filter=108 channel=30
    -1, -6, 0, 4, 5, 0, 6, -7, 1,
    -- filter=108 channel=31
    4, -1, -3, 2, 2, 2, 0, 0, -2,
    -- filter=108 channel=32
    -2, -2, -1, 0, -5, 0, -1, -1, 3,
    -- filter=108 channel=33
    2, 0, 6, -1, -6, -2, 5, -2, 1,
    -- filter=108 channel=34
    -4, 7, -3, -5, -3, -3, 5, 5, -5,
    -- filter=108 channel=35
    -5, -7, 2, 2, -1, -7, -4, -3, 0,
    -- filter=108 channel=36
    4, -3, -5, 4, -3, -3, 4, 5, 7,
    -- filter=108 channel=37
    3, 6, 0, 1, -2, -1, 0, -6, 7,
    -- filter=108 channel=38
    -4, -5, -1, 1, 1, -4, 6, 5, -4,
    -- filter=108 channel=39
    1, 6, -7, 3, -5, 4, 3, 1, 0,
    -- filter=108 channel=40
    1, 3, 2, 0, 3, 1, 3, 6, -3,
    -- filter=108 channel=41
    6, 0, 2, 8, -7, 6, -3, -6, -3,
    -- filter=108 channel=42
    5, 3, -3, -3, 7, -4, -2, -2, 5,
    -- filter=108 channel=43
    -5, 4, -3, -6, -2, 1, 6, -5, 3,
    -- filter=108 channel=44
    0, -4, -2, -4, 6, 4, -6, 6, 1,
    -- filter=108 channel=45
    -2, 5, 0, 4, -1, 3, 1, -6, -4,
    -- filter=108 channel=46
    4, -5, -1, -4, 1, -2, 2, 4, -3,
    -- filter=108 channel=47
    6, -2, 3, -4, -5, -1, 1, 0, -5,
    -- filter=108 channel=48
    -7, 1, 3, 1, -2, 0, 0, 0, 0,
    -- filter=108 channel=49
    -6, 2, 0, 6, 2, 2, -5, -1, -7,
    -- filter=108 channel=50
    0, -1, 6, 1, -5, 2, 0, 0, -5,
    -- filter=108 channel=51
    3, 0, -6, 0, 4, -7, -1, 0, 6,
    -- filter=108 channel=52
    3, 6, -6, -5, 6, -5, 1, -2, -1,
    -- filter=108 channel=53
    0, -1, 0, -5, 3, -1, 7, -5, -1,
    -- filter=108 channel=54
    -5, -4, 4, -4, 2, 1, 5, 1, 0,
    -- filter=108 channel=55
    -4, -1, -4, 0, 1, -7, -2, -6, -6,
    -- filter=108 channel=56
    5, 2, -5, 1, 0, -6, 5, 0, 3,
    -- filter=108 channel=57
    0, 5, 2, -2, 4, 0, -3, 5, -6,
    -- filter=108 channel=58
    -4, 0, -3, -7, -6, -2, -3, -5, -4,
    -- filter=108 channel=59
    -4, -7, -1, -5, -5, 4, 7, 6, 0,
    -- filter=108 channel=60
    2, -1, -2, 5, -2, 0, -2, -6, 0,
    -- filter=108 channel=61
    -2, 3, -2, -6, 1, 0, -2, 5, -2,
    -- filter=108 channel=62
    -7, 3, -1, -1, -5, -3, 4, 1, 1,
    -- filter=108 channel=63
    -6, 0, 8, 7, -4, -4, 4, -4, -2,
    -- filter=108 channel=64
    1, 3, 7, 0, 0, -5, 0, 0, 2,
    -- filter=108 channel=65
    4, -6, 2, 0, 7, -1, -5, 1, 1,
    -- filter=108 channel=66
    5, 0, 4, 7, -7, -1, -1, 1, 7,
    -- filter=108 channel=67
    -2, -3, 5, 6, 0, 5, 0, 0, 5,
    -- filter=108 channel=68
    -5, -1, -6, -6, -4, -6, 6, 1, 0,
    -- filter=108 channel=69
    6, -6, 5, 0, -2, 7, -1, 1, -2,
    -- filter=108 channel=70
    -5, -5, -7, -5, -3, 0, -2, 3, -5,
    -- filter=108 channel=71
    -3, -3, 5, 4, 3, 6, -6, 6, 4,
    -- filter=108 channel=72
    6, -1, 5, -7, 3, -4, 7, 1, -5,
    -- filter=108 channel=73
    -2, -5, 2, -4, 1, 1, -2, 4, -5,
    -- filter=108 channel=74
    -1, -6, -1, -1, -2, 6, -4, 7, 0,
    -- filter=108 channel=75
    4, 0, 8, -5, -6, 2, 0, 5, 5,
    -- filter=108 channel=76
    -5, -6, 1, 3, 5, 7, 3, 2, 2,
    -- filter=108 channel=77
    -4, 6, 4, 0, -4, 5, -1, 2, 0,
    -- filter=108 channel=78
    3, 2, -7, -6, 0, -5, -2, 2, -4,
    -- filter=108 channel=79
    5, -2, 3, -2, -6, 5, 1, -5, 0,
    -- filter=108 channel=80
    -3, 3, -4, -1, -5, -4, 0, -5, 0,
    -- filter=108 channel=81
    4, -3, -6, 2, 6, 0, -3, 3, -7,
    -- filter=108 channel=82
    1, -4, 4, -4, -6, 1, 2, -5, -2,
    -- filter=108 channel=83
    -4, 2, -5, 4, -4, 1, -6, 3, -2,
    -- filter=108 channel=84
    1, -2, -5, 1, -4, 6, -5, -7, 4,
    -- filter=108 channel=85
    -2, -3, 2, -1, -1, -6, -6, 1, 0,
    -- filter=108 channel=86
    4, 3, 0, 1, -3, -5, 2, 3, 5,
    -- filter=108 channel=87
    -7, -2, 0, 7, 1, 2, 2, -4, 1,
    -- filter=108 channel=88
    -6, 0, -2, -3, -2, 3, -2, 7, 0,
    -- filter=108 channel=89
    -1, 4, 6, 3, 1, -6, 2, -2, -6,
    -- filter=108 channel=90
    0, 6, -5, 6, -5, 4, 0, -5, 4,
    -- filter=108 channel=91
    -1, -5, -5, 2, -2, -4, -1, -6, -2,
    -- filter=108 channel=92
    6, 2, 6, 2, -2, 7, -4, -7, 1,
    -- filter=108 channel=93
    5, 6, 2, 2, 0, 1, -6, 2, 3,
    -- filter=108 channel=94
    3, 4, 1, -6, 6, -2, 2, -1, 4,
    -- filter=108 channel=95
    7, -6, -2, 0, -3, 4, -1, -1, 7,
    -- filter=108 channel=96
    -2, 0, -1, -7, -3, 3, -2, 3, -1,
    -- filter=108 channel=97
    2, 7, 0, 1, -3, -1, 7, 2, 3,
    -- filter=108 channel=98
    2, 0, -2, -6, 0, 2, -5, 5, -7,
    -- filter=108 channel=99
    3, 1, 6, 3, -4, -6, 1, -1, 2,
    -- filter=108 channel=100
    -4, 0, 2, 0, -5, -1, 7, 5, 0,
    -- filter=108 channel=101
    -4, -1, 6, -6, 1, -5, -4, 1, 5,
    -- filter=108 channel=102
    0, -7, 1, -4, 0, 5, -4, -6, 3,
    -- filter=108 channel=103
    3, 0, 8, -7, -7, -6, 1, 1, 4,
    -- filter=108 channel=104
    1, -5, -3, -3, 6, -8, 7, 3, 7,
    -- filter=108 channel=105
    -1, 0, -2, 3, 0, 0, 3, -4, -3,
    -- filter=108 channel=106
    -5, 1, -7, -7, -3, 4, -3, -2, -4,
    -- filter=108 channel=107
    0, 0, 2, -6, 0, 2, 5, -2, -1,
    -- filter=108 channel=108
    3, -4, 2, -6, 3, -7, -6, -1, 1,
    -- filter=108 channel=109
    -5, 4, 3, 1, -6, -2, -2, 1, -8,
    -- filter=108 channel=110
    0, 3, 5, -6, 4, -4, 0, -6, 7,
    -- filter=108 channel=111
    -4, 4, -4, -5, 2, -6, -2, 3, -3,
    -- filter=108 channel=112
    4, 5, 4, 5, 0, 6, -4, -7, -4,
    -- filter=108 channel=113
    -2, -3, -3, -1, -1, -2, 5, 0, -6,
    -- filter=108 channel=114
    3, 2, -5, 3, -6, -5, 0, -1, 5,
    -- filter=108 channel=115
    -4, 6, -2, -6, 0, 6, -3, -3, 5,
    -- filter=108 channel=116
    0, 0, 5, 2, 0, 5, 4, -1, 5,
    -- filter=108 channel=117
    -6, 6, -4, 4, -4, -2, 0, 6, -5,
    -- filter=108 channel=118
    3, 3, 5, 4, -7, -3, -6, -6, 3,
    -- filter=108 channel=119
    0, -1, -3, 0, -3, 3, 3, -4, -5,
    -- filter=108 channel=120
    -6, 6, 6, 0, 2, -2, -5, 5, -1,
    -- filter=108 channel=121
    4, 2, 7, 7, 1, 1, 4, 1, -1,
    -- filter=108 channel=122
    -4, 0, -4, -4, -4, 4, 2, 0, -2,
    -- filter=108 channel=123
    4, 2, -1, -2, 6, -3, -6, 5, 7,
    -- filter=108 channel=124
    2, 3, 2, 2, 3, -2, 6, 7, 2,
    -- filter=108 channel=125
    -5, 5, -4, 4, -3, -2, 2, 1, 5,
    -- filter=108 channel=126
    0, 3, -4, -4, 0, -2, -2, 7, -7,
    -- filter=108 channel=127
    -6, 5, -3, 0, -7, 2, -4, 2, -6,
    -- filter=109 channel=0
    -14, 0, 7, -27, -7, 12, -6, -5, 1,
    -- filter=109 channel=1
    -18, 0, 11, -23, -7, 18, -5, -4, 9,
    -- filter=109 channel=2
    -4, -2, -8, 0, 3, 3, 6, -3, 1,
    -- filter=109 channel=3
    0, -4, -1, -13, -18, 1, -4, -2, 15,
    -- filter=109 channel=4
    -1, -5, -11, 1, -13, 7, -10, -10, 6,
    -- filter=109 channel=5
    1, 9, 3, -14, -2, 3, -7, 8, 8,
    -- filter=109 channel=6
    -4, 1, 2, 3, -4, -7, 4, -11, -7,
    -- filter=109 channel=7
    -5, 4, -7, -5, 0, 5, 0, -1, 0,
    -- filter=109 channel=8
    -8, 0, -3, -6, -2, -5, 0, 4, -4,
    -- filter=109 channel=9
    0, 0, 1, 6, 13, -8, -3, 9, 3,
    -- filter=109 channel=10
    -9, 2, -12, -3, 3, -9, 0, 9, -2,
    -- filter=109 channel=11
    14, 2, -3, 10, 0, 0, 0, 0, -1,
    -- filter=109 channel=12
    6, -7, -7, 5, -8, -2, -7, 1, 2,
    -- filter=109 channel=13
    -5, -5, 0, 0, -9, -8, -3, 5, 1,
    -- filter=109 channel=14
    1, -5, -4, -2, 5, 3, 4, 4, -2,
    -- filter=109 channel=15
    7, 0, -7, 4, 0, -2, 3, -4, -6,
    -- filter=109 channel=16
    0, 0, -11, 0, 6, -8, -5, 19, 0,
    -- filter=109 channel=17
    -2, 0, 7, 0, 5, 5, 4, 5, -4,
    -- filter=109 channel=18
    -4, -7, -1, -6, -2, 7, -2, -19, -5,
    -- filter=109 channel=19
    4, 2, -1, -4, 2, 4, 4, 2, 2,
    -- filter=109 channel=20
    18, 20, -2, 7, 5, 0, 0, 4, -13,
    -- filter=109 channel=21
    -8, 0, -24, 3, 19, -7, 4, 18, 4,
    -- filter=109 channel=22
    -5, 4, 6, 0, -10, 4, -4, 2, -4,
    -- filter=109 channel=23
    9, 0, -16, 12, -5, -26, 11, 7, -15,
    -- filter=109 channel=24
    3, 0, -6, -1, -1, 5, -3, -4, 4,
    -- filter=109 channel=25
    -13, -9, -8, -5, 12, -6, -1, 12, 3,
    -- filter=109 channel=26
    -10, 2, -10, 1, 5, -3, 3, 8, -3,
    -- filter=109 channel=27
    -12, 0, -3, 3, 0, -13, 5, 11, 2,
    -- filter=109 channel=28
    -4, -4, 3, -6, 0, 5, 3, 1, 2,
    -- filter=109 channel=29
    14, 12, 2, 8, 10, -8, 7, -1, -3,
    -- filter=109 channel=30
    -7, 4, -3, -4, -1, -5, -1, 9, 7,
    -- filter=109 channel=31
    5, 0, -30, 20, 12, -33, 12, 30, -13,
    -- filter=109 channel=32
    -7, -2, 3, -8, 3, 6, -5, -3, 0,
    -- filter=109 channel=33
    -13, -8, 0, -8, -4, 0, -1, 10, -4,
    -- filter=109 channel=34
    7, -1, 4, -3, -4, 9, 0, 1, 10,
    -- filter=109 channel=35
    6, -6, -4, -4, -1, -3, 4, 6, 0,
    -- filter=109 channel=36
    -2, -3, -10, 15, 6, -12, 1, 9, -8,
    -- filter=109 channel=37
    -7, 1, -5, -16, 5, 10, -8, -3, 0,
    -- filter=109 channel=38
    0, -2, -9, 4, 2, -5, 9, 11, 2,
    -- filter=109 channel=39
    9, 0, -5, 0, -4, -4, 2, -3, -1,
    -- filter=109 channel=40
    6, -4, 1, 6, 2, -9, 3, -8, -9,
    -- filter=109 channel=41
    -13, -15, 10, -9, -14, 10, -10, -11, 17,
    -- filter=109 channel=42
    -9, -2, -3, -7, 5, 10, 4, 6, 0,
    -- filter=109 channel=43
    2, -3, -6, -13, -3, -2, -8, 0, -6,
    -- filter=109 channel=44
    -6, -6, -2, -8, 13, -5, 2, 7, -5,
    -- filter=109 channel=45
    3, 0, 6, -1, 3, 6, -6, -4, 3,
    -- filter=109 channel=46
    -1, -8, 6, 3, -1, 2, -2, -9, -5,
    -- filter=109 channel=47
    -7, 1, -6, 1, 10, -4, 7, 26, 5,
    -- filter=109 channel=48
    -7, -9, -15, 2, 20, -2, 1, 19, 5,
    -- filter=109 channel=49
    1, 4, 2, 4, 3, 2, -3, 0, -4,
    -- filter=109 channel=50
    0, -3, -15, 9, -5, -13, 2, 4, -5,
    -- filter=109 channel=51
    7, -1, 0, -6, -1, 2, 2, 7, 6,
    -- filter=109 channel=52
    0, 3, -10, 1, -2, -9, -2, 3, -5,
    -- filter=109 channel=53
    8, 5, 1, 11, 8, -3, 1, 3, -1,
    -- filter=109 channel=54
    -1, -6, 1, -2, -4, 6, 1, -4, -2,
    -- filter=109 channel=55
    1, -2, -12, 5, 7, -4, 9, -2, -11,
    -- filter=109 channel=56
    -8, 2, -5, -8, 1, -5, 3, -7, 5,
    -- filter=109 channel=57
    -4, -4, 6, 3, -4, 0, -1, 0, 12,
    -- filter=109 channel=58
    -6, 9, -4, -3, -5, 9, -10, 2, 8,
    -- filter=109 channel=59
    -16, -1, -16, 6, 13, -7, 9, 12, -2,
    -- filter=109 channel=60
    3, -3, -2, -7, 5, -4, -6, -1, 7,
    -- filter=109 channel=61
    6, 0, -2, 2, 0, -7, 8, 10, -3,
    -- filter=109 channel=62
    -2, 5, -2, 4, -7, -3, -4, -2, 0,
    -- filter=109 channel=63
    0, 1, -4, -5, 4, 2, 0, 6, 9,
    -- filter=109 channel=64
    4, 1, -9, 4, 4, -6, 1, 7, -5,
    -- filter=109 channel=65
    -6, -5, -7, 2, -1, 6, 0, -4, -2,
    -- filter=109 channel=66
    0, -9, 2, -1, 0, 9, 7, 0, 11,
    -- filter=109 channel=67
    0, 5, -1, -4, -5, 4, -4, -2, 1,
    -- filter=109 channel=68
    2, 3, 3, 2, -5, 0, 1, 0, 5,
    -- filter=109 channel=69
    4, 4, -4, 0, 8, 4, 6, -1, -2,
    -- filter=109 channel=70
    -9, -11, -13, -1, -11, -11, -10, -3, -4,
    -- filter=109 channel=71
    6, -9, -10, -6, -2, -10, 9, 7, 2,
    -- filter=109 channel=72
    -1, -6, -25, 19, 12, -16, 6, 15, -4,
    -- filter=109 channel=73
    6, -3, -8, 9, 5, -8, -3, 1, -11,
    -- filter=109 channel=74
    7, -9, -11, 7, 1, -12, 9, 0, -2,
    -- filter=109 channel=75
    -13, 1, 4, -23, -11, 6, -1, 6, 19,
    -- filter=109 channel=76
    15, 11, 0, 7, 0, -1, 0, -9, 0,
    -- filter=109 channel=77
    0, 0, -3, 0, -1, 2, -2, 3, 6,
    -- filter=109 channel=78
    -2, 0, 1, -8, 1, -3, 0, 6, 1,
    -- filter=109 channel=79
    -7, -2, 0, -19, -17, 2, 0, -14, -6,
    -- filter=109 channel=80
    -7, 3, -12, 13, 13, -11, 12, 24, -4,
    -- filter=109 channel=81
    -6, 1, -3, -1, 5, 3, 4, 0, -5,
    -- filter=109 channel=82
    0, -6, 0, 1, -3, 0, 0, 4, 6,
    -- filter=109 channel=83
    2, 2, -11, 0, 15, -4, -1, 7, 4,
    -- filter=109 channel=84
    2, -3, -2, 3, -5, -2, -1, 3, -5,
    -- filter=109 channel=85
    -3, 3, 1, 1, -5, 6, -4, -6, -1,
    -- filter=109 channel=86
    -2, -2, 0, -5, 0, 1, -2, -7, -1,
    -- filter=109 channel=87
    4, -1, 2, 9, 6, 1, -5, -6, -7,
    -- filter=109 channel=88
    4, -6, -14, 14, 5, -8, 7, 11, -5,
    -- filter=109 channel=89
    -10, -4, -9, -5, 9, -15, 9, 3, 2,
    -- filter=109 channel=90
    2, -3, -9, -4, 0, -14, -1, 12, -11,
    -- filter=109 channel=91
    -2, 4, -11, 3, -1, -2, -3, 2, -8,
    -- filter=109 channel=92
    -5, -6, -4, 3, 2, 1, -6, 7, -3,
    -- filter=109 channel=93
    -4, 2, -5, 4, 15, 7, 1, 13, -6,
    -- filter=109 channel=94
    2, -6, -5, 7, 7, -1, 4, -4, 1,
    -- filter=109 channel=95
    3, -3, 0, 2, -5, 0, 2, 0, -4,
    -- filter=109 channel=96
    0, -3, 4, -3, -2, 6, -4, 3, -7,
    -- filter=109 channel=97
    -3, -5, -5, -6, -1, -12, 0, 7, 3,
    -- filter=109 channel=98
    -10, -11, -2, 3, 14, -10, 16, 14, 12,
    -- filter=109 channel=99
    6, 6, -30, 21, 13, -25, 10, 28, -17,
    -- filter=109 channel=100
    1, 4, 2, 2, -2, 7, 5, -3, 6,
    -- filter=109 channel=101
    -1, 0, -1, 0, -6, -5, 0, -8, -6,
    -- filter=109 channel=102
    1, 4, 2, -2, -2, -1, 2, -2, 0,
    -- filter=109 channel=103
    -9, 0, -4, 0, 7, -10, 9, 16, 6,
    -- filter=109 channel=104
    -6, 0, -23, 18, 23, -19, 3, 14, -4,
    -- filter=109 channel=105
    3, 15, -2, 5, -4, -1, 7, 5, -8,
    -- filter=109 channel=106
    3, -1, -3, -1, -8, 4, 2, 0, -1,
    -- filter=109 channel=107
    -1, -5, 1, 0, -10, -10, -12, -13, -6,
    -- filter=109 channel=108
    0, -2, 3, 0, 4, 9, -6, 7, 1,
    -- filter=109 channel=109
    -12, 0, -4, 13, 5, 0, 7, 12, -8,
    -- filter=109 channel=110
    1, -4, -16, 1, 6, -3, 11, 10, 2,
    -- filter=109 channel=111
    0, 6, 2, 2, 5, -4, -7, -7, -1,
    -- filter=109 channel=112
    4, 0, 4, 2, -4, -5, 0, 3, -2,
    -- filter=109 channel=113
    -10, -1, 0, -11, 0, -11, 3, 16, 1,
    -- filter=109 channel=114
    -12, 1, 8, -16, -16, 5, -10, -21, -7,
    -- filter=109 channel=115
    2, -2, 2, 4, -2, -1, 7, -2, 1,
    -- filter=109 channel=116
    -6, -5, -7, 14, 15, 0, 5, 15, -3,
    -- filter=109 channel=117
    -8, 1, 0, -6, 1, 4, 0, -6, -1,
    -- filter=109 channel=118
    0, 0, 1, -2, 5, -4, 5, 3, 4,
    -- filter=109 channel=119
    0, -10, -5, 5, -7, 7, -8, 6, 7,
    -- filter=109 channel=120
    9, 1, -14, 16, 14, -14, 8, -1, -16,
    -- filter=109 channel=121
    -6, 0, -7, 5, 0, -7, 4, 4, 7,
    -- filter=109 channel=122
    -6, -12, -24, -7, 17, -17, 7, 34, 1,
    -- filter=109 channel=123
    2, -7, -3, 4, 0, 5, 5, 3, 0,
    -- filter=109 channel=124
    8, 0, 1, 6, 5, -5, 0, 3, -5,
    -- filter=109 channel=125
    4, 4, -11, 7, 18, -11, 12, 20, -7,
    -- filter=109 channel=126
    -5, -6, 2, -11, -11, 1, 10, -1, 11,
    -- filter=109 channel=127
    -7, 4, -3, -4, -3, 7, -1, -9, 11,
    -- filter=110 channel=0
    -6, 2, -6, -2, 3, -18, 2, -2, -1,
    -- filter=110 channel=1
    -8, 11, -4, -11, 10, -13, -3, -4, 3,
    -- filter=110 channel=2
    7, -9, -2, -3, -5, -1, -6, -4, 6,
    -- filter=110 channel=3
    -16, 6, -20, -9, 3, -13, 1, -8, -7,
    -- filter=110 channel=4
    6, -13, -4, -14, -3, -10, -6, 22, -12,
    -- filter=110 channel=5
    0, 11, -5, 11, -1, -14, 1, -11, -4,
    -- filter=110 channel=6
    -1, 3, -1, 10, 5, 7, 4, -3, -1,
    -- filter=110 channel=7
    6, -4, 4, -1, 3, 7, -4, 5, 6,
    -- filter=110 channel=8
    6, -2, 10, 12, 4, 8, -3, 3, 0,
    -- filter=110 channel=9
    2, -9, -2, 4, -15, 0, 0, 0, 4,
    -- filter=110 channel=10
    -5, 17, -5, 9, 4, 10, 9, -1, 5,
    -- filter=110 channel=11
    -3, 4, -7, 1, 4, -10, -2, 1, -4,
    -- filter=110 channel=12
    -2, 32, 12, 11, 25, 19, 1, 20, 11,
    -- filter=110 channel=13
    -8, 14, 2, 3, 5, 2, 0, 8, 8,
    -- filter=110 channel=14
    -3, 0, 0, 1, -6, -4, 4, -4, 5,
    -- filter=110 channel=15
    -9, -7, -6, 0, -9, -6, -4, 0, 0,
    -- filter=110 channel=16
    6, 2, 6, 10, 7, 4, 9, -6, 8,
    -- filter=110 channel=17
    2, 6, -6, -5, 4, -2, -3, 0, -3,
    -- filter=110 channel=18
    0, 11, -14, 5, -8, -7, 7, -11, -2,
    -- filter=110 channel=19
    1, 4, -2, 1, -7, 5, -2, -7, 2,
    -- filter=110 channel=20
    0, 4, -1, 4, 3, 0, 1, 6, 3,
    -- filter=110 channel=21
    4, -4, -10, 1, -13, -5, -1, -6, 3,
    -- filter=110 channel=22
    1, -3, 3, 12, -8, 4, -6, 5, -7,
    -- filter=110 channel=23
    8, -13, -3, 13, -42, 17, 0, -12, 7,
    -- filter=110 channel=24
    7, -4, -6, 1, -6, 5, -7, 1, 6,
    -- filter=110 channel=25
    1, 1, 0, 3, -21, 15, -4, 1, 18,
    -- filter=110 channel=26
    10, 0, 4, -2, 1, -2, 0, -1, -6,
    -- filter=110 channel=27
    15, -22, 0, 17, -56, 17, -2, -10, 21,
    -- filter=110 channel=28
    -6, 0, 7, 3, 4, -7, 0, -3, -5,
    -- filter=110 channel=29
    2, 13, -8, 9, 8, -2, 5, 3, 7,
    -- filter=110 channel=30
    3, -8, 3, 10, -24, -5, -8, -7, 4,
    -- filter=110 channel=31
    3, -19, -5, 1, -50, 14, -7, -12, 16,
    -- filter=110 channel=32
    1, 8, -7, 13, -18, 15, -5, 2, 14,
    -- filter=110 channel=33
    1, -5, -1, 12, -20, 0, -1, -19, 9,
    -- filter=110 channel=34
    10, -4, 19, 25, 15, 25, -2, 20, -1,
    -- filter=110 channel=35
    -5, 0, -1, 1, -1, 0, 0, -2, 3,
    -- filter=110 channel=36
    -6, -2, 5, -5, -5, 16, -10, 4, 12,
    -- filter=110 channel=37
    1, 9, 0, 4, -9, -3, -8, 7, -8,
    -- filter=110 channel=38
    5, 1, -7, 3, -23, 11, -1, -15, 1,
    -- filter=110 channel=39
    -10, -6, -12, -6, 7, -6, 1, -6, 2,
    -- filter=110 channel=40
    -8, -11, -14, -5, 3, -8, -11, -12, -2,
    -- filter=110 channel=41
    5, 27, 16, 5, 81, -22, 12, 36, -4,
    -- filter=110 channel=42
    -7, -6, -8, 0, -4, -16, 0, -2, -1,
    -- filter=110 channel=43
    -12, -2, 2, 4, 1, -9, -1, -14, -6,
    -- filter=110 channel=44
    3, 6, -5, 16, -16, -2, 4, -4, 3,
    -- filter=110 channel=45
    -6, -9, -15, -13, -11, -5, -10, -4, -5,
    -- filter=110 channel=46
    4, -1, 6, -2, 7, -11, 2, 0, 0,
    -- filter=110 channel=47
    -1, 1, -16, 6, -9, -15, 0, -4, 1,
    -- filter=110 channel=48
    6, -5, -9, 8, -27, 8, -4, -6, 7,
    -- filter=110 channel=49
    5, -17, 1, -11, -11, -4, -9, 1, 0,
    -- filter=110 channel=50
    1, -26, -3, 1, -40, 5, -11, -16, -2,
    -- filter=110 channel=51
    -4, -1, 5, 6, 3, -4, 0, 1, -1,
    -- filter=110 channel=52
    -2, 3, 8, 8, 6, 28, 0, 15, 1,
    -- filter=110 channel=53
    -1, 9, 1, 2, -1, 4, -4, 2, -2,
    -- filter=110 channel=54
    -3, 0, 6, -6, -1, -1, -2, 3, 0,
    -- filter=110 channel=55
    -8, 0, -7, 11, 0, 16, 1, -2, 14,
    -- filter=110 channel=56
    19, 8, 16, 11, 18, 16, 13, 22, 0,
    -- filter=110 channel=57
    0, 2, 6, -2, 11, -6, 2, 0, -4,
    -- filter=110 channel=58
    0, 10, -6, 7, 18, -11, -1, 10, -7,
    -- filter=110 channel=59
    -4, 5, -3, 8, -13, 6, -7, -10, 4,
    -- filter=110 channel=60
    0, 1, 5, 0, 4, 5, 1, 0, -1,
    -- filter=110 channel=61
    5, 6, 4, -1, -2, 16, 0, 12, 4,
    -- filter=110 channel=62
    5, -2, 0, -1, 9, -6, -5, -3, 4,
    -- filter=110 channel=63
    7, 14, 5, 6, 3, 0, 7, -3, -7,
    -- filter=110 channel=64
    7, 0, -1, 0, 3, 0, -8, 6, -6,
    -- filter=110 channel=65
    4, -4, 1, 1, 2, -2, 2, 4, 6,
    -- filter=110 channel=66
    -5, 24, 14, 12, 29, 29, 8, 22, 16,
    -- filter=110 channel=67
    0, -4, 0, -1, 1, -5, 2, -4, -1,
    -- filter=110 channel=68
    -11, -2, -3, 0, -4, -1, -4, -5, -6,
    -- filter=110 channel=69
    -5, 9, -3, -3, 1, -6, 1, -4, -3,
    -- filter=110 channel=70
    5, -23, -7, 8, -36, 8, -9, -6, 4,
    -- filter=110 channel=71
    -5, 1, -1, -7, -1, -7, -3, -16, -6,
    -- filter=110 channel=72
    -3, 4, -5, 9, -23, 9, -8, -13, 12,
    -- filter=110 channel=73
    3, 3, 2, 8, -12, 3, -2, -4, 1,
    -- filter=110 channel=74
    13, -15, 16, 8, -25, 35, -9, 1, 16,
    -- filter=110 channel=75
    -3, 21, -5, -1, 12, -29, 8, -9, -1,
    -- filter=110 channel=76
    -1, 7, -12, -6, 1, -7, -1, -8, -5,
    -- filter=110 channel=77
    -7, 0, 0, 3, -1, 1, -1, 0, 5,
    -- filter=110 channel=78
    7, 0, -8, 7, -9, -7, 0, 5, 1,
    -- filter=110 channel=79
    0, 1, 1, 9, -8, 0, -4, -12, 5,
    -- filter=110 channel=80
    -2, 5, 0, -1, -23, 3, -10, -3, 11,
    -- filter=110 channel=81
    6, 2, -5, -6, 6, 0, -4, -5, -4,
    -- filter=110 channel=82
    -5, 0, -3, 2, -3, 1, 3, -1, -12,
    -- filter=110 channel=83
    11, -11, -8, -3, -19, 3, 0, -8, -1,
    -- filter=110 channel=84
    5, 0, -2, 9, -12, 6, -7, 8, 7,
    -- filter=110 channel=85
    -5, 6, 0, 2, 6, 0, -1, -4, 0,
    -- filter=110 channel=86
    4, 18, 5, 10, 0, 16, -1, 16, 11,
    -- filter=110 channel=87
    0, 2, 13, 14, 13, 23, 4, 18, 3,
    -- filter=110 channel=88
    2, -12, -1, -3, -12, 21, -9, 3, -2,
    -- filter=110 channel=89
    -8, 17, -12, -1, -11, 4, -2, -13, 19,
    -- filter=110 channel=90
    -1, -15, -3, -4, 0, 7, -11, 2, 0,
    -- filter=110 channel=91
    8, -17, 3, 7, -27, 9, -14, -9, 9,
    -- filter=110 channel=92
    -3, 0, -1, 10, 10, 4, 8, 3, -6,
    -- filter=110 channel=93
    10, 9, 9, 10, -22, -4, 2, 5, 8,
    -- filter=110 channel=94
    -1, -3, 0, 7, 2, 4, 0, 1, -6,
    -- filter=110 channel=95
    -1, 5, 1, -1, 7, 0, 0, -3, 10,
    -- filter=110 channel=96
    -2, -6, -4, -7, 2, -13, -7, 1, -2,
    -- filter=110 channel=97
    -1, -1, -5, -12, 4, -8, -8, -9, -12,
    -- filter=110 channel=98
    1, 10, -3, 9, -27, 4, 4, -10, 20,
    -- filter=110 channel=99
    11, -15, 0, 13, -35, 41, -16, 7, 27,
    -- filter=110 channel=100
    10, 15, 10, 9, 25, -3, 6, 17, 7,
    -- filter=110 channel=101
    -6, -13, -7, -11, -9, 3, -7, -1, -10,
    -- filter=110 channel=102
    4, -2, -5, 2, 4, -3, 1, 2, -1,
    -- filter=110 channel=103
    -3, 7, -17, 14, -17, -16, 3, -12, 8,
    -- filter=110 channel=104
    0, -5, -2, 6, -28, 14, 1, -2, 5,
    -- filter=110 channel=105
    -5, 4, -5, 6, 18, -7, 9, 3, 6,
    -- filter=110 channel=106
    -10, 0, -5, -5, 0, -7, -5, 2, -5,
    -- filter=110 channel=107
    4, 2, -14, 10, -3, 4, 3, -5, 2,
    -- filter=110 channel=108
    4, 5, -6, 0, 27, -6, 0, 4, -11,
    -- filter=110 channel=109
    6, -11, 1, 26, -39, 19, 0, -8, 18,
    -- filter=110 channel=110
    4, 2, 8, 3, 1, 11, 5, 2, 11,
    -- filter=110 channel=111
    4, 5, 3, 0, 8, 3, 5, 6, 4,
    -- filter=110 channel=112
    5, -13, -5, 10, -19, 16, -12, -12, 5,
    -- filter=110 channel=113
    -3, -1, -9, 12, -7, 0, 4, -19, -1,
    -- filter=110 channel=114
    -8, 8, -6, 16, -18, -6, 2, -3, 6,
    -- filter=110 channel=115
    3, -6, -1, -3, 3, 1, -5, 0, 0,
    -- filter=110 channel=116
    4, 2, 4, 0, -26, 3, -9, 0, 16,
    -- filter=110 channel=117
    0, 2, -4, 0, 1, 2, -2, 5, -2,
    -- filter=110 channel=118
    6, -5, -1, -3, -4, -5, 0, 3, -3,
    -- filter=110 channel=119
    29, 8, 20, 30, 30, 13, 10, 28, -3,
    -- filter=110 channel=120
    17, -20, -5, 15, -52, 18, -18, -18, 17,
    -- filter=110 channel=121
    3, 20, 0, 3, 8, 4, 8, 0, 12,
    -- filter=110 channel=122
    13, -8, -6, 3, -22, 9, 9, 1, 11,
    -- filter=110 channel=123
    5, 3, 9, 1, 2, 4, 5, 3, -2,
    -- filter=110 channel=124
    -3, 8, 0, -2, 4, 0, -4, 2, 0,
    -- filter=110 channel=125
    13, 0, -6, 16, -26, 21, -13, 1, 20,
    -- filter=110 channel=126
    -15, 14, -5, 0, 13, -5, 0, -1, 0,
    -- filter=110 channel=127
    3, 6, 7, 8, 10, 3, -1, -2, 6,
    -- filter=111 channel=0
    12, -11, -1, 9, -26, -7, 12, -11, -7,
    -- filter=111 channel=1
    3, -3, -2, 21, -13, 0, 12, 1, 0,
    -- filter=111 channel=2
    0, -4, 3, -1, -9, -1, 0, 7, 2,
    -- filter=111 channel=3
    1, 2, -16, -12, -13, -24, -7, -4, -6,
    -- filter=111 channel=4
    -9, -7, -14, 0, -8, -14, -16, 3, -11,
    -- filter=111 channel=5
    13, 4, 2, 9, -11, -9, 20, -13, -2,
    -- filter=111 channel=6
    6, 0, -1, -2, 0, -3, 0, -1, 6,
    -- filter=111 channel=7
    6, 2, 6, 4, -1, -1, 1, 4, 5,
    -- filter=111 channel=8
    5, 11, -10, 7, 8, -9, -2, 3, 3,
    -- filter=111 channel=9
    -2, 0, 0, 6, -11, 5, 0, -7, 7,
    -- filter=111 channel=10
    -6, 4, 9, 2, -5, 7, 13, -7, 1,
    -- filter=111 channel=11
    -1, 0, 0, 3, -1, -4, -11, 3, 0,
    -- filter=111 channel=12
    5, 2, -9, 18, 7, 4, 1, 12, 3,
    -- filter=111 channel=13
    0, -7, -2, 15, -14, 14, 13, -5, 1,
    -- filter=111 channel=14
    5, -6, -3, -6, 6, 5, -3, -3, 0,
    -- filter=111 channel=15
    -1, 6, -2, 1, -18, 11, 5, -14, 6,
    -- filter=111 channel=16
    0, 3, -9, 8, -11, 2, 18, -2, 8,
    -- filter=111 channel=17
    1, 0, 4, 2, -7, -3, 1, 5, 4,
    -- filter=111 channel=18
    -1, -4, 13, 17, -28, 13, 9, -14, 15,
    -- filter=111 channel=19
    -2, 3, -4, -5, -7, 5, 0, -7, -1,
    -- filter=111 channel=20
    -4, 3, -7, 1, -2, 0, -11, 0, 7,
    -- filter=111 channel=21
    3, -11, 4, 6, -12, 9, 1, 2, 4,
    -- filter=111 channel=22
    0, -2, -1, 3, -10, 8, -1, -1, 5,
    -- filter=111 channel=23
    -9, 12, -1, -8, 0, 0, 13, -14, 21,
    -- filter=111 channel=24
    0, -4, 2, 5, -4, 1, 0, 7, 4,
    -- filter=111 channel=25
    -4, -21, 10, 19, -33, 23, 10, -16, 16,
    -- filter=111 channel=26
    8, -6, 0, 0, -8, -5, 4, 4, -5,
    -- filter=111 channel=27
    -12, -8, 2, 24, -42, 16, 7, -36, 16,
    -- filter=111 channel=28
    -7, 4, 2, 1, 0, -3, -3, -3, 3,
    -- filter=111 channel=29
    -6, 4, 2, 0, 0, 1, -6, 0, -3,
    -- filter=111 channel=30
    -1, -9, 3, 12, -25, 7, 10, -13, 0,
    -- filter=111 channel=31
    -10, -8, -2, -4, -25, 14, 13, -20, 15,
    -- filter=111 channel=32
    0, -13, 3, 18, -37, 18, 16, -10, 11,
    -- filter=111 channel=33
    0, -10, 2, 5, -33, 19, 17, -19, 16,
    -- filter=111 channel=34
    17, 31, -7, 32, 51, -7, 22, 29, 3,
    -- filter=111 channel=35
    -5, 4, 2, -1, 3, 5, -7, -1, 1,
    -- filter=111 channel=36
    0, -6, 1, -4, 5, 3, -1, 4, -13,
    -- filter=111 channel=37
    9, -1, -7, 9, -5, -5, 11, -3, -8,
    -- filter=111 channel=38
    -2, 0, 4, 9, -15, 7, 11, -19, 4,
    -- filter=111 channel=39
    -2, 1, 0, -1, 4, -9, -6, -10, -9,
    -- filter=111 channel=40
    -4, -8, 7, -13, 2, 4, -10, -1, 5,
    -- filter=111 channel=41
    12, 10, 1, 50, 18, 35, 16, 48, 19,
    -- filter=111 channel=42
    -5, -8, -3, -5, -9, 0, -6, 2, -3,
    -- filter=111 channel=43
    -5, 10, -5, -5, 4, -1, 5, -7, 1,
    -- filter=111 channel=44
    0, 0, 1, 12, -14, -2, 6, -11, 6,
    -- filter=111 channel=45
    4, -12, 6, -9, -9, 6, 2, -8, -7,
    -- filter=111 channel=46
    -5, 0, 1, 0, 12, -6, 4, 3, -2,
    -- filter=111 channel=47
    9, -10, 0, 15, -27, -2, 17, -7, 3,
    -- filter=111 channel=48
    3, -17, 1, 10, -40, 6, 14, -10, 4,
    -- filter=111 channel=49
    -8, -4, 10, -2, -25, -6, 6, -4, 0,
    -- filter=111 channel=50
    -13, -12, 10, 0, -17, 11, 2, -20, 10,
    -- filter=111 channel=51
    -6, 0, 2, -6, -6, 0, 0, -6, -3,
    -- filter=111 channel=52
    -3, 17, -1, 5, 11, 2, 5, 5, 4,
    -- filter=111 channel=53
    4, -1, 1, 3, 1, 2, -2, -8, -2,
    -- filter=111 channel=54
    2, 5, -3, 3, 6, -5, -2, 0, 1,
    -- filter=111 channel=55
    -9, 8, 1, 6, -12, 10, 7, -18, 7,
    -- filter=111 channel=56
    5, 12, -1, 17, 27, -4, 11, 12, -1,
    -- filter=111 channel=57
    5, -2, 4, 3, 4, 9, 0, 13, 1,
    -- filter=111 channel=58
    8, 5, -8, 5, -5, -16, 9, -3, 1,
    -- filter=111 channel=59
    0, -21, 9, 14, -34, 26, 11, -14, 8,
    -- filter=111 channel=60
    1, 5, -6, -7, -2, -7, 6, -6, 0,
    -- filter=111 channel=61
    5, 0, -8, 6, 11, 1, 4, 3, 2,
    -- filter=111 channel=62
    -1, 5, -2, -5, 0, -1, -4, 5, -2,
    -- filter=111 channel=63
    6, 0, -3, 9, 5, -5, 3, 2, -6,
    -- filter=111 channel=64
    -4, 9, -8, -6, 15, -4, 3, 12, -7,
    -- filter=111 channel=65
    -1, -6, 0, -1, -5, -1, -5, -1, 5,
    -- filter=111 channel=66
    16, 8, -8, 28, 0, 24, 12, 21, 4,
    -- filter=111 channel=67
    4, 2, -5, -6, 3, 3, -5, -1, -8,
    -- filter=111 channel=68
    -9, -10, -3, 5, 0, -9, -3, -6, -6,
    -- filter=111 channel=69
    5, 1, -4, 0, -8, -6, 0, 3, 1,
    -- filter=111 channel=70
    1, 0, -8, -5, 0, 3, 1, -8, -1,
    -- filter=111 channel=71
    -9, -7, -3, -10, 0, 0, -2, -8, -9,
    -- filter=111 channel=72
    -8, -3, 9, 8, -25, 26, 13, -18, 10,
    -- filter=111 channel=73
    0, -4, -1, 7, -9, 0, 7, -9, -5,
    -- filter=111 channel=74
    1, 8, -13, 14, -3, 0, 5, -14, -1,
    -- filter=111 channel=75
    11, -9, 0, 6, -15, -3, 24, 0, 5,
    -- filter=111 channel=76
    -3, 4, -1, -1, 0, -3, -4, 0, -1,
    -- filter=111 channel=77
    -5, -7, 3, 5, 5, -6, -6, 6, 0,
    -- filter=111 channel=78
    0, 5, 2, 0, 3, -7, 5, 1, -4,
    -- filter=111 channel=79
    6, -3, 10, 19, -33, 17, 13, -31, 17,
    -- filter=111 channel=80
    -2, -20, 11, 10, -42, 26, 16, -23, 1,
    -- filter=111 channel=81
    -1, 3, -6, -4, 4, -2, 0, 7, 3,
    -- filter=111 channel=82
    0, -3, -5, -10, -2, -8, -2, -2, -1,
    -- filter=111 channel=83
    -1, -4, 0, -7, -11, 0, -2, -6, -10,
    -- filter=111 channel=84
    -9, 3, -1, 10, -15, 4, 10, 0, -1,
    -- filter=111 channel=85
    -4, -2, 0, -4, -4, -2, -4, -1, -6,
    -- filter=111 channel=86
    12, 5, -2, 12, -5, -4, 16, 5, -8,
    -- filter=111 channel=87
    6, 13, -12, 4, 5, 2, 6, 6, 0,
    -- filter=111 channel=88
    -11, 0, -7, -11, 1, 0, 0, 3, -10,
    -- filter=111 channel=89
    -4, -17, 1, 15, -31, 11, 12, -19, 13,
    -- filter=111 channel=90
    -14, 11, -16, -4, 16, -12, 5, 10, 2,
    -- filter=111 channel=91
    -13, -5, 1, 6, -20, 6, 2, -19, 2,
    -- filter=111 channel=92
    1, 14, 6, 10, 18, -6, 12, 14, 3,
    -- filter=111 channel=93
    2, -10, 8, 16, -15, 3, 12, -9, -8,
    -- filter=111 channel=94
    5, -1, -6, 6, 0, 1, 4, 5, 3,
    -- filter=111 channel=95
    4, 3, -7, 3, -3, 6, 7, -4, 8,
    -- filter=111 channel=96
    -3, 2, 6, -2, -2, -3, -5, 3, -9,
    -- filter=111 channel=97
    -10, -2, -5, -11, -4, -7, -7, -8, 2,
    -- filter=111 channel=98
    -1, -11, 4, 12, -43, 20, 16, -25, 14,
    -- filter=111 channel=99
    0, 1, 0, 12, -4, 7, 14, -6, 5,
    -- filter=111 channel=100
    2, 9, 5, 7, 33, 0, 1, 28, 7,
    -- filter=111 channel=101
    -15, -8, 0, -1, -8, -8, -3, -8, -13,
    -- filter=111 channel=102
    1, -1, -2, -1, 7, -5, 4, 7, -3,
    -- filter=111 channel=103
    3, -11, 6, 11, -28, -1, 19, -23, -3,
    -- filter=111 channel=104
    -7, -5, 15, 10, -21, 12, 4, -6, -2,
    -- filter=111 channel=105
    0, 3, -6, 2, 10, -8, 0, 0, 3,
    -- filter=111 channel=106
    0, 1, -1, -5, 7, -1, -11, 0, -1,
    -- filter=111 channel=107
    2, 4, -5, -9, -2, 0, 2, -8, -2,
    -- filter=111 channel=108
    5, 7, 2, 5, -1, 6, 0, 4, 1,
    -- filter=111 channel=109
    -9, -9, 10, 12, -34, 20, 19, -25, 13,
    -- filter=111 channel=110
    6, -1, 4, 1, 6, 7, -1, 6, 10,
    -- filter=111 channel=111
    1, 1, -3, 0, -5, 9, 3, 3, -6,
    -- filter=111 channel=112
    -12, -6, -1, 9, -8, 4, 3, -19, 5,
    -- filter=111 channel=113
    4, -8, 0, 6, -17, 5, 10, -18, 7,
    -- filter=111 channel=114
    13, -16, 11, 17, -44, 2, 11, -15, 2,
    -- filter=111 channel=115
    5, 2, -3, -4, 2, 6, 0, -5, -4,
    -- filter=111 channel=116
    -2, -8, 7, 16, -31, 11, 11, -6, 4,
    -- filter=111 channel=117
    -2, -5, 8, 0, -12, 9, -5, 0, 7,
    -- filter=111 channel=118
    -2, 0, 0, -7, -6, 0, -7, 0, 0,
    -- filter=111 channel=119
    9, 31, -8, 15, 44, -6, 23, 36, -3,
    -- filter=111 channel=120
    -15, -2, -8, 11, -22, -5, 10, -35, 3,
    -- filter=111 channel=121
    2, 3, -8, 12, 0, 14, 9, 6, 3,
    -- filter=111 channel=122
    0, -8, -13, 15, -27, 9, 24, -8, 3,
    -- filter=111 channel=123
    9, 11, 0, 12, 24, -5, 14, 5, 1,
    -- filter=111 channel=124
    -4, 6, 0, -1, -6, -2, -2, -9, -2,
    -- filter=111 channel=125
    -3, -2, -1, 15, -20, 11, 15, -20, 0,
    -- filter=111 channel=126
    3, -6, -3, 10, -9, 14, 10, -4, 1,
    -- filter=111 channel=127
    1, 8, -3, 7, 12, 13, 1, 0, 12,
    -- filter=112 channel=0
    -13, 3, 6, -10, 29, 16, -10, 5, 7,
    -- filter=112 channel=1
    -9, 8, -2, 3, 33, 11, -4, 8, -4,
    -- filter=112 channel=2
    1, -3, 3, 0, -7, -8, -7, -8, -4,
    -- filter=112 channel=3
    1, 10, -1, -3, 0, 7, -1, 0, 2,
    -- filter=112 channel=4
    0, 0, 2, -6, -7, -4, -3, 2, -2,
    -- filter=112 channel=5
    -3, 13, -4, -5, 30, 15, -14, 9, -4,
    -- filter=112 channel=6
    6, 8, -4, -1, 5, 3, -6, -6, -4,
    -- filter=112 channel=7
    -6, -6, 0, -6, 5, 2, 1, -5, -5,
    -- filter=112 channel=8
    0, -5, -4, 3, 4, 1, -3, -3, -4,
    -- filter=112 channel=9
    5, 4, 0, 4, 10, 6, -5, 6, -3,
    -- filter=112 channel=10
    7, -6, -8, 3, -6, -1, 0, 2, -8,
    -- filter=112 channel=11
    4, -2, -4, 6, -8, -1, 0, -1, 9,
    -- filter=112 channel=12
    0, 1, 6, -7, -6, 5, 6, 0, 5,
    -- filter=112 channel=13
    4, -12, 3, 5, -4, 0, -5, -5, 0,
    -- filter=112 channel=14
    1, 4, -1, -1, 3, -7, -3, 4, 2,
    -- filter=112 channel=15
    -7, 3, -8, 7, -5, -4, 2, -8, 1,
    -- filter=112 channel=16
    0, 1, 0, 10, 9, -3, -1, 2, -10,
    -- filter=112 channel=17
    -1, 1, 2, -3, -7, -4, -4, 2, 2,
    -- filter=112 channel=18
    -3, 0, 4, 7, 7, 5, -3, -3, -11,
    -- filter=112 channel=19
    4, -2, -2, 1, -2, 3, -2, -1, 0,
    -- filter=112 channel=20
    7, 2, 0, 9, -3, 0, 5, 4, 6,
    -- filter=112 channel=21
    4, -2, -5, 12, 0, -10, 4, -4, -3,
    -- filter=112 channel=22
    3, 7, 2, 0, 11, -1, 4, -3, -7,
    -- filter=112 channel=23
    4, -8, -1, 10, -12, -3, 2, 0, 0,
    -- filter=112 channel=24
    2, -6, 1, -5, 0, -6, -7, 2, -1,
    -- filter=112 channel=25
    6, -5, -7, -3, 2, 5, 0, 3, -7,
    -- filter=112 channel=26
    5, 7, 0, 9, 1, 8, -7, -4, 0,
    -- filter=112 channel=27
    -1, 4, -3, 3, 4, 8, -8, -1, -10,
    -- filter=112 channel=28
    3, -6, -4, 3, -1, -6, -6, -2, 4,
    -- filter=112 channel=29
    10, -4, 2, 5, -5, -5, 11, -5, 0,
    -- filter=112 channel=30
    -9, 5, -4, -6, 9, 11, -12, 6, 2,
    -- filter=112 channel=31
    6, -19, -18, -2, -15, -8, -7, -7, -2,
    -- filter=112 channel=32
    -2, 2, 2, -1, 7, 7, -3, -1, -3,
    -- filter=112 channel=33
    -3, -3, -8, 7, 2, 2, -3, -2, -8,
    -- filter=112 channel=34
    5, 6, 5, 7, -6, 1, 9, -1, 6,
    -- filter=112 channel=35
    6, 0, -1, 2, 5, 3, 0, 0, 4,
    -- filter=112 channel=36
    9, -9, 4, 0, -14, -8, -5, -9, 4,
    -- filter=112 channel=37
    -7, 10, 12, 3, 32, 25, -6, -2, -7,
    -- filter=112 channel=38
    6, 4, -10, 3, -6, -3, -2, -1, -1,
    -- filter=112 channel=39
    11, 3, 5, -5, 1, -2, 5, 6, 6,
    -- filter=112 channel=40
    2, -6, -4, 5, 2, -7, 6, -3, 6,
    -- filter=112 channel=41
    11, -4, 4, 5, -11, -15, 10, 1, -3,
    -- filter=112 channel=42
    -6, 0, -2, 0, 13, 11, -12, -2, 5,
    -- filter=112 channel=43
    0, 2, 0, 0, -8, -7, 8, 1, 7,
    -- filter=112 channel=44
    -7, 5, 3, 4, 20, 1, -12, -1, -2,
    -- filter=112 channel=45
    4, 4, -3, -6, 0, 10, 5, 0, 0,
    -- filter=112 channel=46
    4, 3, 2, 6, 10, -3, 1, -2, -5,
    -- filter=112 channel=47
    0, 8, -2, 8, 11, 0, 5, 9, 0,
    -- filter=112 channel=48
    -4, -1, 4, 3, 14, 8, -5, -8, -15,
    -- filter=112 channel=49
    -4, 3, -3, 5, 5, 3, -6, -2, -3,
    -- filter=112 channel=50
    -8, -3, 0, -5, -7, 2, -8, -5, -3,
    -- filter=112 channel=51
    7, 3, -2, 6, -2, -1, -4, 7, 2,
    -- filter=112 channel=52
    13, -5, -7, 10, -5, 3, 1, -5, 3,
    -- filter=112 channel=53
    1, -2, 3, 0, -5, -3, 7, 6, 4,
    -- filter=112 channel=54
    -6, 0, 5, -2, -6, -6, 0, 4, -1,
    -- filter=112 channel=55
    2, -11, -13, 8, -9, -14, -1, -9, 0,
    -- filter=112 channel=56
    3, -5, -8, 2, -7, 4, 7, 5, -4,
    -- filter=112 channel=57
    7, -2, -4, 3, 1, -8, 0, -3, 2,
    -- filter=112 channel=58
    -11, 9, 1, 3, 21, 14, -1, 11, 9,
    -- filter=112 channel=59
    -5, 2, -11, 7, 0, 0, -9, 0, -2,
    -- filter=112 channel=60
    -2, 0, -4, 0, 4, -6, 0, 3, 5,
    -- filter=112 channel=61
    6, -5, -2, 1, -1, -4, -4, -1, -8,
    -- filter=112 channel=62
    7, -6, -4, -6, -6, 5, 4, 0, 3,
    -- filter=112 channel=63
    -2, 6, -4, -2, 4, 9, -10, 7, -2,
    -- filter=112 channel=64
    -1, -6, -4, 6, -2, 0, 5, -6, 5,
    -- filter=112 channel=65
    -2, 4, -2, -1, -3, 1, -4, 7, 5,
    -- filter=112 channel=66
    2, -2, 0, 0, -10, -10, 6, -8, -8,
    -- filter=112 channel=67
    5, -3, -3, 2, 1, -7, 7, -2, 6,
    -- filter=112 channel=68
    -3, -4, -1, -2, -1, 3, 1, -2, 7,
    -- filter=112 channel=69
    -2, 5, -3, 6, 0, 6, -4, -3, -7,
    -- filter=112 channel=70
    -2, 0, 0, 2, -1, 6, -4, -10, 0,
    -- filter=112 channel=71
    -1, 6, -1, -3, -1, -9, -3, 5, 8,
    -- filter=112 channel=72
    -4, -7, -10, 6, -16, -11, 2, -2, -3,
    -- filter=112 channel=73
    2, -9, -5, 2, -8, -4, 0, 1, -2,
    -- filter=112 channel=74
    2, -3, 3, 6, -12, -1, 5, -10, 0,
    -- filter=112 channel=75
    -19, 5, 0, -3, 36, 18, -13, 18, -9,
    -- filter=112 channel=76
    13, 0, -4, 12, -10, -7, 5, -4, 11,
    -- filter=112 channel=77
    -1, 0, -5, -5, -6, -6, 2, -4, -7,
    -- filter=112 channel=78
    -1, 8, 5, -3, 8, 7, -8, -5, -7,
    -- filter=112 channel=79
    0, 3, 0, -1, -1, 12, 0, -6, -5,
    -- filter=112 channel=80
    6, -3, -16, 10, 3, 1, -5, -5, -16,
    -- filter=112 channel=81
    6, 5, 1, 2, 7, 0, -7, 5, -5,
    -- filter=112 channel=82
    0, -3, -6, 4, 4, 5, 1, -3, 6,
    -- filter=112 channel=83
    6, 6, -5, -1, -1, -1, 2, 4, 1,
    -- filter=112 channel=84
    -5, 0, -1, 4, -1, -4, -8, 2, -7,
    -- filter=112 channel=85
    -3, 5, -3, -3, -3, 1, 5, -3, 2,
    -- filter=112 channel=86
    -2, 6, 6, -8, 12, 2, 2, 7, 3,
    -- filter=112 channel=87
    9, -6, 0, 5, -4, -6, 0, 6, 2,
    -- filter=112 channel=88
    11, 0, 0, 2, -10, -12, -1, 0, -2,
    -- filter=112 channel=89
    8, -2, -9, -5, -17, -11, -9, -16, -10,
    -- filter=112 channel=90
    14, 0, -6, 9, -12, -9, 10, 1, 1,
    -- filter=112 channel=91
    1, -5, -2, 0, -3, 0, -6, -1, 1,
    -- filter=112 channel=92
    -6, 0, 1, -3, 3, -7, 5, -6, 1,
    -- filter=112 channel=93
    -2, 3, -1, -1, 15, 12, -7, -7, -10,
    -- filter=112 channel=94
    5, -4, -2, 3, 6, 4, 0, -2, -1,
    -- filter=112 channel=95
    7, -2, 1, 0, 5, 1, 4, -1, -6,
    -- filter=112 channel=96
    -8, 4, -3, -6, -3, 4, 2, 2, 6,
    -- filter=112 channel=97
    -1, 7, -2, -5, 5, 0, 1, 11, 7,
    -- filter=112 channel=98
    0, -2, -6, 3, 10, 9, 2, -6, -3,
    -- filter=112 channel=99
    15, -14, -14, 5, -21, -10, 1, -16, -9,
    -- filter=112 channel=100
    3, 0, 0, 3, 2, 4, 7, 0, -8,
    -- filter=112 channel=101
    12, 5, 3, -3, 2, -6, -4, -1, -6,
    -- filter=112 channel=102
    3, 3, 7, -4, -7, -7, 0, 1, 6,
    -- filter=112 channel=103
    2, 0, -4, 8, 20, 7, 0, 5, 1,
    -- filter=112 channel=104
    10, 0, -8, 0, 2, -12, -7, -10, -10,
    -- filter=112 channel=105
    10, 0, -2, 10, -1, -3, 8, 4, 5,
    -- filter=112 channel=106
    -1, -1, -3, 7, 1, 2, 3, -1, 3,
    -- filter=112 channel=107
    2, 0, 2, 4, -9, 8, 5, -6, 7,
    -- filter=112 channel=108
    3, 10, 5, -4, -2, -5, 1, 9, -3,
    -- filter=112 channel=109
    6, 3, -4, 3, 3, -7, -9, -10, -13,
    -- filter=112 channel=110
    7, -5, 0, -4, -12, -10, 0, -6, 6,
    -- filter=112 channel=111
    3, 1, -4, -3, -1, -10, 1, 7, -2,
    -- filter=112 channel=112
    3, 6, 0, -3, 5, 3, 4, -1, -4,
    -- filter=112 channel=113
    -2, -9, -10, 8, 4, -5, 5, -1, 1,
    -- filter=112 channel=114
    -12, 2, 4, 5, 17, 20, -14, -7, -1,
    -- filter=112 channel=115
    2, -6, 0, -5, 6, 2, 2, 2, -5,
    -- filter=112 channel=116
    6, -4, -12, 1, -8, 1, -11, -12, -2,
    -- filter=112 channel=117
    -4, -6, -1, -6, 4, 4, -8, -8, -1,
    -- filter=112 channel=118
    6, 3, 0, -5, 6, 4, -5, -4, 6,
    -- filter=112 channel=119
    1, -5, 4, 9, 0, -6, 4, -3, 2,
    -- filter=112 channel=120
    1, -8, -2, 5, -1, -1, -3, -6, -2,
    -- filter=112 channel=121
    -3, -5, 0, -2, 2, -10, 7, -6, -3,
    -- filter=112 channel=122
    18, 4, -2, 18, 11, 0, 11, 1, -2,
    -- filter=112 channel=123
    8, -2, -3, 5, -4, -8, 5, 0, 5,
    -- filter=112 channel=124
    3, -4, 4, 9, 1, -6, 0, 0, 1,
    -- filter=112 channel=125
    3, -12, -11, 1, -5, -1, -5, -11, -9,
    -- filter=112 channel=126
    -4, -5, -9, 4, 5, -4, -3, -3, -10,
    -- filter=112 channel=127
    0, -2, 2, 8, -8, 2, 6, -5, 2,
    -- filter=113 channel=0
    -6, -13, 20, -19, -17, 21, -15, -16, 10,
    -- filter=113 channel=1
    -3, -2, 16, -4, 0, 9, -18, -3, 10,
    -- filter=113 channel=2
    0, -4, 5, -5, -3, -8, -6, 0, 0,
    -- filter=113 channel=3
    -10, -1, 1, 4, 3, 0, 3, 0, 4,
    -- filter=113 channel=4
    -5, 1, -1, -12, -3, -9, 0, -9, 5,
    -- filter=113 channel=5
    -1, 0, 6, -4, -1, 12, -18, -4, 0,
    -- filter=113 channel=6
    -6, -2, 2, -3, -3, -3, -7, -5, 4,
    -- filter=113 channel=7
    6, 6, -2, 6, -1, 4, 6, -4, -3,
    -- filter=113 channel=8
    4, 8, -5, 7, 2, 2, -4, -4, -8,
    -- filter=113 channel=9
    2, -5, -3, -5, 6, 3, 1, 1, 1,
    -- filter=113 channel=10
    1, 12, -10, 9, 15, -9, -1, -3, -9,
    -- filter=113 channel=11
    5, -1, -9, 9, -3, -9, -2, -4, 1,
    -- filter=113 channel=12
    6, 0, -2, -1, 0, 7, 7, 7, 1,
    -- filter=113 channel=13
    -1, 8, 1, 4, 2, 0, 9, 5, -3,
    -- filter=113 channel=14
    6, -2, 4, -4, 0, -3, 4, -1, -4,
    -- filter=113 channel=15
    4, 0, 13, 6, 0, 7, -7, -1, 0,
    -- filter=113 channel=16
    -4, 7, -3, 2, 17, -2, 1, 1, 5,
    -- filter=113 channel=17
    0, 0, 5, -4, -7, -4, -2, 3, 4,
    -- filter=113 channel=18
    0, 0, 14, -7, -11, 3, -14, -17, 1,
    -- filter=113 channel=19
    -3, 1, -2, -6, -4, 3, -5, 4, 7,
    -- filter=113 channel=20
    6, 7, 0, 11, 4, -8, 10, 4, 0,
    -- filter=113 channel=21
    9, 14, -19, 4, 12, -13, 4, 5, 4,
    -- filter=113 channel=22
    2, -8, 12, 1, -6, 5, -6, -1, -1,
    -- filter=113 channel=23
    7, 1, 11, 9, -5, 2, 5, -4, 0,
    -- filter=113 channel=24
    3, -6, -1, -4, 6, 5, -1, 0, -1,
    -- filter=113 channel=25
    4, 0, -3, -4, 3, -3, -10, -9, -2,
    -- filter=113 channel=26
    -1, 2, 1, -8, 1, -11, -1, 4, 6,
    -- filter=113 channel=27
    0, -3, 9, 0, -5, 15, -7, -20, 7,
    -- filter=113 channel=28
    -3, 7, -5, -3, 4, -6, -3, 7, 5,
    -- filter=113 channel=29
    -4, -2, -4, 7, 0, -7, -4, -6, -13,
    -- filter=113 channel=30
    -5, -4, 8, 4, -8, -1, 0, 0, 0,
    -- filter=113 channel=31
    13, 7, -17, 19, 9, -12, 0, -2, -7,
    -- filter=113 channel=32
    -1, -2, 7, 1, -10, 14, -9, -14, -2,
    -- filter=113 channel=33
    -2, -6, 16, -2, -9, 20, -8, -2, 8,
    -- filter=113 channel=34
    5, 2, 1, 21, 0, -7, 12, 6, -1,
    -- filter=113 channel=35
    1, -6, 0, -7, 4, -6, -5, 1, 2,
    -- filter=113 channel=36
    13, 12, -13, 15, 14, -9, 17, 6, -8,
    -- filter=113 channel=37
    1, 0, 6, -14, 0, 14, -13, -11, 7,
    -- filter=113 channel=38
    3, -3, 3, 2, 5, 1, -3, -6, 0,
    -- filter=113 channel=39
    5, 4, 1, -2, -3, -7, 4, -6, 1,
    -- filter=113 channel=40
    5, 8, 0, 2, 4, 8, -3, 0, 8,
    -- filter=113 channel=41
    6, 3, 5, 8, 12, -17, 8, 2, -7,
    -- filter=113 channel=42
    1, 0, 4, -7, 5, -3, -7, -7, 7,
    -- filter=113 channel=43
    0, 2, 6, -5, 2, 10, -9, -4, -5,
    -- filter=113 channel=44
    0, 5, 2, -2, 1, 2, 0, -7, 3,
    -- filter=113 channel=45
    -5, 5, 8, -2, -1, 1, 4, -3, 9,
    -- filter=113 channel=46
    -1, 9, 5, -1, 0, -3, -6, 4, 0,
    -- filter=113 channel=47
    -2, 1, -12, -1, 17, -1, -4, 9, 1,
    -- filter=113 channel=48
    3, 8, 2, 0, 6, -4, -7, 0, 3,
    -- filter=113 channel=49
    -2, 3, 5, -16, -17, -3, -9, -15, 0,
    -- filter=113 channel=50
    7, -4, 0, 9, -11, 0, 5, -8, -4,
    -- filter=113 channel=51
    -5, -5, 7, 3, -2, 0, 4, 7, 0,
    -- filter=113 channel=52
    6, 6, 2, 13, -5, 1, 0, 2, 5,
    -- filter=113 channel=53
    -4, -1, 3, -3, -1, -5, -3, 3, -6,
    -- filter=113 channel=54
    2, 0, 6, 6, 0, 5, 0, 0, 2,
    -- filter=113 channel=55
    11, 2, 1, 15, 0, -8, 5, -10, -13,
    -- filter=113 channel=56
    7, 5, 1, 7, 10, -6, -3, 2, 4,
    -- filter=113 channel=57
    2, -2, 0, 5, 4, 2, 0, 1, 2,
    -- filter=113 channel=58
    -8, -5, -2, -8, 5, -4, -11, -6, 6,
    -- filter=113 channel=59
    3, 6, 1, -1, 12, 3, -12, 0, -2,
    -- filter=113 channel=60
    -1, 2, -7, -1, 6, -5, 2, 0, 1,
    -- filter=113 channel=61
    9, 4, 0, 2, 3, -3, 9, 8, -7,
    -- filter=113 channel=62
    -7, 6, 1, 2, -3, -1, 1, 0, 0,
    -- filter=113 channel=63
    -1, 2, -10, -7, -5, -7, -4, 3, -4,
    -- filter=113 channel=64
    7, 6, -3, 0, 10, -7, 1, 11, -9,
    -- filter=113 channel=65
    6, 1, 5, 5, -3, 0, 2, 0, -1,
    -- filter=113 channel=66
    4, 8, 5, 2, 5, 4, 9, -1, 0,
    -- filter=113 channel=67
    0, 0, -6, -1, -2, -7, -2, 8, 2,
    -- filter=113 channel=68
    0, 7, -8, -6, -2, 0, 6, -8, 5,
    -- filter=113 channel=69
    -1, -1, 0, -5, 2, 3, 0, 0, -4,
    -- filter=113 channel=70
    9, 3, 16, 5, -8, 14, -7, -8, 9,
    -- filter=113 channel=71
    4, 1, 6, 6, 5, 0, -2, -1, -3,
    -- filter=113 channel=72
    9, -1, -11, 14, 6, -19, -1, 4, -15,
    -- filter=113 channel=73
    0, 2, 2, -3, -6, 5, 5, -11, -12,
    -- filter=113 channel=74
    11, -4, 11, 15, -4, -7, -3, -8, -6,
    -- filter=113 channel=75
    1, -1, 12, -5, -3, 22, -17, 0, 4,
    -- filter=113 channel=76
    8, 11, 8, 0, 7, 0, 11, 1, 6,
    -- filter=113 channel=77
    4, -5, -1, 0, -6, -7, -3, 4, 0,
    -- filter=113 channel=78
    -7, 1, -6, 6, 2, 0, 1, 1, 2,
    -- filter=113 channel=79
    -9, 0, 16, -5, -13, 25, -22, -20, 3,
    -- filter=113 channel=80
    1, 2, -22, 1, 7, -18, -8, 6, -6,
    -- filter=113 channel=81
    4, 2, -4, 7, 6, 1, -3, 2, -1,
    -- filter=113 channel=82
    -6, 6, 5, -2, 5, 7, -2, 5, -1,
    -- filter=113 channel=83
    -6, 0, 1, -8, 2, 2, -7, 2, 2,
    -- filter=113 channel=84
    -1, -5, 1, -9, 0, -3, 0, -12, -1,
    -- filter=113 channel=85
    -3, 5, -7, 5, -3, 5, -7, 6, 2,
    -- filter=113 channel=86
    -3, -3, 0, -2, 1, 5, 2, 5, 8,
    -- filter=113 channel=87
    8, -5, 7, 9, 0, 5, 9, -5, 0,
    -- filter=113 channel=88
    13, 9, -9, 12, 13, -7, 16, 3, -2,
    -- filter=113 channel=89
    0, -7, -11, 7, 8, -10, -4, -11, -5,
    -- filter=113 channel=90
    4, 15, -12, 24, 11, -9, 17, 19, -6,
    -- filter=113 channel=91
    -3, -4, 11, 1, -3, 4, -5, -16, -5,
    -- filter=113 channel=92
    -2, 4, 6, 0, 6, 6, 3, -3, 5,
    -- filter=113 channel=93
    3, -5, -7, -10, 1, -3, -6, 0, 4,
    -- filter=113 channel=94
    5, -4, 7, -6, 0, -5, -7, -2, 7,
    -- filter=113 channel=95
    4, -4, -6, -3, 6, 1, 0, -2, 4,
    -- filter=113 channel=96
    -7, 0, 4, -5, -4, 2, -4, -4, 0,
    -- filter=113 channel=97
    5, 1, 1, 6, -1, 0, 1, 9, -4,
    -- filter=113 channel=98
    0, -6, 0, 6, -11, -7, -8, -4, -10,
    -- filter=113 channel=99
    4, -2, -16, 23, 3, -17, 13, 0, -15,
    -- filter=113 channel=100
    8, 9, -1, -4, 12, -1, 1, 8, 1,
    -- filter=113 channel=101
    -3, -6, -8, 2, -6, -10, 0, -8, 3,
    -- filter=113 channel=102
    0, -4, -4, 4, 6, 3, 0, 0, -1,
    -- filter=113 channel=103
    0, 7, -8, 4, 8, -9, -10, -2, 2,
    -- filter=113 channel=104
    9, 5, -21, 2, 12, -15, -7, 1, -5,
    -- filter=113 channel=105
    -6, -4, -3, 0, 8, 0, 6, -3, 4,
    -- filter=113 channel=106
    0, 7, 0, 7, 1, 2, 4, 11, 1,
    -- filter=113 channel=107
    2, 4, 7, -6, -2, 4, -2, 0, 3,
    -- filter=113 channel=108
    -7, 7, 3, -8, 0, 4, 5, 7, -9,
    -- filter=113 channel=109
    -3, -1, 11, 0, -3, 6, -6, -12, -3,
    -- filter=113 channel=110
    8, -2, -6, 15, 9, -8, 1, 0, -7,
    -- filter=113 channel=111
    -2, 7, -4, -5, -1, -1, 5, 6, 4,
    -- filter=113 channel=112
    -5, -5, 8, -3, -8, 1, -12, -8, -1,
    -- filter=113 channel=113
    5, -1, 5, 1, 7, 2, -8, -2, 0,
    -- filter=113 channel=114
    -19, -19, 24, -26, -30, 17, -31, -31, 3,
    -- filter=113 channel=115
    -2, -3, -7, 7, -3, -4, 2, -2, 6,
    -- filter=113 channel=116
    -4, 4, 1, 2, -8, -11, 0, -4, -10,
    -- filter=113 channel=117
    6, 5, 3, 0, 1, -4, -2, 4, 0,
    -- filter=113 channel=118
    -2, 1, 1, -5, -1, -2, 3, -3, 4,
    -- filter=113 channel=119
    5, 0, 11, 8, 10, -1, 5, 3, 8,
    -- filter=113 channel=120
    2, 0, 0, 2, -17, -3, -8, -9, -14,
    -- filter=113 channel=121
    5, 0, -10, 3, 8, 0, 4, 0, -1,
    -- filter=113 channel=122
    1, 9, -13, 13, 27, -16, 3, 17, -5,
    -- filter=113 channel=123
    10, -1, 9, 14, 4, -7, 8, 3, 4,
    -- filter=113 channel=124
    4, -2, 4, 0, 4, 0, 5, 6, 2,
    -- filter=113 channel=125
    -3, 6, -11, 0, 6, -11, 4, -4, -14,
    -- filter=113 channel=126
    0, -7, -4, 2, -1, -9, -4, -2, -8,
    -- filter=113 channel=127
    2, 1, 6, -4, 1, -4, 9, 8, -4,
    -- filter=114 channel=0
    4, -4, 1, 4, 3, -4, 8, 5, -3,
    -- filter=114 channel=1
    -1, -8, 2, -11, -6, -12, -4, 0, -8,
    -- filter=114 channel=2
    7, -4, -3, -5, 7, 3, -8, 2, 0,
    -- filter=114 channel=3
    0, 0, 9, 6, 1, 8, 2, 0, 0,
    -- filter=114 channel=4
    1, -3, -1, -11, -10, -7, -6, -4, 6,
    -- filter=114 channel=5
    -5, -3, -5, 0, -7, -10, 0, 2, -7,
    -- filter=114 channel=6
    8, 4, -1, 5, -5, 2, 6, 0, -2,
    -- filter=114 channel=7
    0, -4, 2, 2, -2, -5, -2, 5, 0,
    -- filter=114 channel=8
    4, 7, 0, 2, -2, 2, -7, -8, 3,
    -- filter=114 channel=9
    -5, -5, 6, -9, 0, 5, -10, 4, -1,
    -- filter=114 channel=10
    -2, -8, 5, 1, 4, -2, -4, 2, -2,
    -- filter=114 channel=11
    -2, 4, 8, -4, 3, 0, 1, 2, 11,
    -- filter=114 channel=12
    0, 4, -5, -3, 7, 5, -2, -2, 0,
    -- filter=114 channel=13
    -3, 1, 0, -7, 10, -4, -19, -7, -5,
    -- filter=114 channel=14
    -6, 5, 2, 1, 2, 0, 4, 0, 1,
    -- filter=114 channel=15
    -6, 4, 2, 2, 5, 0, -17, -2, -4,
    -- filter=114 channel=16
    1, 2, 2, 0, 8, 7, -1, 3, -5,
    -- filter=114 channel=17
    -6, 2, -3, -5, 5, 3, -5, 2, 6,
    -- filter=114 channel=18
    -17, -5, 7, -10, -4, 0, -25, -12, -6,
    -- filter=114 channel=19
    -4, -3, 3, 4, 2, 0, 5, 2, 2,
    -- filter=114 channel=20
    8, 7, 14, 14, 11, 12, 9, 11, 9,
    -- filter=114 channel=21
    3, 0, 6, -6, 10, 0, 3, 2, 0,
    -- filter=114 channel=22
    2, -3, 3, 0, 2, -7, 0, 0, -4,
    -- filter=114 channel=23
    -4, 10, 5, 13, 7, 2, -7, 10, -8,
    -- filter=114 channel=24
    6, -2, 1, 0, -6, -3, 6, -1, 7,
    -- filter=114 channel=25
    0, 0, 4, -8, 11, -1, -21, -14, -9,
    -- filter=114 channel=26
    8, 2, 5, -1, 7, -5, 9, 0, 9,
    -- filter=114 channel=27
    -10, 11, 4, -12, 4, -8, -34, -18, -16,
    -- filter=114 channel=28
    -1, -2, 6, 1, 5, 0, 0, 1, 6,
    -- filter=114 channel=29
    0, 11, 12, -4, 13, 8, -3, 6, 5,
    -- filter=114 channel=30
    0, 7, 3, 0, 3, -2, -6, -7, -8,
    -- filter=114 channel=31
    3, 9, 11, 5, 17, 0, -11, 10, 0,
    -- filter=114 channel=32
    -9, -3, -5, -14, 8, -5, -25, -7, -3,
    -- filter=114 channel=33
    -7, 5, -3, -3, 10, -1, -20, 1, -7,
    -- filter=114 channel=34
    6, 2, -2, 7, 5, -4, -4, 8, 4,
    -- filter=114 channel=35
    6, 1, 3, 0, 6, 3, 5, 6, 4,
    -- filter=114 channel=36
    2, 8, 2, 2, 7, 0, 6, 6, 7,
    -- filter=114 channel=37
    7, 3, -7, -3, 2, -12, -9, -14, 0,
    -- filter=114 channel=38
    -4, 5, 5, 0, 3, 4, -1, 0, -6,
    -- filter=114 channel=39
    -3, 2, 8, 0, 11, 8, 4, 9, 8,
    -- filter=114 channel=40
    1, 0, 12, 2, 9, 0, 10, 13, 5,
    -- filter=114 channel=41
    -4, -7, 3, -10, -5, 1, -2, -12, 4,
    -- filter=114 channel=42
    -7, 0, -6, 3, 0, -6, -8, 2, 0,
    -- filter=114 channel=43
    6, 0, 9, 4, 0, -2, -1, 10, 0,
    -- filter=114 channel=44
    0, -2, -1, 2, 0, -11, -13, 3, -10,
    -- filter=114 channel=45
    0, -2, 6, -1, 9, 7, 3, -3, 9,
    -- filter=114 channel=46
    0, 4, 7, 0, 2, 2, -4, 4, 6,
    -- filter=114 channel=47
    -9, -5, 5, -12, -2, 5, -6, 2, -7,
    -- filter=114 channel=48
    0, 2, 0, -5, 9, -3, -23, -2, -11,
    -- filter=114 channel=49
    1, 0, -1, -3, -8, -8, -13, -3, -11,
    -- filter=114 channel=50
    0, 5, 2, 0, -2, 0, -6, -7, -3,
    -- filter=114 channel=51
    -7, 3, -2, -6, 5, 5, 2, -5, 5,
    -- filter=114 channel=52
    0, 3, -2, 7, 5, -4, 4, 4, 4,
    -- filter=114 channel=53
    -6, 4, 5, 0, -1, -1, 3, 0, -1,
    -- filter=114 channel=54
    3, -3, -7, 6, 4, -4, 6, 5, -6,
    -- filter=114 channel=55
    -10, 5, -1, -8, 2, 8, -18, -4, -4,
    -- filter=114 channel=56
    -3, -3, -2, 2, 5, 6, -7, 5, -2,
    -- filter=114 channel=57
    4, 1, -4, -2, -4, -6, -5, -1, -3,
    -- filter=114 channel=58
    3, 7, -7, 2, -5, -3, 0, 7, -7,
    -- filter=114 channel=59
    -10, 6, 9, -12, 11, -3, -26, -12, -10,
    -- filter=114 channel=60
    -2, 0, 7, -6, 6, 1, 1, 2, 5,
    -- filter=114 channel=61
    4, 0, 2, 8, 9, -5, -5, 9, 7,
    -- filter=114 channel=62
    -6, 2, 6, -2, -2, -4, -4, 0, -3,
    -- filter=114 channel=63
    -1, -4, 2, 2, 7, 0, 0, -4, 0,
    -- filter=114 channel=64
    -4, -3, 3, 5, 10, 2, 2, 6, 4,
    -- filter=114 channel=65
    -5, -3, 3, -2, -5, 0, 2, 0, -5,
    -- filter=114 channel=66
    -2, -8, 7, 5, 5, -5, -9, 5, -1,
    -- filter=114 channel=67
    -2, 6, 0, 0, 8, 7, 6, -1, -4,
    -- filter=114 channel=68
    0, 1, 0, 6, 4, 6, -2, -1, 3,
    -- filter=114 channel=69
    -6, -3, -7, -4, 5, 0, 5, 0, 1,
    -- filter=114 channel=70
    -5, 3, -5, 6, 5, -1, -10, -7, -2,
    -- filter=114 channel=71
    -3, -4, 0, 7, 8, 10, 9, 4, 5,
    -- filter=114 channel=72
    -3, 7, 0, -6, 8, 8, -20, 7, 2,
    -- filter=114 channel=73
    -12, 3, 1, -1, 9, -11, -20, -14, -2,
    -- filter=114 channel=74
    0, 12, 2, 4, 7, 0, -3, 6, -11,
    -- filter=114 channel=75
    -8, -3, -2, -4, -2, -11, -14, -11, -10,
    -- filter=114 channel=76
    6, 11, 3, 2, 16, 12, 5, 14, 2,
    -- filter=114 channel=77
    0, 1, 1, 1, -7, -2, 6, 5, -2,
    -- filter=114 channel=78
    -3, 4, 3, 8, 4, -1, -4, 1, 4,
    -- filter=114 channel=79
    -15, -7, -1, -19, -1, -4, -31, -6, -9,
    -- filter=114 channel=80
    -8, 7, 5, -10, 10, 4, -23, -1, -1,
    -- filter=114 channel=81
    7, 4, -6, -3, 6, -3, -2, 3, -5,
    -- filter=114 channel=82
    -1, -4, 5, 7, 8, -5, 1, 3, 5,
    -- filter=114 channel=83
    -4, 4, -1, -8, -1, 0, -7, 0, 0,
    -- filter=114 channel=84
    -7, -6, -6, -3, -4, -1, -8, -5, -11,
    -- filter=114 channel=85
    -3, -2, 0, -7, 6, 3, -4, 6, -3,
    -- filter=114 channel=86
    -6, -5, 6, 1, -4, 0, -1, 7, -4,
    -- filter=114 channel=87
    7, 0, 7, 14, 11, 0, 3, 12, 1,
    -- filter=114 channel=88
    10, 15, 6, 14, 16, 6, 1, 4, 2,
    -- filter=114 channel=89
    -18, 2, 1, -7, 7, 6, -25, -7, -11,
    -- filter=114 channel=90
    1, 14, -1, 19, 17, 1, 12, 17, 12,
    -- filter=114 channel=91
    0, 9, -2, -10, -2, -11, -22, -18, -16,
    -- filter=114 channel=92
    0, 6, -2, 6, 2, 3, 6, 4, 4,
    -- filter=114 channel=93
    -2, -3, 2, 0, -6, -11, -13, -4, -12,
    -- filter=114 channel=94
    3, -1, -1, 5, -4, -2, 2, -5, -4,
    -- filter=114 channel=95
    -4, 1, 5, -6, 0, -2, -6, -5, 0,
    -- filter=114 channel=96
    -5, 0, 2, -4, 6, 3, -7, -4, -2,
    -- filter=114 channel=97
    9, -3, 2, 6, 7, 0, 5, 1, 8,
    -- filter=114 channel=98
    -16, 1, 1, -3, 6, 1, -20, -2, -10,
    -- filter=114 channel=99
    -4, 8, 0, 4, 17, 1, -2, 12, 0,
    -- filter=114 channel=100
    2, 4, 2, 3, -7, 0, 4, 3, 0,
    -- filter=114 channel=101
    8, 6, 4, 2, -1, -2, -3, 0, 5,
    -- filter=114 channel=102
    6, -1, 6, -1, -6, -2, 3, -1, 2,
    -- filter=114 channel=103
    2, 0, -1, -6, -4, 4, -16, 7, -1,
    -- filter=114 channel=104
    -6, 2, 11, -10, 15, -2, -8, 7, 3,
    -- filter=114 channel=105
    9, -1, 3, -1, 7, 2, 7, 13, 4,
    -- filter=114 channel=106
    0, 0, 1, -3, -4, 9, -1, 7, -2,
    -- filter=114 channel=107
    -1, 11, 3, 14, -2, 5, 1, 8, 8,
    -- filter=114 channel=108
    4, -6, 0, -5, 3, 7, -2, -3, 0,
    -- filter=114 channel=109
    -16, -2, -3, -5, 8, -10, -28, -11, -12,
    -- filter=114 channel=110
    -3, 0, 6, 8, 1, -4, 2, 6, 3,
    -- filter=114 channel=111
    -7, -5, 1, 0, 0, 1, -2, -1, -4,
    -- filter=114 channel=112
    5, 0, 4, -6, -4, -9, -6, -7, -10,
    -- filter=114 channel=113
    -6, 0, 1, -6, 5, 6, -7, -1, 4,
    -- filter=114 channel=114
    -8, -9, -4, -19, -3, -16, -17, -14, -7,
    -- filter=114 channel=115
    -5, -7, 0, 4, 6, 4, 6, -1, 0,
    -- filter=114 channel=116
    -5, 0, 7, -11, -1, -8, -24, -9, -1,
    -- filter=114 channel=117
    6, 6, 0, -5, -2, 2, -6, -4, 7,
    -- filter=114 channel=118
    -4, 2, 0, 3, -2, -7, 4, 0, 0,
    -- filter=114 channel=119
    4, 0, -6, 2, 3, 6, 6, 6, 5,
    -- filter=114 channel=120
    -1, 15, -5, 2, 13, -10, -21, -1, -5,
    -- filter=114 channel=121
    1, 0, 8, 0, 5, -1, -3, 2, 4,
    -- filter=114 channel=122
    2, 7, -2, 0, 9, -3, -14, 7, -9,
    -- filter=114 channel=123
    -4, 0, 3, 1, 7, 1, 4, 4, 4,
    -- filter=114 channel=124
    4, 2, -3, 4, 7, 4, -1, -3, 1,
    -- filter=114 channel=125
    -2, 7, 2, -13, 14, 6, -14, -2, -9,
    -- filter=114 channel=126
    -10, -5, 9, -5, 3, -1, 0, -1, -2,
    -- filter=114 channel=127
    1, -6, 6, -1, -6, 7, -4, 0, 5,
    -- filter=115 channel=0
    -5, -20, -6, -19, -13, -9, -9, -13, 8,
    -- filter=115 channel=1
    -4, -22, -10, -23, -19, 0, -7, -11, 3,
    -- filter=115 channel=2
    -1, -4, 4, -2, 4, 8, -2, -3, 11,
    -- filter=115 channel=3
    -8, -4, 0, -18, -5, -8, -17, -4, 1,
    -- filter=115 channel=4
    -5, -2, -5, -7, -3, 1, -1, -6, 7,
    -- filter=115 channel=5
    -7, -4, 10, -16, -9, 7, 0, -2, 13,
    -- filter=115 channel=6
    4, 0, -5, 6, 5, 3, -5, 2, -4,
    -- filter=115 channel=7
    0, -2, 5, -2, -2, -7, -5, -2, -3,
    -- filter=115 channel=8
    3, -12, -2, 6, -5, -1, -3, -3, 4,
    -- filter=115 channel=9
    0, -7, 4, 0, -5, 9, 5, 5, 4,
    -- filter=115 channel=10
    0, 6, -4, 1, 0, -7, 0, 1, 0,
    -- filter=115 channel=11
    2, 9, -6, 11, 12, 3, -1, -4, -9,
    -- filter=115 channel=12
    -1, -6, -2, -5, -1, 0, 6, -9, -3,
    -- filter=115 channel=13
    -4, 4, -10, -7, 6, -4, 6, 0, -8,
    -- filter=115 channel=14
    7, -2, 4, 0, 5, 3, 3, -3, 5,
    -- filter=115 channel=15
    -3, 0, -8, 6, 15, -10, 6, -5, -10,
    -- filter=115 channel=16
    -6, -6, 4, -9, -7, 5, -4, 0, 7,
    -- filter=115 channel=17
    -5, 4, 3, -2, 5, 0, 0, -4, -3,
    -- filter=115 channel=18
    7, 6, -19, 9, 10, -10, 0, 7, -15,
    -- filter=115 channel=19
    7, 5, 0, -1, 4, 5, 0, -7, -7,
    -- filter=115 channel=20
    -4, 15, -2, 13, 23, 0, -8, -10, -9,
    -- filter=115 channel=21
    -11, -2, 11, -14, 0, 15, -6, 0, 22,
    -- filter=115 channel=22
    3, -1, 0, -3, -2, 0, 3, -5, -1,
    -- filter=115 channel=23
    9, -7, -9, 9, 8, -13, 7, 0, -4,
    -- filter=115 channel=24
    -7, -2, -5, -1, -2, 7, -1, -1, -6,
    -- filter=115 channel=25
    1, -9, -2, -5, 0, -9, 1, 10, 7,
    -- filter=115 channel=26
    0, -4, 0, -12, 0, 4, -7, 1, 2,
    -- filter=115 channel=27
    -2, 0, -18, 10, -2, -7, 15, 8, 11,
    -- filter=115 channel=28
    -6, -2, 3, -4, 3, -1, 0, 5, -2,
    -- filter=115 channel=29
    7, 22, 4, 13, 21, -5, -4, 0, -13,
    -- filter=115 channel=30
    -2, -4, 1, -3, 0, -3, 5, 1, 5,
    -- filter=115 channel=31
    -2, -1, -8, -3, 1, 5, 3, 11, 12,
    -- filter=115 channel=32
    -4, -1, -13, 0, 12, -7, 4, 10, -11,
    -- filter=115 channel=33
    8, -2, -7, -3, 0, -12, -4, 4, 0,
    -- filter=115 channel=34
    0, -8, -8, 3, -10, -14, -3, -4, -6,
    -- filter=115 channel=35
    1, 4, 2, -4, 0, 1, -7, 1, -3,
    -- filter=115 channel=36
    -2, 7, 5, -3, -1, 7, -3, 4, -2,
    -- filter=115 channel=37
    -13, -12, 2, -23, -21, -7, -4, -8, 9,
    -- filter=115 channel=38
    1, 0, 1, 1, 8, 3, 5, 6, 3,
    -- filter=115 channel=39
    0, 9, -6, 9, 7, 0, -4, 4, -8,
    -- filter=115 channel=40
    -4, -3, 4, 0, 0, 0, -3, -1, -5,
    -- filter=115 channel=41
    -1, -2, -6, -1, -8, -8, -1, -9, -11,
    -- filter=115 channel=42
    4, -3, -1, -6, -1, -4, 3, 2, 4,
    -- filter=115 channel=43
    2, 2, -6, 4, -8, -12, -7, 0, 1,
    -- filter=115 channel=44
    -16, -2, 6, -16, -16, 4, -5, 6, 10,
    -- filter=115 channel=45
    3, 0, 2, 2, 6, 2, 3, 2, 4,
    -- filter=115 channel=46
    5, 0, -3, -2, -1, -3, 2, -1, 3,
    -- filter=115 channel=47
    -6, -4, 8, -11, -13, 3, -1, 10, 25,
    -- filter=115 channel=48
    -1, -3, -3, -7, -11, 8, 13, 14, 19,
    -- filter=115 channel=49
    1, 1, -14, 7, 4, 0, 3, 13, 6,
    -- filter=115 channel=50
    6, 0, -2, 2, -1, -4, 8, 7, 6,
    -- filter=115 channel=51
    -7, 0, -7, -5, 4, 0, 2, 3, 7,
    -- filter=115 channel=52
    -6, -2, 0, 0, -1, -6, -8, -1, -10,
    -- filter=115 channel=53
    -2, 4, 2, 0, 4, -1, -2, -6, -1,
    -- filter=115 channel=54
    -2, -6, 5, 2, -2, -6, -2, 5, 7,
    -- filter=115 channel=55
    0, 3, -7, 14, 11, -17, -4, 5, -12,
    -- filter=115 channel=56
    2, -9, -8, 4, -2, -3, 3, -1, 0,
    -- filter=115 channel=57
    5, 5, 2, 4, -2, -7, -6, -6, 2,
    -- filter=115 channel=58
    4, 0, -2, -9, -11, 3, 0, -5, 5,
    -- filter=115 channel=59
    0, -8, -3, 3, -2, 7, 5, 0, 1,
    -- filter=115 channel=60
    -3, 1, 0, 1, -3, 3, 0, 0, 5,
    -- filter=115 channel=61
    -8, 4, 5, 0, 0, -5, 4, -9, 0,
    -- filter=115 channel=62
    -4, 6, 4, 6, 3, -2, -8, -5, -5,
    -- filter=115 channel=63
    3, 5, 1, -3, 6, -3, 5, 3, 9,
    -- filter=115 channel=64
    5, 5, -3, 1, -5, -3, -4, -2, -6,
    -- filter=115 channel=65
    -6, 4, 0, 5, -1, 4, 4, -1, 5,
    -- filter=115 channel=66
    -6, -3, 2, -13, 3, -7, 0, -1, -8,
    -- filter=115 channel=67
    1, 0, -4, -2, -6, 1, 0, 1, -2,
    -- filter=115 channel=68
    6, 7, -2, -3, -4, -2, -2, 4, 7,
    -- filter=115 channel=69
    5, -5, 0, -7, 1, 2, 0, -5, 0,
    -- filter=115 channel=70
    -1, -11, -17, 5, 3, -11, 0, 3, -1,
    -- filter=115 channel=71
    -1, -3, -5, 2, 2, 5, 0, 3, 0,
    -- filter=115 channel=72
    0, 2, 4, -3, 10, 4, 0, 3, 12,
    -- filter=115 channel=73
    5, 8, -7, 13, 10, -8, 4, -4, -6,
    -- filter=115 channel=74
    -3, 0, -9, 0, -10, -12, 8, 2, -8,
    -- filter=115 channel=75
    -7, -19, -4, -27, -22, -9, -2, 0, 1,
    -- filter=115 channel=76
    -7, 7, 0, 9, 13, 0, -14, -9, -10,
    -- filter=115 channel=77
    -2, 2, 1, -4, 0, 1, 4, 3, 4,
    -- filter=115 channel=78
    -2, -6, -2, 6, -7, -3, 6, -5, 11,
    -- filter=115 channel=79
    9, 3, -21, 8, 8, -22, -1, 11, -13,
    -- filter=115 channel=80
    1, -2, 0, -2, -4, 0, 5, 17, 10,
    -- filter=115 channel=81
    6, 7, 0, 3, 5, 4, -1, -4, 3,
    -- filter=115 channel=82
    6, -3, -2, 0, 0, -7, 3, 1, 0,
    -- filter=115 channel=83
    3, 2, 6, 6, 0, 9, -3, 3, 0,
    -- filter=115 channel=84
    3, 2, -11, 2, 9, -1, 1, 1, -4,
    -- filter=115 channel=85
    -3, -1, 0, 2, 4, 2, 0, 0, -7,
    -- filter=115 channel=86
    -8, 1, 2, 0, -7, -6, -2, -11, -1,
    -- filter=115 channel=87
    -4, 6, -8, 3, 7, -5, -5, 2, -12,
    -- filter=115 channel=88
    -9, -4, -5, -5, -2, 7, 6, -4, -1,
    -- filter=115 channel=89
    0, 3, -8, 6, 15, -6, 3, 6, 1,
    -- filter=115 channel=90
    -4, -6, -4, 2, -5, 5, -8, -11, 4,
    -- filter=115 channel=91
    -3, -1, -8, 2, 14, -9, 9, 11, 1,
    -- filter=115 channel=92
    0, -2, 0, -4, -9, -6, 0, -8, -1,
    -- filter=115 channel=93
    -7, -11, 4, -17, -16, 0, -2, 5, 20,
    -- filter=115 channel=94
    -3, 4, -1, -3, -3, 0, -2, 6, -4,
    -- filter=115 channel=95
    1, -2, -8, 0, 3, -9, 3, -2, -8,
    -- filter=115 channel=96
    -5, 6, -3, 7, 0, -4, 6, 8, -1,
    -- filter=115 channel=97
    -1, -9, -1, -10, 0, -2, -4, 2, 1,
    -- filter=115 channel=98
    3, 5, -3, -4, 10, -11, 3, 13, 6,
    -- filter=115 channel=99
    5, 0, -9, 8, -1, 2, 4, 7, -1,
    -- filter=115 channel=100
    7, -8, -10, 2, -6, -5, 10, 2, 0,
    -- filter=115 channel=101
    3, 1, -2, -11, 4, 6, -1, 4, 12,
    -- filter=115 channel=102
    -5, -4, -5, 3, -5, -4, -3, -4, -2,
    -- filter=115 channel=103
    -3, 3, 14, -18, -11, 11, -4, 0, 22,
    -- filter=115 channel=104
    0, -4, 9, -8, 2, 6, 1, 6, 17,
    -- filter=115 channel=105
    -6, 11, -6, 3, 5, 1, 2, 2, -13,
    -- filter=115 channel=106
    -5, 0, -5, -1, 0, -2, 5, 2, -1,
    -- filter=115 channel=107
    -8, 0, -6, -1, 9, -8, -3, -6, -13,
    -- filter=115 channel=108
    -3, -1, 6, 0, 3, -2, 3, -7, 5,
    -- filter=115 channel=109
    2, -1, -10, 12, 0, -2, 13, 15, 7,
    -- filter=115 channel=110
    2, 2, 3, 0, -4, -8, -1, 0, 5,
    -- filter=115 channel=111
    3, 0, 6, 6, 5, -7, -3, 5, -8,
    -- filter=115 channel=112
    8, -8, -8, 2, 0, -5, -1, 2, 9,
    -- filter=115 channel=113
    3, -8, -6, 5, 0, -8, 0, -4, 0,
    -- filter=115 channel=114
    5, -3, -10, 7, -1, -11, 2, 6, 1,
    -- filter=115 channel=115
    7, -4, 0, 3, 5, -3, 2, -6, -5,
    -- filter=115 channel=116
    8, 7, -6, 2, 11, 0, 14, 2, 6,
    -- filter=115 channel=117
    -7, 4, -1, 0, -1, 0, 0, 0, -5,
    -- filter=115 channel=118
    3, -6, 3, -1, -4, -6, 3, 0, 5,
    -- filter=115 channel=119
    -4, -10, 0, 3, -9, -6, 6, -4, 0,
    -- filter=115 channel=120
    8, 3, -11, 7, 2, -1, 3, 1, 1,
    -- filter=115 channel=121
    2, -4, 3, -1, -6, -3, 6, -1, -3,
    -- filter=115 channel=122
    -17, -4, 10, -23, -13, 16, -8, 0, 31,
    -- filter=115 channel=123
    -4, 0, 3, -4, -9, 4, 4, 1, 4,
    -- filter=115 channel=124
    5, 5, -7, 6, -2, -10, -6, -5, -12,
    -- filter=115 channel=125
    5, 6, -13, -2, 13, -6, 2, 12, 2,
    -- filter=115 channel=126
    8, 7, -7, 7, 3, -10, 5, 4, 2,
    -- filter=115 channel=127
    4, 0, 0, -2, 0, 1, -2, 2, -5,
    -- filter=116 channel=0
    0, 4, 12, -1, -14, 0, 0, 4, 1,
    -- filter=116 channel=1
    0, -2, 1, 6, -13, -15, -2, 1, -9,
    -- filter=116 channel=2
    5, 1, 1, 4, 20, 4, 8, -2, 0,
    -- filter=116 channel=3
    10, 42, 24, 12, 27, -1, 24, 41, 12,
    -- filter=116 channel=4
    21, 24, 13, 33, 66, 36, 15, 14, 8,
    -- filter=116 channel=5
    2, 3, -2, 5, 3, -1, -1, -4, 0,
    -- filter=116 channel=6
    2, 4, -4, -6, -2, 3, 6, -1, 6,
    -- filter=116 channel=7
    -7, 3, -2, 0, 2, 2, 1, -6, 7,
    -- filter=116 channel=8
    11, -4, -1, 2, 12, 6, 7, 5, 5,
    -- filter=116 channel=9
    4, 11, 7, -16, -18, -4, 7, 15, 5,
    -- filter=116 channel=10
    0, 15, 9, -18, -18, -19, 17, 25, 8,
    -- filter=116 channel=11
    5, 3, -9, -3, -2, -6, 5, 7, -4,
    -- filter=116 channel=12
    1, -2, 2, 0, -9, -3, 1, -4, 7,
    -- filter=116 channel=13
    6, 18, 15, -16, -33, -24, 12, 9, 18,
    -- filter=116 channel=14
    -5, 0, -6, 0, 4, 2, 1, 0, -1,
    -- filter=116 channel=15
    0, 10, 3, -15, -33, -22, 6, 21, 15,
    -- filter=116 channel=16
    0, 1, 4, -9, -6, -13, 9, 5, 2,
    -- filter=116 channel=17
    6, 1, -3, -4, 1, -3, -6, 0, -4,
    -- filter=116 channel=18
    3, 15, 8, -15, -32, -22, 4, 9, 13,
    -- filter=116 channel=19
    1, 0, 0, -3, 1, 3, -1, 5, -4,
    -- filter=116 channel=20
    6, 2, -7, -14, -11, -11, 6, 9, -3,
    -- filter=116 channel=21
    -5, -2, 0, -12, -15, -13, 0, 11, 5,
    -- filter=116 channel=22
    10, 11, -1, -6, -7, -7, 6, -3, -1,
    -- filter=116 channel=23
    11, 28, 16, -49, -48, -36, 28, 36, 7,
    -- filter=116 channel=24
    -1, -6, 4, 5, 0, -3, 0, 6, 7,
    -- filter=116 channel=25
    5, 19, 9, -28, -49, -25, 11, 8, 20,
    -- filter=116 channel=26
    0, -11, -3, 10, 10, 9, -5, 4, 8,
    -- filter=116 channel=27
    15, 22, 15, -48, -68, -34, 17, 30, 20,
    -- filter=116 channel=28
    0, -2, -4, -4, -2, -2, 7, 7, 4,
    -- filter=116 channel=29
    -2, -1, -1, 1, -6, -1, 9, 15, 4,
    -- filter=116 channel=30
    6, 18, 6, -21, -28, -10, 8, 7, 1,
    -- filter=116 channel=31
    0, 21, 9, -26, -39, -30, 22, 38, 18,
    -- filter=116 channel=32
    12, 21, 8, -26, -38, -30, 14, 16, 10,
    -- filter=116 channel=33
    7, 11, 19, -12, -37, -32, 15, 29, 15,
    -- filter=116 channel=34
    11, 2, -8, -11, -18, -9, 9, -6, -4,
    -- filter=116 channel=35
    -6, -5, 3, -2, 5, 6, 0, 4, -3,
    -- filter=116 channel=36
    2, -9, -3, -1, 4, -7, 6, 5, 6,
    -- filter=116 channel=37
    -8, -5, -4, 4, 5, 6, 2, -2, -3,
    -- filter=116 channel=38
    5, 7, 5, -15, -18, -13, 2, 18, 12,
    -- filter=116 channel=39
    0, 4, -2, -11, -1, 0, 1, 11, 5,
    -- filter=116 channel=40
    -8, -4, -1, -5, -15, -10, -7, 7, -3,
    -- filter=116 channel=41
    -3, -1, -4, 19, -5, -31, -9, -13, 6,
    -- filter=116 channel=42
    -4, -2, 3, -7, -10, -8, 2, 9, 5,
    -- filter=116 channel=43
    7, 17, 8, 11, 1, -5, 12, 20, 11,
    -- filter=116 channel=44
    1, 9, -6, -8, -15, -4, -1, 9, -2,
    -- filter=116 channel=45
    -8, -8, 4, 0, 6, 11, -3, 2, -1,
    -- filter=116 channel=46
    -3, 4, -4, 4, -2, -6, -5, 1, 4,
    -- filter=116 channel=47
    4, 1, 2, -8, -9, -15, 0, 18, 5,
    -- filter=116 channel=48
    12, 17, -9, -9, -23, -7, 10, 17, 17,
    -- filter=116 channel=49
    9, 0, 6, -4, 6, 9, 6, 10, 5,
    -- filter=116 channel=50
    -2, 18, 2, -24, -32, -11, -1, 20, 6,
    -- filter=116 channel=51
    -1, 4, 1, -3, -6, 2, -1, -6, 0,
    -- filter=116 channel=52
    11, 2, -9, 0, -13, -1, -3, 2, 3,
    -- filter=116 channel=53
    0, -1, 5, 0, -9, -5, 4, 6, 5,
    -- filter=116 channel=54
    6, 1, -1, 2, -1, -3, -6, 3, 3,
    -- filter=116 channel=55
    7, 6, 7, -20, -38, -26, 14, 20, 10,
    -- filter=116 channel=56
    6, -6, -7, -6, -9, -1, 0, -5, 2,
    -- filter=116 channel=57
    -5, 3, -3, -2, 8, -3, 5, 2, 1,
    -- filter=116 channel=58
    3, 3, 2, 4, 3, -6, 0, -2, 0,
    -- filter=116 channel=59
    -5, 8, 5, -18, -33, -24, 4, 15, 8,
    -- filter=116 channel=60
    -1, -7, -1, -5, -4, 4, 4, 2, -4,
    -- filter=116 channel=61
    3, -10, -4, -2, -1, 4, -4, -8, -5,
    -- filter=116 channel=62
    -6, -2, 1, -3, 2, -2, 2, 1, 1,
    -- filter=116 channel=63
    -6, 0, -8, 2, 6, 0, -6, -1, -7,
    -- filter=116 channel=64
    -2, 0, -1, -4, -4, 1, -5, 6, -5,
    -- filter=116 channel=65
    7, -2, -5, 6, -4, -1, -4, -5, -5,
    -- filter=116 channel=66
    4, -5, 0, 2, -20, -13, -4, -13, 2,
    -- filter=116 channel=67
    -2, 0, -3, 4, 3, 4, 4, -4, -2,
    -- filter=116 channel=68
    2, 0, 5, -5, 9, 6, 4, -7, 5,
    -- filter=116 channel=69
    2, 2, 0, 4, -4, 3, -7, 0, 5,
    -- filter=116 channel=70
    9, 5, 9, -20, -24, -7, 3, 14, 10,
    -- filter=116 channel=71
    1, 7, 2, 2, 14, 0, 3, 18, 6,
    -- filter=116 channel=72
    -7, 7, 8, -21, -35, -16, 5, 23, 11,
    -- filter=116 channel=73
    0, 1, 0, -12, -4, -7, 0, 2, 0,
    -- filter=116 channel=74
    9, -6, -4, -7, -20, -4, -1, 2, 9,
    -- filter=116 channel=75
    10, 11, 13, 6, -19, -20, 4, 11, 0,
    -- filter=116 channel=76
    5, 3, 6, -15, -20, -9, 3, 12, 9,
    -- filter=116 channel=77
    2, 2, 1, -5, -2, 5, -5, -1, -7,
    -- filter=116 channel=78
    1, 1, 4, -1, -2, 1, 6, 4, -1,
    -- filter=116 channel=79
    13, 20, 15, -31, -53, -40, 20, 27, 18,
    -- filter=116 channel=80
    5, 18, 8, -27, -51, -37, 11, 22, 18,
    -- filter=116 channel=81
    -4, -5, 6, -6, 6, 6, -1, -7, 4,
    -- filter=116 channel=82
    -4, 4, -3, 2, -7, 5, 0, -3, -6,
    -- filter=116 channel=83
    -7, -8, -3, 5, 5, 1, -3, 4, -5,
    -- filter=116 channel=84
    -4, 2, -6, -12, -10, 0, 0, 2, 5,
    -- filter=116 channel=85
    0, -4, 2, -7, -3, -1, 7, -5, -7,
    -- filter=116 channel=86
    2, -7, -3, -10, -12, 2, -2, 0, 5,
    -- filter=116 channel=87
    14, 3, -9, -12, -10, 0, 8, 9, -1,
    -- filter=116 channel=88
    -3, -5, -10, -9, -12, -6, 0, 4, 1,
    -- filter=116 channel=89
    4, 16, 16, -21, -45, -32, 19, 34, 14,
    -- filter=116 channel=90
    10, -5, 3, -2, 1, -3, 5, -9, -4,
    -- filter=116 channel=91
    15, 7, -3, -13, -20, -13, 1, 11, 3,
    -- filter=116 channel=92
    3, 10, 4, -7, 0, 0, 6, 5, 2,
    -- filter=116 channel=93
    1, 10, 0, -1, -11, -11, -4, 6, 14,
    -- filter=116 channel=94
    -4, -1, 1, 6, 4, -1, 0, 2, 7,
    -- filter=116 channel=95
    0, -1, 5, 4, -5, 6, -2, 3, 3,
    -- filter=116 channel=96
    6, 0, 3, -5, 8, -3, -7, 3, 8,
    -- filter=116 channel=97
    1, 17, 9, 2, 17, 2, 4, 8, 1,
    -- filter=116 channel=98
    13, 28, 12, -35, -47, -25, 16, 28, 23,
    -- filter=116 channel=99
    2, 18, -8, -31, -44, -19, 30, 31, 5,
    -- filter=116 channel=100
    8, -1, 2, -3, -13, -2, 0, -1, -9,
    -- filter=116 channel=101
    6, 15, 9, 25, 46, 16, 12, 14, 15,
    -- filter=116 channel=102
    0, -3, 0, 5, 3, 5, -5, 2, 0,
    -- filter=116 channel=103
    -6, 6, 6, -6, -9, -9, 9, 13, 8,
    -- filter=116 channel=104
    -3, -7, -6, -8, -19, -6, 11, 17, 10,
    -- filter=116 channel=105
    -5, 11, 3, 0, 0, -10, 5, 1, 2,
    -- filter=116 channel=106
    -2, 6, -5, -9, -1, -3, 0, -3, -3,
    -- filter=116 channel=107
    0, 5, 0, -8, -14, 10, 12, -2, -8,
    -- filter=116 channel=108
    -1, 0, 0, 7, 1, -4, -4, -8, 6,
    -- filter=116 channel=109
    12, 8, 0, -21, -42, -23, 3, 19, 16,
    -- filter=116 channel=110
    -6, 13, -1, -4, -8, -6, 7, 19, 12,
    -- filter=116 channel=111
    7, 0, -4, -2, 3, -4, 5, -8, 0,
    -- filter=116 channel=112
    10, 7, -1, -7, -11, -10, 1, 9, 5,
    -- filter=116 channel=113
    7, 17, 10, -17, -28, -10, 18, 22, 9,
    -- filter=116 channel=114
    8, 10, 2, -14, -30, -13, 16, 7, 10,
    -- filter=116 channel=115
    1, 2, -5, 2, 0, -1, 4, -6, 4,
    -- filter=116 channel=116
    13, 13, 2, -16, -23, -22, 16, 22, 16,
    -- filter=116 channel=117
    -2, 4, 7, -3, -7, -11, 5, 1, 2,
    -- filter=116 channel=118
    0, 1, 4, -4, 7, 0, 4, 3, -6,
    -- filter=116 channel=119
    3, -10, -5, -22, -14, -4, 3, -14, -6,
    -- filter=116 channel=120
    19, 14, -14, -34, -19, -1, 11, 15, 5,
    -- filter=116 channel=121
    -2, 12, 0, 3, -21, -21, 3, 15, 3,
    -- filter=116 channel=122
    -8, 10, 5, -4, -15, -7, -4, 16, 11,
    -- filter=116 channel=123
    2, -6, 7, -3, -11, 4, 9, -3, -3,
    -- filter=116 channel=124
    4, -3, -2, -1, -4, 2, -2, 13, -3,
    -- filter=116 channel=125
    1, 4, -3, -16, -28, -18, 7, 16, 6,
    -- filter=116 channel=126
    9, 18, 16, -12, -18, -11, 5, 11, 8,
    -- filter=116 channel=127
    -4, 6, 0, -1, -8, -4, 5, 1, -7,
    -- filter=117 channel=0
    11, 14, -12, 4, -2, -29, 0, -12, -21,
    -- filter=117 channel=1
    19, 11, -17, 9, -6, -18, -2, -13, -26,
    -- filter=117 channel=2
    1, 1, -7, -7, 0, 5, 1, 2, 6,
    -- filter=117 channel=3
    -10, 3, 5, 0, 5, -6, -6, -4, -1,
    -- filter=117 channel=4
    11, -4, 1, 1, 0, -2, 4, 4, 7,
    -- filter=117 channel=5
    14, 7, -4, 12, -4, -10, 3, 3, -12,
    -- filter=117 channel=6
    -6, -10, -6, 0, -5, -3, -3, -6, -2,
    -- filter=117 channel=7
    5, 5, -4, 0, -3, 0, 4, 0, 5,
    -- filter=117 channel=8
    -1, 0, 1, -2, 4, -8, 6, -1, -10,
    -- filter=117 channel=9
    1, 10, 1, 6, 1, -4, 3, 1, -4,
    -- filter=117 channel=10
    1, -3, 8, 7, 1, 9, 4, 6, 1,
    -- filter=117 channel=11
    -11, -16, -2, -5, -2, 6, 0, 9, 6,
    -- filter=117 channel=12
    7, -3, -5, 0, -2, -1, 6, 1, -4,
    -- filter=117 channel=13
    -1, -9, 0, 2, 5, 6, 0, 7, 0,
    -- filter=117 channel=14
    3, -1, -5, -3, 0, 3, 2, -2, -4,
    -- filter=117 channel=15
    -8, -13, -1, 4, 6, 1, 7, 1, 8,
    -- filter=117 channel=16
    -4, -2, -2, 7, 7, -14, -3, -5, -12,
    -- filter=117 channel=17
    -5, 5, 0, -6, 6, 5, 1, 3, -6,
    -- filter=117 channel=18
    9, -6, -7, 4, 0, 7, 7, -4, 1,
    -- filter=117 channel=19
    7, 6, 0, 2, 3, 6, -2, -6, -5,
    -- filter=117 channel=20
    -14, -20, 6, -14, 0, 17, -2, 3, 16,
    -- filter=117 channel=21
    -7, 6, 7, -5, 0, -2, 1, 2, -7,
    -- filter=117 channel=22
    11, -6, -7, 3, -7, -6, 9, 1, -16,
    -- filter=117 channel=23
    -2, -11, -16, 2, 1, -9, 7, 3, -9,
    -- filter=117 channel=24
    0, 0, 1, 2, 0, 5, 4, 0, 7,
    -- filter=117 channel=25
    7, 5, -5, 10, 2, -15, 7, -1, -13,
    -- filter=117 channel=26
    3, 4, 2, 2, 0, -8, 1, -8, -4,
    -- filter=117 channel=27
    11, 6, -17, 17, 8, -14, 6, 3, -14,
    -- filter=117 channel=28
    6, -2, 2, 0, 5, 6, 2, 0, -1,
    -- filter=117 channel=29
    -7, -19, 0, 0, 11, 25, -5, 1, 20,
    -- filter=117 channel=30
    11, 12, -7, 1, 5, -5, 0, -2, -12,
    -- filter=117 channel=31
    -10, 14, -4, -3, -2, -8, -2, -2, -12,
    -- filter=117 channel=32
    9, -6, -11, 0, -3, -8, 4, -2, -7,
    -- filter=117 channel=33
    0, -1, -6, 0, -2, 0, 1, 1, -7,
    -- filter=117 channel=34
    13, 6, -12, 5, -8, -8, 12, 10, -18,
    -- filter=117 channel=35
    5, 0, 2, 4, 6, 4, 0, -5, -1,
    -- filter=117 channel=36
    0, -8, -2, 3, 0, 4, 1, 0, 11,
    -- filter=117 channel=37
    4, 0, -7, 4, 2, -23, 4, -14, -20,
    -- filter=117 channel=38
    -3, 6, -1, -5, 0, 0, 4, -4, 4,
    -- filter=117 channel=39
    -3, -4, 5, -2, -2, 10, -2, 8, 16,
    -- filter=117 channel=40
    0, -4, 4, 0, 0, 1, -3, 4, 2,
    -- filter=117 channel=41
    6, -2, -3, 14, 16, -1, 4, 15, 7,
    -- filter=117 channel=42
    -3, -1, -5, 6, 0, 0, -5, -5, 0,
    -- filter=117 channel=43
    -3, -4, -6, -1, 0, -2, 9, -6, -6,
    -- filter=117 channel=44
    0, 6, -2, 8, -2, -12, -3, -9, -17,
    -- filter=117 channel=45
    -2, 5, 6, -6, -5, -5, -5, 0, 2,
    -- filter=117 channel=46
    9, 0, 0, 3, -3, -4, -3, 6, -9,
    -- filter=117 channel=47
    2, 1, -6, -3, 0, -9, -3, -13, -16,
    -- filter=117 channel=48
    9, 12, -5, 8, 6, -8, 6, -5, -8,
    -- filter=117 channel=49
    7, 0, -2, -2, 0, 0, 1, 0, 5,
    -- filter=117 channel=50
    -3, 3, -10, 0, -4, -15, 2, -7, -9,
    -- filter=117 channel=51
    5, -2, -1, 5, 2, -3, 3, -2, 3,
    -- filter=117 channel=52
    -6, -7, -5, -2, 1, 2, -2, 5, -1,
    -- filter=117 channel=53
    -9, -10, 0, -5, 7, 10, -3, -2, 5,
    -- filter=117 channel=54
    6, 4, 6, 5, -1, -4, 0, 2, 1,
    -- filter=117 channel=55
    -11, -7, 5, -2, 7, 15, 7, 11, 12,
    -- filter=117 channel=56
    3, -8, -9, 0, -3, -7, 8, -1, 0,
    -- filter=117 channel=57
    -2, 0, -1, 1, 6, -3, 6, 4, 2,
    -- filter=117 channel=58
    5, 11, -4, 0, 0, 0, 1, -4, -7,
    -- filter=117 channel=59
    -4, 5, 1, 9, 5, -11, -5, 3, -12,
    -- filter=117 channel=60
    4, 0, -6, 6, -6, -2, 3, 1, 7,
    -- filter=117 channel=61
    4, 1, 6, 2, 0, 4, -7, -5, 0,
    -- filter=117 channel=62
    5, 0, 0, 6, 6, -3, 4, -2, 5,
    -- filter=117 channel=63
    1, 7, 3, -3, 8, -2, -4, -1, -4,
    -- filter=117 channel=64
    -9, -3, 1, 3, -3, 7, -4, 5, 5,
    -- filter=117 channel=65
    -3, -6, 2, 1, 1, 0, 1, 5, -6,
    -- filter=117 channel=66
    4, 5, 1, 11, -1, 8, 0, 5, 4,
    -- filter=117 channel=67
    4, 5, -5, 0, -6, 4, 2, 7, -4,
    -- filter=117 channel=68
    5, -9, 5, 4, -6, 0, 5, -1, 6,
    -- filter=117 channel=69
    5, -4, -2, 0, -6, 0, 5, 3, -3,
    -- filter=117 channel=70
    5, -7, -18, 7, -1, -16, 4, -9, -22,
    -- filter=117 channel=71
    -2, 5, 5, 1, 0, 2, 5, -4, 0,
    -- filter=117 channel=72
    0, 3, 3, 3, 10, 6, -3, 3, -4,
    -- filter=117 channel=73
    -1, 1, 1, 7, -5, 1, 0, -1, -3,
    -- filter=117 channel=74
    11, 1, -15, 3, -7, -11, 5, 5, -19,
    -- filter=117 channel=75
    12, 9, -10, 14, -3, -25, 2, -12, -19,
    -- filter=117 channel=76
    -18, -20, 12, -2, -2, 15, -4, 13, 15,
    -- filter=117 channel=77
    -5, 7, 8, 1, 2, 1, -7, 4, 7,
    -- filter=117 channel=78
    -5, 0, -1, 8, 5, 4, 3, 7, 0,
    -- filter=117 channel=79
    -1, 0, 1, 10, 5, 3, 0, 5, -1,
    -- filter=117 channel=80
    3, 7, 7, 1, 0, -3, 3, 0, 0,
    -- filter=117 channel=81
    1, 5, -2, 5, 0, -7, -6, -4, 4,
    -- filter=117 channel=82
    -7, 0, 0, 3, -1, 0, 6, 5, 5,
    -- filter=117 channel=83
    7, 4, -1, -4, -1, -11, 2, -6, 0,
    -- filter=117 channel=84
    1, -4, -1, 3, 3, -5, 5, -4, 1,
    -- filter=117 channel=85
    6, 2, 0, -4, 4, -6, 3, -4, -4,
    -- filter=117 channel=86
    3, 3, 0, 0, 4, -12, 2, 7, -6,
    -- filter=117 channel=87
    1, -14, 0, 3, 4, 0, -3, 2, -1,
    -- filter=117 channel=88
    -5, 2, 4, -4, 1, 4, -2, 3, -3,
    -- filter=117 channel=89
    -11, 2, 0, 6, 6, 13, -1, 6, 3,
    -- filter=117 channel=90
    -10, -5, -5, -9, -10, -8, 3, 0, 1,
    -- filter=117 channel=91
    -2, -4, -3, 8, 0, -10, -4, 2, -6,
    -- filter=117 channel=92
    -3, 3, 0, 4, 3, -7, 5, 6, -5,
    -- filter=117 channel=93
    15, 13, 0, 2, -4, -22, -8, -2, -10,
    -- filter=117 channel=94
    0, -2, 0, 6, -1, 7, -5, -5, -1,
    -- filter=117 channel=95
    2, -2, 3, 6, -1, -1, -3, 0, 3,
    -- filter=117 channel=96
    0, 5, 0, -6, 0, -4, 3, -2, -1,
    -- filter=117 channel=97
    -4, -1, -2, -8, 1, 1, 6, -8, 4,
    -- filter=117 channel=98
    0, 13, -2, 2, 6, 2, -3, 0, 2,
    -- filter=117 channel=99
    -10, -5, -2, -1, -6, -12, -3, 8, -4,
    -- filter=117 channel=100
    -5, 0, 1, 0, 6, 6, -2, 0, 0,
    -- filter=117 channel=101
    -4, 4, 6, -8, -3, 5, 0, 1, 9,
    -- filter=117 channel=102
    3, -5, -2, 6, -2, 6, -4, 6, -1,
    -- filter=117 channel=103
    3, 9, -10, -1, -7, -11, -9, 0, -17,
    -- filter=117 channel=104
    -7, 0, 0, 2, 2, -5, -6, -2, -8,
    -- filter=117 channel=105
    -5, -10, 6, -2, 0, 22, -3, 0, 18,
    -- filter=117 channel=106
    0, -4, 7, -3, 5, 14, 7, 8, 11,
    -- filter=117 channel=107
    -7, -17, -8, 4, -4, 0, -6, -5, -1,
    -- filter=117 channel=108
    0, -4, 6, 10, 2, -3, 8, -1, -5,
    -- filter=117 channel=109
    12, 5, -13, 5, 7, -6, 10, -7, -14,
    -- filter=117 channel=110
    -2, 4, 8, 5, 0, 5, 0, 8, 0,
    -- filter=117 channel=111
    4, -3, -1, -1, 0, -6, 1, 6, 8,
    -- filter=117 channel=112
    8, 9, -7, 11, 3, -18, 7, -5, -18,
    -- filter=117 channel=113
    -4, 0, -7, 6, -3, -6, 2, -1, 1,
    -- filter=117 channel=114
    9, 3, -4, 16, 6, -21, 10, 2, -5,
    -- filter=117 channel=115
    0, -3, 2, 6, 2, -5, 2, 4, 5,
    -- filter=117 channel=116
    3, -2, 1, -4, 1, 0, 4, 0, 0,
    -- filter=117 channel=117
    3, -7, 8, 7, 0, -1, 4, 3, 2,
    -- filter=117 channel=118
    -1, -4, -5, 5, -4, 1, -4, 0, -5,
    -- filter=117 channel=119
    13, 6, -13, 7, 6, -17, 5, 0, -13,
    -- filter=117 channel=120
    -2, -5, -4, 2, -7, -13, 7, 3, -21,
    -- filter=117 channel=121
    6, 0, -2, 1, -2, 3, 9, -3, 4,
    -- filter=117 channel=122
    1, 11, -12, -4, -8, -19, -10, -16, -24,
    -- filter=117 channel=123
    -1, -4, -3, 5, -7, -11, 0, -6, -6,
    -- filter=117 channel=124
    -8, -15, 2, 0, 2, 13, 5, -3, 8,
    -- filter=117 channel=125
    -7, 9, 5, 7, -3, -10, -1, 0, -1,
    -- filter=117 channel=126
    2, -6, 8, 1, 8, 10, 9, 5, 6,
    -- filter=117 channel=127
    4, -6, -3, 0, 4, 0, 4, 3, 6,
    -- filter=118 channel=0
    2, -5, 0, 2, 2, 9, 0, 1, 6,
    -- filter=118 channel=1
    -5, -8, -1, 14, 0, 2, 0, -5, 0,
    -- filter=118 channel=2
    1, -6, 0, 7, 0, -7, 0, 4, 4,
    -- filter=118 channel=3
    -1, -1, -9, -1, -6, -7, 2, 14, -6,
    -- filter=118 channel=4
    7, -3, -1, 18, 7, -12, 10, 9, 1,
    -- filter=118 channel=5
    -7, -3, 4, -4, -5, 8, -4, -4, -7,
    -- filter=118 channel=6
    -3, -7, -3, -4, 2, 2, 9, 0, 9,
    -- filter=118 channel=7
    -2, -7, -3, 5, 4, 5, 0, -1, -7,
    -- filter=118 channel=8
    2, 8, 7, 11, 0, -2, 1, 2, -1,
    -- filter=118 channel=9
    -3, -1, -7, 7, -2, -6, 0, -6, -9,
    -- filter=118 channel=10
    -8, -15, -10, -14, -3, 0, 11, 13, 1,
    -- filter=118 channel=11
    -19, -19, -12, -2, -2, 7, 18, 2, 8,
    -- filter=118 channel=12
    0, 0, 7, 0, -5, 1, -6, 4, -4,
    -- filter=118 channel=13
    -5, -21, 0, -1, 0, -2, 7, 25, 11,
    -- filter=118 channel=14
    -5, 4, -1, -4, -5, -4, 0, 0, 0,
    -- filter=118 channel=15
    -19, -28, -12, 1, -9, -7, 24, 26, 4,
    -- filter=118 channel=16
    3, 15, -1, 3, -1, 3, -10, -1, -3,
    -- filter=118 channel=17
    6, -7, -6, 5, 3, 1, -3, -6, -4,
    -- filter=118 channel=18
    -21, -36, -18, -3, 0, -2, 25, 25, 5,
    -- filter=118 channel=19
    -4, -5, 7, 3, -3, 3, 2, -2, 1,
    -- filter=118 channel=20
    -12, -15, -12, 4, 3, 3, 18, 20, 12,
    -- filter=118 channel=21
    10, 11, 7, 0, 1, 6, -4, -12, -4,
    -- filter=118 channel=22
    -3, -3, 2, -4, -11, 1, -1, 8, 9,
    -- filter=118 channel=23
    -20, -34, -10, -8, -17, -7, 25, 25, 6,
    -- filter=118 channel=24
    1, -6, -6, 3, 5, 0, 0, 0, 7,
    -- filter=118 channel=25
    -7, -19, 2, -1, 9, 2, -2, 6, 4,
    -- filter=118 channel=26
    11, 8, 10, 6, 6, 2, 5, -7, 1,
    -- filter=118 channel=27
    -28, -24, -6, 10, 4, -6, 15, 20, 6,
    -- filter=118 channel=28
    -6, 5, 0, 5, -1, 0, -6, 0, 5,
    -- filter=118 channel=29
    -22, -20, -4, 3, -3, 5, 25, 18, 8,
    -- filter=118 channel=30
    -10, 0, -7, 6, 13, 3, -1, -7, 0,
    -- filter=118 channel=31
    -13, -4, 11, 4, -2, 0, 8, -1, -5,
    -- filter=118 channel=32
    -18, -32, -8, -6, -7, 6, 12, 19, 9,
    -- filter=118 channel=33
    -15, -22, -12, 0, -10, 0, 3, 11, 1,
    -- filter=118 channel=34
    -6, -2, 4, -11, 3, -7, 0, 4, 1,
    -- filter=118 channel=35
    0, 5, -4, 3, 7, 6, 0, -1, 6,
    -- filter=118 channel=36
    2, 3, -1, 3, 12, 5, -2, -1, 4,
    -- filter=118 channel=37
    3, 1, 8, 13, 7, 2, -5, -3, -2,
    -- filter=118 channel=38
    0, -7, 2, 0, 2, 3, 8, 7, 0,
    -- filter=118 channel=39
    -8, -16, -7, 1, 1, -5, 5, 10, 5,
    -- filter=118 channel=40
    2, -5, -4, -11, -7, 4, 7, 3, -2,
    -- filter=118 channel=41
    12, -14, 0, -1, 3, -1, 2, 14, 9,
    -- filter=118 channel=42
    2, -8, 3, -5, 0, 2, 0, -2, -3,
    -- filter=118 channel=43
    -7, -6, -12, -8, 0, -5, 3, 15, 2,
    -- filter=118 channel=44
    -10, 9, 9, 5, 3, 2, 0, -15, -12,
    -- filter=118 channel=45
    1, 1, 4, -3, -9, -1, 6, 6, -3,
    -- filter=118 channel=46
    0, 0, -6, -5, 5, -5, 0, -4, 3,
    -- filter=118 channel=47
    1, 6, 14, 2, 2, 6, -14, -4, -14,
    -- filter=118 channel=48
    -11, 3, 9, 6, 17, -3, -7, -3, -6,
    -- filter=118 channel=49
    -6, -18, -2, 6, 11, 0, 0, 7, 4,
    -- filter=118 channel=50
    -5, -12, -3, 6, -5, 3, 6, 6, -6,
    -- filter=118 channel=51
    0, 0, -6, -6, 7, -5, 1, 6, -4,
    -- filter=118 channel=52
    -3, -11, 0, 2, -2, 4, 0, 0, 0,
    -- filter=118 channel=53
    -7, -14, -4, 1, 2, 7, 6, 13, -1,
    -- filter=118 channel=54
    3, -4, 4, -1, -2, -1, 3, 2, 1,
    -- filter=118 channel=55
    -19, -33, -14, -11, 3, -5, 25, 33, 17,
    -- filter=118 channel=56
    -2, -3, 0, 6, -5, -1, 5, 2, 0,
    -- filter=118 channel=57
    3, -2, -5, -1, 0, -1, 8, 4, -3,
    -- filter=118 channel=58
    7, 11, 9, -1, -1, 0, 0, 0, 3,
    -- filter=118 channel=59
    -14, -15, -6, 5, 2, 1, -6, 3, -2,
    -- filter=118 channel=60
    5, 6, -1, 0, -2, 2, 3, 0, 1,
    -- filter=118 channel=61
    -8, 3, 5, 9, 8, -6, -3, 3, -6,
    -- filter=118 channel=62
    -2, -5, 2, 1, -1, -5, -2, 5, 7,
    -- filter=118 channel=63
    -1, 0, 0, 0, 4, 0, 0, -15, 0,
    -- filter=118 channel=64
    -1, 0, 7, 2, 2, 0, 9, -2, 3,
    -- filter=118 channel=65
    -2, -1, -6, 0, 0, 6, -5, 0, 1,
    -- filter=118 channel=66
    8, -10, 0, 1, 4, 1, -6, 12, 4,
    -- filter=118 channel=67
    -3, 6, 3, 1, 0, 6, 0, 5, 1,
    -- filter=118 channel=68
    2, -3, -4, 2, 9, 0, -6, 2, -6,
    -- filter=118 channel=69
    -5, 4, 2, -5, -9, 0, -5, -6, -2,
    -- filter=118 channel=70
    -25, -17, 1, -4, -9, -7, 11, 10, 0,
    -- filter=118 channel=71
    0, 3, -4, 2, -2, 0, -5, 6, 1,
    -- filter=118 channel=72
    -15, -7, -2, 6, 9, 5, 5, 2, -6,
    -- filter=118 channel=73
    -7, -16, 0, 8, 9, -3, 12, 19, -1,
    -- filter=118 channel=74
    -5, -5, 4, 0, 9, 0, 6, -6, -2,
    -- filter=118 channel=75
    -13, -12, -9, 0, -18, -10, -2, -2, 3,
    -- filter=118 channel=76
    -7, -23, 0, -11, 0, -1, 16, 13, 5,
    -- filter=118 channel=77
    0, 0, 1, 0, -5, -2, -2, 7, -1,
    -- filter=118 channel=78
    3, 7, 11, -8, 5, 2, 3, 2, -5,
    -- filter=118 channel=79
    -24, -36, -15, -3, 0, 2, 26, 33, 9,
    -- filter=118 channel=80
    -5, -4, -3, -4, 1, -4, 0, -5, -11,
    -- filter=118 channel=81
    0, 1, -3, -4, -1, -1, 2, -2, -5,
    -- filter=118 channel=82
    -5, -9, -3, -8, -10, -3, -4, 6, 0,
    -- filter=118 channel=83
    2, 2, -1, -1, 7, 0, -6, -2, -4,
    -- filter=118 channel=84
    -11, -16, -6, 12, 11, 0, 14, 10, 8,
    -- filter=118 channel=85
    1, -1, 0, -4, 5, -2, 2, -1, 1,
    -- filter=118 channel=86
    -6, 3, 2, -5, 0, -4, 0, 3, 0,
    -- filter=118 channel=87
    0, -9, 5, 4, -7, 6, 14, 3, 0,
    -- filter=118 channel=88
    -7, 7, 6, 8, 7, 7, 0, -2, -7,
    -- filter=118 channel=89
    -18, -28, -10, -12, -7, 3, 21, 17, 5,
    -- filter=118 channel=90
    1, 4, 7, 2, -1, 3, 4, -3, -2,
    -- filter=118 channel=91
    -15, -19, -1, 13, 15, -6, 7, 5, 9,
    -- filter=118 channel=92
    1, 1, -7, -2, -7, -8, -1, -2, 1,
    -- filter=118 channel=93
    6, 7, 8, 13, 13, 0, -5, 0, 0,
    -- filter=118 channel=94
    -4, 2, 1, 5, -2, 6, -4, 6, 2,
    -- filter=118 channel=95
    -3, -4, -3, 0, -3, 0, 5, 3, 2,
    -- filter=118 channel=96
    3, 0, 0, -5, -3, -7, 0, 3, 5,
    -- filter=118 channel=97
    -2, -8, -10, -12, -13, -1, -3, 1, 4,
    -- filter=118 channel=98
    -8, -18, -1, 2, -1, 2, 11, 13, -4,
    -- filter=118 channel=99
    -15, -20, 1, 4, 7, -4, 15, 9, 0,
    -- filter=118 channel=100
    0, -3, 4, -8, -4, -3, -5, 9, -1,
    -- filter=118 channel=101
    1, 0, -8, 5, 6, 2, 14, 11, -1,
    -- filter=118 channel=102
    2, -4, 2, 7, 1, -4, 5, -6, 6,
    -- filter=118 channel=103
    -9, -2, -6, -1, 1, -3, -1, -12, -11,
    -- filter=118 channel=104
    0, -4, 9, 6, 11, 0, 1, -6, -10,
    -- filter=118 channel=105
    -3, -12, -8, 0, 3, 7, 14, 11, 9,
    -- filter=118 channel=106
    -6, -2, -2, 3, 2, 5, 11, 8, 7,
    -- filter=118 channel=107
    -19, -13, 0, -7, -2, 6, 9, 10, 15,
    -- filter=118 channel=108
    3, -3, -5, -6, 2, -3, 1, -5, -5,
    -- filter=118 channel=109
    -16, -17, -13, 4, 12, 1, 7, 22, 7,
    -- filter=118 channel=110
    -10, -12, 4, -5, 1, 3, 12, 2, 6,
    -- filter=118 channel=111
    5, -3, 4, -2, -3, -6, 7, 6, 0,
    -- filter=118 channel=112
    -1, -3, 2, 6, 4, -8, -1, 4, -7,
    -- filter=118 channel=113
    -16, -14, -16, -5, -9, 0, -2, 4, -5,
    -- filter=118 channel=114
    -23, -44, -21, 11, 1, -4, 19, 20, 6,
    -- filter=118 channel=115
    2, 0, -1, -5, -1, 0, 0, -4, -2,
    -- filter=118 channel=116
    -10, -13, -6, 18, 14, 2, 10, 4, 0,
    -- filter=118 channel=117
    -1, -9, 2, 5, -3, 2, -3, 4, -7,
    -- filter=118 channel=118
    6, -5, 3, -1, 8, 0, 5, 7, -2,
    -- filter=118 channel=119
    -8, -5, 9, 0, 3, -2, 8, -1, -5,
    -- filter=118 channel=120
    -28, -33, 0, 14, 15, 4, 19, 11, 5,
    -- filter=118 channel=121
    5, -8, -10, -8, 0, -1, 4, 2, -4,
    -- filter=118 channel=122
    4, 34, 20, 10, 15, 4, -20, -15, -23,
    -- filter=118 channel=123
    -1, -6, -3, 0, 2, -5, -1, 7, 4,
    -- filter=118 channel=124
    0, -6, -3, 2, 3, -4, 14, 14, 5,
    -- filter=118 channel=125
    -11, -9, -2, 5, 10, 0, 4, 7, 0,
    -- filter=118 channel=126
    0, -15, -7, -13, -10, 0, 8, 19, 2,
    -- filter=118 channel=127
    7, 0, 3, -3, 6, -5, -3, 0, 1,
    -- filter=119 channel=0
    -7, 7, 0, 3, 5, -2, -5, 1, -7,
    -- filter=119 channel=1
    0, 7, 3, -5, -2, -2, -4, -2, -7,
    -- filter=119 channel=2
    0, 2, 4, 2, 7, -5, -4, -5, 7,
    -- filter=119 channel=3
    2, -5, -1, -4, -7, -1, 2, 1, 3,
    -- filter=119 channel=4
    4, -6, 3, -3, -2, 4, -2, -1, -1,
    -- filter=119 channel=5
    6, 6, -1, 0, 6, -1, 1, 5, -3,
    -- filter=119 channel=6
    -1, -6, -4, 7, 7, -6, 2, 4, -1,
    -- filter=119 channel=7
    6, -2, -2, -7, -3, 7, -3, 4, 1,
    -- filter=119 channel=8
    -5, 1, 6, 6, 2, -2, 0, 4, 5,
    -- filter=119 channel=9
    7, 0, 1, 2, -5, 1, 4, -4, -5,
    -- filter=119 channel=10
    -1, -1, 1, -3, 5, 2, -6, -5, -3,
    -- filter=119 channel=11
    -2, -3, 3, -1, -1, 2, -4, 0, 3,
    -- filter=119 channel=12
    -5, -4, 3, -4, 5, 4, -1, 1, 0,
    -- filter=119 channel=13
    3, 5, -3, 0, -5, -3, 1, 4, -6,
    -- filter=119 channel=14
    6, -1, -2, -5, -3, 4, 0, 0, 0,
    -- filter=119 channel=15
    0, 5, 8, 5, 3, -6, 4, 0, 5,
    -- filter=119 channel=16
    2, -2, 0, 0, -6, -1, 5, 5, 2,
    -- filter=119 channel=17
    -6, 0, -5, 0, -6, 7, -2, -1, 5,
    -- filter=119 channel=18
    2, -1, -6, 5, -6, 2, 8, -5, -1,
    -- filter=119 channel=19
    -5, 7, 5, -5, 4, 1, 2, 6, -6,
    -- filter=119 channel=20
    6, -1, 0, 0, 0, 6, 8, 1, 3,
    -- filter=119 channel=21
    1, -2, 3, 0, -1, 0, 4, -7, 5,
    -- filter=119 channel=22
    1, 0, 7, 4, 7, 0, 7, 2, 6,
    -- filter=119 channel=23
    -1, 4, 0, 2, 6, -4, -3, 0, 3,
    -- filter=119 channel=24
    -4, -6, 4, 1, -2, 0, 3, -2, 1,
    -- filter=119 channel=25
    -8, -5, 2, 3, 0, -6, -4, -4, 0,
    -- filter=119 channel=26
    7, 2, -2, 0, -1, 4, -3, 7, 5,
    -- filter=119 channel=27
    -2, -5, 0, 1, -4, -5, -2, -7, -1,
    -- filter=119 channel=28
    -4, 5, 3, 4, 5, 6, -2, -1, -2,
    -- filter=119 channel=29
    4, -6, 0, 1, -5, 1, 9, -5, 7,
    -- filter=119 channel=30
    -2, -5, -6, -1, 1, -3, 2, 0, -6,
    -- filter=119 channel=31
    -7, -5, 0, -5, -3, -7, -5, -1, 4,
    -- filter=119 channel=32
    2, -1, -6, -1, -6, -1, -5, -3, 1,
    -- filter=119 channel=33
    6, 2, -5, 1, -4, 0, 2, 4, 1,
    -- filter=119 channel=34
    -4, -5, 3, 5, -3, -1, 1, -4, 1,
    -- filter=119 channel=35
    -4, -4, 5, 0, 5, -2, -6, -3, 0,
    -- filter=119 channel=36
    -1, -3, 4, 1, 0, -6, -4, 3, 5,
    -- filter=119 channel=37
    -4, 1, -5, -6, 0, 6, 3, 7, 2,
    -- filter=119 channel=38
    0, -7, 2, -5, -7, 0, -3, -5, -3,
    -- filter=119 channel=39
    -4, 0, 0, 4, 1, 1, 1, -1, 0,
    -- filter=119 channel=40
    2, 4, 4, 0, -5, 5, -3, -2, 3,
    -- filter=119 channel=41
    -6, -3, -2, 0, -2, -2, 0, 6, 1,
    -- filter=119 channel=42
    -4, 4, 1, 6, -2, -5, -6, -1, -2,
    -- filter=119 channel=43
    -2, -2, 7, 0, -4, -3, -5, 6, -4,
    -- filter=119 channel=44
    -6, 0, -5, -4, 4, 2, 0, 2, -2,
    -- filter=119 channel=45
    3, 3, 6, 5, -6, 4, -2, 0, 5,
    -- filter=119 channel=46
    7, 6, -6, -5, -7, -4, 1, -5, -1,
    -- filter=119 channel=47
    -5, 5, 1, 1, -2, 1, -3, 1, -7,
    -- filter=119 channel=48
    -3, -1, -7, 1, 0, 0, -7, 6, 4,
    -- filter=119 channel=49
    -6, -2, 5, -7, 2, -6, 3, -5, 3,
    -- filter=119 channel=50
    1, -2, 0, -6, -7, -6, 6, 3, 6,
    -- filter=119 channel=51
    -2, -2, 3, 6, -7, 7, -4, -5, -3,
    -- filter=119 channel=52
    1, 0, -1, 3, 1, 3, -2, -7, -1,
    -- filter=119 channel=53
    -1, -1, -4, -6, -5, -2, 0, 6, -1,
    -- filter=119 channel=54
    -3, 7, 6, 6, -2, 3, 1, -3, 3,
    -- filter=119 channel=55
    3, -3, 4, -5, -3, -1, 6, -4, -4,
    -- filter=119 channel=56
    -4, 1, 4, -4, 2, -4, 4, -2, 6,
    -- filter=119 channel=57
    -1, -1, 2, 6, -6, 2, 4, 7, 0,
    -- filter=119 channel=58
    -1, -1, -6, 1, -5, 5, -7, -3, 2,
    -- filter=119 channel=59
    3, 0, -6, 2, -1, 5, -4, 3, 0,
    -- filter=119 channel=60
    3, -4, 0, 3, -2, -2, 1, 6, 5,
    -- filter=119 channel=61
    -5, 3, 6, 1, 6, 0, 5, 4, -4,
    -- filter=119 channel=62
    7, 3, -5, 0, 0, 3, 1, 1, 6,
    -- filter=119 channel=63
    -1, -1, 7, 5, 4, -6, 2, -3, -7,
    -- filter=119 channel=64
    4, 4, -1, 6, 0, 1, 1, 2, -6,
    -- filter=119 channel=65
    -5, 0, 2, 7, -2, 4, 0, 6, 0,
    -- filter=119 channel=66
    -7, 7, -5, 3, 7, -4, 4, 5, -6,
    -- filter=119 channel=67
    -2, 4, 0, 3, 5, -5, -6, 0, -2,
    -- filter=119 channel=68
    -1, -1, 4, 0, -3, 4, 0, -3, 5,
    -- filter=119 channel=69
    6, -4, 1, -3, -4, 6, -6, 5, 0,
    -- filter=119 channel=70
    -6, -5, 5, 3, -1, -2, 6, 6, -4,
    -- filter=119 channel=71
    -1, -5, -5, 0, 0, 6, -2, 0, -3,
    -- filter=119 channel=72
    0, -6, -7, 4, 5, -1, -1, -3, -3,
    -- filter=119 channel=73
    -2, -5, 2, -2, -2, 3, -5, 0, 7,
    -- filter=119 channel=74
    -4, -2, 0, 1, 4, -1, 0, 3, 4,
    -- filter=119 channel=75
    4, 1, 0, 0, 5, 2, -4, -1, 1,
    -- filter=119 channel=76
    3, 2, 2, 1, -2, 0, 8, 2, 0,
    -- filter=119 channel=77
    -6, -5, 6, 4, -3, -1, 0, 7, -2,
    -- filter=119 channel=78
    -7, 5, 6, -5, 2, 0, 0, 7, -5,
    -- filter=119 channel=79
    6, 1, 5, 1, 4, 3, -2, -3, 5,
    -- filter=119 channel=80
    2, 6, 5, -8, 0, -2, 3, 6, 5,
    -- filter=119 channel=81
    -3, -6, 5, 7, -5, 0, 6, 4, -6,
    -- filter=119 channel=82
    1, 4, 4, -2, 2, 0, 2, 0, 0,
    -- filter=119 channel=83
    3, -4, -3, 3, 5, -7, -6, 5, 0,
    -- filter=119 channel=84
    6, 4, -5, 7, 1, -1, 1, -6, 5,
    -- filter=119 channel=85
    1, 6, -3, 5, -4, 7, 4, -4, -5,
    -- filter=119 channel=86
    0, 2, 3, 4, -3, 2, 5, 0, 4,
    -- filter=119 channel=87
    5, 0, 0, 5, -6, 6, 0, 5, 7,
    -- filter=119 channel=88
    2, -3, 2, 2, 0, 7, 6, -4, 5,
    -- filter=119 channel=89
    -1, -1, 0, -6, 2, -5, 1, 2, 4,
    -- filter=119 channel=90
    -6, 0, -3, -4, -4, 0, -1, 0, 6,
    -- filter=119 channel=91
    6, 1, -2, 3, -1, -5, 0, -6, 0,
    -- filter=119 channel=92
    -4, 0, 4, -6, -3, -4, 0, 2, 2,
    -- filter=119 channel=93
    6, 5, -2, 0, 2, 7, 1, -3, -7,
    -- filter=119 channel=94
    -5, 0, 6, -1, -3, 4, -5, -3, 0,
    -- filter=119 channel=95
    -7, 0, 0, 0, 1, 5, 6, 5, -5,
    -- filter=119 channel=96
    1, 0, -4, 6, 7, 5, 3, -5, 1,
    -- filter=119 channel=97
    2, -7, -6, 3, 5, -1, -7, 0, 0,
    -- filter=119 channel=98
    -6, -1, -5, -6, 2, -5, 5, -5, -1,
    -- filter=119 channel=99
    0, 2, 5, 4, -8, -1, -1, -2, 6,
    -- filter=119 channel=100
    -5, 4, -2, 5, -7, 6, 2, -4, 2,
    -- filter=119 channel=101
    0, -5, -5, 0, 1, -2, 0, -5, 3,
    -- filter=119 channel=102
    6, 6, 4, -4, 7, 3, -3, -3, -1,
    -- filter=119 channel=103
    -1, 3, -6, 6, 0, -7, -8, 2, 6,
    -- filter=119 channel=104
    0, -2, 4, 4, 5, -4, -7, -3, -5,
    -- filter=119 channel=105
    -5, -4, 6, 5, -6, 6, 0, 0, 3,
    -- filter=119 channel=106
    1, -4, 2, -6, 5, -3, -6, -4, 0,
    -- filter=119 channel=107
    -3, 2, 6, 3, 7, -2, -1, -6, 5,
    -- filter=119 channel=108
    -2, 1, -1, -3, -5, 0, 5, -2, 4,
    -- filter=119 channel=109
    5, 3, 2, 5, -2, -2, 0, 4, -4,
    -- filter=119 channel=110
    -3, -5, 3, -2, -5, -7, 3, -2, 3,
    -- filter=119 channel=111
    -1, -3, -6, 2, 5, 0, 0, -7, -7,
    -- filter=119 channel=112
    -4, 0, 4, -7, 1, 0, 3, 4, -2,
    -- filter=119 channel=113
    -3, -6, -1, -6, -4, 0, -4, -2, 0,
    -- filter=119 channel=114
    -5, -3, -3, -1, -5, -3, 5, -4, 5,
    -- filter=119 channel=115
    -6, 6, -6, 1, 5, -1, 5, -5, 6,
    -- filter=119 channel=116
    -1, -7, 3, -3, 1, -5, -7, 3, 4,
    -- filter=119 channel=117
    -6, 3, 6, -3, 5, 5, -2, -5, 1,
    -- filter=119 channel=118
    -1, 0, 0, -4, 0, -4, 0, -2, 0,
    -- filter=119 channel=119
    3, 7, -2, -3, 6, 0, 0, 4, -1,
    -- filter=119 channel=120
    7, 0, -5, 1, 0, -2, 2, -6, 0,
    -- filter=119 channel=121
    7, -2, -6, -1, 0, -6, 3, -4, 0,
    -- filter=119 channel=122
    -3, -6, -5, -6, 4, 5, 0, 0, -2,
    -- filter=119 channel=123
    -1, -2, 2, -7, -1, 5, 3, 3, 4,
    -- filter=119 channel=124
    8, 3, 2, 3, -4, -6, -2, -4, -6,
    -- filter=119 channel=125
    0, 0, -4, -3, 3, 0, -7, -3, 0,
    -- filter=119 channel=126
    7, 0, -1, 1, 3, 5, 4, -3, 2,
    -- filter=119 channel=127
    -3, 3, 5, -4, -6, 5, -1, 6, 0,
    -- filter=120 channel=0
    14, 10, -9, 3, 3, -2, 9, 6, 3,
    -- filter=120 channel=1
    0, 5, 5, -2, -8, 10, 8, 7, 2,
    -- filter=120 channel=2
    -1, -3, -4, 3, -10, 4, 0, -7, -5,
    -- filter=120 channel=3
    14, 20, 2, 8, 5, -11, 8, 11, 5,
    -- filter=120 channel=4
    12, 10, 6, 14, 2, 0, 10, 0, -7,
    -- filter=120 channel=5
    11, 0, 0, 4, -10, -1, -5, -6, 7,
    -- filter=120 channel=6
    2, -3, -2, -1, -4, -1, 4, 4, 5,
    -- filter=120 channel=7
    3, 3, 3, -5, -3, 0, 0, 2, 4,
    -- filter=120 channel=8
    2, 5, 5, -4, 0, 4, 0, 1, 2,
    -- filter=120 channel=9
    3, -1, 7, -5, 0, 6, -7, 0, -5,
    -- filter=120 channel=10
    -7, 2, 9, -11, -11, 2, -3, -4, -2,
    -- filter=120 channel=11
    -7, -5, 0, -8, -5, 6, 1, -5, 0,
    -- filter=120 channel=12
    -7, 7, 11, -2, -2, 13, -3, -7, 10,
    -- filter=120 channel=13
    0, 13, 5, -9, -10, 5, 2, -8, -1,
    -- filter=120 channel=14
    -4, 0, 2, 1, 1, -5, 2, 1, 1,
    -- filter=120 channel=15
    0, 11, -11, 2, 10, 6, 3, -5, 8,
    -- filter=120 channel=16
    -2, 0, 1, -9, -4, 14, 3, -12, 5,
    -- filter=120 channel=17
    -4, -5, -4, -1, 1, -1, -7, -2, 0,
    -- filter=120 channel=18
    1, 5, -12, -7, 0, 7, 4, -7, 0,
    -- filter=120 channel=19
    -3, -3, 0, 0, 5, 0, 0, 0, -2,
    -- filter=120 channel=20
    -7, 3, -8, -7, 8, 4, 0, 1, 11,
    -- filter=120 channel=21
    -10, 0, 10, -14, -14, 11, -15, -22, 3,
    -- filter=120 channel=22
    5, 0, -4, 4, 12, 6, 6, 9, 3,
    -- filter=120 channel=23
    3, 11, -3, -11, 10, 3, 0, -5, 4,
    -- filter=120 channel=24
    0, -7, 0, 3, 0, 3, 6, 4, -5,
    -- filter=120 channel=25
    1, 7, -3, -16, -12, 11, 5, -6, 6,
    -- filter=120 channel=26
    0, 1, -3, -1, -5, 7, 0, -12, 0,
    -- filter=120 channel=27
    11, 6, -6, -22, -1, 13, 0, 0, -1,
    -- filter=120 channel=28
    -5, -6, 6, 4, -4, -7, -2, 6, 5,
    -- filter=120 channel=29
    -8, 1, -5, -6, 4, 0, 2, -3, 5,
    -- filter=120 channel=30
    11, 12, 2, -6, 0, 9, 6, -8, -3,
    -- filter=120 channel=31
    -7, 12, -2, -34, -13, 14, -8, -18, 12,
    -- filter=120 channel=32
    3, 9, 0, -5, 2, 9, 6, -5, -4,
    -- filter=120 channel=33
    6, 20, -1, -9, 3, 2, -7, -9, 1,
    -- filter=120 channel=34
    9, 0, 0, 0, 13, 8, 5, 2, 11,
    -- filter=120 channel=35
    4, -1, -1, 3, -2, -6, -2, 2, 5,
    -- filter=120 channel=36
    -1, 4, 3, -4, -10, 2, -2, -5, 1,
    -- filter=120 channel=37
    14, 7, 7, -4, -8, 5, 1, -2, 6,
    -- filter=120 channel=38
    0, 0, -4, -11, 5, -2, 0, -6, 2,
    -- filter=120 channel=39
    -4, -8, -4, -6, -5, 8, 0, -2, -3,
    -- filter=120 channel=40
    0, -3, -7, 4, 4, -5, -2, 4, 1,
    -- filter=120 channel=41
    -20, -8, 12, -10, -9, 9, -4, 6, 3,
    -- filter=120 channel=42
    0, 3, -3, -5, -9, -6, -3, -7, 0,
    -- filter=120 channel=43
    4, 11, -8, 10, 15, -1, 0, 6, 7,
    -- filter=120 channel=44
    0, 9, 5, -9, 3, 4, 5, 0, 5,
    -- filter=120 channel=45
    11, 2, 0, 3, -4, -8, 4, -5, -5,
    -- filter=120 channel=46
    -2, -4, 7, -6, -7, 4, 2, -1, -3,
    -- filter=120 channel=47
    1, 11, 19, -8, -6, 15, -9, -20, -1,
    -- filter=120 channel=48
    1, 1, 7, -19, -8, 10, -9, 0, 0,
    -- filter=120 channel=49
    10, 8, -1, 3, 0, 7, 7, -2, 0,
    -- filter=120 channel=50
    1, 0, 5, -13, 4, 4, -1, -11, 8,
    -- filter=120 channel=51
    5, -6, 3, -6, -2, -2, -5, 3, 7,
    -- filter=120 channel=52
    5, -2, 3, -1, 12, 0, 1, -5, 0,
    -- filter=120 channel=53
    -6, -1, 0, -6, -2, -1, -5, 0, -1,
    -- filter=120 channel=54
    0, -7, -4, -3, 4, -4, 7, 6, 0,
    -- filter=120 channel=55
    -9, 5, -1, -12, -1, 1, -9, -4, 1,
    -- filter=120 channel=56
    1, -9, 8, -7, -1, 2, -4, -3, 6,
    -- filter=120 channel=57
    -3, 1, 5, 7, -6, 3, -7, 0, -5,
    -- filter=120 channel=58
    11, -7, -6, 8, -6, -1, 7, -1, -7,
    -- filter=120 channel=59
    -14, 8, 11, -12, -13, 16, -3, -12, 7,
    -- filter=120 channel=60
    -3, -7, 0, -5, 3, 5, -2, 2, 5,
    -- filter=120 channel=61
    0, -9, -8, 2, -2, 2, 0, -6, -2,
    -- filter=120 channel=62
    0, 1, -7, 2, 5, -2, 1, -4, -1,
    -- filter=120 channel=63
    2, -3, -6, -2, -8, 2, 4, 2, 6,
    -- filter=120 channel=64
    -6, -3, -1, 0, -2, 3, 5, -8, 8,
    -- filter=120 channel=65
    -4, -5, 0, 7, 4, 6, -3, 0, -4,
    -- filter=120 channel=66
    -5, 7, -1, -9, -7, 14, -6, 6, 14,
    -- filter=120 channel=67
    4, 0, -1, -8, 8, -1, -9, 7, -1,
    -- filter=120 channel=68
    2, 0, 8, -3, -1, -4, -5, 6, -6,
    -- filter=120 channel=69
    0, -6, 10, -5, -4, 2, -1, 4, 8,
    -- filter=120 channel=70
    9, 14, 4, -2, 14, 6, 3, 0, 3,
    -- filter=120 channel=71
    11, 2, -2, 6, -2, -7, 0, 4, 5,
    -- filter=120 channel=72
    -16, 2, 11, -27, -5, 17, -16, -15, -1,
    -- filter=120 channel=73
    -5, 8, -3, -11, -8, -2, -10, -4, 5,
    -- filter=120 channel=74
    2, -4, -6, -10, 8, 14, -9, 0, 13,
    -- filter=120 channel=75
    9, 11, 1, -2, 2, -5, 9, -2, 5,
    -- filter=120 channel=76
    -6, 4, -2, -3, -1, 1, 3, -7, 0,
    -- filter=120 channel=77
    5, -5, 8, -4, -1, 7, -3, 7, -3,
    -- filter=120 channel=78
    1, -9, 0, 3, -10, 6, -7, -6, -2,
    -- filter=120 channel=79
    -4, 17, -4, -3, -1, 13, 3, 0, 8,
    -- filter=120 channel=80
    0, 7, 9, -34, -15, 19, -15, -19, 5,
    -- filter=120 channel=81
    -6, 0, 1, 5, -3, 5, 0, 6, -1,
    -- filter=120 channel=82
    4, -3, -6, -1, 0, -2, 5, 0, 5,
    -- filter=120 channel=83
    -8, 3, 3, -3, -8, -4, -3, -4, -11,
    -- filter=120 channel=84
    6, -3, -1, -4, -5, 3, 3, 2, -8,
    -- filter=120 channel=85
    -1, -4, 1, 3, 1, -6, -6, 5, 7,
    -- filter=120 channel=86
    5, 6, 1, 2, -1, -2, 10, 2, 2,
    -- filter=120 channel=87
    5, 1, -11, -5, -2, 5, 9, 8, 7,
    -- filter=120 channel=88
    -10, -2, 6, -10, 2, 4, -12, 3, 10,
    -- filter=120 channel=89
    -6, 3, -1, -22, -18, 9, -17, -19, 5,
    -- filter=120 channel=90
    4, -12, 2, 0, -4, 2, -7, -9, 6,
    -- filter=120 channel=91
    6, 13, -7, -14, -1, 14, 4, -2, -1,
    -- filter=120 channel=92
    11, 2, 3, -3, 7, 8, -3, 2, 1,
    -- filter=120 channel=93
    17, 6, 12, -6, -19, 0, 3, -10, -6,
    -- filter=120 channel=94
    4, 5, -1, -1, -5, 2, -6, 1, 5,
    -- filter=120 channel=95
    -4, 3, 0, 7, -3, -1, -1, -1, -1,
    -- filter=120 channel=96
    -3, 3, -2, -6, -4, -3, 3, -7, 4,
    -- filter=120 channel=97
    1, 10, -5, -1, 3, 1, -5, 4, 5,
    -- filter=120 channel=98
    0, 3, 8, -16, -10, 11, -4, -6, 4,
    -- filter=120 channel=99
    -5, 1, -14, -27, -6, 14, -23, -13, 12,
    -- filter=120 channel=100
    -9, -9, -2, -6, 2, -1, 0, 6, -2,
    -- filter=120 channel=101
    5, 5, 0, 6, -1, -5, 5, 8, -4,
    -- filter=120 channel=102
    0, 3, -1, -5, 6, 5, -4, -1, -1,
    -- filter=120 channel=103
    1, 8, 4, -16, -9, 19, -7, -10, 6,
    -- filter=120 channel=104
    0, -4, 13, -27, -15, 10, -6, -18, 5,
    -- filter=120 channel=105
    0, 4, 4, 4, -3, -1, 3, 2, 8,
    -- filter=120 channel=106
    -6, -6, -6, 3, 4, -6, -8, 8, 0,
    -- filter=120 channel=107
    11, 7, -5, 16, 11, 2, 11, 12, 0,
    -- filter=120 channel=108
    0, 4, 4, -11, -7, -1, -4, 2, 4,
    -- filter=120 channel=109
    3, 8, -2, -24, -2, 9, -9, -14, 2,
    -- filter=120 channel=110
    4, -4, 5, -14, -7, -1, -1, -4, 2,
    -- filter=120 channel=111
    -8, 0, -3, -1, 1, -5, -1, -7, 3,
    -- filter=120 channel=112
    0, 11, 4, -8, 7, 10, -1, -4, 8,
    -- filter=120 channel=113
    4, 6, -3, -7, 4, 11, 0, 0, 2,
    -- filter=120 channel=114
    8, 11, -17, -2, 0, -4, 0, -3, -11,
    -- filter=120 channel=115
    5, 3, 0, -8, 1, -5, 5, 3, -6,
    -- filter=120 channel=116
    -8, 7, 2, -13, -19, 4, -4, -13, 0,
    -- filter=120 channel=117
    1, -1, 5, -1, -9, -2, -3, 4, 3,
    -- filter=120 channel=118
    -1, 0, 6, -7, -6, 0, 1, -6, -5,
    -- filter=120 channel=119
    -3, -8, 13, -8, 0, 8, -11, 10, 18,
    -- filter=120 channel=120
    8, 7, -15, -24, 5, 18, -8, 2, 5,
    -- filter=120 channel=121
    -6, -4, -5, -1, -1, 3, -10, -12, 8,
    -- filter=120 channel=122
    2, 5, 21, -21, -19, 16, -4, -25, 13,
    -- filter=120 channel=123
    0, -4, 3, 5, 2, 5, -2, 8, 14,
    -- filter=120 channel=124
    7, -5, 1, -1, -1, -4, 1, -3, -1,
    -- filter=120 channel=125
    -8, 9, 2, -26, -11, 19, -15, -8, 2,
    -- filter=120 channel=126
    -14, -4, 4, -10, -6, -3, -14, -12, 8,
    -- filter=120 channel=127
    1, 0, 6, 1, 0, 0, -3, 3, 9,
    -- filter=121 channel=0
    4, 5, -3, -14, 2, 18, -4, -4, 10,
    -- filter=121 channel=1
    0, 0, 12, -14, -10, 12, -7, 2, 11,
    -- filter=121 channel=2
    -5, -4, 0, 2, -6, -2, 3, 0, -6,
    -- filter=121 channel=3
    7, -9, -6, -9, -4, -7, 1, -2, 5,
    -- filter=121 channel=4
    -1, 4, 5, -2, -9, -3, -5, -2, -3,
    -- filter=121 channel=5
    0, 3, -9, -9, 10, 6, 0, 4, -1,
    -- filter=121 channel=6
    -4, 1, -1, -1, -1, -2, -8, -9, 8,
    -- filter=121 channel=7
    -3, -5, 0, -5, 4, 5, -3, 6, 2,
    -- filter=121 channel=8
    -7, 9, 1, 0, -5, 2, 4, 3, 3,
    -- filter=121 channel=9
    -1, 4, -8, 3, 9, 6, -5, 2, -8,
    -- filter=121 channel=10
    -3, -1, -6, -13, 4, 9, -12, -1, 9,
    -- filter=121 channel=11
    -5, 0, 3, 7, -3, -3, 0, -5, 4,
    -- filter=121 channel=12
    -6, 2, 8, -9, 0, 2, -10, -4, 1,
    -- filter=121 channel=13
    -17, -8, 6, -21, -3, 17, -16, -3, 11,
    -- filter=121 channel=14
    1, -1, 5, -6, 0, 4, -5, 5, 3,
    -- filter=121 channel=15
    -8, -7, 0, -18, -5, 8, -7, -1, 6,
    -- filter=121 channel=16
    -4, 7, -1, -12, 11, 3, -12, 9, 3,
    -- filter=121 channel=17
    -6, 0, -5, 2, 0, -4, -3, -3, -5,
    -- filter=121 channel=18
    -17, -14, 4, -27, -17, 10, -12, -10, 11,
    -- filter=121 channel=19
    -2, 5, 6, -4, -4, 0, 2, -5, -3,
    -- filter=121 channel=20
    -3, -5, 1, 4, -2, -5, -8, 0, 6,
    -- filter=121 channel=21
    -2, 7, -10, -11, 9, -10, -12, 10, -6,
    -- filter=121 channel=22
    -4, -3, 4, -5, -6, 7, -7, 0, 2,
    -- filter=121 channel=23
    -14, 0, -3, -8, 9, 7, -12, 3, 8,
    -- filter=121 channel=24
    0, 6, 2, -5, -4, 1, -4, -6, -4,
    -- filter=121 channel=25
    -16, 3, 4, -27, 9, 18, -16, -5, 7,
    -- filter=121 channel=26
    3, 9, 5, 7, 10, 0, 0, 0, 3,
    -- filter=121 channel=27
    -19, 5, 3, -18, 11, 17, -10, -5, 8,
    -- filter=121 channel=28
    -3, -1, 1, -6, 4, -3, 0, -4, -2,
    -- filter=121 channel=29
    -6, -6, 10, -5, -7, 5, 1, -14, 3,
    -- filter=121 channel=30
    1, 2, -4, -3, 5, 5, 4, 5, 4,
    -- filter=121 channel=31
    -6, 11, -7, -4, 24, -3, -14, 18, 0,
    -- filter=121 channel=32
    -16, 2, 9, -29, 0, 16, -17, -10, 6,
    -- filter=121 channel=33
    -12, -3, 3, -21, 7, 18, -19, -4, 12,
    -- filter=121 channel=34
    -12, 0, 16, 5, 5, 16, -7, 0, 15,
    -- filter=121 channel=35
    -1, 6, -1, 5, 5, -3, -5, 5, 3,
    -- filter=121 channel=36
    0, -1, 0, 6, -2, -1, -8, -7, -4,
    -- filter=121 channel=37
    -6, -2, 10, -17, 7, 18, -9, 0, 2,
    -- filter=121 channel=38
    0, -4, -5, -1, 4, 7, -9, 3, -1,
    -- filter=121 channel=39
    0, -6, -2, 5, -11, -3, -1, -3, 3,
    -- filter=121 channel=40
    -2, 0, 4, -3, -4, 3, -7, -9, 4,
    -- filter=121 channel=41
    -14, -1, 10, -36, -18, 21, -26, -9, 10,
    -- filter=121 channel=42
    -1, 0, 7, -8, 1, 2, 2, 0, 3,
    -- filter=121 channel=43
    -1, 3, 1, -1, -5, -5, 0, -1, 1,
    -- filter=121 channel=44
    -8, 8, -1, -6, 9, 15, 2, 14, 9,
    -- filter=121 channel=45
    9, -2, -4, 7, 0, 0, -3, -5, 1,
    -- filter=121 channel=46
    -6, 4, 3, -8, 4, -2, 5, 2, 6,
    -- filter=121 channel=47
    -15, -4, -1, -12, 19, 2, -16, 7, -2,
    -- filter=121 channel=48
    -12, 6, 9, -11, 6, 13, -8, -1, -8,
    -- filter=121 channel=49
    -14, -4, 12, -6, -13, -2, 0, -5, 3,
    -- filter=121 channel=50
    0, -3, -4, 1, 2, 9, 3, 0, 0,
    -- filter=121 channel=51
    5, 3, -2, -3, 5, -5, -3, -2, 5,
    -- filter=121 channel=52
    3, 5, 1, 0, -4, 8, -8, 1, 4,
    -- filter=121 channel=53
    3, 1, -1, -4, -5, 6, 1, 4, 3,
    -- filter=121 channel=54
    6, -4, 6, -1, 4, 0, -3, 7, 1,
    -- filter=121 channel=55
    -15, -1, 0, -11, -9, 3, -15, 0, 2,
    -- filter=121 channel=56
    -3, 0, 5, 4, -2, 8, 0, 0, 5,
    -- filter=121 channel=57
    -2, -3, 5, 0, -4, 5, -2, 5, 8,
    -- filter=121 channel=58
    9, 7, 0, -5, 0, 3, 1, 1, 1,
    -- filter=121 channel=59
    -13, 4, 0, -23, 14, 11, -21, -5, -2,
    -- filter=121 channel=60
    3, 2, -4, 0, 0, -2, -4, 5, -5,
    -- filter=121 channel=61
    -7, 4, 0, 5, 8, -3, 4, 4, -7,
    -- filter=121 channel=62
    1, -7, -2, -4, -7, -1, -7, -5, -5,
    -- filter=121 channel=63
    3, -4, -4, 0, -1, -6, -5, 0, 3,
    -- filter=121 channel=64
    2, -3, 4, 8, -5, -11, -6, 1, -6,
    -- filter=121 channel=65
    4, 1, -1, 2, 0, -6, -1, -3, 0,
    -- filter=121 channel=66
    -14, -8, 2, -13, 2, 11, -17, 0, 12,
    -- filter=121 channel=67
    -5, -2, 7, -4, -4, 1, -1, -4, -3,
    -- filter=121 channel=68
    -1, -3, 6, -3, -3, -7, 7, -8, -4,
    -- filter=121 channel=69
    -6, 3, -6, -10, -6, 4, -2, 2, 1,
    -- filter=121 channel=70
    -14, -2, 4, -12, -1, 17, -11, 5, 12,
    -- filter=121 channel=71
    1, 0, -5, 3, 3, 0, -10, 0, 0,
    -- filter=121 channel=72
    -9, 0, 0, -5, 14, -5, -8, 4, -1,
    -- filter=121 channel=73
    -6, -10, 3, -14, -4, 0, -1, 0, -3,
    -- filter=121 channel=74
    -5, 6, 4, 5, 9, 10, -11, 9, 7,
    -- filter=121 channel=75
    -7, -7, -7, -18, -7, 20, -15, 5, 20,
    -- filter=121 channel=76
    -2, -9, 9, 0, -9, 2, -8, -12, 2,
    -- filter=121 channel=77
    -3, 0, 5, 1, 2, -5, 6, 4, 0,
    -- filter=121 channel=78
    1, -4, 0, 4, 4, 1, -5, 8, -2,
    -- filter=121 channel=79
    -13, -8, 13, -35, -12, 20, -19, -9, 13,
    -- filter=121 channel=80
    -6, 11, -16, -16, 20, 4, -14, 6, -4,
    -- filter=121 channel=81
    6, 5, 4, 3, -5, 3, 5, -5, 6,
    -- filter=121 channel=82
    0, 0, 1, -1, -5, -3, 3, 2, -4,
    -- filter=121 channel=83
    -3, 1, 5, -1, 8, -6, 0, 6, -6,
    -- filter=121 channel=84
    -6, 1, 6, -7, -6, 16, -4, -7, -1,
    -- filter=121 channel=85
    -4, 0, 3, -4, -6, -3, 5, -4, -3,
    -- filter=121 channel=86
    1, -2, 3, -2, 2, 0, 0, 1, 7,
    -- filter=121 channel=87
    -3, -4, -2, -9, -9, 6, -11, 0, -4,
    -- filter=121 channel=88
    5, 6, -4, 1, 14, -6, 6, -2, -3,
    -- filter=121 channel=89
    -14, -5, 6, -16, -5, 2, -19, 6, -2,
    -- filter=121 channel=90
    5, 0, -3, 2, 3, 0, 4, 4, 5,
    -- filter=121 channel=91
    -12, -4, 9, -22, 8, 12, -6, -2, -4,
    -- filter=121 channel=92
    0, 4, 6, -2, -4, 9, -1, 5, 5,
    -- filter=121 channel=93
    -1, 10, 6, -15, 15, 13, 4, 0, 1,
    -- filter=121 channel=94
    2, 2, 1, 0, -2, 2, 0, 5, 6,
    -- filter=121 channel=95
    1, 0, 2, 0, 4, 5, -3, 1, 1,
    -- filter=121 channel=96
    2, -2, 2, -8, -7, 5, -7, -9, 3,
    -- filter=121 channel=97
    -1, 6, -6, 0, -3, 0, -4, 2, 7,
    -- filter=121 channel=98
    -12, -5, 4, -14, 3, 15, -18, 7, 12,
    -- filter=121 channel=99
    -9, 3, -2, -9, 23, 9, -3, 5, 1,
    -- filter=121 channel=100
    -6, -3, -2, -2, 0, 6, 0, -6, 6,
    -- filter=121 channel=101
    -3, 0, 4, -4, -9, 2, 7, -7, -4,
    -- filter=121 channel=102
    2, -7, -1, 4, 3, 3, 4, 2, 6,
    -- filter=121 channel=103
    -1, -4, -10, -4, 20, 10, -13, 13, 0,
    -- filter=121 channel=104
    -15, 0, -7, -12, 15, -3, -5, 10, -8,
    -- filter=121 channel=105
    5, -6, 0, -5, -7, -1, -5, -6, -4,
    -- filter=121 channel=106
    -5, 0, -7, -2, -1, -7, -5, -8, 2,
    -- filter=121 channel=107
    -9, -5, 6, -5, -9, 7, 4, 0, 8,
    -- filter=121 channel=108
    -9, -9, 0, -4, -8, 5, -1, -7, 1,
    -- filter=121 channel=109
    -13, 1, 6, -23, 3, 21, -20, -1, 1,
    -- filter=121 channel=110
    -10, -3, -2, -10, 12, -2, -7, 6, 3,
    -- filter=121 channel=111
    0, 3, 6, 2, -3, 5, 0, -5, 4,
    -- filter=121 channel=112
    -9, 9, 7, 0, 4, 10, -12, 7, 5,
    -- filter=121 channel=113
    -7, 1, -11, -4, 5, 12, -10, 5, 10,
    -- filter=121 channel=114
    -20, -10, 6, -31, -7, 20, -18, -1, 9,
    -- filter=121 channel=115
    0, 1, -3, -7, -7, 3, -3, -3, -2,
    -- filter=121 channel=116
    -6, 1, 11, -24, 0, 11, -13, -4, -7,
    -- filter=121 channel=117
    0, -1, 6, -13, -7, -3, 3, 1, 0,
    -- filter=121 channel=118
    -1, -3, 0, 4, 0, -3, 0, 4, 0,
    -- filter=121 channel=119
    4, 7, 7, 1, 6, 17, 0, -3, 13,
    -- filter=121 channel=120
    -13, -2, 9, -13, 5, 18, -11, 3, 5,
    -- filter=121 channel=121
    -12, 3, -7, -11, -7, 8, -15, 1, 2,
    -- filter=121 channel=122
    -11, 9, -15, -6, 25, 4, -8, 11, 6,
    -- filter=121 channel=123
    0, -4, 0, 11, -2, 9, -1, 5, 0,
    -- filter=121 channel=124
    5, 1, -5, 3, 4, 3, -7, -7, -1,
    -- filter=121 channel=125
    -16, 8, 2, -10, 17, 8, -12, 7, 0,
    -- filter=121 channel=126
    -15, -3, 6, -20, -7, 1, -9, -7, 7,
    -- filter=121 channel=127
    2, 0, 8, -4, 3, -1, -7, -8, 4,
    -- filter=122 channel=0
    4, 5, -5, 13, -1, 2, 5, 3, -11,
    -- filter=122 channel=1
    14, 1, -7, 15, 2, 2, 9, -3, -1,
    -- filter=122 channel=2
    1, 4, -2, 0, -5, -1, 4, -5, -3,
    -- filter=122 channel=3
    11, 6, 5, 8, 0, -7, 11, 11, 3,
    -- filter=122 channel=4
    2, 9, 0, 8, 9, 7, 1, 0, 9,
    -- filter=122 channel=5
    -4, -5, -8, 10, -7, -3, 8, -5, -5,
    -- filter=122 channel=6
    -6, -4, 2, 6, 6, -1, 1, -5, 1,
    -- filter=122 channel=7
    -7, 4, -7, 5, -1, -4, -5, -3, 5,
    -- filter=122 channel=8
    0, 2, 9, 4, 0, 5, 6, 1, 2,
    -- filter=122 channel=9
    4, -7, -1, -3, -5, -2, 3, 5, -7,
    -- filter=122 channel=10
    -7, -8, -5, -5, 3, -4, -5, -4, 0,
    -- filter=122 channel=11
    2, 0, -6, -7, 5, -7, -8, 3, 4,
    -- filter=122 channel=12
    5, 7, 5, 7, 2, 1, 0, 0, 0,
    -- filter=122 channel=13
    4, -5, -2, -5, -4, 11, -6, 7, 11,
    -- filter=122 channel=14
    -4, -2, 0, 1, -1, 0, 6, 0, -6,
    -- filter=122 channel=15
    -3, -5, -2, -5, 6, -6, 5, -5, 0,
    -- filter=122 channel=16
    5, -8, 4, 1, 2, 0, 2, 6, 5,
    -- filter=122 channel=17
    7, 4, 1, -6, 6, -6, 5, -4, -5,
    -- filter=122 channel=18
    1, -6, -2, -2, 0, 9, 0, 1, 1,
    -- filter=122 channel=19
    3, -5, 5, 4, 4, 0, 0, -2, 4,
    -- filter=122 channel=20
    -3, 2, -3, 0, -6, -4, -5, 2, -4,
    -- filter=122 channel=21
    3, -1, 5, -10, 0, 0, -5, 1, 11,
    -- filter=122 channel=22
    -1, -3, 0, 3, -1, -4, -2, 0, -6,
    -- filter=122 channel=23
    2, -10, 3, -1, 2, -4, -6, 3, 8,
    -- filter=122 channel=24
    2, -6, 4, 4, 2, 4, -4, 2, -4,
    -- filter=122 channel=25
    3, -12, -2, -2, -6, 1, -10, 6, 2,
    -- filter=122 channel=26
    1, -5, 0, -1, 1, -1, 5, 0, 0,
    -- filter=122 channel=27
    1, -8, 0, -6, -6, 4, -4, 2, -2,
    -- filter=122 channel=28
    7, 0, 7, -3, 3, -3, -2, -5, -2,
    -- filter=122 channel=29
    4, 1, 1, -6, -8, -4, -5, 3, 0,
    -- filter=122 channel=30
    5, 4, -10, 3, 6, -4, -3, 7, 3,
    -- filter=122 channel=31
    -8, -4, -13, -14, 5, 5, 0, 16, 6,
    -- filter=122 channel=32
    0, -5, -7, -6, -8, 0, -7, -4, 4,
    -- filter=122 channel=33
    1, -3, -9, -6, -2, -4, -3, -3, 6,
    -- filter=122 channel=34
    -3, 3, 6, 2, -1, 0, -1, 10, 0,
    -- filter=122 channel=35
    0, 0, -6, -6, 1, 3, -7, 6, -6,
    -- filter=122 channel=36
    -6, 6, 1, 0, 3, 14, 6, 4, 6,
    -- filter=122 channel=37
    0, 0, 4, 15, 4, -7, 13, 8, -6,
    -- filter=122 channel=38
    -3, -6, -7, 2, 2, 0, -5, -5, 8,
    -- filter=122 channel=39
    -5, -7, -1, 5, -2, -1, -3, 4, -1,
    -- filter=122 channel=40
    8, 9, -1, 0, -3, -1, 1, 2, 1,
    -- filter=122 channel=41
    9, 0, 4, -5, 5, 11, 4, -6, 4,
    -- filter=122 channel=42
    -3, 4, 1, 1, -6, 2, -6, -6, -6,
    -- filter=122 channel=43
    -2, 6, 0, -1, -2, 0, 0, 5, -3,
    -- filter=122 channel=44
    0, -10, 1, 7, 7, -7, 2, 4, 0,
    -- filter=122 channel=45
    5, 0, -4, 0, 5, -5, 0, -6, -2,
    -- filter=122 channel=46
    -4, -1, 5, 6, 4, 3, 0, 0, -3,
    -- filter=122 channel=47
    0, -12, 0, -4, -9, -2, -2, 1, 5,
    -- filter=122 channel=48
    3, -2, -7, -11, 2, 3, -1, -4, 0,
    -- filter=122 channel=49
    6, 6, 0, -6, -1, 4, -6, -5, -2,
    -- filter=122 channel=50
    -6, -5, -5, -4, -4, -7, -1, 0, 6,
    -- filter=122 channel=51
    5, 3, 1, -4, -3, 0, -6, -7, -3,
    -- filter=122 channel=52
    5, -2, 0, -4, 9, 6, -2, 3, 6,
    -- filter=122 channel=53
    1, 0, -4, -6, -2, 4, -7, -5, -5,
    -- filter=122 channel=54
    -1, -5, -1, -5, 4, -2, 4, 7, 0,
    -- filter=122 channel=55
    -5, 0, 0, 0, -1, 8, -10, 7, 2,
    -- filter=122 channel=56
    3, -1, 3, 3, 1, -4, 6, 4, 2,
    -- filter=122 channel=57
    1, 1, 0, -2, 1, 0, 1, 0, -4,
    -- filter=122 channel=58
    -1, -5, 1, 10, -1, 1, 5, 4, -5,
    -- filter=122 channel=59
    5, -12, -8, -10, -8, 4, 0, 1, 0,
    -- filter=122 channel=60
    5, 6, 1, -1, 5, 3, -1, 2, -6,
    -- filter=122 channel=61
    -3, -6, 0, -4, 2, -2, -6, 0, 7,
    -- filter=122 channel=62
    -2, 4, 3, 6, 0, -6, 0, 6, -1,
    -- filter=122 channel=63
    0, 2, -6, 0, 1, 0, 6, -3, -5,
    -- filter=122 channel=64
    5, 6, 5, -3, -4, 5, 5, -5, -3,
    -- filter=122 channel=65
    2, -7, -4, -2, 4, 4, 3, -1, 5,
    -- filter=122 channel=66
    6, 0, 3, -6, 7, 12, 4, 7, 6,
    -- filter=122 channel=67
    -6, 6, 0, 2, -5, -6, -3, -2, -7,
    -- filter=122 channel=68
    -2, -3, -4, -5, -4, 10, 0, 7, 1,
    -- filter=122 channel=69
    7, 0, 5, -2, 0, 6, 0, -1, 7,
    -- filter=122 channel=70
    5, -6, 1, 8, 3, 0, 3, -3, -3,
    -- filter=122 channel=71
    6, 1, 3, 3, 5, 6, 2, 3, 8,
    -- filter=122 channel=72
    -9, -7, -11, -7, 0, 8, -6, 3, 2,
    -- filter=122 channel=73
    1, 3, -7, 0, -8, 8, -8, -1, 2,
    -- filter=122 channel=74
    3, 2, 6, 3, 4, 0, 6, 0, 2,
    -- filter=122 channel=75
    5, -7, -14, 10, -3, -9, 1, 0, -4,
    -- filter=122 channel=76
    -1, 9, 0, -2, -3, -1, -5, 2, -2,
    -- filter=122 channel=77
    7, 4, 1, -6, 7, 0, -1, -7, -6,
    -- filter=122 channel=78
    3, 2, 0, 6, -2, -3, -4, -6, -3,
    -- filter=122 channel=79
    1, 0, -2, -3, -7, 7, 1, -4, 3,
    -- filter=122 channel=80
    -8, -9, -11, -11, -2, 7, -10, 1, 12,
    -- filter=122 channel=81
    -1, 1, 6, 1, -7, -2, 4, 0, -2,
    -- filter=122 channel=82
    1, -2, 0, 7, 5, -7, 7, -3, -1,
    -- filter=122 channel=83
    -6, -2, -5, 0, -7, -4, -6, 4, 1,
    -- filter=122 channel=84
    2, -1, -2, 0, 4, -2, -6, 7, 1,
    -- filter=122 channel=85
    -2, -2, 2, -7, -6, -6, -1, -5, 3,
    -- filter=122 channel=86
    -4, -2, 4, 0, -3, -6, 1, 9, 1,
    -- filter=122 channel=87
    -1, -1, 5, 5, 1, -4, -1, 7, 3,
    -- filter=122 channel=88
    -8, 1, -1, -4, -3, 8, 4, 12, 2,
    -- filter=122 channel=89
    0, -4, -3, -1, -11, 9, -10, 4, 8,
    -- filter=122 channel=90
    0, 0, 3, 1, 0, 0, -1, 10, 7,
    -- filter=122 channel=91
    6, -4, -3, -5, -4, 0, -4, -6, 7,
    -- filter=122 channel=92
    -2, 3, 7, 3, 0, 4, 1, -5, 1,
    -- filter=122 channel=93
    6, -7, -9, -5, 2, 5, -4, 7, 5,
    -- filter=122 channel=94
    0, 3, 5, 1, 2, -6, 5, 0, -3,
    -- filter=122 channel=95
    0, 0, 7, -3, 2, 1, -5, -5, 4,
    -- filter=122 channel=96
    2, -4, -1, -7, 3, 1, -6, 2, 3,
    -- filter=122 channel=97
    -2, -4, -6, 6, -6, -5, 8, -1, 1,
    -- filter=122 channel=98
    2, -7, -14, -6, -8, 1, -2, -7, 8,
    -- filter=122 channel=99
    -13, -15, -10, -4, 4, -1, -9, 14, -1,
    -- filter=122 channel=100
    -4, 0, -3, 5, 0, -5, 6, -2, -4,
    -- filter=122 channel=101
    9, 3, 9, -2, 8, -2, 1, 11, 7,
    -- filter=122 channel=102
    0, 3, 6, -6, -3, -3, -5, 1, -2,
    -- filter=122 channel=103
    4, -9, -2, 2, -2, 0, 3, 3, -1,
    -- filter=122 channel=104
    -9, -14, 1, -1, 0, -2, -7, 0, 1,
    -- filter=122 channel=105
    1, 4, -1, 0, 3, 0, -2, 5, 0,
    -- filter=122 channel=106
    -5, 8, 0, -5, 5, -4, 2, 0, -2,
    -- filter=122 channel=107
    6, 4, -5, 11, 5, 7, 4, 0, -2,
    -- filter=122 channel=108
    0, 6, 0, 2, 4, 5, -1, -7, 6,
    -- filter=122 channel=109
    4, -7, -2, -9, -2, 6, -2, 1, 2,
    -- filter=122 channel=110
    -9, -7, -3, -3, 2, 4, -7, 4, 10,
    -- filter=122 channel=111
    4, -1, -1, -8, 5, 3, -6, -7, 1,
    -- filter=122 channel=112
    -6, -1, -5, 0, -3, -1, 0, -4, -4,
    -- filter=122 channel=113
    -1, -9, 1, 3, -4, 6, -7, 8, 8,
    -- filter=122 channel=114
    10, -2, -6, 0, 5, -3, -1, -8, -7,
    -- filter=122 channel=115
    6, 2, 0, 1, 1, -1, -6, -6, -7,
    -- filter=122 channel=116
    -4, -11, -3, -11, -1, 1, -7, 7, 0,
    -- filter=122 channel=117
    -6, 4, 7, -1, -3, 8, -7, 5, 6,
    -- filter=122 channel=118
    -7, 2, -6, -4, 3, -1, 5, -3, 2,
    -- filter=122 channel=119
    0, 0, 6, -5, -2, 3, -3, 7, 0,
    -- filter=122 channel=120
    5, -5, 2, 1, -2, 0, -5, -3, -7,
    -- filter=122 channel=121
    -3, -1, -3, -5, 8, 6, -3, 3, 0,
    -- filter=122 channel=122
    0, -14, -2, -5, 0, 12, -5, 11, 14,
    -- filter=122 channel=123
    -7, 3, -1, 4, 1, -4, 8, 1, 5,
    -- filter=122 channel=124
    -4, 6, -5, -3, 6, -3, 0, -1, 1,
    -- filter=122 channel=125
    0, -6, -7, -6, -8, 1, -11, 4, 0,
    -- filter=122 channel=126
    -2, -6, -8, -4, -7, -5, -1, 6, 0,
    -- filter=122 channel=127
    3, 3, 7, -7, 2, 0, -6, 4, 2,
    -- filter=123 channel=0
    -5, -3, -5, 2, 10, 3, 2, 17, 16,
    -- filter=123 channel=1
    -2, -4, 4, 5, 9, 6, 0, 10, 6,
    -- filter=123 channel=2
    -4, 1, 5, -4, -3, 1, -4, 0, 4,
    -- filter=123 channel=3
    0, 3, -1, 7, -3, 2, 0, -5, 2,
    -- filter=123 channel=4
    5, -1, 3, 9, 2, -7, 7, 3, 2,
    -- filter=123 channel=5
    -5, 6, 3, 1, 17, 15, 9, 15, 7,
    -- filter=123 channel=6
    0, 0, 0, -2, -6, -6, 1, -5, 4,
    -- filter=123 channel=7
    -3, 0, -6, -7, 4, 2, 2, -1, 0,
    -- filter=123 channel=8
    0, -1, 3, 0, 6, -5, 4, -5, -5,
    -- filter=123 channel=9
    -1, 0, -2, -9, 3, -1, 2, 3, -2,
    -- filter=123 channel=10
    -9, -4, 2, -13, -1, 2, -11, -11, 2,
    -- filter=123 channel=11
    -6, 4, -7, 4, 1, -1, -5, -5, 0,
    -- filter=123 channel=12
    -1, 6, -3, -7, -3, -3, 0, 4, -5,
    -- filter=123 channel=13
    -13, -4, -4, -18, -6, -9, -8, -4, -12,
    -- filter=123 channel=14
    4, -5, -2, 0, 4, -6, -7, 1, -6,
    -- filter=123 channel=15
    -12, 0, -8, -8, -2, -6, 1, -11, -5,
    -- filter=123 channel=16
    -6, 2, 9, -1, 0, 4, 2, 3, 3,
    -- filter=123 channel=17
    1, 3, -5, -4, -6, 0, 2, -2, 6,
    -- filter=123 channel=18
    -17, -10, -7, -14, -9, -16, -6, -6, -16,
    -- filter=123 channel=19
    4, 1, -1, 5, 1, 4, -2, 0, 2,
    -- filter=123 channel=20
    -4, 1, -8, -5, -5, -9, 5, -11, -3,
    -- filter=123 channel=21
    -2, 1, 11, -9, -2, 4, -8, -1, 10,
    -- filter=123 channel=22
    8, -1, -8, -4, 3, 0, -3, -3, 3,
    -- filter=123 channel=23
    -5, 8, -11, -12, -13, -6, -6, -4, -17,
    -- filter=123 channel=24
    -1, 0, -5, 4, 5, 7, -1, 0, 6,
    -- filter=123 channel=25
    -14, 10, 4, -19, -1, -1, -16, 0, -7,
    -- filter=123 channel=26
    5, 2, 1, 1, 10, 1, 7, 7, 1,
    -- filter=123 channel=27
    -14, 3, -8, -22, -4, -6, -8, 1, 0,
    -- filter=123 channel=28
    3, 5, -3, 6, -1, -3, 0, 3, -1,
    -- filter=123 channel=29
    -6, -7, -3, -5, 2, 4, -3, 1, -6,
    -- filter=123 channel=30
    -6, 8, 7, -3, 0, -4, -3, 10, 0,
    -- filter=123 channel=31
    -6, 5, 3, -8, 0, 6, -13, 1, -4,
    -- filter=123 channel=32
    -7, 2, -3, -14, -11, -13, -10, -6, -6,
    -- filter=123 channel=33
    -9, 7, -7, -12, -4, 0, -7, -10, -7,
    -- filter=123 channel=34
    10, 5, 3, -2, 3, 2, -4, 8, 1,
    -- filter=123 channel=35
    5, -4, 3, -1, -3, -1, 1, -4, -1,
    -- filter=123 channel=36
    -1, 3, 3, -10, -8, -7, -6, -5, 5,
    -- filter=123 channel=37
    -3, 8, 6, 2, 15, 4, 7, 13, 12,
    -- filter=123 channel=38
    1, 11, -5, -12, 4, -4, -8, 4, 1,
    -- filter=123 channel=39
    -1, 4, -8, 2, 0, 0, -6, -7, -9,
    -- filter=123 channel=40
    -4, 5, -5, -2, 0, -1, 7, -7, -3,
    -- filter=123 channel=41
    -5, -7, 8, -8, -16, -2, -11, -9, 4,
    -- filter=123 channel=42
    -8, 1, -1, -3, -7, -4, 0, 0, 3,
    -- filter=123 channel=43
    0, 0, 3, 9, 3, -5, 5, 4, 2,
    -- filter=123 channel=44
    -4, 9, 10, 0, -1, -1, -11, 10, 8,
    -- filter=123 channel=45
    -3, -6, 5, -3, -6, -6, 5, -3, -6,
    -- filter=123 channel=46
    3, 5, 7, 2, 0, -5, 1, -7, 7,
    -- filter=123 channel=47
    0, 4, 17, -4, 14, 17, -6, 8, 9,
    -- filter=123 channel=48
    -10, 3, 5, -19, -3, 4, -15, -5, 4,
    -- filter=123 channel=49
    -6, 0, -1, -8, -4, -8, -6, 3, -5,
    -- filter=123 channel=50
    -8, 5, 1, -16, -2, 0, -11, -7, -9,
    -- filter=123 channel=51
    1, 3, -2, 2, 7, -7, 3, 0, 0,
    -- filter=123 channel=52
    2, 2, -2, -5, 3, 3, -4, 2, -8,
    -- filter=123 channel=53
    0, -4, -8, -9, -8, -8, -3, -3, -6,
    -- filter=123 channel=54
    3, 6, -7, -6, -3, 6, -3, 3, -2,
    -- filter=123 channel=55
    -1, 4, -1, -6, -5, -9, -7, -14, -12,
    -- filter=123 channel=56
    -6, -1, -1, -2, -7, 4, 1, -1, -8,
    -- filter=123 channel=57
    -7, 4, 0, -4, -3, 6, -1, -6, -4,
    -- filter=123 channel=58
    1, -3, 8, 1, 14, 4, 6, 0, 3,
    -- filter=123 channel=59
    -15, 3, 1, -19, -5, 5, -24, -2, -8,
    -- filter=123 channel=60
    -3, 0, 4, -3, -2, 0, 0, 0, 0,
    -- filter=123 channel=61
    -6, 1, -2, -3, -4, -7, 0, 1, -6,
    -- filter=123 channel=62
    2, -2, -1, -5, 2, 1, -1, 6, -4,
    -- filter=123 channel=63
    9, 7, 11, 0, 11, 5, 3, 13, 4,
    -- filter=123 channel=64
    -6, 4, 1, -2, 5, 3, 3, -7, -8,
    -- filter=123 channel=65
    -2, 7, -7, 5, 0, 5, 1, -2, -5,
    -- filter=123 channel=66
    -2, -1, 0, 2, -4, -6, -4, 2, -6,
    -- filter=123 channel=67
    5, 0, 3, -1, 4, -3, 2, -5, 0,
    -- filter=123 channel=68
    -7, -1, 5, 3, -4, -3, -2, 4, -7,
    -- filter=123 channel=69
    0, -4, -2, -8, -1, -6, 0, 0, 6,
    -- filter=123 channel=70
    3, 6, -3, -17, -5, -8, -4, -1, -8,
    -- filter=123 channel=71
    8, 0, -6, -1, 1, 5, 1, -4, -7,
    -- filter=123 channel=72
    -16, 1, 0, -18, -2, -2, -7, -11, -9,
    -- filter=123 channel=73
    0, -8, -1, -11, 2, -6, -3, 0, -8,
    -- filter=123 channel=74
    1, 7, 4, -6, 5, 2, 4, 4, -2,
    -- filter=123 channel=75
    2, 5, 0, -6, 14, 9, -12, 13, 12,
    -- filter=123 channel=76
    -1, 4, -5, 3, 1, -4, -1, -9, -3,
    -- filter=123 channel=77
    -6, -4, -5, -2, -3, -4, 5, -4, 3,
    -- filter=123 channel=78
    2, -1, 4, -5, -1, 5, -7, 10, 8,
    -- filter=123 channel=79
    -19, -10, -16, -13, -7, -12, -20, -6, -9,
    -- filter=123 channel=80
    -21, 12, 11, -26, -9, 1, -20, 0, -3,
    -- filter=123 channel=81
    -2, -2, -1, -1, -6, 1, -3, 2, 3,
    -- filter=123 channel=82
    7, 1, 5, 3, 3, 6, 5, 3, -3,
    -- filter=123 channel=83
    1, -2, -2, -3, -6, 0, -9, -4, -3,
    -- filter=123 channel=84
    1, 5, 0, 1, -4, -4, -9, 1, -4,
    -- filter=123 channel=85
    -3, 2, 0, 0, 6, 4, -5, 1, 1,
    -- filter=123 channel=86
    2, 0, -5, 3, 13, -1, 9, 0, 3,
    -- filter=123 channel=87
    -4, 5, 0, 1, 4, 5, 6, 4, 1,
    -- filter=123 channel=88
    -6, -2, 1, -3, -5, 0, -5, -7, -5,
    -- filter=123 channel=89
    -14, -6, 3, -12, -5, -8, -17, -14, -5,
    -- filter=123 channel=90
    -1, 0, 4, 6, -1, 1, -2, 4, 3,
    -- filter=123 channel=91
    -13, -2, 3, -7, 0, 0, 0, -3, 1,
    -- filter=123 channel=92
    8, 2, 4, 0, 0, -1, 4, 1, -6,
    -- filter=123 channel=93
    -4, 1, 0, -2, 5, 8, 1, 2, 13,
    -- filter=123 channel=94
    -2, 2, 5, -2, -2, -3, -7, 2, 5,
    -- filter=123 channel=95
    -7, -2, -3, -4, -5, 7, 6, 3, -5,
    -- filter=123 channel=96
    3, 4, -6, -4, -5, 3, -10, 1, -1,
    -- filter=123 channel=97
    6, -3, 4, 0, -2, 9, -4, 1, 4,
    -- filter=123 channel=98
    -7, 9, 3, -11, -9, 7, -11, 1, -5,
    -- filter=123 channel=99
    0, 14, 0, -11, -2, 0, -4, -9, -8,
    -- filter=123 channel=100
    2, 1, -3, -3, -4, 1, -1, -1, 0,
    -- filter=123 channel=101
    -7, -3, 2, 6, -5, 0, -1, -3, 1,
    -- filter=123 channel=102
    6, 7, -1, -6, 2, -5, 7, -1, -7,
    -- filter=123 channel=103
    -1, 11, 7, -15, 12, 12, -11, 6, 13,
    -- filter=123 channel=104
    -16, 9, 9, -13, 3, 3, -8, 4, 8,
    -- filter=123 channel=105
    5, 1, 0, -3, 3, -8, -7, -1, 0,
    -- filter=123 channel=106
    0, -3, -5, -4, -8, 5, 1, -6, 2,
    -- filter=123 channel=107
    -3, -2, 0, 5, 1, 0, -4, 4, 0,
    -- filter=123 channel=108
    -6, -1, 5, 1, 0, 0, 0, -2, -1,
    -- filter=123 channel=109
    -18, 7, -4, -15, -7, -10, -18, -1, 1,
    -- filter=123 channel=110
    0, -1, 5, -12, 4, 0, -12, -8, 5,
    -- filter=123 channel=111
    0, -7, -5, -7, 3, 1, 3, 1, 7,
    -- filter=123 channel=112
    0, -4, -3, 0, 5, -1, -2, 0, 5,
    -- filter=123 channel=113
    -9, 1, -1, -5, 4, 1, -11, 3, -4,
    -- filter=123 channel=114
    -3, -1, -9, -2, 2, -9, -8, 2, -2,
    -- filter=123 channel=115
    4, 0, -6, -8, -7, 5, 2, 0, -7,
    -- filter=123 channel=116
    -16, 0, 5, -11, -11, -9, -7, -3, 3,
    -- filter=123 channel=117
    -5, 3, -1, -5, 0, 5, 1, -8, -8,
    -- filter=123 channel=118
    -3, 0, 4, -4, -2, -3, 6, 0, 3,
    -- filter=123 channel=119
    3, 5, 0, 3, -3, -4, 8, 3, 3,
    -- filter=123 channel=120
    0, -6, -11, -7, -9, -6, 4, 1, -7,
    -- filter=123 channel=121
    -12, 1, 0, -4, -5, -5, -2, -7, -4,
    -- filter=123 channel=122
    0, 19, 23, -17, 15, 16, -8, 1, 15,
    -- filter=123 channel=123
    -4, 4, 0, 0, 2, 4, 1, 3, 0,
    -- filter=123 channel=124
    -7, -4, -2, 2, 1, -4, -1, 4, -3,
    -- filter=123 channel=125
    -11, 10, 7, -6, -1, 2, -15, -7, -2,
    -- filter=123 channel=126
    -1, 4, -6, -11, -11, -6, -14, -7, 0,
    -- filter=123 channel=127
    4, 0, -6, -2, -3, 0, 2, -1, -6,
    -- filter=124 channel=0
    4, -5, -13, 10, 2, -15, 11, -4, -4,
    -- filter=124 channel=1
    0, 3, 3, 13, 10, 2, 0, 7, -1,
    -- filter=124 channel=2
    -6, 1, 5, -5, -8, 0, -2, 1, -2,
    -- filter=124 channel=3
    8, 6, 0, 3, -7, -4, -2, -1, -5,
    -- filter=124 channel=4
    0, -4, 3, -11, 3, 0, 3, -4, 0,
    -- filter=124 channel=5
    4, -1, 0, 14, 3, 0, 5, 1, -10,
    -- filter=124 channel=6
    -12, -11, -4, -11, -3, 2, -2, -11, -9,
    -- filter=124 channel=7
    -5, 3, -4, 4, -5, 2, -1, -2, 1,
    -- filter=124 channel=8
    8, 1, 3, 0, -4, 1, 1, -2, -1,
    -- filter=124 channel=9
    5, 6, -6, -3, 0, -1, 0, 1, 2,
    -- filter=124 channel=10
    5, 7, 4, 2, 6, -8, 0, -6, -10,
    -- filter=124 channel=11
    -13, -5, -10, -7, -3, -9, -10, -8, -10,
    -- filter=124 channel=12
    1, 5, 6, -6, 0, -9, -7, 0, -5,
    -- filter=124 channel=13
    -7, 2, 4, -7, 6, 2, 2, 5, 7,
    -- filter=124 channel=14
    5, 0, -1, 0, 2, 1, 7, 0, 1,
    -- filter=124 channel=15
    -4, -11, -12, -4, -9, -10, 0, 4, 0,
    -- filter=124 channel=16
    5, 12, 8, 9, 2, 7, -3, -6, 5,
    -- filter=124 channel=17
    5, 5, -3, 3, -4, -6, -4, 4, -1,
    -- filter=124 channel=18
    -4, 5, -7, -12, -9, -6, -6, -6, -10,
    -- filter=124 channel=19
    4, -1, -5, -7, 0, 3, -1, -2, -5,
    -- filter=124 channel=20
    -10, -6, -11, -7, -13, -3, -7, -9, -3,
    -- filter=124 channel=21
    -4, 8, 0, 12, 1, 6, -10, 1, -1,
    -- filter=124 channel=22
    5, -4, 2, -4, -4, -2, -5, 4, 2,
    -- filter=124 channel=23
    8, 5, -2, -2, -9, -7, 4, -7, 0,
    -- filter=124 channel=24
    3, 0, 0, 0, -7, -6, 1, -2, -7,
    -- filter=124 channel=25
    -4, 5, -6, 0, 8, 4, -5, 1, -1,
    -- filter=124 channel=26
    7, 1, 0, 9, 3, -4, 1, 0, -6,
    -- filter=124 channel=27
    11, -1, -13, 3, 4, -9, 0, 0, -4,
    -- filter=124 channel=28
    -7, 2, 5, -3, 2, -1, -2, 2, -6,
    -- filter=124 channel=29
    -10, -10, -5, -6, -1, -14, -3, 2, -5,
    -- filter=124 channel=30
    -2, -7, -11, 15, -5, -6, 3, 5, -8,
    -- filter=124 channel=31
    0, 1, -4, 8, -8, 0, -13, -5, -4,
    -- filter=124 channel=32
    -3, 10, -2, 0, -6, -5, -12, 3, -9,
    -- filter=124 channel=33
    1, 9, 0, -1, 1, -3, -2, 4, -1,
    -- filter=124 channel=34
    2, -2, 1, 13, -7, -8, -3, -9, -6,
    -- filter=124 channel=35
    0, -3, -1, -5, 2, 2, -3, 1, 2,
    -- filter=124 channel=36
    1, 1, -2, 0, 3, 3, -8, -7, 6,
    -- filter=124 channel=37
    1, 5, -5, 12, 12, 4, 9, -1, -3,
    -- filter=124 channel=38
    2, 3, 0, -4, 2, -9, -5, 4, -2,
    -- filter=124 channel=39
    0, -1, -3, 0, -3, 1, -2, 0, 2,
    -- filter=124 channel=40
    -2, 0, -6, -7, 0, -5, 1, -2, -3,
    -- filter=124 channel=41
    4, 7, 13, -6, 0, -3, -8, -6, 1,
    -- filter=124 channel=42
    -3, -3, 1, 0, -2, 5, -2, 6, 5,
    -- filter=124 channel=43
    -7, -11, 4, -12, -5, -13, -9, -1, -3,
    -- filter=124 channel=44
    12, 11, 0, 15, 10, 4, 0, 5, -6,
    -- filter=124 channel=45
    2, -10, -7, -7, 0, -3, 0, -8, -8,
    -- filter=124 channel=46
    0, -2, 3, 4, 5, 3, -2, 2, -2,
    -- filter=124 channel=47
    3, 14, 2, 12, 10, 4, 0, -5, 0,
    -- filter=124 channel=48
    7, 8, 1, 11, 9, -3, 0, 7, 3,
    -- filter=124 channel=49
    -11, -2, 0, -9, -3, -5, -1, 0, 0,
    -- filter=124 channel=50
    0, -6, -8, 5, 6, 4, 8, 1, -4,
    -- filter=124 channel=51
    2, 5, 5, 6, 6, 0, -1, -2, 3,
    -- filter=124 channel=52
    0, 6, -4, -6, -3, -8, -3, 2, 5,
    -- filter=124 channel=53
    -6, -3, -1, 0, -2, 1, 2, -5, -8,
    -- filter=124 channel=54
    -3, 4, -1, -5, 1, 5, 4, 0, 0,
    -- filter=124 channel=55
    -14, -12, -14, -12, -14, -19, -8, -1, -8,
    -- filter=124 channel=56
    0, -11, 8, -2, -1, -5, 0, -6, -6,
    -- filter=124 channel=57
    4, 0, 4, 0, -3, 0, 2, -6, 4,
    -- filter=124 channel=58
    4, 0, -9, 1, -8, -10, -2, -8, -12,
    -- filter=124 channel=59
    4, 11, -4, -5, 9, -6, -9, 8, -6,
    -- filter=124 channel=60
    -6, 5, 0, -5, -4, 3, 6, 2, -1,
    -- filter=124 channel=61
    -8, 0, -1, -9, -5, 3, 0, -3, 5,
    -- filter=124 channel=62
    7, 5, -6, -5, 0, 0, 0, 4, 5,
    -- filter=124 channel=63
    -2, -9, -10, 6, -10, -4, 5, -11, -4,
    -- filter=124 channel=64
    -7, 0, -1, -5, 3, -5, -5, 0, -1,
    -- filter=124 channel=65
    -3, -3, -7, 7, -5, 3, -6, -4, -3,
    -- filter=124 channel=66
    -9, 0, -3, 1, -2, 5, 0, -7, 1,
    -- filter=124 channel=67
    -4, 2, 7, 0, -7, 3, 7, 3, -5,
    -- filter=124 channel=68
    -2, 0, -2, -3, 3, 5, 0, -4, 8,
    -- filter=124 channel=69
    4, -2, -7, 3, -4, -6, -8, -1, -8,
    -- filter=124 channel=70
    0, 7, 2, 8, 1, 2, 8, 2, -3,
    -- filter=124 channel=71
    -1, 8, 0, 6, 5, 3, -1, 1, 5,
    -- filter=124 channel=72
    -9, 3, 0, -5, -6, -9, -3, 0, 1,
    -- filter=124 channel=73
    -8, 2, -1, -2, -8, -10, 2, -1, -1,
    -- filter=124 channel=74
    12, -2, -4, 11, -9, -6, -1, 0, -1,
    -- filter=124 channel=75
    12, 11, -6, 7, 10, -3, 8, 8, -12,
    -- filter=124 channel=76
    -14, -5, -10, -14, -2, -10, -10, -10, -9,
    -- filter=124 channel=77
    -5, 3, -2, 6, 0, -6, 1, 7, -5,
    -- filter=124 channel=78
    0, -1, -4, 0, -3, -3, 4, 0, -11,
    -- filter=124 channel=79
    -8, 10, -2, -10, 4, -17, -2, 6, -10,
    -- filter=124 channel=80
    2, 9, 1, 10, 5, -4, -15, -2, -5,
    -- filter=124 channel=81
    0, -5, -5, 2, 6, -5, 0, 3, -5,
    -- filter=124 channel=82
    0, -2, 5, -7, 4, 0, 3, -5, -4,
    -- filter=124 channel=83
    4, 4, 1, 6, 5, -1, 3, 0, 0,
    -- filter=124 channel=84
    -5, 0, -10, 1, -9, -1, -8, 0, -7,
    -- filter=124 channel=85
    6, 0, 3, 0, -6, 5, 0, 5, 3,
    -- filter=124 channel=86
    -2, 4, -8, 9, -9, -4, 6, -3, 0,
    -- filter=124 channel=87
    2, 1, 0, -6, -8, 0, -10, 0, -10,
    -- filter=124 channel=88
    -8, -5, 1, -4, 0, 2, -8, -2, -2,
    -- filter=124 channel=89
    -5, 10, 3, -4, -5, -1, -3, 0, -9,
    -- filter=124 channel=90
    0, -3, 7, -6, -8, 2, -4, 0, 2,
    -- filter=124 channel=91
    -1, 4, -10, -5, -2, -1, 6, 6, 0,
    -- filter=124 channel=92
    2, -5, 7, 5, -2, -6, 5, -8, 4,
    -- filter=124 channel=93
    12, 5, -3, 16, 10, -1, 7, 9, 0,
    -- filter=124 channel=94
    -2, 0, 2, -2, 6, 3, 2, 7, 4,
    -- filter=124 channel=95
    -3, 1, -5, -8, 3, 6, 0, 6, 5,
    -- filter=124 channel=96
    6, -1, 0, 2, -1, -4, 4, -2, 1,
    -- filter=124 channel=97
    0, 0, 3, -4, 10, 0, 2, 6, 1,
    -- filter=124 channel=98
    -2, 5, 1, 8, 8, 1, -2, 0, 1,
    -- filter=124 channel=99
    -2, -11, -5, -1, -10, -5, -8, -14, 2,
    -- filter=124 channel=100
    -1, -4, 6, 2, 0, -3, -4, -6, 1,
    -- filter=124 channel=101
    -5, 7, -7, 2, -6, -2, -5, -2, -3,
    -- filter=124 channel=102
    4, 1, -1, 4, 0, -5, -3, -2, 5,
    -- filter=124 channel=103
    9, 7, 0, 6, 13, 5, -3, 5, -8,
    -- filter=124 channel=104
    3, 4, -7, 0, 3, -5, -13, 1, 0,
    -- filter=124 channel=105
    -6, -8, -2, -7, -6, 3, -7, -7, -5,
    -- filter=124 channel=106
    4, -2, 0, -8, -8, 4, 6, -8, 2,
    -- filter=124 channel=107
    -3, -8, -2, -5, -19, -3, -8, -13, -12,
    -- filter=124 channel=108
    -5, 5, 6, -1, -2, -7, -3, 0, 0,
    -- filter=124 channel=109
    7, -2, -9, 6, -6, -1, -6, 8, -3,
    -- filter=124 channel=110
    3, 5, 3, -2, 3, 0, 0, -6, -8,
    -- filter=124 channel=111
    -7, 1, -6, -5, -6, 3, -7, -5, 4,
    -- filter=124 channel=112
    0, 2, 6, 2, -2, -5, 2, 3, 0,
    -- filter=124 channel=113
    4, 5, 1, 7, 6, -3, -7, 2, -6,
    -- filter=124 channel=114
    -7, -8, -15, 2, -13, -21, -9, -4, -7,
    -- filter=124 channel=115
    1, -5, 2, -4, 6, -1, 0, 0, -4,
    -- filter=124 channel=116
    -4, 2, 0, 0, -4, -8, -4, 6, 1,
    -- filter=124 channel=117
    -5, -1, -6, -1, 7, -5, 1, -5, 3,
    -- filter=124 channel=118
    2, 4, -6, -4, -3, 0, -5, 0, 4,
    -- filter=124 channel=119
    8, -5, -2, 1, -14, -7, -5, 1, 6,
    -- filter=124 channel=120
    -7, -5, -11, 0, -17, -10, 6, 4, -1,
    -- filter=124 channel=121
    3, 6, 2, -1, 11, 0, -2, -5, 1,
    -- filter=124 channel=122
    15, 13, 1, 20, 19, 13, -3, 0, -4,
    -- filter=124 channel=123
    7, -2, 0, 0, 2, 4, 3, -3, -7,
    -- filter=124 channel=124
    -2, -1, -3, 1, 0, -6, 0, -7, 3,
    -- filter=124 channel=125
    0, -3, -12, 2, -4, -2, -1, -7, 0,
    -- filter=124 channel=126
    7, 4, 9, 1, 1, -4, 0, -3, 2,
    -- filter=124 channel=127
    1, 2, -2, -9, 7, 2, 3, 5, 0,
    -- filter=125 channel=0
    -4, 4, -4, 7, -2, -1, 0, -1, 1,
    -- filter=125 channel=1
    4, -3, 3, 1, -4, 5, -1, 0, -7,
    -- filter=125 channel=2
    -6, 0, -7, -5, 7, -3, -4, 3, 4,
    -- filter=125 channel=3
    -5, 5, 5, 0, -6, -5, -4, 0, -3,
    -- filter=125 channel=4
    2, 4, 1, 0, -4, 0, 0, 0, -4,
    -- filter=125 channel=5
    5, 0, 0, 7, 0, 8, -1, 5, 0,
    -- filter=125 channel=6
    -7, -1, 6, -5, 6, -6, -6, -5, 1,
    -- filter=125 channel=7
    6, 0, 5, -1, -2, -4, -4, -4, 6,
    -- filter=125 channel=8
    -2, 5, -1, 6, 3, -2, 0, 2, 4,
    -- filter=125 channel=9
    1, -1, 4, -2, -2, -2, -1, 4, 5,
    -- filter=125 channel=10
    -4, 0, 4, -6, 0, 0, -1, 0, -4,
    -- filter=125 channel=11
    0, 4, 0, 2, 4, -3, -4, 4, 0,
    -- filter=125 channel=12
    3, -3, -3, -3, 0, 3, -7, 0, 4,
    -- filter=125 channel=13
    2, -3, 5, 0, 0, -5, 3, 0, 1,
    -- filter=125 channel=14
    3, 5, 0, 3, 5, 4, -7, -5, 6,
    -- filter=125 channel=15
    4, -5, 3, -4, 0, 2, -3, 7, -2,
    -- filter=125 channel=16
    -4, -3, 1, 3, 2, 5, 6, -2, -7,
    -- filter=125 channel=17
    -4, -5, 1, 0, 1, 4, -1, 7, -4,
    -- filter=125 channel=18
    3, 0, 3, -1, 8, 1, -2, 2, -3,
    -- filter=125 channel=19
    -1, 1, -6, -3, 6, -7, 1, -6, -4,
    -- filter=125 channel=20
    -3, 6, 2, -3, 1, 0, -6, 6, 0,
    -- filter=125 channel=21
    -5, 0, 3, -6, 3, 5, 3, -8, 1,
    -- filter=125 channel=22
    -7, -3, 7, 5, -6, -3, -4, 7, -2,
    -- filter=125 channel=23
    0, -4, 6, -6, -7, 2, -3, 0, -6,
    -- filter=125 channel=24
    -5, 7, -6, -3, -4, -2, -4, 3, 6,
    -- filter=125 channel=25
    -6, 1, -2, 0, -3, -5, 3, 0, -8,
    -- filter=125 channel=26
    4, -3, -5, 3, 6, -5, 4, 5, -5,
    -- filter=125 channel=27
    -5, -1, 8, 4, -5, 6, 7, -6, 0,
    -- filter=125 channel=28
    -3, 4, -6, 2, 6, -6, 0, -5, -6,
    -- filter=125 channel=29
    5, 7, 1, -7, -4, 1, 6, -4, 6,
    -- filter=125 channel=30
    -5, -3, 0, 7, -6, 5, 0, 0, 3,
    -- filter=125 channel=31
    2, 7, 4, 7, -9, 4, 7, -3, -6,
    -- filter=125 channel=32
    1, -3, 2, 6, 4, 0, -1, 1, 0,
    -- filter=125 channel=33
    -5, 7, 8, 0, -3, 5, -2, 3, -7,
    -- filter=125 channel=34
    1, -1, 6, -4, -3, 3, -1, 0, 0,
    -- filter=125 channel=35
    5, 4, -2, 4, -3, -6, 4, 6, -2,
    -- filter=125 channel=36
    3, -5, -6, -6, 2, 0, -4, -7, 6,
    -- filter=125 channel=37
    -5, -3, -2, 6, 4, -4, 0, 2, -7,
    -- filter=125 channel=38
    -2, 6, -3, 6, -4, 4, -4, 6, 2,
    -- filter=125 channel=39
    1, -6, 5, 3, 6, 0, -5, 4, 2,
    -- filter=125 channel=40
    -4, 2, 7, 2, -4, 1, 1, 7, 1,
    -- filter=125 channel=41
    -3, 2, -6, 10, 1, -4, 6, 8, -5,
    -- filter=125 channel=42
    6, -6, 3, 6, 0, 0, -2, -2, -7,
    -- filter=125 channel=43
    4, 0, -2, -1, 2, 7, -6, 5, -6,
    -- filter=125 channel=44
    1, 2, 2, 2, -5, 6, 2, -7, -6,
    -- filter=125 channel=45
    -5, 7, -6, 0, 4, -3, -2, -6, 1,
    -- filter=125 channel=46
    0, -6, 5, 0, -4, 1, -4, -5, 0,
    -- filter=125 channel=47
    -3, 2, 8, 1, -8, 5, 6, -8, 3,
    -- filter=125 channel=48
    1, 4, 3, -1, 2, 1, 1, 0, -4,
    -- filter=125 channel=49
    -2, -4, 1, 3, -4, 2, 6, 6, -1,
    -- filter=125 channel=50
    2, 7, -3, -2, 0, -3, 4, 0, -6,
    -- filter=125 channel=51
    3, -3, 3, 0, 2, -6, 3, 5, 0,
    -- filter=125 channel=52
    4, -5, 4, 4, -7, -2, 1, -6, 0,
    -- filter=125 channel=53
    1, 3, 1, 2, -2, -1, 0, -5, 1,
    -- filter=125 channel=54
    -5, 4, 6, -5, 5, 6, -2, 4, 0,
    -- filter=125 channel=55
    0, -2, 1, 2, -3, -5, -3, -3, -1,
    -- filter=125 channel=56
    5, -5, 1, 0, 0, -2, 2, -3, 5,
    -- filter=125 channel=57
    6, -2, 6, -3, -3, -3, -3, 8, -1,
    -- filter=125 channel=58
    -3, -6, 8, -2, -3, -5, 1, -6, 3,
    -- filter=125 channel=59
    -4, -4, 6, -1, -4, -5, 0, 0, 5,
    -- filter=125 channel=60
    0, 3, 6, 1, -6, -3, -5, 6, 4,
    -- filter=125 channel=61
    -2, -2, 2, 0, 6, 1, -8, -4, 7,
    -- filter=125 channel=62
    0, 3, 6, -3, 0, -3, -4, -3, 0,
    -- filter=125 channel=63
    3, 2, 1, -3, -7, -3, -1, -4, -2,
    -- filter=125 channel=64
    -2, 4, 3, 2, -2, 3, 0, 7, 2,
    -- filter=125 channel=65
    7, 4, -7, -5, 0, 0, -6, -6, 5,
    -- filter=125 channel=66
    -4, -7, 0, 7, 5, 1, -6, 6, 0,
    -- filter=125 channel=67
    6, 5, -1, -3, 1, 0, 7, -6, 5,
    -- filter=125 channel=68
    2, 0, 1, -1, -5, 5, 6, 3, 6,
    -- filter=125 channel=69
    6, 6, 3, 5, 0, 1, -2, 2, 0,
    -- filter=125 channel=70
    -3, 3, 7, 4, 0, 6, -1, 4, 6,
    -- filter=125 channel=71
    -1, 2, -4, 6, 4, 0, -4, 0, -3,
    -- filter=125 channel=72
    -7, 6, -5, -7, 4, 3, -4, -5, -4,
    -- filter=125 channel=73
    -7, -4, -5, 2, -2, 5, -3, -6, 4,
    -- filter=125 channel=74
    -5, 1, -4, 1, 6, -1, 4, 1, -3,
    -- filter=125 channel=75
    -4, -6, -4, -3, -6, 8, 3, -4, -3,
    -- filter=125 channel=76
    -7, -6, -5, 5, -1, -5, 4, 3, 6,
    -- filter=125 channel=77
    1, 3, 5, 1, -6, 0, 0, -5, -6,
    -- filter=125 channel=78
    1, 0, 4, 1, 6, -4, -1, 6, 2,
    -- filter=125 channel=79
    -2, -1, 0, 0, -1, -5, -3, 7, -7,
    -- filter=125 channel=80
    6, -1, -1, 3, 5, 2, 0, 0, -2,
    -- filter=125 channel=81
    -3, -2, 3, 6, -1, 4, -7, -4, 4,
    -- filter=125 channel=82
    4, 0, 0, 0, 6, 0, 2, 4, 3,
    -- filter=125 channel=83
    -2, 1, -2, -5, 3, 0, 5, -1, -3,
    -- filter=125 channel=84
    -6, 6, 0, 3, 0, 6, 3, 6, -5,
    -- filter=125 channel=85
    6, 6, 7, -5, 4, -4, 2, 6, -3,
    -- filter=125 channel=86
    3, -5, 3, 6, 7, -5, 7, 6, -1,
    -- filter=125 channel=87
    4, 6, -2, -2, -6, -1, 0, -6, -6,
    -- filter=125 channel=88
    0, 1, -1, 1, -8, 5, 0, 0, 0,
    -- filter=125 channel=89
    1, -4, -4, -3, -2, -3, 0, 3, -3,
    -- filter=125 channel=90
    -4, -1, 6, -6, -5, -4, -3, 1, 5,
    -- filter=125 channel=91
    -3, 3, -5, -5, -2, -5, -6, -2, 5,
    -- filter=125 channel=92
    0, 1, -5, -4, 1, -6, -1, 3, -4,
    -- filter=125 channel=93
    -5, 0, 0, -4, -5, 1, -5, 0, -4,
    -- filter=125 channel=94
    -1, -7, -2, 6, 0, 2, -4, 7, 0,
    -- filter=125 channel=95
    -1, 1, 4, 6, 5, 4, -2, -2, 0,
    -- filter=125 channel=96
    4, -5, -4, -4, 2, -1, -5, 0, -7,
    -- filter=125 channel=97
    4, 3, 6, 5, 1, 0, 7, 3, -5,
    -- filter=125 channel=98
    -1, -4, 2, 6, 2, 0, 5, -2, -6,
    -- filter=125 channel=99
    -2, 1, 6, -4, 0, 0, 5, -2, -7,
    -- filter=125 channel=100
    5, -2, -1, 2, -3, 5, 6, -3, 5,
    -- filter=125 channel=101
    0, 4, -4, -4, 6, -5, 0, -5, -2,
    -- filter=125 channel=102
    0, -3, 0, -7, 5, 0, 0, -1, -6,
    -- filter=125 channel=103
    -1, -3, 4, -5, 0, 5, 5, -8, 1,
    -- filter=125 channel=104
    3, -6, 6, -2, -6, 6, 4, 5, -3,
    -- filter=125 channel=105
    -6, 7, 7, 2, 7, 6, -4, -5, 2,
    -- filter=125 channel=106
    -1, -6, -7, -5, -6, -3, -6, -5, 3,
    -- filter=125 channel=107
    -1, -5, 0, -3, -4, -5, 6, 6, 7,
    -- filter=125 channel=108
    2, -6, -5, -2, -6, 5, -2, 1, 7,
    -- filter=125 channel=109
    1, -6, -1, 5, -5, 0, 0, -2, 6,
    -- filter=125 channel=110
    4, 3, -2, 5, 4, 5, 0, -7, 2,
    -- filter=125 channel=111
    3, 6, -4, -3, 4, 5, 1, 1, -4,
    -- filter=125 channel=112
    -4, -1, -5, 0, 5, 3, 2, 2, -1,
    -- filter=125 channel=113
    4, 4, 0, 6, 2, -1, 7, -7, 3,
    -- filter=125 channel=114
    0, -5, 0, 1, -2, 0, -3, -2, 6,
    -- filter=125 channel=115
    1, 2, 7, -5, 2, -3, 0, 1, 1,
    -- filter=125 channel=116
    -4, -3, -2, 2, 0, -8, -1, 0, -8,
    -- filter=125 channel=117
    3, -4, 0, -1, 5, -3, -5, -5, 1,
    -- filter=125 channel=118
    4, -2, -2, 3, -4, 3, -7, 4, 4,
    -- filter=125 channel=119
    -8, 4, 0, 2, -4, 2, 2, -1, 5,
    -- filter=125 channel=120
    1, 2, 0, -6, -5, -4, 8, -7, -3,
    -- filter=125 channel=121
    -3, -6, 4, -3, 5, 2, 4, 0, -7,
    -- filter=125 channel=122
    -3, -2, 0, 1, -9, -2, 9, -8, -8,
    -- filter=125 channel=123
    1, 1, 2, 4, -5, -3, 6, 0, 1,
    -- filter=125 channel=124
    -3, 6, 0, -1, -2, 0, -6, 2, 7,
    -- filter=125 channel=125
    2, 3, -3, 5, -2, 5, -1, -6, 4,
    -- filter=125 channel=126
    -5, -4, -4, 0, 2, -2, -6, -5, -6,
    -- filter=125 channel=127
    -6, 0, 4, -5, -2, 0, -2, 6, -4,
    -- filter=126 channel=0
    -6, 0, -3, 1, 2, 6, 5, -3, -3,
    -- filter=126 channel=1
    -7, -1, -4, 2, 6, -2, 0, -6, 1,
    -- filter=126 channel=2
    6, 0, 3, 3, 4, 7, -6, 0, 3,
    -- filter=126 channel=3
    5, 4, 4, -2, 1, -5, -1, 5, 6,
    -- filter=126 channel=4
    -4, -5, 5, -5, -3, -2, 5, -2, -2,
    -- filter=126 channel=5
    6, 0, 4, -1, -6, 8, 0, 5, 4,
    -- filter=126 channel=6
    -6, 2, 0, -2, 1, 1, 1, 1, -3,
    -- filter=126 channel=7
    -2, 6, 7, 5, 0, 6, 7, 1, 6,
    -- filter=126 channel=8
    -4, 2, 1, -1, 5, 0, 4, 4, -3,
    -- filter=126 channel=9
    -7, -3, 2, -7, 5, 5, 4, 6, -6,
    -- filter=126 channel=10
    -3, 0, 3, 5, -2, 3, 7, 0, 2,
    -- filter=126 channel=11
    -7, 2, -4, 5, 5, 0, 0, 2, -4,
    -- filter=126 channel=12
    6, 5, 8, 0, -4, 2, 0, 2, 1,
    -- filter=126 channel=13
    -6, 2, 6, 1, -9, -1, -3, 1, 7,
    -- filter=126 channel=14
    2, 1, 5, 7, -4, 0, -2, 2, -4,
    -- filter=126 channel=15
    3, -5, -2, -1, 4, 2, 3, -6, -4,
    -- filter=126 channel=16
    -4, 0, 0, 5, -3, 7, 1, 0, -6,
    -- filter=126 channel=17
    6, -2, 4, 7, 6, 5, 2, 7, 0,
    -- filter=126 channel=18
    -9, 3, 1, 4, 0, -7, -7, -5, -6,
    -- filter=126 channel=19
    -5, 2, 4, 7, -5, 2, -4, 4, 4,
    -- filter=126 channel=20
    -2, 6, 3, 5, 0, -7, 3, 3, 4,
    -- filter=126 channel=21
    -5, -3, 6, 0, -2, -1, -2, 1, -6,
    -- filter=126 channel=22
    0, 2, -5, -6, -4, 0, 0, 6, 5,
    -- filter=126 channel=23
    0, -2, 6, 0, -5, -3, -2, -1, 6,
    -- filter=126 channel=24
    -7, 0, -5, 0, -6, -6, -5, -2, 6,
    -- filter=126 channel=25
    -1, -7, 6, -7, -8, 3, -7, 5, -2,
    -- filter=126 channel=26
    4, -3, 0, -6, 3, -3, 2, -3, 3,
    -- filter=126 channel=27
    1, -8, 7, -6, 0, -4, -2, -1, -2,
    -- filter=126 channel=28
    2, -2, 4, -2, 0, 5, -7, -6, -7,
    -- filter=126 channel=29
    -1, 1, 2, -5, 4, 1, 3, -6, 0,
    -- filter=126 channel=30
    -7, -1, 1, 3, -4, 5, -2, -5, 0,
    -- filter=126 channel=31
    -2, 0, -5, 0, -1, 4, 1, 5, -6,
    -- filter=126 channel=32
    -8, 3, 7, 1, -1, -1, -3, 2, 6,
    -- filter=126 channel=33
    -1, -1, 4, -8, 0, -5, 3, 3, 7,
    -- filter=126 channel=34
    1, 7, 0, -6, -4, -5, 5, 7, 0,
    -- filter=126 channel=35
    6, -6, 7, 2, -6, 0, 2, 0, -5,
    -- filter=126 channel=36
    -6, 5, 1, 6, -1, -4, 3, -3, -2,
    -- filter=126 channel=37
    -1, 3, 5, 8, 2, -3, 2, -7, 2,
    -- filter=126 channel=38
    1, 0, 3, 3, -5, 3, -6, 4, -2,
    -- filter=126 channel=39
    5, 6, -4, -4, -2, -1, -3, 5, 3,
    -- filter=126 channel=40
    0, -5, -4, 2, -6, 2, 3, -4, -3,
    -- filter=126 channel=41
    2, 2, -2, 4, 0, -4, 4, 0, -7,
    -- filter=126 channel=42
    3, 0, 1, -3, -6, -3, -5, 2, -3,
    -- filter=126 channel=43
    -5, 8, 0, 0, 5, 5, 0, 0, -5,
    -- filter=126 channel=44
    6, 4, 5, 1, -4, -1, -2, 6, -5,
    -- filter=126 channel=45
    1, -4, 1, 0, -2, 7, 6, 1, 4,
    -- filter=126 channel=46
    -5, 6, 3, 6, -2, 2, 4, 0, -2,
    -- filter=126 channel=47
    -2, -2, -3, 5, 5, -3, 5, 0, 3,
    -- filter=126 channel=48
    2, 0, -3, 1, -3, -3, -5, 2, -2,
    -- filter=126 channel=49
    -3, -2, 1, 4, 4, -6, -2, -3, -3,
    -- filter=126 channel=50
    6, -7, -2, 2, -1, 1, 6, -2, 4,
    -- filter=126 channel=51
    0, 1, -1, 5, -2, -5, 0, -5, 3,
    -- filter=126 channel=52
    0, -4, -2, 6, -3, -6, -7, -3, 7,
    -- filter=126 channel=53
    -5, -7, 3, -6, 2, -6, -7, -3, -5,
    -- filter=126 channel=54
    -2, -4, 0, 0, -6, 5, 3, -4, 7,
    -- filter=126 channel=55
    -2, -7, -6, -3, -2, 0, 3, 6, -1,
    -- filter=126 channel=56
    1, -5, 3, -7, -1, 6, 0, 3, 1,
    -- filter=126 channel=57
    2, -6, -7, -4, -4, -4, 3, -1, -6,
    -- filter=126 channel=58
    5, 6, -2, -3, -1, 7, -1, -3, -1,
    -- filter=126 channel=59
    -8, -2, 5, -2, -7, 2, -6, -1, 7,
    -- filter=126 channel=60
    -5, 6, 5, 6, 1, 0, 0, 0, 2,
    -- filter=126 channel=61
    6, -1, 0, -2, 0, -4, 0, -4, 1,
    -- filter=126 channel=62
    -3, -5, -2, -5, 4, 1, -5, -2, -5,
    -- filter=126 channel=63
    -4, 1, 5, -5, 1, -4, -2, 1, -6,
    -- filter=126 channel=64
    -6, -3, 2, 4, 3, 5, -3, 2, -1,
    -- filter=126 channel=65
    1, 0, 6, 1, -3, -3, -2, -6, 6,
    -- filter=126 channel=66
    -5, 2, 5, -7, -5, 7, -5, 3, -2,
    -- filter=126 channel=67
    -4, -3, -7, 4, -3, -7, 0, -1, -3,
    -- filter=126 channel=68
    -3, 4, 0, 3, -2, 2, -5, 0, 0,
    -- filter=126 channel=69
    0, 3, 6, -4, 1, 5, 7, 2, -1,
    -- filter=126 channel=70
    -1, 7, -6, 5, 6, 3, -5, 3, 5,
    -- filter=126 channel=71
    -2, -5, 0, 1, 6, -5, -3, 5, 6,
    -- filter=126 channel=72
    5, 5, -3, 3, -8, -6, -4, -2, 2,
    -- filter=126 channel=73
    -2, -3, 4, -4, 3, -6, 5, -3, -2,
    -- filter=126 channel=74
    -5, 1, 0, -6, -1, 6, -2, 0, 5,
    -- filter=126 channel=75
    -7, 4, 7, 4, 2, -3, 3, -3, 2,
    -- filter=126 channel=76
    2, -6, 5, -6, 3, -1, 4, -4, 5,
    -- filter=126 channel=77
    -2, -5, -1, -5, 0, 2, 2, 7, -1,
    -- filter=126 channel=78
    -2, 0, -2, 0, -4, -3, -4, 5, 4,
    -- filter=126 channel=79
    -9, 2, 7, 3, -6, 0, -7, 3, -6,
    -- filter=126 channel=80
    -4, -5, 4, -6, -6, 1, -4, 5, 5,
    -- filter=126 channel=81
    5, 1, -6, -2, -2, 2, 1, -5, -4,
    -- filter=126 channel=82
    -6, 0, 3, 0, -3, 3, 7, 5, -2,
    -- filter=126 channel=83
    4, -5, 0, 3, 5, 0, 0, -1, 3,
    -- filter=126 channel=84
    3, 3, -1, 5, -4, 0, 6, 4, 0,
    -- filter=126 channel=85
    -2, 5, -1, 0, 7, 0, -2, -6, -4,
    -- filter=126 channel=86
    -6, 2, 6, -4, -3, 2, -2, 6, 6,
    -- filter=126 channel=87
    3, 8, -5, 4, -3, 6, 0, 2, -3,
    -- filter=126 channel=88
    -3, 2, -7, 3, -3, 3, -4, 2, 1,
    -- filter=126 channel=89
    -7, 0, 2, 1, -6, -2, -1, -3, 1,
    -- filter=126 channel=90
    -5, 4, 1, 6, -3, -3, 2, 0, 2,
    -- filter=126 channel=91
    2, -1, 1, 6, -6, 6, 2, -4, 3,
    -- filter=126 channel=92
    4, 3, -1, 3, 5, 4, 3, -1, 0,
    -- filter=126 channel=93
    0, 3, -2, 0, 3, -6, -6, -6, -7,
    -- filter=126 channel=94
    -6, 0, 3, -2, 0, -1, 0, -2, 1,
    -- filter=126 channel=95
    -2, -1, 6, 6, 2, -3, 2, 5, 3,
    -- filter=126 channel=96
    4, -2, 4, -3, -7, -1, 0, -5, 6,
    -- filter=126 channel=97
    0, -5, -3, -7, -7, -6, -4, 8, -2,
    -- filter=126 channel=98
    -1, 2, 5, 0, -1, -7, 2, 4, 0,
    -- filter=126 channel=99
    0, 0, -6, -5, 0, -6, 3, 5, 1,
    -- filter=126 channel=100
    -6, -4, 1, -5, -6, 3, 3, 0, -4,
    -- filter=126 channel=101
    1, 6, -2, 8, 7, 7, -6, 0, -1,
    -- filter=126 channel=102
    1, -7, -7, 3, 1, 0, -5, 6, 6,
    -- filter=126 channel=103
    -5, 0, 8, -4, -6, -3, 7, 3, -5,
    -- filter=126 channel=104
    3, 4, -7, -4, -5, 7, -7, -5, -5,
    -- filter=126 channel=105
    -3, 5, 6, 4, 0, -1, 5, 2, 0,
    -- filter=126 channel=106
    2, 7, 2, 3, 2, 0, 0, 5, -3,
    -- filter=126 channel=107
    -3, -1, 0, -6, 0, 3, 6, 0, 0,
    -- filter=126 channel=108
    4, 0, -6, -2, -6, -1, -1, -4, 0,
    -- filter=126 channel=109
    0, 4, -6, -4, -6, -3, -1, 0, 3,
    -- filter=126 channel=110
    1, 5, 4, 0, -1, 4, 4, 1, 3,
    -- filter=126 channel=111
    -5, -4, 3, 1, 0, -7, 4, 6, -4,
    -- filter=126 channel=112
    5, 7, -2, -5, -5, -2, -1, -2, 5,
    -- filter=126 channel=113
    -3, -3, 7, 0, -2, -3, 1, -2, 1,
    -- filter=126 channel=114
    -8, -4, 6, -1, 6, -1, -4, -5, -3,
    -- filter=126 channel=115
    -3, 4, -1, 2, 4, -2, -4, 0, -2,
    -- filter=126 channel=116
    -4, -2, 4, -5, -6, 3, 3, 1, -5,
    -- filter=126 channel=117
    -7, -6, -6, 5, 0, 7, -1, 5, 2,
    -- filter=126 channel=118
    -4, 0, 1, 4, 1, 6, -1, 1, -1,
    -- filter=126 channel=119
    -4, 7, -5, -1, 7, -3, -2, 0, 5,
    -- filter=126 channel=120
    -1, -3, -2, 5, 2, -1, -1, -7, 1,
    -- filter=126 channel=121
    2, 0, -3, 1, 0, 1, -2, -1, 3,
    -- filter=126 channel=122
    -6, -3, 2, -2, 0, -2, 2, 1, -5,
    -- filter=126 channel=123
    6, 0, -6, -4, -7, -5, 0, 6, -3,
    -- filter=126 channel=124
    -7, 3, -1, 3, 0, -6, -5, -3, -1,
    -- filter=126 channel=125
    -1, 0, -3, 1, 5, -2, -4, -1, 6,
    -- filter=126 channel=126
    -3, -4, 0, -5, 0, -2, -2, -2, 3,
    -- filter=126 channel=127
    2, -6, 1, -3, 0, 0, 3, 5, 2,
    -- filter=127 channel=0
    2, 3, 9, 3, -1, -1, 0, -2, -11,
    -- filter=127 channel=1
    1, 3, 2, 8, -1, 1, 0, -3, -4,
    -- filter=127 channel=2
    2, -8, 5, -2, 1, 3, 1, -3, 1,
    -- filter=127 channel=3
    7, -2, -5, 0, -6, 2, 2, 3, -3,
    -- filter=127 channel=4
    5, 8, 14, 5, 8, 7, 1, 6, 2,
    -- filter=127 channel=5
    2, 9, 5, -1, 4, -4, 5, -8, -9,
    -- filter=127 channel=6
    0, -4, 7, -1, -2, 3, -7, -1, 0,
    -- filter=127 channel=7
    5, -7, 3, -5, 4, 6, 0, -2, -2,
    -- filter=127 channel=8
    0, 3, 3, -5, 6, 2, 2, 0, 9,
    -- filter=127 channel=9
    2, -7, -7, 5, 0, 5, -1, 0, 3,
    -- filter=127 channel=10
    -12, -13, -16, -10, 0, -5, 11, 4, -1,
    -- filter=127 channel=11
    2, -3, -2, -4, 0, 9, 6, 6, 11,
    -- filter=127 channel=12
    3, -11, 0, 5, 0, 1, 2, -9, -3,
    -- filter=127 channel=13
    5, -14, -11, -9, -13, -6, 2, 1, 0,
    -- filter=127 channel=14
    5, -7, 0, 0, 2, 1, 2, 1, 6,
    -- filter=127 channel=15
    -11, -13, 0, -17, -19, 4, 0, -2, 1,
    -- filter=127 channel=16
    7, 1, -9, 14, 12, -7, 6, 0, 2,
    -- filter=127 channel=17
    6, 0, 2, 0, 6, -1, 6, -5, 5,
    -- filter=127 channel=18
    -4, -19, -15, -11, -11, -6, -7, -1, 10,
    -- filter=127 channel=19
    -7, -4, 6, 6, 7, -2, 7, 4, -4,
    -- filter=127 channel=20
    2, -9, 7, -16, -8, 9, -2, 10, 12,
    -- filter=127 channel=21
    5, 3, -13, 14, 3, 1, 21, 4, 1,
    -- filter=127 channel=22
    2, -6, 5, -4, -11, -1, -8, 0, -1,
    -- filter=127 channel=23
    -17, -27, -5, -27, -14, 10, 0, -7, 10,
    -- filter=127 channel=24
    0, 1, 1, 2, -5, 5, 4, 6, 7,
    -- filter=127 channel=25
    1, -19, -15, 5, -1, -5, 11, -4, -4,
    -- filter=127 channel=26
    2, 11, 8, 12, 10, 0, 4, 8, -6,
    -- filter=127 channel=27
    -12, -23, -6, -7, -6, 11, 8, 3, 6,
    -- filter=127 channel=28
    7, 4, -3, -1, 2, -1, 5, -4, -1,
    -- filter=127 channel=29
    -8, -7, -1, -12, -8, -2, -4, 11, 16,
    -- filter=127 channel=30
    -7, -3, -5, -1, 1, 0, 7, -4, 2,
    -- filter=127 channel=31
    -14, -33, -14, 8, -9, -2, 18, 11, 11,
    -- filter=127 channel=32
    -5, -22, -4, -15, -11, 7, -9, -3, -1,
    -- filter=127 channel=33
    1, -21, -10, 0, -16, 1, 6, -5, -1,
    -- filter=127 channel=34
    -5, -3, 3, -5, -8, 2, -11, -3, 7,
    -- filter=127 channel=35
    -5, 0, 5, 5, 2, -3, -6, 4, 5,
    -- filter=127 channel=36
    -1, -4, -7, 1, 7, 11, 3, 16, 1,
    -- filter=127 channel=37
    7, 4, 1, 5, 7, 12, 0, -9, -5,
    -- filter=127 channel=38
    -8, -15, -4, -1, -7, -3, 9, -6, -4,
    -- filter=127 channel=39
    5, -7, -1, -5, -1, 10, 5, 3, 0,
    -- filter=127 channel=40
    0, -6, 3, -1, -9, -4, -2, -3, 6,
    -- filter=127 channel=41
    7, -8, -15, -6, 3, -18, 2, -3, -5,
    -- filter=127 channel=42
    -5, -6, -6, 0, -2, -3, 0, 0, 5,
    -- filter=127 channel=43
    2, -7, -6, 0, -11, 0, 2, 5, 6,
    -- filter=127 channel=44
    8, -6, 6, 1, -1, 5, 6, 5, -8,
    -- filter=127 channel=45
    9, 6, 7, -1, -3, 4, 8, -3, 4,
    -- filter=127 channel=46
    -2, 1, -5, 8, 5, -5, 4, -3, -5,
    -- filter=127 channel=47
    9, 1, -13, 20, 6, -10, 11, -2, -5,
    -- filter=127 channel=48
    3, -10, -8, 14, 14, 0, 15, 11, 2,
    -- filter=127 channel=49
    -8, 2, -1, -7, 5, 11, 0, 2, 13,
    -- filter=127 channel=50
    -4, -4, -6, 5, -10, 3, -1, 1, 2,
    -- filter=127 channel=51
    -3, 5, 4, 2, 0, 4, 4, 0, 6,
    -- filter=127 channel=52
    1, -1, 0, -9, -7, 10, -8, -4, 6,
    -- filter=127 channel=53
    -5, -8, 1, -6, -7, -4, 1, 0, 1,
    -- filter=127 channel=54
    -2, 2, 6, 4, 0, 3, 5, -2, -3,
    -- filter=127 channel=55
    -17, -24, -9, -10, -12, 0, 2, 7, 12,
    -- filter=127 channel=56
    2, -5, -1, 0, -7, 7, -7, -3, 4,
    -- filter=127 channel=57
    -7, 6, 2, 1, -6, 5, -5, 1, 1,
    -- filter=127 channel=58
    4, 3, 1, 0, 10, -5, 0, -1, -2,
    -- filter=127 channel=59
    -2, -21, -6, 5, 1, -4, 15, 3, -3,
    -- filter=127 channel=60
    8, 1, 3, -4, 3, 0, -4, -2, -4,
    -- filter=127 channel=61
    -5, 0, 0, -7, 5, -5, -5, 1, 4,
    -- filter=127 channel=62
    0, -4, 6, -5, 0, 6, 4, 0, 6,
    -- filter=127 channel=63
    -1, 0, 5, 7, 1, -4, 6, -6, -8,
    -- filter=127 channel=64
    -8, -4, -5, 5, 1, 0, 8, 11, 0,
    -- filter=127 channel=65
    0, 3, 2, -1, 0, -1, 4, 2, 4,
    -- filter=127 channel=66
    1, -1, 2, 3, -12, -7, -3, -8, -3,
    -- filter=127 channel=67
    0, -3, 1, 1, -1, -1, 5, 4, -5,
    -- filter=127 channel=68
    3, -3, 2, 1, -3, 8, 2, 9, 0,
    -- filter=127 channel=69
    8, -4, -4, 1, -2, 3, 4, -2, -2,
    -- filter=127 channel=70
    -12, -14, 0, -17, -8, 13, 0, -8, 7,
    -- filter=127 channel=71
    1, -7, -1, 1, 9, 1, 5, 1, 4,
    -- filter=127 channel=72
    -2, -26, -7, -2, -11, -2, 20, 4, 6,
    -- filter=127 channel=73
    -2, -15, -1, -8, -3, 2, -3, 11, 5,
    -- filter=127 channel=74
    -14, -6, 8, 2, 1, 13, 4, 4, -1,
    -- filter=127 channel=75
    9, -5, -11, -5, -9, -12, -1, -13, -19,
    -- filter=127 channel=76
    4, 1, 3, -1, -5, 6, 5, 2, 10,
    -- filter=127 channel=77
    0, 7, -4, -3, 6, -7, 0, -5, 4,
    -- filter=127 channel=78
    -8, -6, 1, -6, 6, -1, 5, 0, 0,
    -- filter=127 channel=79
    -10, -20, -17, -11, -13, 3, -6, 0, 0,
    -- filter=127 channel=80
    1, -17, -24, 17, 2, 0, 19, 7, 6,
    -- filter=127 channel=81
    -6, -2, -6, 3, -3, -3, 3, 1, 4,
    -- filter=127 channel=82
    -2, 5, 0, 6, 3, 2, 0, -5, -2,
    -- filter=127 channel=83
    -6, -5, 1, 0, 9, -2, 10, 4, -1,
    -- filter=127 channel=84
    -9, -5, -7, -12, -4, 0, 2, 9, 3,
    -- filter=127 channel=85
    7, 4, 4, 5, -7, -6, 0, 0, 0,
    -- filter=127 channel=86
    -3, 3, -1, -5, -1, 7, -5, -1, -9,
    -- filter=127 channel=87
    1, -5, 0, -14, -11, 9, -1, -2, 7,
    -- filter=127 channel=88
    -3, -5, 2, 10, 10, 0, 8, 4, 11,
    -- filter=127 channel=89
    -4, -14, -13, -2, -8, -3, -1, 9, 13,
    -- filter=127 channel=90
    0, 1, 4, -5, 8, 2, 0, 0, 2,
    -- filter=127 channel=91
    0, -13, -4, -8, 0, 17, -1, 1, 13,
    -- filter=127 channel=92
    0, 1, -4, 1, 2, 5, 1, 4, 0,
    -- filter=127 channel=93
    8, -2, -6, 15, 6, 5, 10, 9, 0,
    -- filter=127 channel=94
    5, 1, 3, 7, 5, -4, 4, 0, -4,
    -- filter=127 channel=95
    3, 3, 4, -6, 2, 6, 7, 6, 5,
    -- filter=127 channel=96
    8, -2, -2, 1, 6, 1, 2, -2, 1,
    -- filter=127 channel=97
    8, -2, 4, 0, 7, -5, 5, -2, -2,
    -- filter=127 channel=98
    -1, -19, -13, 6, -4, 0, 8, 4, -3,
    -- filter=127 channel=99
    -10, -30, -7, -1, -10, 0, 16, 7, 7,
    -- filter=127 channel=100
    -6, 4, 2, 0, -8, 5, 1, 1, -6,
    -- filter=127 channel=101
    -5, 7, 0, 3, 11, 12, -2, 7, 0,
    -- filter=127 channel=102
    -6, 0, 2, -4, 3, 0, -3, -3, 5,
    -- filter=127 channel=103
    11, -10, -2, 12, 9, -3, 15, -1, 0,
    -- filter=127 channel=104
    -3, -13, -12, 4, 4, -4, 12, 13, 3,
    -- filter=127 channel=105
    1, 5, -4, 0, -1, -1, -2, 1, 2,
    -- filter=127 channel=106
    2, 0, -4, -3, 6, -2, 1, 8, 0,
    -- filter=127 channel=107
    -7, -8, 3, -6, -11, 4, 3, -5, 5,
    -- filter=127 channel=108
    0, 3, -1, -5, -2, -1, 0, 0, -9,
    -- filter=127 channel=109
    -3, -19, -14, -4, -9, 8, 9, 7, 5,
    -- filter=127 channel=110
    -3, -5, -6, -8, -5, 3, 3, 3, 0,
    -- filter=127 channel=111
    7, 1, -6, -5, -3, -2, 1, -3, -7,
    -- filter=127 channel=112
    -4, -11, 2, -10, -10, 10, 5, 0, 6,
    -- filter=127 channel=113
    0, -18, -8, 0, -6, -2, -3, 0, 9,
    -- filter=127 channel=114
    -1, -10, 4, -14, -7, 11, -5, -1, 7,
    -- filter=127 channel=115
    1, 1, 3, -4, 7, 0, -7, -1, -1,
    -- filter=127 channel=116
    -8, -14, -19, 2, -5, -2, 14, 14, 6,
    -- filter=127 channel=117
    3, 1, -1, -1, -5, 2, 1, 6, 0,
    -- filter=127 channel=118
    6, 0, -6, 0, 7, 3, 4, -5, -1,
    -- filter=127 channel=119
    -3, -7, 12, -4, 1, -4, -2, -7, 8,
    -- filter=127 channel=120
    -21, -19, 5, -11, -3, 17, 9, 14, 18,
    -- filter=127 channel=121
    -1, -15, -5, -7, -3, -10, 8, -7, 0,
    -- filter=127 channel=122
    13, -7, -11, 29, 24, 0, 26, 17, -10,
    -- filter=127 channel=123
    1, 1, -3, 1, -9, -3, 0, 3, -1,
    -- filter=127 channel=124
    0, -6, -5, -8, -3, 4, -2, 5, 0,
    -- filter=127 channel=125
    -1, -16, -11, 6, -10, 9, 16, 14, 0,
    -- filter=127 channel=126
    4, -4, -7, -7, -8, -7, -1, -1, 4,
    -- filter=127 channel=127
    5, 1, -7, -4, 6, 0, -3, 0, 0,
    -- filter=128 channel=0
    -3, 0, -1, 2, 0, -6, 0, 3, -2,
    -- filter=128 channel=1
    5, 3, -2, -2, 4, 2, 0, 6, -1,
    -- filter=128 channel=2
    -6, 1, 0, 1, -2, -2, 2, 5, 7,
    -- filter=128 channel=3
    -5, -9, -7, -4, 7, 4, 1, -1, -5,
    -- filter=128 channel=4
    -4, -7, -3, 3, 5, 1, 2, 6, -3,
    -- filter=128 channel=5
    -2, -4, -2, -4, -9, 6, 8, -9, -1,
    -- filter=128 channel=6
    3, -1, -3, -1, 3, 0, -5, 3, 5,
    -- filter=128 channel=7
    -2, -6, -1, -2, 5, -3, 0, 2, 4,
    -- filter=128 channel=8
    -1, -2, -4, 6, -3, -4, 3, 4, 0,
    -- filter=128 channel=9
    -1, 0, 2, 0, -8, -1, -4, -5, -1,
    -- filter=128 channel=10
    4, -6, -1, 2, 4, 1, -5, 0, 1,
    -- filter=128 channel=11
    -2, -5, -3, -3, -4, -5, 5, 3, 1,
    -- filter=128 channel=12
    0, 3, 2, -5, 6, -1, 0, 6, 3,
    -- filter=128 channel=13
    1, -1, -6, 8, 7, -4, 1, 0, -8,
    -- filter=128 channel=14
    -2, -2, -3, -6, -7, 0, -6, -1, 2,
    -- filter=128 channel=15
    -6, -7, 0, -5, 0, 1, 0, 6, 4,
    -- filter=128 channel=16
    4, -8, 4, 6, -7, -4, 8, -8, 6,
    -- filter=128 channel=17
    -2, 0, 2, -5, 1, 6, -5, 0, -6,
    -- filter=128 channel=18
    2, -7, 2, 5, 3, 0, -7, 2, -7,
    -- filter=128 channel=19
    0, 5, 6, -5, -5, 4, -7, -7, -6,
    -- filter=128 channel=20
    2, -5, -4, -2, 4, 2, -5, -5, 4,
    -- filter=128 channel=21
    -3, 7, 8, -2, 6, 3, 8, 5, -2,
    -- filter=128 channel=22
    3, 0, -1, 5, 1, 1, 5, 2, 4,
    -- filter=128 channel=23
    -5, -8, -1, 2, -12, -10, 6, 3, 5,
    -- filter=128 channel=24
    5, -2, 7, -4, 4, 4, -3, 3, -6,
    -- filter=128 channel=25
    5, -4, -7, 8, -3, 0, 9, 2, -3,
    -- filter=128 channel=26
    5, 2, -3, -3, 2, 8, -6, 4, 2,
    -- filter=128 channel=27
    2, -10, -7, -2, -8, -6, 10, -7, 5,
    -- filter=128 channel=28
    0, 0, 6, -2, -4, 7, -5, 0, 0,
    -- filter=128 channel=29
    0, -2, 0, 5, 2, 1, -8, -3, 4,
    -- filter=128 channel=30
    -7, -7, 0, 6, 0, 0, 0, -2, -2,
    -- filter=128 channel=31
    -3, -4, 4, -1, -1, 4, 8, -10, 5,
    -- filter=128 channel=32
    -3, -4, 1, 1, 2, -5, 8, 6, -2,
    -- filter=128 channel=33
    2, -7, -9, -2, -3, -3, -5, 4, -8,
    -- filter=128 channel=34
    -6, 1, 1, 0, -6, 2, -7, 1, 1,
    -- filter=128 channel=35
    2, 1, -4, -1, -3, -5, 3, -3, -4,
    -- filter=128 channel=36
    9, 5, 4, 5, -4, 3, -1, 5, 3,
    -- filter=128 channel=37
    -1, -10, -8, 9, -5, -2, 0, -8, 7,
    -- filter=128 channel=38
    -7, -3, 0, 2, 0, 0, -1, -6, -3,
    -- filter=128 channel=39
    6, -4, 0, -5, 6, -4, -4, 4, -3,
    -- filter=128 channel=40
    0, 5, -6, 3, 4, 3, -5, -5, -2,
    -- filter=128 channel=41
    9, 15, 1, 6, 10, -1, 2, 15, 3,
    -- filter=128 channel=42
    2, 0, -2, -5, 1, -3, 0, 2, 6,
    -- filter=128 channel=43
    -7, 5, -5, -4, 0, -4, 0, 2, 1,
    -- filter=128 channel=44
    5, -10, -6, 9, -3, -6, 9, -9, -5,
    -- filter=128 channel=45
    3, -1, -2, 3, 2, 0, 6, -2, -3,
    -- filter=128 channel=46
    -1, -5, 1, 0, -5, 6, 0, 5, -2,
    -- filter=128 channel=47
    2, -5, -1, 9, -10, -7, -2, -5, -6,
    -- filter=128 channel=48
    10, 6, 0, 9, -4, -7, 1, -5, 3,
    -- filter=128 channel=49
    -4, -5, -7, -4, -7, -5, -3, -4, 1,
    -- filter=128 channel=50
    2, -8, -8, 2, -5, 0, 0, 1, 4,
    -- filter=128 channel=51
    6, -1, 1, -2, -6, 2, 7, -1, -1,
    -- filter=128 channel=52
    1, -3, -6, 4, -7, -2, -5, 0, -6,
    -- filter=128 channel=53
    0, -7, 3, -5, -3, 3, 5, -1, -6,
    -- filter=128 channel=54
    2, -1, -1, 0, 4, -7, -3, -3, -5,
    -- filter=128 channel=55
    8, -6, -10, -1, -5, -5, -5, 0, 0,
    -- filter=128 channel=56
    1, -6, -3, 3, -1, 0, -5, 6, -1,
    -- filter=128 channel=57
    5, 0, -2, 0, 7, 6, 0, 0, 1,
    -- filter=128 channel=58
    -6, -8, 0, -4, -9, -5, 7, 3, -2,
    -- filter=128 channel=59
    -4, 5, -6, -4, 0, -3, 0, 8, 1,
    -- filter=128 channel=60
    -6, 0, -1, 7, 3, -5, 4, -6, 7,
    -- filter=128 channel=61
    1, -2, 5, 4, -1, 7, -7, 4, 3,
    -- filter=128 channel=62
    -4, 0, -5, 7, -6, 1, 7, -5, 3,
    -- filter=128 channel=63
    -7, -8, 6, -8, -1, 1, 0, 3, 3,
    -- filter=128 channel=64
    -4, 2, 0, -2, 0, 1, 2, -3, -1,
    -- filter=128 channel=65
    7, 0, -6, -1, 2, 0, -7, -1, -3,
    -- filter=128 channel=66
    3, 4, 6, 4, 3, -1, -6, 5, 6,
    -- filter=128 channel=67
    -6, 3, -3, 0, 5, 0, 0, 3, 0,
    -- filter=128 channel=68
    -3, -4, -6, -6, -1, 3, -3, 2, 3,
    -- filter=128 channel=69
    2, -4, -4, 5, 0, 4, -6, -4, 0,
    -- filter=128 channel=70
    0, -3, -2, 0, -3, -3, 8, -1, 3,
    -- filter=128 channel=71
    1, 7, -2, -6, 6, -4, 0, 4, -5,
    -- filter=128 channel=72
    10, -3, -3, 7, -4, 3, 0, 4, -6,
    -- filter=128 channel=73
    8, -2, -4, -3, 2, -4, 1, 7, -5,
    -- filter=128 channel=74
    -6, -9, -3, 3, -5, 0, -2, 4, -4,
    -- filter=128 channel=75
    3, -2, -5, -4, 0, 0, 2, -8, 0,
    -- filter=128 channel=76
    4, -5, -2, -3, 0, -1, 4, -3, -3,
    -- filter=128 channel=77
    4, -3, -2, 6, 4, 1, -1, 3, -3,
    -- filter=128 channel=78
    -8, 4, -7, 0, -7, -7, 3, 6, 1,
    -- filter=128 channel=79
    2, -10, -5, 2, 0, -5, 3, 2, 2,
    -- filter=128 channel=80
    3, 6, 1, 11, 5, -7, -1, 2, 0,
    -- filter=128 channel=81
    6, 4, -6, -6, 4, 6, -4, -5, -6,
    -- filter=128 channel=82
    1, -5, -5, 4, 0, 0, 0, -5, 0,
    -- filter=128 channel=83
    0, 0, -3, -4, -3, -7, -4, -3, -2,
    -- filter=128 channel=84
    -6, -3, -7, 5, 4, -5, 5, -2, 5,
    -- filter=128 channel=85
    -1, -2, 6, -4, 0, 0, -4, 4, -7,
    -- filter=128 channel=86
    5, -5, -4, 7, -8, -7, -4, 0, 3,
    -- filter=128 channel=87
    -4, 5, 0, 1, -2, 4, -7, -3, 5,
    -- filter=128 channel=88
    -4, 0, -4, -5, 0, 9, 0, -7, -4,
    -- filter=128 channel=89
    0, 7, -5, -3, 3, 3, -3, 3, 3,
    -- filter=128 channel=90
    3, 7, 6, 3, 6, 0, 1, -7, -4,
    -- filter=128 channel=91
    -1, 4, 1, -1, -8, -5, 3, 5, -5,
    -- filter=128 channel=92
    0, -3, -7, -2, -2, 0, 3, -7, -5,
    -- filter=128 channel=93
    6, -1, 3, 8, 0, 0, 8, 2, 8,
    -- filter=128 channel=94
    2, 0, 2, 0, -3, 7, -2, -5, 6,
    -- filter=128 channel=95
    -4, 0, 6, -2, -2, -3, -2, -4, 2,
    -- filter=128 channel=96
    0, -6, 1, 3, -2, -4, 6, 6, 3,
    -- filter=128 channel=97
    5, 0, 3, -7, -3, -4, 7, 0, 4,
    -- filter=128 channel=98
    1, 0, 0, 8, -2, -2, -2, -7, 4,
    -- filter=128 channel=99
    1, -6, -1, 8, -7, -9, 6, 0, 7,
    -- filter=128 channel=100
    -7, -4, 1, 5, -3, -2, -5, -1, 1,
    -- filter=128 channel=101
    -2, -4, 4, 1, 5, 2, 1, -3, -1,
    -- filter=128 channel=102
    -6, 4, -6, 2, 0, 0, -3, -7, 0,
    -- filter=128 channel=103
    -6, 0, -5, 1, -8, 4, 2, 3, -5,
    -- filter=128 channel=104
    1, -5, 7, 9, 4, -1, 2, 0, -6,
    -- filter=128 channel=105
    5, -1, -4, 5, -7, 3, 2, -4, -6,
    -- filter=128 channel=106
    8, 7, 1, 4, 10, 0, -7, -4, 6,
    -- filter=128 channel=107
    0, 3, -7, -7, 1, -4, -7, 6, -5,
    -- filter=128 channel=108
    -6, -3, 2, 1, 8, 0, -7, -2, 4,
    -- filter=128 channel=109
    0, -4, -8, 1, -3, -9, 0, 3, -5,
    -- filter=128 channel=110
    -2, 1, 2, 0, -4, -7, 5, -3, 0,
    -- filter=128 channel=111
    -6, 8, 7, -3, 1, -4, -1, -1, 0,
    -- filter=128 channel=112
    0, -9, -4, -4, 3, -5, 8, -7, -6,
    -- filter=128 channel=113
    4, -5, -6, 0, 1, 2, -1, -7, 1,
    -- filter=128 channel=114
    -7, 0, -10, 1, -10, -11, 5, -4, 6,
    -- filter=128 channel=115
    2, -7, -4, 6, 2, 5, 4, 3, 0,
    -- filter=128 channel=116
    0, 1, -4, -3, -6, -9, 1, 3, 7,
    -- filter=128 channel=117
    0, 7, -2, -5, 8, -7, -1, 0, 6,
    -- filter=128 channel=118
    -6, -2, -6, 3, 1, 3, -5, 4, 0,
    -- filter=128 channel=119
    0, 3, 2, 3, -5, 5, -1, 0, -2,
    -- filter=128 channel=120
    7, -11, -2, 1, -2, 1, 7, -3, 6,
    -- filter=128 channel=121
    -3, -2, -5, 6, 9, 0, 2, 3, -7,
    -- filter=128 channel=122
    6, -3, 7, 3, -5, 4, 0, -9, -1,
    -- filter=128 channel=123
    -6, -7, -4, -2, 0, 3, 3, 5, -4,
    -- filter=128 channel=124
    -1, -2, 5, 6, 3, 5, -7, -7, 7,
    -- filter=128 channel=125
    7, -5, -5, 4, -9, 6, 2, 6, 7,
    -- filter=128 channel=126
    -6, -6, -3, 0, 4, -1, 0, -4, -7,
    -- filter=128 channel=127
    4, 6, 2, -4, -3, -6, 0, 9, 1,
    -- filter=129 channel=0
    -6, -4, -4, 4, 10, 6, -18, -7, -5,
    -- filter=129 channel=1
    14, -3, -15, 9, 14, -2, 0, -12, 0,
    -- filter=129 channel=2
    9, 5, -1, -2, 4, 2, 6, 1, 2,
    -- filter=129 channel=3
    5, 12, 11, 42, 42, 15, -10, 4, 6,
    -- filter=129 channel=4
    12, 15, 4, 17, 28, 19, 28, 25, 1,
    -- filter=129 channel=5
    -12, 1, 8, 6, 0, -5, -10, 0, 3,
    -- filter=129 channel=6
    2, -7, 5, 10, 3, 3, -4, -8, 3,
    -- filter=129 channel=7
    -5, -3, 1, 3, 3, -7, -5, 0, -1,
    -- filter=129 channel=8
    9, 10, -3, -6, -3, -1, 4, -2, -5,
    -- filter=129 channel=9
    -9, -7, 1, 15, 5, 0, -13, 2, 5,
    -- filter=129 channel=10
    -7, -12, -10, 10, 20, 3, -5, -4, -3,
    -- filter=129 channel=11
    1, -2, 1, 8, 2, 0, -6, -5, -1,
    -- filter=129 channel=12
    -7, 0, -3, -8, 5, -11, -4, 0, -10,
    -- filter=129 channel=13
    -8, -23, -14, 18, 32, 7, -10, -5, -8,
    -- filter=129 channel=14
    -2, -7, -2, 0, 0, 5, 5, 5, 6,
    -- filter=129 channel=15
    -9, -11, -5, 22, 34, 7, -6, -10, 0,
    -- filter=129 channel=16
    0, -6, -8, 6, 13, -11, -2, -4, -5,
    -- filter=129 channel=17
    -5, -6, 0, 3, -7, 6, 0, -6, 5,
    -- filter=129 channel=18
    -5, -17, -16, 17, 25, 10, -28, -19, 1,
    -- filter=129 channel=19
    3, -6, -7, 1, 1, 6, 0, 4, -3,
    -- filter=129 channel=20
    -3, -4, 8, 14, 20, 7, -11, 0, 0,
    -- filter=129 channel=21
    -5, -4, -3, 7, 10, 1, -5, 5, 6,
    -- filter=129 channel=22
    -8, -4, 0, 10, 0, -3, -8, 1, 0,
    -- filter=129 channel=23
    -19, -20, -10, 50, 45, 3, -31, -18, -2,
    -- filter=129 channel=24
    -5, 4, -4, 0, -7, -4, -3, 5, 1,
    -- filter=129 channel=25
    -5, -29, -6, 25, 33, 1, -14, -23, -4,
    -- filter=129 channel=26
    8, -3, -7, -9, -1, -8, 7, -8, -7,
    -- filter=129 channel=27
    -18, -37, -18, 50, 48, 17, -33, -23, -1,
    -- filter=129 channel=28
    5, 6, -2, -2, 5, 2, 7, 2, 3,
    -- filter=129 channel=29
    -4, -1, -2, 14, 5, 5, -4, -14, 2,
    -- filter=129 channel=30
    -12, -22, -8, 26, 33, 15, -14, -10, -7,
    -- filter=129 channel=31
    -29, -30, -16, 33, 26, 0, -6, -5, 5,
    -- filter=129 channel=32
    -6, -18, -9, 39, 33, 17, -26, -23, -3,
    -- filter=129 channel=33
    -17, -14, -9, 33, 37, 9, -18, -12, 2,
    -- filter=129 channel=34
    -6, -1, -4, 4, -14, -15, -8, -5, -6,
    -- filter=129 channel=35
    -2, 4, 0, -1, 6, 5, -5, -4, 5,
    -- filter=129 channel=36
    -5, 0, -6, -2, -6, 1, 15, 0, -9,
    -- filter=129 channel=37
    10, 6, 5, 4, 2, -6, -1, -9, -3,
    -- filter=129 channel=38
    -8, -7, -9, 15, 21, 0, -11, -11, 1,
    -- filter=129 channel=39
    2, 0, -4, 0, 13, 6, -9, -3, 0,
    -- filter=129 channel=40
    -11, -3, 2, 0, 8, 0, 0, -9, -4,
    -- filter=129 channel=41
    15, 3, -15, -21, 0, 6, 12, -14, -14,
    -- filter=129 channel=42
    0, -1, 0, 7, 15, 1, -6, -5, 5,
    -- filter=129 channel=43
    -2, 7, 9, 15, 21, 2, -1, -8, -4,
    -- filter=129 channel=44
    -8, 4, 7, 9, 12, 0, -5, -4, 5,
    -- filter=129 channel=45
    -5, 4, -3, 7, 0, -6, -9, 6, 0,
    -- filter=129 channel=46
    1, 6, 6, 3, -2, -1, 1, -4, 1,
    -- filter=129 channel=47
    -8, -7, -7, 13, 24, 1, -7, -2, 0,
    -- filter=129 channel=48
    -5, -9, -5, 18, 18, 10, -8, 0, -11,
    -- filter=129 channel=49
    5, -6, -8, 9, 16, 15, 10, -8, 3,
    -- filter=129 channel=50
    -10, -17, -10, 18, 16, -1, -2, -12, 6,
    -- filter=129 channel=51
    0, 6, 0, -5, 2, -3, 2, -1, 3,
    -- filter=129 channel=52
    7, 5, 3, 6, -5, -3, 3, 7, 4,
    -- filter=129 channel=53
    4, -8, 4, 0, 8, 0, -6, -1, -1,
    -- filter=129 channel=54
    -3, 4, 7, -7, 6, 0, -1, -6, 0,
    -- filter=129 channel=55
    -7, -8, -7, 25, 19, 3, -17, -12, -5,
    -- filter=129 channel=56
    0, 1, -7, -1, -7, -8, -3, -5, -4,
    -- filter=129 channel=57
    8, 10, 2, 6, 7, 4, 0, 2, 1,
    -- filter=129 channel=58
    3, 1, 1, -7, 1, -1, -9, -12, -3,
    -- filter=129 channel=59
    -7, -19, -13, 18, 17, 5, -1, -13, -7,
    -- filter=129 channel=60
    1, -5, 3, 4, -2, 1, 0, 3, 1,
    -- filter=129 channel=61
    3, -1, -5, -9, 0, -5, 4, -4, 3,
    -- filter=129 channel=62
    8, -4, -3, -2, 0, 1, -3, 3, -5,
    -- filter=129 channel=63
    5, -2, -2, -11, -11, -4, -1, -4, -7,
    -- filter=129 channel=64
    -6, -1, -4, 1, 2, 10, 1, -4, 1,
    -- filter=129 channel=65
    -3, -3, -1, -4, 7, 1, 5, 1, -5,
    -- filter=129 channel=66
    9, -3, -4, -11, -4, 0, 5, -8, -3,
    -- filter=129 channel=67
    -1, 1, 6, 6, -1, 0, 8, -6, 6,
    -- filter=129 channel=68
    -2, 3, -7, 0, 1, 7, 11, 1, -2,
    -- filter=129 channel=69
    6, -5, -3, -9, -6, 5, -7, -8, -5,
    -- filter=129 channel=70
    -1, -6, 2, 26, 21, 11, -2, -4, 7,
    -- filter=129 channel=71
    -6, 11, 3, 15, 15, 0, -3, 8, 0,
    -- filter=129 channel=72
    -12, -24, -11, 17, 20, -5, -8, -10, -3,
    -- filter=129 channel=73
    1, 0, -1, 18, 7, 3, 2, 1, 3,
    -- filter=129 channel=74
    -5, -10, 1, 0, -4, 0, -4, -2, 4,
    -- filter=129 channel=75
    -4, -16, -2, 21, 22, 11, -21, -13, -6,
    -- filter=129 channel=76
    1, -8, 0, 7, 7, 9, -12, -2, 3,
    -- filter=129 channel=77
    4, 4, -6, 6, -1, -1, 3, 5, -9,
    -- filter=129 channel=78
    -9, 3, 0, -1, 5, -6, 4, 3, -6,
    -- filter=129 channel=79
    -17, -33, -17, 40, 54, 21, -31, -28, -10,
    -- filter=129 channel=80
    -8, -27, -16, 26, 23, 8, -10, -16, -8,
    -- filter=129 channel=81
    -1, -5, 4, -6, 5, 2, -2, 0, -5,
    -- filter=129 channel=82
    -6, -5, 7, 2, 1, 0, -3, 7, 0,
    -- filter=129 channel=83
    10, -2, 0, 0, 0, -1, 1, 7, -5,
    -- filter=129 channel=84
    7, -2, -12, 9, 17, 3, 4, -7, -8,
    -- filter=129 channel=85
    -7, -4, -6, 6, 7, 6, 5, -4, -2,
    -- filter=129 channel=86
    -2, 3, 5, -5, 2, -9, -2, 4, -5,
    -- filter=129 channel=87
    0, -2, 2, 10, 9, 1, 2, 1, 2,
    -- filter=129 channel=88
    -9, -8, -6, -1, -9, -7, 0, -5, 1,
    -- filter=129 channel=89
    -12, -24, -4, 37, 39, 2, -26, -21, 0,
    -- filter=129 channel=90
    -3, 6, 8, 10, -7, -14, 4, 10, -3,
    -- filter=129 channel=91
    0, -20, -9, 13, 18, 6, -4, -15, 1,
    -- filter=129 channel=92
    2, 0, 5, 9, -1, 1, 5, 11, 0,
    -- filter=129 channel=93
    2, -3, -1, 13, 19, 12, -11, 0, -2,
    -- filter=129 channel=94
    -4, -1, 2, 1, -1, 3, 1, -2, -7,
    -- filter=129 channel=95
    -3, 6, 4, 8, 4, -1, -4, -3, -2,
    -- filter=129 channel=96
    0, 4, -3, 5, -1, -4, 1, 6, -2,
    -- filter=129 channel=97
    -2, 11, 10, 11, 9, 0, 0, 9, 12,
    -- filter=129 channel=98
    -15, -25, -6, 43, 36, 9, -32, -11, -7,
    -- filter=129 channel=99
    -19, -24, -16, 13, 11, -5, -10, -2, 3,
    -- filter=129 channel=100
    9, 0, 7, 0, -9, 8, -5, 0, 7,
    -- filter=129 channel=101
    17, 16, 0, 12, 22, 11, 23, 18, 4,
    -- filter=129 channel=102
    -1, -2, 2, -4, 6, -1, -7, 2, 1,
    -- filter=129 channel=103
    -4, 0, 3, 9, 18, -3, -2, 2, 3,
    -- filter=129 channel=104
    -6, -17, -6, 3, 11, 6, -2, -6, 4,
    -- filter=129 channel=105
    1, 1, 8, 0, 2, 12, -6, 1, -5,
    -- filter=129 channel=106
    -2, -1, 3, 7, -1, 5, -4, 7, 0,
    -- filter=129 channel=107
    -1, -7, 2, 7, 5, 0, -11, 0, -2,
    -- filter=129 channel=108
    7, 5, 4, -10, 1, 7, -1, -8, 4,
    -- filter=129 channel=109
    -6, -29, -15, 22, 32, 13, -17, -24, -7,
    -- filter=129 channel=110
    -13, -7, 2, 12, 5, -4, -2, -8, 3,
    -- filter=129 channel=111
    -1, 3, 2, -5, -2, -2, 3, -5, -10,
    -- filter=129 channel=112
    -10, -13, 0, 19, 3, -2, -4, -6, 0,
    -- filter=129 channel=113
    -14, -3, -2, 27, 18, 7, -8, -4, 9,
    -- filter=129 channel=114
    2, -32, -19, 18, 34, 20, -21, -22, -2,
    -- filter=129 channel=115
    1, 7, 1, -1, 2, -4, -1, -4, 1,
    -- filter=129 channel=116
    3, -31, -18, 16, 31, 15, -5, -14, -10,
    -- filter=129 channel=117
    -7, -8, -9, 0, 5, -1, -2, -5, 0,
    -- filter=129 channel=118
    -2, 0, -4, 6, -1, 2, 3, -2, -2,
    -- filter=129 channel=119
    5, -5, 3, -2, -8, -9, 1, -9, -7,
    -- filter=129 channel=120
    -16, -20, -11, 19, 8, 9, -18, -20, -8,
    -- filter=129 channel=121
    2, -11, 0, 17, 12, -1, 3, -13, -1,
    -- filter=129 channel=122
    -10, -4, 0, 14, 13, -9, -2, -5, 8,
    -- filter=129 channel=123
    -1, 2, 6, 11, -5, 1, 8, 6, 9,
    -- filter=129 channel=124
    -5, -2, 7, 2, 8, 4, -5, 1, -3,
    -- filter=129 channel=125
    -7, -24, -12, 8, 17, -4, -13, -4, -5,
    -- filter=129 channel=126
    -13, -18, -7, 18, 12, 15, -9, -13, -2,
    -- filter=129 channel=127
    0, 5, -8, 0, -1, -5, -2, -7, -2,
    -- filter=130 channel=0
    7, 5, 9, -5, 2, 3, -2, 10, 10,
    -- filter=130 channel=1
    5, -5, 12, -3, 3, 3, -5, 2, 10,
    -- filter=130 channel=2
    -2, 3, 1, 5, -8, 7, -1, 4, 6,
    -- filter=130 channel=3
    3, 5, 8, 4, 2, 8, 0, -4, 10,
    -- filter=130 channel=4
    0, -6, -3, -7, -3, 8, -2, 9, 2,
    -- filter=130 channel=5
    2, 2, 5, 0, 6, 12, 2, 11, 2,
    -- filter=130 channel=6
    4, 3, 0, 1, 1, 1, 6, 3, 8,
    -- filter=130 channel=7
    -2, 1, -3, -1, 6, -3, 0, -1, 4,
    -- filter=130 channel=8
    5, 3, -2, 2, -6, 0, -5, -7, -6,
    -- filter=130 channel=9
    -5, 1, 1, 2, -10, -3, 4, -3, -5,
    -- filter=130 channel=10
    10, 5, 3, 5, -7, -7, 0, -13, 0,
    -- filter=130 channel=11
    -4, -1, 0, 5, 10, 1, 3, 0, 9,
    -- filter=130 channel=12
    1, -6, 1, 1, -10, 2, 6, -2, 2,
    -- filter=130 channel=13
    -1, 1, 0, 7, -2, -3, 0, -13, -9,
    -- filter=130 channel=14
    3, 6, -5, -6, 2, 3, 7, 0, -6,
    -- filter=130 channel=15
    -8, 3, -1, -3, 2, -1, -10, 1, -8,
    -- filter=130 channel=16
    -7, -12, -3, -10, -2, -1, 0, -13, 5,
    -- filter=130 channel=17
    -3, 2, -5, -4, 5, -2, 0, 1, 0,
    -- filter=130 channel=18
    5, 2, -9, 6, 18, 4, -9, 8, -8,
    -- filter=130 channel=19
    -1, -3, 1, -6, 0, 3, -4, 1, 5,
    -- filter=130 channel=20
    0, -4, -4, 15, 23, -1, -4, 15, 9,
    -- filter=130 channel=21
    -10, -7, -2, -7, -18, -8, -16, -16, -6,
    -- filter=130 channel=22
    -2, 9, -3, 1, 5, 3, -4, 0, 0,
    -- filter=130 channel=23
    5, 4, -9, 9, 4, -2, -1, -5, 9,
    -- filter=130 channel=24
    -4, -3, -5, 5, -5, 6, 7, 1, 4,
    -- filter=130 channel=25
    -4, -1, -5, -9, -4, -2, -7, -5, -10,
    -- filter=130 channel=26
    -6, 6, 6, 2, 5, 10, -4, 6, 3,
    -- filter=130 channel=27
    3, -6, 0, -5, -5, -3, -8, -8, 0,
    -- filter=130 channel=28
    1, -4, -6, -1, 0, 4, -4, -2, -4,
    -- filter=130 channel=29
    5, 13, -11, 14, 22, -2, -4, 11, 9,
    -- filter=130 channel=30
    -3, -1, 0, -1, 0, 0, -4, 0, 4,
    -- filter=130 channel=31
    -11, -7, -3, -14, -21, 4, -14, -15, 7,
    -- filter=130 channel=32
    3, 7, 1, 0, 8, 3, -12, 3, 1,
    -- filter=130 channel=33
    3, 0, 1, 0, 2, -2, -11, -2, 6,
    -- filter=130 channel=34
    7, -4, -1, 4, -9, 1, 1, -4, 2,
    -- filter=130 channel=35
    -1, 3, 5, 7, -5, 0, -6, 0, 6,
    -- filter=130 channel=36
    -5, -2, -5, -1, -8, 5, -1, -2, 5,
    -- filter=130 channel=37
    -3, -5, 10, -10, 3, 2, 5, 5, 7,
    -- filter=130 channel=38
    4, -6, -8, 6, 2, 5, -7, -4, 0,
    -- filter=130 channel=39
    4, 5, 0, 0, 0, 2, -2, 3, -6,
    -- filter=130 channel=40
    0, -6, -7, 6, 4, -5, -5, 4, 3,
    -- filter=130 channel=41
    7, -2, -1, 12, 0, -5, 7, -4, -1,
    -- filter=130 channel=42
    -2, -7, -2, -7, -6, -2, -8, 2, 6,
    -- filter=130 channel=43
    6, 8, 2, 7, 15, 5, 8, -1, 5,
    -- filter=130 channel=44
    -7, -8, 4, -12, -4, 7, -3, -14, -8,
    -- filter=130 channel=45
    -8, 3, 0, -8, 3, 2, -6, 0, -4,
    -- filter=130 channel=46
    2, 8, -6, 8, 3, 2, 2, 3, -6,
    -- filter=130 channel=47
    -6, -8, 0, -18, -13, -6, -2, -8, -2,
    -- filter=130 channel=48
    -8, -9, -9, -14, -22, -4, -5, -13, -2,
    -- filter=130 channel=49
    2, 6, -4, -5, -2, -4, -3, 8, 1,
    -- filter=130 channel=50
    0, -1, -4, -6, -10, -1, -6, 0, -9,
    -- filter=130 channel=51
    -5, 1, -6, 4, 5, 2, 1, 4, 5,
    -- filter=130 channel=52
    2, -6, -4, 1, 6, -4, 5, -7, 4,
    -- filter=130 channel=53
    -4, 1, -9, 5, 10, -3, 4, 0, 7,
    -- filter=130 channel=54
    2, -4, -6, -5, -4, -7, -1, -2, -2,
    -- filter=130 channel=55
    -1, -4, -2, 11, 9, -6, -3, -3, 3,
    -- filter=130 channel=56
    7, 0, -3, -3, -6, 6, 0, 7, 5,
    -- filter=130 channel=57
    -1, 5, -2, -4, -3, -6, 6, 3, 0,
    -- filter=130 channel=58
    6, 2, 8, 5, 0, 2, 8, 0, 12,
    -- filter=130 channel=59
    -7, -1, -11, -5, -18, -6, -1, -17, -3,
    -- filter=130 channel=60
    0, -7, 7, 4, 7, 3, -4, 1, 3,
    -- filter=130 channel=61
    7, 5, 0, -2, 0, 4, 1, 0, 0,
    -- filter=130 channel=62
    7, -2, 3, -3, 8, -4, 6, 4, -6,
    -- filter=130 channel=63
    1, 0, 0, -1, 0, 13, 1, 0, 8,
    -- filter=130 channel=64
    1, -7, 0, -3, 0, -6, -4, 3, 5,
    -- filter=130 channel=65
    -7, -2, 4, 4, -2, -1, -5, 0, 3,
    -- filter=130 channel=66
    0, -5, -10, 0, 0, 2, 5, 2, -4,
    -- filter=130 channel=67
    -1, 3, 5, -4, -3, 1, 3, -5, -5,
    -- filter=130 channel=68
    -4, -8, -5, 0, -6, -5, 6, 7, -4,
    -- filter=130 channel=69
    3, 5, 6, 0, 0, -5, 1, 0, 1,
    -- filter=130 channel=70
    6, 0, 0, 3, -2, 3, -4, -7, -3,
    -- filter=130 channel=71
    5, 3, -1, -4, 0, 7, 1, 2, 7,
    -- filter=130 channel=72
    -5, -4, -4, -7, -11, 1, 0, -5, 3,
    -- filter=130 channel=73
    -7, -2, -6, -2, -4, 0, -3, 4, 1,
    -- filter=130 channel=74
    0, -5, 1, 6, -8, 5, 7, 1, -8,
    -- filter=130 channel=75
    0, 7, 6, -6, -4, 2, 2, -5, 2,
    -- filter=130 channel=76
    -2, 8, -10, 6, 23, 4, -8, 0, 2,
    -- filter=130 channel=77
    -4, 2, 7, 2, 4, 5, 4, -4, 0,
    -- filter=130 channel=78
    2, -4, 0, -4, -5, -2, 4, 2, 6,
    -- filter=130 channel=79
    8, 5, -3, 3, 7, -9, -11, 7, -5,
    -- filter=130 channel=80
    -5, -18, -6, -18, -25, 2, -8, -17, -5,
    -- filter=130 channel=81
    1, 1, -5, 6, 0, -5, 2, 0, 2,
    -- filter=130 channel=82
    -1, -5, -6, -5, -5, 3, -4, -5, 4,
    -- filter=130 channel=83
    4, -7, 5, 0, -8, 1, -8, 4, -1,
    -- filter=130 channel=84
    1, 1, -9, -4, 9, 4, -10, 1, -7,
    -- filter=130 channel=85
    -3, 0, 1, 6, 1, 1, 6, 4, -2,
    -- filter=130 channel=86
    7, 2, 0, 7, -3, 5, 9, 5, -4,
    -- filter=130 channel=87
    6, 6, 3, 13, 9, -1, 4, 9, 1,
    -- filter=130 channel=88
    8, 5, -6, 7, -5, -4, -6, 5, 6,
    -- filter=130 channel=89
    -1, 2, -3, 1, 0, -4, -14, -1, -8,
    -- filter=130 channel=90
    -1, -11, 0, -6, -6, 6, -4, -10, -7,
    -- filter=130 channel=91
    3, 4, -10, -5, 0, -5, -7, 3, 0,
    -- filter=130 channel=92
    -6, 2, -3, -2, -1, 0, 2, 1, 0,
    -- filter=130 channel=93
    0, -1, 0, -6, -15, 1, -4, -10, 4,
    -- filter=130 channel=94
    4, -7, 0, -5, 1, 0, 1, 0, -5,
    -- filter=130 channel=95
    6, 1, 0, 5, 0, 6, -5, -3, 4,
    -- filter=130 channel=96
    0, 1, 2, 4, 4, 1, -8, -2, 4,
    -- filter=130 channel=97
    2, 0, -4, -9, -2, 8, 5, 5, 0,
    -- filter=130 channel=98
    7, 2, -6, -6, -13, -11, -12, -10, -3,
    -- filter=130 channel=99
    6, -4, -12, 0, -6, -5, -9, -4, 0,
    -- filter=130 channel=100
    4, 2, -5, 5, 0, 0, 0, -5, -6,
    -- filter=130 channel=101
    8, -1, 2, -10, -7, 5, -1, -3, 10,
    -- filter=130 channel=102
    6, 0, 6, -1, 2, 5, 4, -1, 4,
    -- filter=130 channel=103
    -3, -3, -12, -10, -17, 0, -17, -12, 0,
    -- filter=130 channel=104
    -7, -7, -2, -11, -7, -5, -3, -16, 0,
    -- filter=130 channel=105
    2, 5, 2, 3, 18, -6, -6, 9, -2,
    -- filter=130 channel=106
    6, 2, -3, 3, 8, 0, 2, 4, -7,
    -- filter=130 channel=107
    1, 3, 0, 8, 17, 8, -6, 5, 8,
    -- filter=130 channel=108
    -2, 7, 1, 0, 8, 8, 2, -3, 2,
    -- filter=130 channel=109
    -4, -1, -8, 0, 2, 0, -12, -4, -2,
    -- filter=130 channel=110
    -2, 2, -1, -1, -3, -2, 2, 0, -1,
    -- filter=130 channel=111
    7, -4, 8, -4, 7, 2, 8, -6, 3,
    -- filter=130 channel=112
    -6, 0, -1, 0, -10, 3, -8, -4, 3,
    -- filter=130 channel=113
    9, -2, -1, 4, -7, -6, -3, -3, -7,
    -- filter=130 channel=114
    2, 7, 7, 7, 18, 12, -11, 6, 12,
    -- filter=130 channel=115
    -1, -7, 1, 4, 4, 6, -5, 1, 0,
    -- filter=130 channel=116
    7, 0, -6, -1, 0, -4, -9, 1, -5,
    -- filter=130 channel=117
    -5, 0, 1, 0, -7, 1, 0, -5, 3,
    -- filter=130 channel=118
    -7, 2, 5, -5, -1, 4, 1, 1, 3,
    -- filter=130 channel=119
    5, 6, -6, 3, -1, 3, -5, -7, -4,
    -- filter=130 channel=120
    3, 7, -10, -4, -2, 0, -2, -3, 6,
    -- filter=130 channel=121
    0, 4, -3, 4, -10, -8, -1, -6, 5,
    -- filter=130 channel=122
    -10, -26, -9, -11, -20, -4, -21, -23, -17,
    -- filter=130 channel=123
    -4, 2, 2, -6, 1, -3, -7, -9, 5,
    -- filter=130 channel=124
    -3, 0, -4, 10, 5, 8, -2, 8, -6,
    -- filter=130 channel=125
    8, 1, 1, -11, -2, 1, -11, 0, -6,
    -- filter=130 channel=126
    8, 8, 5, -7, -4, 3, -4, 6, 0,
    -- filter=130 channel=127
    2, 2, 0, 2, -3, 1, -2, 5, 4,
    -- filter=131 channel=0
    8, 5, 8, 1, 6, -1, -2, 5, 8,
    -- filter=131 channel=1
    10, -1, 0, 0, -1, -7, 7, 0, -1,
    -- filter=131 channel=2
    -1, 0, 0, -1, 0, 1, -5, -4, -6,
    -- filter=131 channel=3
    6, 12, 23, 3, -5, 4, 3, -9, 0,
    -- filter=131 channel=4
    -3, -10, 8, -7, -8, 3, 0, 9, 5,
    -- filter=131 channel=5
    0, 15, 12, -3, 11, 11, 1, 2, 0,
    -- filter=131 channel=6
    7, 1, -1, -2, 9, -4, 0, 8, 6,
    -- filter=131 channel=7
    -4, -3, 4, 2, 7, 6, -2, -5, -2,
    -- filter=131 channel=8
    0, 5, -4, 2, -3, -2, 5, -6, -4,
    -- filter=131 channel=9
    -9, -2, 2, -8, 3, 5, 0, 3, 0,
    -- filter=131 channel=10
    8, 0, 2, -4, -11, 0, -1, -12, -11,
    -- filter=131 channel=11
    4, 4, 4, 1, -9, 2, -2, 4, -1,
    -- filter=131 channel=12
    -3, -7, 1, -3, -13, 2, 1, -1, -8,
    -- filter=131 channel=13
    0, -10, -5, 4, -19, -12, 0, -14, -15,
    -- filter=131 channel=14
    -2, 6, -6, 5, -4, 4, -4, 1, 3,
    -- filter=131 channel=15
    9, 8, 11, 0, -15, -9, 2, -2, -3,
    -- filter=131 channel=16
    10, 0, 11, 4, 3, 10, -4, 7, 2,
    -- filter=131 channel=17
    -7, 2, 7, 6, -3, -2, -1, 5, 2,
    -- filter=131 channel=18
    -1, -5, 8, -4, -12, -9, 7, -6, -5,
    -- filter=131 channel=19
    5, 5, 2, -4, -2, -4, 4, -4, 2,
    -- filter=131 channel=20
    0, 8, 4, 4, 7, 14, 15, 3, 9,
    -- filter=131 channel=21
    0, 7, -1, 6, 8, 4, 5, 0, 2,
    -- filter=131 channel=22
    -2, 10, 6, -1, 4, -1, -5, 0, -7,
    -- filter=131 channel=23
    -5, 11, 32, -12, -20, -1, -10, -11, -11,
    -- filter=131 channel=24
    3, 2, 4, 2, -6, -6, 0, -2, 4,
    -- filter=131 channel=25
    -9, -2, -4, 3, -16, -15, 6, -4, -2,
    -- filter=131 channel=26
    2, 0, -4, 5, 9, 3, 10, 15, 13,
    -- filter=131 channel=27
    -12, -2, 20, -17, -20, -13, 0, -15, -19,
    -- filter=131 channel=28
    3, -3, -3, 6, 3, 2, -2, -7, -2,
    -- filter=131 channel=29
    0, -7, 5, -3, 2, 6, 12, -1, 6,
    -- filter=131 channel=30
    0, -9, 7, 0, -2, -10, -2, -3, -9,
    -- filter=131 channel=31
    -7, 8, 20, -12, -12, 0, -2, -8, -5,
    -- filter=131 channel=32
    1, -11, 4, -12, -20, -5, -6, -3, -10,
    -- filter=131 channel=33
    0, 2, 10, -8, -11, 1, -9, -17, -10,
    -- filter=131 channel=34
    -10, 12, 14, -3, -2, 2, 4, -9, 4,
    -- filter=131 channel=35
    -4, 3, -3, -4, 3, -4, 4, -6, 7,
    -- filter=131 channel=36
    0, -2, 3, 0, 6, -2, 13, 5, 9,
    -- filter=131 channel=37
    -5, 4, 7, -9, 5, 0, -4, 5, 1,
    -- filter=131 channel=38
    -8, -1, 13, -9, -3, -1, -7, -11, -3,
    -- filter=131 channel=39
    6, -5, 8, -2, 1, 2, 9, 0, 6,
    -- filter=131 channel=40
    12, 9, 14, 9, -2, 2, 3, 7, -1,
    -- filter=131 channel=41
    17, -15, -13, 11, -3, -14, 6, -8, -14,
    -- filter=131 channel=42
    -3, -2, 0, 4, -7, 2, -9, -1, 5,
    -- filter=131 channel=43
    3, 10, 15, 2, 5, 10, -1, -6, 6,
    -- filter=131 channel=44
    0, -2, 1, 0, -9, -6, -1, -8, -1,
    -- filter=131 channel=45
    9, -1, 8, -4, 10, 11, 4, 10, 1,
    -- filter=131 channel=46
    3, 7, 6, -2, -6, -3, 7, 4, 5,
    -- filter=131 channel=47
    5, 5, 10, 1, -6, 6, -9, 2, -2,
    -- filter=131 channel=48
    -10, -14, 4, -1, -3, -3, 0, 6, -11,
    -- filter=131 channel=49
    1, 2, 3, -5, -13, 1, 1, 0, -1,
    -- filter=131 channel=50
    -2, 1, 0, -8, -3, -6, -7, -3, -10,
    -- filter=131 channel=51
    7, 5, 3, -1, 0, 1, -3, -4, -6,
    -- filter=131 channel=52
    -1, 6, 10, -8, 3, 6, 1, -6, -3,
    -- filter=131 channel=53
    -7, 3, 9, 5, -8, -5, -2, 1, 2,
    -- filter=131 channel=54
    1, -3, 1, -6, -3, 4, -1, -3, 1,
    -- filter=131 channel=55
    -1, 1, 3, 3, -18, -10, 2, -1, -13,
    -- filter=131 channel=56
    1, -7, -5, 1, 0, 2, -1, -9, -1,
    -- filter=131 channel=57
    -5, -6, 0, -4, -5, -4, -1, -5, -4,
    -- filter=131 channel=58
    -1, 7, 7, -4, 5, 2, -1, 6, 8,
    -- filter=131 channel=59
    6, -2, -4, -1, -10, -13, 2, 0, -9,
    -- filter=131 channel=60
    4, -4, 0, 5, -1, -6, -3, 0, 8,
    -- filter=131 channel=61
    -4, 4, 4, 3, 0, 1, 4, 6, 3,
    -- filter=131 channel=62
    1, 0, 6, 7, 2, -5, -6, 4, 2,
    -- filter=131 channel=63
    5, 4, -1, 9, 8, 11, 9, 10, 12,
    -- filter=131 channel=64
    5, -3, 7, -4, 2, -4, 8, 5, 8,
    -- filter=131 channel=65
    -4, -6, -5, -7, -4, 6, -1, -3, 5,
    -- filter=131 channel=66
    1, -12, -6, -1, -6, -12, 10, -12, -7,
    -- filter=131 channel=67
    1, -2, 8, 5, 5, -4, 8, 5, 0,
    -- filter=131 channel=68
    1, 0, 0, -2, 0, -5, -2, 5, 3,
    -- filter=131 channel=69
    -4, 0, 0, 6, -7, 1, 2, -1, 5,
    -- filter=131 channel=70
    -1, -3, 16, -15, -9, -7, -6, -17, -11,
    -- filter=131 channel=71
    1, 13, 16, 5, 1, 2, -4, -4, 2,
    -- filter=131 channel=72
    -1, -10, 7, 4, -6, -4, -5, -8, -9,
    -- filter=131 channel=73
    -5, -1, 0, -7, -6, -7, -4, 1, -6,
    -- filter=131 channel=74
    -3, 6, 18, -3, -9, 8, -1, -11, -2,
    -- filter=131 channel=75
    5, 0, 10, 1, -7, 0, -7, -2, -3,
    -- filter=131 channel=76
    13, 0, 12, 4, 2, 0, 2, -2, 3,
    -- filter=131 channel=77
    7, -2, 4, 6, 0, -3, 4, -3, 1,
    -- filter=131 channel=78
    5, 11, 1, -8, 9, 5, -2, -4, 11,
    -- filter=131 channel=79
    4, 3, 15, 0, -20, -10, 0, -13, -21,
    -- filter=131 channel=80
    2, -1, 6, -6, -10, 0, 1, -3, -5,
    -- filter=131 channel=81
    0, -5, -1, -6, 2, 1, 0, 0, -5,
    -- filter=131 channel=82
    -4, -1, 12, 4, 8, 0, -5, -7, -2,
    -- filter=131 channel=83
    3, 2, -6, 2, -5, 0, 1, 4, -4,
    -- filter=131 channel=84
    -6, -6, 8, 0, -5, -5, -6, 3, -11,
    -- filter=131 channel=85
    3, -7, 0, 6, 5, 3, -2, 7, 6,
    -- filter=131 channel=86
    -4, 4, 3, -9, -3, 2, 6, 3, 4,
    -- filter=131 channel=87
    2, 0, 0, 6, -3, 0, -4, 0, 7,
    -- filter=131 channel=88
    2, 0, -2, -3, -2, -1, 11, 8, 9,
    -- filter=131 channel=89
    5, -2, 8, 3, -10, -3, -3, -5, -11,
    -- filter=131 channel=90
    9, 15, 6, 0, 8, 15, 1, 6, 0,
    -- filter=131 channel=91
    -9, -12, 2, 0, -14, -14, -3, -9, -12,
    -- filter=131 channel=92
    0, -1, 4, -4, 3, 3, 1, -2, 2,
    -- filter=131 channel=93
    -1, -9, 4, -5, 0, -6, 3, 6, 7,
    -- filter=131 channel=94
    -6, 1, 4, -1, -3, -7, 0, 1, -5,
    -- filter=131 channel=95
    7, 3, 6, 0, -5, 3, 2, -7, 4,
    -- filter=131 channel=96
    -2, -7, 7, 6, 6, 0, -4, -1, -7,
    -- filter=131 channel=97
    7, 8, 9, 4, 0, 6, 2, 1, -6,
    -- filter=131 channel=98
    0, -9, 3, -1, -18, -10, -6, -4, -14,
    -- filter=131 channel=99
    -10, -5, 18, 0, -17, -4, 0, -6, -10,
    -- filter=131 channel=100
    -7, 4, 2, -3, -1, -6, 3, 0, -4,
    -- filter=131 channel=101
    3, 1, 9, 0, 3, 2, 7, -1, 0,
    -- filter=131 channel=102
    -7, -7, 4, -2, 0, 0, 3, 7, 4,
    -- filter=131 channel=103
    -3, 6, 8, -9, 0, 7, -8, -2, 2,
    -- filter=131 channel=104
    -1, -10, 7, 2, -12, -6, 6, -4, -7,
    -- filter=131 channel=105
    9, -1, 9, 3, 5, 6, 0, 6, 4,
    -- filter=131 channel=106
    6, 7, -5, 9, 7, 4, 3, 2, 5,
    -- filter=131 channel=107
    7, 6, 9, 7, -2, 12, 0, -2, -2,
    -- filter=131 channel=108
    3, 2, 0, 8, 4, -6, 6, -2, 2,
    -- filter=131 channel=109
    0, -12, 4, -8, -11, -18, -4, -12, -3,
    -- filter=131 channel=110
    -1, 6, 3, 0, 0, 1, -3, -6, 0,
    -- filter=131 channel=111
    6, -6, 0, 10, 3, -8, -2, 10, 0,
    -- filter=131 channel=112
    -10, 8, 9, -6, 0, -4, -9, -1, -4,
    -- filter=131 channel=113
    0, 11, 13, -1, -13, 0, -2, -8, -14,
    -- filter=131 channel=114
    5, -8, 5, -10, -18, -11, 8, 0, -12,
    -- filter=131 channel=115
    4, 6, 6, -1, 7, -2, 7, -6, -3,
    -- filter=131 channel=116
    -1, -6, -2, 4, -4, -6, 2, -5, -1,
    -- filter=131 channel=117
    0, -7, 0, 6, -7, -8, 5, 1, -1,
    -- filter=131 channel=118
    0, 6, 2, 4, -3, 0, -1, -5, -5,
    -- filter=131 channel=119
    -6, 1, 8, -5, -4, 3, -2, -7, -4,
    -- filter=131 channel=120
    -8, 4, 13, -4, -10, -7, 6, 2, -4,
    -- filter=131 channel=121
    3, -8, -4, -2, -3, -12, 7, -2, -6,
    -- filter=131 channel=122
    1, 10, 4, 8, 5, 4, -2, 10, 14,
    -- filter=131 channel=123
    1, 5, 10, -3, 6, -1, 1, -8, 1,
    -- filter=131 channel=124
    -5, -3, 10, 6, -1, -2, 5, 2, 9,
    -- filter=131 channel=125
    -4, -4, -4, -9, -12, -14, 0, 3, -8,
    -- filter=131 channel=126
    5, -4, 7, -1, -6, -3, -5, 0, 0,
    -- filter=131 channel=127
    -1, 1, -6, -2, 5, -5, 5, 2, -8,
    -- filter=132 channel=0
    -5, -5, 2, -5, -14, -2, 5, -9, 0,
    -- filter=132 channel=1
    5, -8, -6, 5, -4, -1, -1, 0, -3,
    -- filter=132 channel=2
    4, 2, 0, 5, -4, -1, 0, -3, -3,
    -- filter=132 channel=3
    -3, -8, -5, 2, -1, 4, 2, -6, 2,
    -- filter=132 channel=4
    9, -3, -6, -5, 1, 0, 2, 7, 1,
    -- filter=132 channel=5
    -9, 1, 5, -14, -10, 3, -4, 1, 16,
    -- filter=132 channel=6
    3, -4, -7, 8, -7, -1, -2, 0, -9,
    -- filter=132 channel=7
    4, 2, 2, 0, -3, 0, -6, 3, 5,
    -- filter=132 channel=8
    -5, 2, 2, -9, -5, -10, 5, -3, 0,
    -- filter=132 channel=9
    -5, 2, 4, 4, -7, -3, 1, 4, 6,
    -- filter=132 channel=10
    14, 0, -2, 16, -2, 0, 7, 2, -4,
    -- filter=132 channel=11
    5, -5, 1, 6, 6, 0, -3, -4, -9,
    -- filter=132 channel=12
    -1, -1, -3, -6, -7, 3, 3, 1, 0,
    -- filter=132 channel=13
    20, 0, -15, 19, -14, -11, 13, 2, -2,
    -- filter=132 channel=14
    0, -2, 0, -4, 0, 0, -4, 2, -6,
    -- filter=132 channel=15
    20, -11, -10, 18, -9, -16, 3, -19, -15,
    -- filter=132 channel=16
    -12, 4, 5, -9, -4, 11, -1, 9, 10,
    -- filter=132 channel=17
    7, 5, 7, 0, 1, -2, 1, -1, -1,
    -- filter=132 channel=18
    25, -8, -13, 18, -7, -27, 7, -18, -13,
    -- filter=132 channel=19
    0, -4, -5, 4, -5, -6, -7, 5, 4,
    -- filter=132 channel=20
    17, 9, -8, 16, 0, -6, 4, -2, -2,
    -- filter=132 channel=21
    -12, -4, 15, -8, 11, 22, 6, 3, 10,
    -- filter=132 channel=22
    -5, -8, -11, 5, -1, -2, 5, -10, -8,
    -- filter=132 channel=23
    9, -17, -24, 8, -15, -17, -4, -21, -21,
    -- filter=132 channel=24
    -4, 0, 0, -2, -6, 0, 0, -5, -3,
    -- filter=132 channel=25
    4, -3, 0, 5, -7, -3, 1, 3, -7,
    -- filter=132 channel=26
    -1, -3, 9, -12, 4, 2, 3, 2, 12,
    -- filter=132 channel=27
    16, -19, -12, 0, -24, -24, 2, -17, -14,
    -- filter=132 channel=28
    -6, -6, -3, -4, 3, -3, 5, -5, 7,
    -- filter=132 channel=29
    21, 3, -7, 12, 2, -8, 3, 2, -10,
    -- filter=132 channel=30
    -4, -3, 0, -3, -13, 3, -7, 3, 3,
    -- filter=132 channel=31
    -15, -2, 8, -6, -2, 0, 0, 13, 12,
    -- filter=132 channel=32
    23, -10, -10, 7, -10, -20, 8, -13, -10,
    -- filter=132 channel=33
    9, -10, -14, 6, -12, -13, 0, -9, -3,
    -- filter=132 channel=34
    -3, -6, -5, -12, -9, -7, -9, -12, -9,
    -- filter=132 channel=35
    -5, -4, 1, 0, 6, 2, 5, 4, -7,
    -- filter=132 channel=36
    3, 8, -2, -4, 3, 1, 6, 3, 7,
    -- filter=132 channel=37
    -10, -12, 11, -10, -12, 5, -8, -4, 14,
    -- filter=132 channel=38
    7, -8, -6, 7, -5, -6, -2, -4, 3,
    -- filter=132 channel=39
    8, 8, 1, 12, -3, 3, 0, -7, 4,
    -- filter=132 channel=40
    -2, 3, 4, 0, 4, 1, 5, -1, -8,
    -- filter=132 channel=41
    26, 0, -10, 20, 4, -6, 14, 2, -10,
    -- filter=132 channel=42
    -4, 2, 0, 5, -1, -3, 2, 3, -6,
    -- filter=132 channel=43
    3, 0, -10, 8, 2, -13, -2, -9, -1,
    -- filter=132 channel=44
    -4, -10, 10, -15, -10, -2, 3, 6, 8,
    -- filter=132 channel=45
    0, -2, 1, 4, 0, 7, -6, 0, -2,
    -- filter=132 channel=46
    2, -3, -7, -2, 5, -7, -3, 0, -5,
    -- filter=132 channel=47
    -8, 0, 4, -10, 3, 17, 6, 2, 6,
    -- filter=132 channel=48
    -3, 0, 3, -4, -4, -6, 3, 11, 0,
    -- filter=132 channel=49
    3, -8, -3, 5, -13, -9, 2, -3, -7,
    -- filter=132 channel=50
    6, -12, -8, -3, -8, 1, 2, 3, -8,
    -- filter=132 channel=51
    6, 2, -4, -7, -1, -3, 6, 2, 7,
    -- filter=132 channel=52
    1, 2, -8, -5, -5, 0, -5, -5, 0,
    -- filter=132 channel=53
    8, 4, 1, 0, 3, 2, 5, -4, -11,
    -- filter=132 channel=54
    -5, 6, 6, 0, 5, 7, 4, -4, 6,
    -- filter=132 channel=55
    28, -8, -22, 19, -11, -17, 8, -10, -13,
    -- filter=132 channel=56
    -6, 4, -8, 6, 5, -11, 3, 5, -7,
    -- filter=132 channel=57
    -2, -3, -7, -3, 3, -7, -2, 0, -2,
    -- filter=132 channel=58
    -3, 3, -1, -8, 0, 8, 5, 0, 1,
    -- filter=132 channel=59
    15, -1, -8, 9, 0, -3, 3, 4, -2,
    -- filter=132 channel=60
    -1, -4, -1, -2, 0, 5, 4, 6, -4,
    -- filter=132 channel=61
    -3, -6, 0, -3, -2, 4, -5, 3, -1,
    -- filter=132 channel=62
    5, -2, -1, 0, 3, -4, -2, 6, -5,
    -- filter=132 channel=63
    1, 0, 12, -8, -6, 12, -2, 9, 7,
    -- filter=132 channel=64
    0, 0, -3, -2, 7, 0, 4, 7, 1,
    -- filter=132 channel=65
    -1, 4, -2, -2, -4, 1, 3, 4, -1,
    -- filter=132 channel=66
    7, -5, -6, -4, -8, -1, 0, 0, -1,
    -- filter=132 channel=67
    -1, -4, 5, 3, 0, -2, -4, -3, -6,
    -- filter=132 channel=68
    6, 0, -2, 3, -3, -2, 0, 6, -1,
    -- filter=132 channel=69
    0, 1, 7, -1, 5, 4, 8, 3, -3,
    -- filter=132 channel=70
    7, -19, -17, 6, -20, -20, -2, -5, -16,
    -- filter=132 channel=71
    2, 6, 0, -1, 8, 0, 8, -3, -1,
    -- filter=132 channel=72
    5, -4, 4, 2, 9, 1, 7, 7, 6,
    -- filter=132 channel=73
    11, -5, -7, 14, -2, -16, 1, -13, -2,
    -- filter=132 channel=74
    -5, -10, -12, -14, -17, -2, -3, -8, -9,
    -- filter=132 channel=75
    -4, -4, -7, 2, -4, 4, 6, -8, -1,
    -- filter=132 channel=76
    10, -1, -12, 22, 3, -8, 8, -10, -13,
    -- filter=132 channel=77
    -1, 1, -5, 0, -2, 6, 1, -6, -1,
    -- filter=132 channel=78
    0, 0, 4, -4, 4, 1, -2, 6, 0,
    -- filter=132 channel=79
    19, -3, -23, 26, -21, -24, 6, -21, -25,
    -- filter=132 channel=80
    0, -3, 10, 8, -7, 6, 12, 4, 1,
    -- filter=132 channel=81
    -3, 5, -7, 0, 5, -1, 1, 6, 0,
    -- filter=132 channel=82
    3, -4, -7, 0, -7, 4, -6, 6, 0,
    -- filter=132 channel=83
    2, -5, 4, -6, -5, -1, -1, 0, 2,
    -- filter=132 channel=84
    9, 0, -13, 9, -3, -18, 4, -1, -4,
    -- filter=132 channel=85
    -3, 0, -5, -1, 0, -2, 7, 7, -1,
    -- filter=132 channel=86
    -12, -8, -10, -7, -12, 0, -9, -5, -3,
    -- filter=132 channel=87
    1, 0, -4, -3, 1, -2, -10, -8, -4,
    -- filter=132 channel=88
    -5, 5, 10, -9, 0, 4, -3, 9, 11,
    -- filter=132 channel=89
    19, 2, -11, 17, -6, -15, 19, 2, -17,
    -- filter=132 channel=90
    -8, -8, 5, -4, 8, 4, 0, -1, 6,
    -- filter=132 channel=91
    14, -5, -13, 0, -6, -13, 0, -1, -13,
    -- filter=132 channel=92
    -1, 2, -7, -4, 3, -4, -2, -7, -3,
    -- filter=132 channel=93
    -12, -2, 4, -9, -11, 9, 5, -2, 2,
    -- filter=132 channel=94
    5, -1, 6, -2, 4, 4, -7, 3, -5,
    -- filter=132 channel=95
    4, -6, 0, 5, -1, -3, -6, 0, -8,
    -- filter=132 channel=96
    7, 2, -5, -4, -1, -3, 6, 3, 2,
    -- filter=132 channel=97
    0, 8, 5, -5, 0, 3, 5, 7, -8,
    -- filter=132 channel=98
    15, -1, -2, 16, -11, -13, 9, -9, 2,
    -- filter=132 channel=99
    1, -2, -12, -5, -7, -6, -4, -1, 1,
    -- filter=132 channel=100
    0, 4, 0, -2, 8, 1, 7, -7, -10,
    -- filter=132 channel=101
    0, 0, 2, 5, 2, -6, -6, 7, 4,
    -- filter=132 channel=102
    7, -3, 0, -4, -1, 6, 3, 0, -2,
    -- filter=132 channel=103
    -11, -4, -2, -12, 3, 9, 0, 8, 19,
    -- filter=132 channel=104
    -2, 5, 0, 0, 2, 5, 8, -1, 12,
    -- filter=132 channel=105
    13, 7, -9, 5, 7, -12, -2, -8, 0,
    -- filter=132 channel=106
    6, 3, 0, 4, 1, -4, -1, 1, -3,
    -- filter=132 channel=107
    0, -8, -8, 5, -3, -5, -12, -17, -6,
    -- filter=132 channel=108
    0, 7, 0, 4, -2, -6, 5, 6, -3,
    -- filter=132 channel=109
    8, -4, -5, 9, -20, -12, 8, -14, -5,
    -- filter=132 channel=110
    -4, -3, -1, 0, 6, 4, -2, 6, -6,
    -- filter=132 channel=111
    8, 7, 7, 1, 2, -1, -1, 5, 0,
    -- filter=132 channel=112
    -7, -6, -2, -5, -1, -4, -8, -12, 4,
    -- filter=132 channel=113
    7, -9, -10, 10, 2, -7, 6, 3, -9,
    -- filter=132 channel=114
    18, -5, -21, 3, -14, -18, -2, -10, -16,
    -- filter=132 channel=115
    0, -4, 1, -2, -1, 2, -3, 5, 0,
    -- filter=132 channel=116
    19, 6, 1, 14, -4, -7, 1, -1, -4,
    -- filter=132 channel=117
    1, 7, 3, -5, 0, -6, 0, 0, -3,
    -- filter=132 channel=118
    2, 1, -1, -1, 0, 0, 6, -6, 7,
    -- filter=132 channel=119
    0, 1, -6, 1, -8, -11, -2, -11, -3,
    -- filter=132 channel=120
    6, -10, -17, 4, -14, -13, -1, -9, -18,
    -- filter=132 channel=121
    14, 6, -9, 9, 2, -9, 3, -1, 0,
    -- filter=132 channel=122
    -23, 2, 24, -27, 7, 32, -1, 19, 31,
    -- filter=132 channel=123
    2, -2, 2, -7, -3, -9, 0, -4, -4,
    -- filter=132 channel=124
    3, 6, 0, -2, 5, -8, -6, 3, -7,
    -- filter=132 channel=125
    10, -5, 5, 6, -13, 0, 5, 0, 0,
    -- filter=132 channel=126
    9, 7, -8, 23, -2, -12, 6, -4, 2,
    -- filter=132 channel=127
    0, -4, 4, 10, 4, -6, -4, -3, -5,
    -- filter=133 channel=0
    -8, 6, -4, -18, 10, -2, -15, 1, 2,
    -- filter=133 channel=1
    -7, 15, -6, -13, 8, -10, -2, -3, -7,
    -- filter=133 channel=2
    -8, -2, -4, -8, -6, 0, 0, 3, 4,
    -- filter=133 channel=3
    5, -14, 0, 3, -9, -16, -13, -14, -21,
    -- filter=133 channel=4
    2, -14, 4, -8, -4, -4, -8, -26, -8,
    -- filter=133 channel=5
    6, 4, 3, 2, 0, -5, -10, 9, 7,
    -- filter=133 channel=6
    -1, -1, -6, 1, -5, -2, 0, 1, -6,
    -- filter=133 channel=7
    0, -1, -5, 1, -1, 6, -2, -1, -7,
    -- filter=133 channel=8
    -7, -3, 3, 3, 7, -7, -9, -2, -8,
    -- filter=133 channel=9
    -6, 4, -1, -14, 6, 0, -8, -2, 9,
    -- filter=133 channel=10
    2, -3, -8, -1, 4, -6, -11, 10, 0,
    -- filter=133 channel=11
    -2, -2, -3, 8, -7, -2, 0, 0, 6,
    -- filter=133 channel=12
    0, 3, -5, 0, 11, -1, 5, 11, 1,
    -- filter=133 channel=13
    5, -2, -8, -14, 15, -6, -4, 5, -2,
    -- filter=133 channel=14
    -6, -3, -4, 4, 4, -4, -5, -3, -4,
    -- filter=133 channel=15
    8, 3, -2, -3, 6, -13, -4, 13, -8,
    -- filter=133 channel=16
    3, 3, -7, -6, 8, 1, -1, 10, -3,
    -- filter=133 channel=17
    1, 3, 6, -1, 0, -1, -5, 1, 2,
    -- filter=133 channel=18
    3, 11, -15, -2, 9, -8, 0, 2, 0,
    -- filter=133 channel=19
    -2, -1, 5, 0, -2, 6, 5, 2, -5,
    -- filter=133 channel=20
    3, -13, 5, 5, -3, -10, -1, 7, -9,
    -- filter=133 channel=21
    -8, 5, -2, -18, 6, 0, 1, 7, -1,
    -- filter=133 channel=22
    -2, -3, 0, 5, 7, -14, 3, 2, -2,
    -- filter=133 channel=23
    4, -9, 0, 4, 20, -18, -16, 22, -20,
    -- filter=133 channel=24
    7, 4, 6, -2, -1, -3, -6, -4, 5,
    -- filter=133 channel=25
    -1, 20, -2, -19, 31, 1, -21, 13, -5,
    -- filter=133 channel=26
    6, 1, -3, -4, 1, 0, -2, -4, 0,
    -- filter=133 channel=27
    0, 20, -14, -29, 47, -12, -29, 31, -3,
    -- filter=133 channel=28
    0, -1, -2, -4, -4, 2, -6, -5, 3,
    -- filter=133 channel=29
    6, 1, 0, 5, 3, 2, -5, 5, -2,
    -- filter=133 channel=30
    5, 2, -9, -15, 14, -1, -16, 10, 3,
    -- filter=133 channel=31
    -10, 0, -2, -30, 12, 1, -29, 21, 2,
    -- filter=133 channel=32
    3, 15, -6, -18, 32, -16, -7, 16, -13,
    -- filter=133 channel=33
    -3, 14, -2, -13, 15, 0, -15, 19, -9,
    -- filter=133 channel=34
    12, -2, -4, 11, 24, -2, 0, 26, -19,
    -- filter=133 channel=35
    0, 5, 4, -1, 1, -5, -2, -7, -1,
    -- filter=133 channel=36
    -4, -3, -2, 1, -3, 3, 5, -5, -4,
    -- filter=133 channel=37
    2, 13, -7, -13, 2, -5, -6, 7, -10,
    -- filter=133 channel=38
    6, 7, -6, -10, 11, 2, -10, 15, -8,
    -- filter=133 channel=39
    0, -9, 4, 2, 2, -3, -7, 2, 4,
    -- filter=133 channel=40
    -6, -5, -2, 6, 3, -7, -3, 5, -11,
    -- filter=133 channel=41
    4, 13, -21, 9, 24, -16, 23, 15, 1,
    -- filter=133 channel=42
    -8, 4, 10, -4, -4, 14, -6, -12, 11,
    -- filter=133 channel=43
    -1, -4, -7, 9, 5, -13, -6, 6, -14,
    -- filter=133 channel=44
    -7, 8, -4, -19, 10, 2, -7, 14, -6,
    -- filter=133 channel=45
    5, 1, -4, 3, -6, -2, -7, -1, 2,
    -- filter=133 channel=46
    2, 0, -6, 2, -6, 1, 8, -3, 0,
    -- filter=133 channel=47
    9, -1, -10, -18, 14, 7, -10, 7, 8,
    -- filter=133 channel=48
    0, 6, -7, -29, 8, 8, -18, -2, 8,
    -- filter=133 channel=49
    -4, 5, 5, -8, 10, -9, -4, -4, 0,
    -- filter=133 channel=50
    -3, 5, -7, -7, 18, -4, -16, 4, 0,
    -- filter=133 channel=51
    1, -2, 5, 4, -1, 0, 3, -3, 1,
    -- filter=133 channel=52
    -1, 1, -10, 6, 14, -16, -3, 19, -3,
    -- filter=133 channel=53
    4, -2, 6, 7, 7, -6, -2, 4, -6,
    -- filter=133 channel=54
    -3, 4, 1, -5, -6, -5, -2, 1, 0,
    -- filter=133 channel=55
    10, 5, -1, 1, 6, -3, 0, 4, -5,
    -- filter=133 channel=56
    2, 2, 3, 8, 8, 2, 11, 1, 0,
    -- filter=133 channel=57
    7, 5, -5, 4, -2, -4, 8, -1, -3,
    -- filter=133 channel=58
    10, 0, -6, -3, -2, 3, 5, -5, 0,
    -- filter=133 channel=59
    -10, 13, -1, -17, 20, 4, -9, 5, 1,
    -- filter=133 channel=60
    -2, -1, 5, 4, -3, 6, 5, -1, 5,
    -- filter=133 channel=61
    -7, 1, -1, 0, 13, -3, 5, -1, -6,
    -- filter=133 channel=62
    2, -9, -5, 6, -7, -4, 5, 4, 1,
    -- filter=133 channel=63
    6, 0, 7, 4, -2, 2, 3, 0, -1,
    -- filter=133 channel=64
    6, 2, -7, -1, -9, -3, -1, 4, 4,
    -- filter=133 channel=65
    1, -5, 1, 0, 5, 0, -3, 7, 5,
    -- filter=133 channel=66
    12, 4, -2, 2, 13, -11, 9, 24, -9,
    -- filter=133 channel=67
    -2, 1, -4, -1, -6, -3, -2, -4, -7,
    -- filter=133 channel=68
    -1, -1, 4, -4, -6, 5, -4, -8, -3,
    -- filter=133 channel=69
    -1, 4, 6, -1, 0, -2, -1, 0, 4,
    -- filter=133 channel=70
    0, 0, -4, -11, 6, -14, -20, 8, -3,
    -- filter=133 channel=71
    -1, 2, 0, -3, -1, 1, -12, -6, -5,
    -- filter=133 channel=72
    2, 0, -5, -12, 12, 7, -11, 14, 4,
    -- filter=133 channel=73
    0, 0, -3, 0, 13, 1, -6, 5, -5,
    -- filter=133 channel=74
    -4, 4, -18, -10, 26, -13, -17, 31, -16,
    -- filter=133 channel=75
    0, 11, -4, -7, 13, -6, -1, -1, -2,
    -- filter=133 channel=76
    5, -8, -4, 8, -8, -3, 4, -9, -2,
    -- filter=133 channel=77
    2, -4, 3, 0, -6, 4, 6, 4, 5,
    -- filter=133 channel=78
    -4, -3, 6, -4, 3, -7, 6, 0, -4,
    -- filter=133 channel=79
    -4, 17, -4, -21, 32, -15, -18, 10, -3,
    -- filter=133 channel=80
    -7, 15, -6, -32, 27, 11, -20, 3, 20,
    -- filter=133 channel=81
    -1, 6, 7, -6, -7, -5, -5, 4, 2,
    -- filter=133 channel=82
    5, -8, -6, 9, -2, 0, -2, -6, 2,
    -- filter=133 channel=83
    -5, -1, 6, -7, 8, 2, -9, -7, 13,
    -- filter=133 channel=84
    -4, 11, -9, -5, 17, -14, -3, 7, -5,
    -- filter=133 channel=85
    5, -3, -3, -7, -1, -5, 4, 1, -5,
    -- filter=133 channel=86
    7, 11, -8, -6, 10, -4, 1, 21, -6,
    -- filter=133 channel=87
    0, 3, -3, -2, 0, -7, -4, 5, -10,
    -- filter=133 channel=88
    1, -4, -10, -6, -2, -1, 1, -1, 1,
    -- filter=133 channel=89
    -8, 7, 2, -18, 10, -4, -13, 8, 6,
    -- filter=133 channel=90
    -7, -6, -7, 7, -3, -10, 2, 0, -6,
    -- filter=133 channel=91
    -4, 0, 0, -11, 14, -13, -15, 10, 6,
    -- filter=133 channel=92
    5, 3, 0, 12, 4, 5, -4, 0, -3,
    -- filter=133 channel=93
    -1, 1, 2, -4, 1, 3, -9, -7, 0,
    -- filter=133 channel=94
    -6, 2, 6, 6, -1, 1, 6, 6, -4,
    -- filter=133 channel=95
    -6, -7, 2, 1, -2, -4, -6, 1, 5,
    -- filter=133 channel=96
    -4, 3, 6, -8, 2, 0, 0, -3, -2,
    -- filter=133 channel=97
    8, -9, -5, -3, -2, -2, -7, -2, 0,
    -- filter=133 channel=98
    -9, 6, 2, -28, 20, 5, -26, 18, 2,
    -- filter=133 channel=99
    -6, 0, -6, -14, 30, -19, -21, 27, -13,
    -- filter=133 channel=100
    4, -1, -4, 1, -2, 8, 1, 2, 2,
    -- filter=133 channel=101
    2, -5, 3, -10, -5, -13, -4, -10, -13,
    -- filter=133 channel=102
    4, 6, -4, 4, -3, 2, -6, 1, 7,
    -- filter=133 channel=103
    1, 13, -2, -17, 2, -3, -6, 10, -5,
    -- filter=133 channel=104
    -8, 4, -7, -19, 7, 0, -7, 10, 5,
    -- filter=133 channel=105
    9, -1, 7, 1, -11, -6, 10, 4, -4,
    -- filter=133 channel=106
    3, -6, -1, -1, -2, 5, 5, -13, -6,
    -- filter=133 channel=107
    0, 0, -6, -3, -2, -14, -3, 10, -10,
    -- filter=133 channel=108
    7, -1, 0, 0, 5, -5, 6, -5, 3,
    -- filter=133 channel=109
    0, 18, -4, -11, 33, 0, -15, 25, -2,
    -- filter=133 channel=110
    -1, -2, 2, 0, 8, -8, 1, 0, 3,
    -- filter=133 channel=111
    -4, -2, -7, -3, -2, -5, 8, -2, -1,
    -- filter=133 channel=112
    0, 0, 1, -7, 14, -9, -17, 15, 1,
    -- filter=133 channel=113
    8, 10, -6, -12, 8, 0, -17, 16, 2,
    -- filter=133 channel=114
    -4, 24, -18, -14, 27, -9, -11, 18, -2,
    -- filter=133 channel=115
    6, 0, -7, 6, 0, -2, -4, -2, -2,
    -- filter=133 channel=116
    -1, 5, -4, -8, 25, 9, -13, -3, 15,
    -- filter=133 channel=117
    -3, 0, -6, -5, 0, 6, -2, -6, -1,
    -- filter=133 channel=118
    3, -2, 5, 6, 6, -1, 1, 1, 6,
    -- filter=133 channel=119
    12, 0, -11, 20, 14, -9, 7, 23, -12,
    -- filter=133 channel=120
    1, 8, -13, -20, 29, -9, -16, 22, -5,
    -- filter=133 channel=121
    -5, 7, -2, -5, 6, -9, 4, 0, -7,
    -- filter=133 channel=122
    1, 1, -2, -10, 8, -8, -8, 4, -6,
    -- filter=133 channel=123
    6, -2, 1, 16, 0, 0, -1, 8, -6,
    -- filter=133 channel=124
    0, -1, 5, -1, -1, -5, -4, 0, 2,
    -- filter=133 channel=125
    -8, 4, -5, -21, 19, 0, -19, 17, 3,
    -- filter=133 channel=126
    -3, 0, -4, -4, 12, 2, 0, 1, 1,
    -- filter=133 channel=127
    3, 8, 0, 8, 8, 4, -2, 6, 2,
    -- filter=134 channel=0
    -4, 12, 8, 12, 11, -7, -6, -14, 0,
    -- filter=134 channel=1
    7, 20, 13, 14, 5, 0, -7, -2, -9,
    -- filter=134 channel=2
    2, -5, 1, 0, 0, 3, -7, 3, 5,
    -- filter=134 channel=3
    -3, -3, -1, 1, 0, 3, 0, 6, 3,
    -- filter=134 channel=4
    6, 0, 11, 0, 7, 1, 1, 6, 19,
    -- filter=134 channel=5
    0, 6, -4, 3, -3, 1, -13, -17, -13,
    -- filter=134 channel=6
    0, 2, -9, 2, 0, -4, 5, 6, -4,
    -- filter=134 channel=7
    -4, 0, 0, -1, 2, 0, 5, -2, -4,
    -- filter=134 channel=8
    3, 1, 8, 3, 3, 4, -1, 0, 2,
    -- filter=134 channel=9
    3, -5, -9, 1, 4, -1, -9, -11, 2,
    -- filter=134 channel=10
    -3, -4, 0, 0, -2, -3, 5, 0, -1,
    -- filter=134 channel=11
    -10, -13, -15, 4, 2, -4, 4, 1, 2,
    -- filter=134 channel=12
    8, 9, 5, 8, 9, -5, 9, -2, -1,
    -- filter=134 channel=13
    -4, -3, 7, 10, 12, -1, 9, 2, 8,
    -- filter=134 channel=14
    -2, -1, 2, 2, -1, -1, 5, 1, -6,
    -- filter=134 channel=15
    -1, -11, -3, 1, 4, -7, 2, 12, -3,
    -- filter=134 channel=16
    5, 9, 0, 2, 5, 7, -6, -4, -4,
    -- filter=134 channel=17
    1, 4, 0, 4, -4, 3, -1, -1, 6,
    -- filter=134 channel=18
    -7, 0, -3, 8, 7, 1, -5, -6, 0,
    -- filter=134 channel=19
    -6, -6, 4, -7, 1, 4, 3, -3, -2,
    -- filter=134 channel=20
    -4, -19, -11, -5, 0, 0, 12, 12, -1,
    -- filter=134 channel=21
    9, 2, -1, 3, -6, -4, -2, -6, -5,
    -- filter=134 channel=22
    0, 8, -5, -2, -2, -6, -1, 1, 6,
    -- filter=134 channel=23
    -10, -12, 2, -2, 1, -7, -3, 15, 5,
    -- filter=134 channel=24
    -5, -2, 3, 4, -3, 0, -3, 0, 1,
    -- filter=134 channel=25
    0, -2, 8, -4, 10, -11, -14, -6, 8,
    -- filter=134 channel=26
    -2, 9, 4, -1, 3, -3, -1, 2, 2,
    -- filter=134 channel=27
    5, 0, 6, 8, 4, -4, -7, -3, 9,
    -- filter=134 channel=28
    -1, 6, -5, 5, -4, -1, 0, 2, 5,
    -- filter=134 channel=29
    -8, -6, -14, 2, -3, -3, 10, 11, 7,
    -- filter=134 channel=30
    -4, 5, 2, 7, -2, -6, -5, 0, 0,
    -- filter=134 channel=31
    5, -4, -2, 1, 2, -1, -8, -11, 11,
    -- filter=134 channel=32
    -4, -6, -7, 4, 7, -9, 3, 6, 8,
    -- filter=134 channel=33
    -4, 5, 1, 0, -1, -6, -5, 2, -9,
    -- filter=134 channel=34
    -3, 8, 12, -7, 5, 4, -3, 8, 7,
    -- filter=134 channel=35
    7, 3, -3, 0, 2, 0, -2, -2, 5,
    -- filter=134 channel=36
    5, -2, 2, 0, -2, 5, 2, 0, 0,
    -- filter=134 channel=37
    6, 8, 8, 12, 11, -1, -7, -4, 2,
    -- filter=134 channel=38
    -7, 0, 0, 0, 1, -2, 2, -3, 2,
    -- filter=134 channel=39
    -5, -4, -4, 0, -2, -7, -2, -2, 0,
    -- filter=134 channel=40
    4, -5, 4, -3, 5, 4, 5, 5, 1,
    -- filter=134 channel=41
    2, 8, 13, 3, -2, 8, 1, -9, 2,
    -- filter=134 channel=42
    -6, -3, 0, 3, -2, -7, -5, -2, -6,
    -- filter=134 channel=43
    -1, 5, 8, 3, 4, 3, 6, 9, 0,
    -- filter=134 channel=44
    11, 15, 8, 3, 0, 3, -4, -5, 0,
    -- filter=134 channel=45
    6, 4, -9, 1, -7, -8, 4, 3, -6,
    -- filter=134 channel=46
    7, 0, 2, -3, -6, 3, 0, 0, 1,
    -- filter=134 channel=47
    3, 15, -1, 9, 4, -5, -15, -16, 0,
    -- filter=134 channel=48
    9, 4, 5, -3, 1, -2, -17, -16, 0,
    -- filter=134 channel=49
    -8, 0, -10, -4, 2, 0, -2, 0, 11,
    -- filter=134 channel=50
    -1, 0, -8, -1, 0, -1, -11, -5, 7,
    -- filter=134 channel=51
    1, 0, -3, -6, -5, 6, 0, 4, 5,
    -- filter=134 channel=52
    2, -1, 0, 2, 9, -1, 3, 7, 8,
    -- filter=134 channel=53
    0, 0, -11, 8, 0, 2, -1, 6, 0,
    -- filter=134 channel=54
    -1, -5, 4, 6, 0, 1, 4, -2, 5,
    -- filter=134 channel=55
    -2, -12, -14, -3, -3, -9, 0, 8, -1,
    -- filter=134 channel=56
    9, 6, 7, 6, 3, 0, -7, 3, 2,
    -- filter=134 channel=57
    -3, 6, -6, -2, -2, 1, 0, 0, 0,
    -- filter=134 channel=58
    -3, -1, 0, 0, 0, 3, -4, -8, -10,
    -- filter=134 channel=59
    -1, 7, 0, 6, -4, -3, -7, -9, 0,
    -- filter=134 channel=60
    3, 0, -7, -4, 4, 1, 2, -5, 3,
    -- filter=134 channel=61
    5, 0, -5, 5, 5, 1, -2, -1, 4,
    -- filter=134 channel=62
    5, -2, 1, 3, -3, 2, 3, 6, 6,
    -- filter=134 channel=63
    0, -2, -2, 2, 2, 2, -2, -13, 0,
    -- filter=134 channel=64
    -3, 2, 1, -2, -1, 8, 2, 1, -4,
    -- filter=134 channel=65
    -1, -4, 1, 3, 5, 0, 2, -6, 6,
    -- filter=134 channel=66
    10, -1, 4, -2, 4, 2, -2, -3, 2,
    -- filter=134 channel=67
    4, -7, 2, -6, -2, -5, 7, 3, 6,
    -- filter=134 channel=68
    1, 1, 0, -2, -5, 2, 1, 6, -2,
    -- filter=134 channel=69
    6, 7, -4, -1, 7, -7, 4, -1, -1,
    -- filter=134 channel=70
    -6, 4, 0, -2, -3, -2, -4, -2, 8,
    -- filter=134 channel=71
    -4, 8, 4, -2, 7, -5, -6, 7, -6,
    -- filter=134 channel=72
    -7, -7, -8, -1, -3, -5, 0, -9, 3,
    -- filter=134 channel=73
    -1, -4, -3, 0, 2, -9, -5, -6, 9,
    -- filter=134 channel=74
    -5, 8, -4, -1, 3, -5, -7, -5, 4,
    -- filter=134 channel=75
    7, 7, 1, 15, 0, -2, -6, -5, -9,
    -- filter=134 channel=76
    -12, -17, 0, 3, -6, 3, 4, 14, 3,
    -- filter=134 channel=77
    2, -4, -2, 6, -1, 0, -7, -2, -5,
    -- filter=134 channel=78
    4, -5, -5, 0, 0, -3, -2, -8, -8,
    -- filter=134 channel=79
    1, -1, 0, 4, 5, -12, 2, 7, -7,
    -- filter=134 channel=80
    0, 5, 1, 0, 6, -3, -14, -13, 2,
    -- filter=134 channel=81
    -1, 5, 0, -2, -7, 0, -5, -5, 1,
    -- filter=134 channel=82
    3, 6, 3, -6, 0, -3, -7, -3, 5,
    -- filter=134 channel=83
    1, -4, -5, -3, 0, -8, 0, -5, 8,
    -- filter=134 channel=84
    -2, -3, -2, 7, 8, -2, 4, -5, 5,
    -- filter=134 channel=85
    4, 4, 3, 5, -6, 4, -7, 0, -2,
    -- filter=134 channel=86
    -5, 7, 5, 3, 8, 6, 5, 0, -1,
    -- filter=134 channel=87
    4, 3, 6, 0, 5, -2, 7, 3, 11,
    -- filter=134 channel=88
    2, -3, -2, 1, 6, 0, 2, 7, 0,
    -- filter=134 channel=89
    1, -5, -4, 6, 3, 0, -6, 3, -6,
    -- filter=134 channel=90
    -3, 5, -4, 0, 0, 9, 3, 7, 3,
    -- filter=134 channel=91
    0, 0, -6, -4, 2, -8, -10, 3, 14,
    -- filter=134 channel=92
    -1, 0, -2, 4, 2, -3, 0, 7, -2,
    -- filter=134 channel=93
    5, 13, 0, 6, 0, -5, -9, -9, 9,
    -- filter=134 channel=94
    0, 4, 7, -6, 0, -1, -2, 0, 5,
    -- filter=134 channel=95
    -1, -3, 1, 0, 3, -5, -4, 4, 5,
    -- filter=134 channel=96
    6, 0, 3, -4, 2, -6, 3, 1, -6,
    -- filter=134 channel=97
    2, -5, -3, 4, 1, -2, -6, -4, -9,
    -- filter=134 channel=98
    1, 2, -3, 5, -3, -5, -10, -11, -3,
    -- filter=134 channel=99
    -1, -4, -5, 5, 0, -13, -9, 9, 4,
    -- filter=134 channel=100
    8, -1, 0, 3, 6, 9, -6, 6, 7,
    -- filter=134 channel=101
    0, 2, 5, -4, 0, 6, -1, 11, 13,
    -- filter=134 channel=102
    2, 5, -1, -2, -5, -1, -3, -2, 0,
    -- filter=134 channel=103
    3, 9, -12, 1, -4, -5, -13, -10, -7,
    -- filter=134 channel=104
    5, 8, -9, 3, -1, -2, -5, 0, -1,
    -- filter=134 channel=105
    -9, -9, -3, 0, -3, 5, -1, 13, 0,
    -- filter=134 channel=106
    3, -8, -5, 0, -6, -1, 9, 8, -1,
    -- filter=134 channel=107
    5, -2, -11, 1, 8, 1, 5, 13, 8,
    -- filter=134 channel=108
    -6, 6, 0, 3, 0, -1, -6, 1, -7,
    -- filter=134 channel=109
    2, -6, 1, 8, -4, -3, -14, 1, 6,
    -- filter=134 channel=110
    5, 4, 0, -3, 6, 0, 1, -5, 0,
    -- filter=134 channel=111
    -7, 4, 6, 5, -6, 7, 5, -2, 0,
    -- filter=134 channel=112
    0, 2, 2, 4, -5, -6, 2, -6, 1,
    -- filter=134 channel=113
    5, -5, 2, 4, 7, 0, -2, -4, 5,
    -- filter=134 channel=114
    5, -8, 0, 2, 0, -4, 0, -1, -6,
    -- filter=134 channel=115
    6, 5, 3, 5, -5, -5, 4, 3, 0,
    -- filter=134 channel=116
    1, 0, -5, 0, -2, -13, -4, 0, 2,
    -- filter=134 channel=117
    7, -4, -4, 6, -5, -6, 2, 0, 0,
    -- filter=134 channel=118
    -7, -5, 7, -5, -5, -1, 6, 0, -4,
    -- filter=134 channel=119
    10, -5, -1, 4, 0, -1, -6, 2, -2,
    -- filter=134 channel=120
    -3, -5, -1, 8, -5, -12, -7, -9, 14,
    -- filter=134 channel=121
    5, 9, 9, -3, 3, 0, 5, 5, 3,
    -- filter=134 channel=122
    23, 17, -1, 3, 9, 7, -8, -13, -1,
    -- filter=134 channel=123
    0, 1, 2, -2, -5, 0, 3, 8, 5,
    -- filter=134 channel=124
    -7, -11, 1, 5, 2, -7, 6, 11, 3,
    -- filter=134 channel=125
    0, 3, 2, 0, 1, -8, -10, -4, 12,
    -- filter=134 channel=126
    3, 3, 5, 5, -3, 2, -3, 0, -7,
    -- filter=134 channel=127
    -5, -5, -1, 3, 1, 1, 0, -3, 0,
    -- filter=135 channel=0
    -4, -2, -4, -7, 3, 0, -4, 1, -3,
    -- filter=135 channel=1
    0, -2, 2, -1, 2, 6, -7, -7, -6,
    -- filter=135 channel=2
    -4, -5, 0, 2, -5, -2, -1, 0, 1,
    -- filter=135 channel=3
    1, -1, -3, 0, 4, -6, 2, -4, -5,
    -- filter=135 channel=4
    -3, 0, 0, -4, 0, 3, 7, 4, 6,
    -- filter=135 channel=5
    0, 7, 3, -4, -5, -2, 0, -2, -6,
    -- filter=135 channel=6
    1, 5, -6, 4, 2, 7, 0, -1, -2,
    -- filter=135 channel=7
    -7, 5, 4, 6, -1, -6, 1, 0, 0,
    -- filter=135 channel=8
    -4, -1, 3, -5, 0, 0, -6, 0, 4,
    -- filter=135 channel=9
    -2, 4, -6, -3, 7, 3, -4, 7, 4,
    -- filter=135 channel=10
    -7, -5, -2, -7, -5, -5, -5, 0, 1,
    -- filter=135 channel=11
    0, 4, -7, -3, 2, 4, 1, -7, -2,
    -- filter=135 channel=12
    -4, 4, -6, 7, 7, 1, 0, 1, 0,
    -- filter=135 channel=13
    0, -3, 6, -6, -3, -2, 0, -1, 0,
    -- filter=135 channel=14
    6, 0, -6, 4, 3, 4, 3, 0, 0,
    -- filter=135 channel=15
    5, -4, 6, -5, -6, -4, 5, 0, 2,
    -- filter=135 channel=16
    6, -1, 5, 0, 0, 0, 0, -1, -1,
    -- filter=135 channel=17
    -1, 3, -2, 3, -1, 2, -3, -6, -5,
    -- filter=135 channel=18
    0, 5, 4, 5, 5, 2, -2, 1, 6,
    -- filter=135 channel=19
    3, 4, 6, -2, -3, -2, 4, -1, -2,
    -- filter=135 channel=20
    0, -5, -4, 0, 6, -4, -6, -1, -5,
    -- filter=135 channel=21
    5, 4, 4, 1, 5, 1, 0, -7, 4,
    -- filter=135 channel=22
    -1, -1, -6, 4, -6, 0, 3, 4, 0,
    -- filter=135 channel=23
    0, -6, 1, 0, -3, -7, 0, -3, -1,
    -- filter=135 channel=24
    3, 6, -5, -2, 3, 3, -6, -2, 0,
    -- filter=135 channel=25
    -4, 0, 6, -6, 1, -5, 1, -5, -3,
    -- filter=135 channel=26
    -1, -7, 5, 2, -1, 3, 3, 2, -7,
    -- filter=135 channel=27
    4, -7, -5, -6, 3, -1, -4, 2, -3,
    -- filter=135 channel=28
    -3, 1, 5, 2, 1, 7, 4, 4, 2,
    -- filter=135 channel=29
    -4, -7, -3, -3, 6, 5, -6, -3, -7,
    -- filter=135 channel=30
    -6, -4, 2, 0, 4, 3, 6, -1, 5,
    -- filter=135 channel=31
    -4, -3, -3, -5, 2, 6, 0, -6, 2,
    -- filter=135 channel=32
    -1, -1, 2, 1, 5, -5, 6, 6, 0,
    -- filter=135 channel=33
    1, -6, -5, -7, -5, -5, -4, -5, -1,
    -- filter=135 channel=34
    -1, -3, 3, -6, -6, -4, -6, 4, 4,
    -- filter=135 channel=35
    2, 7, 0, 6, -3, 0, -1, 7, 7,
    -- filter=135 channel=36
    -5, -7, -3, -3, -6, -4, 3, 5, -2,
    -- filter=135 channel=37
    -2, 6, -1, -5, 6, -3, -1, 0, 6,
    -- filter=135 channel=38
    4, -6, 1, 0, 1, 6, 0, 0, -5,
    -- filter=135 channel=39
    0, -1, -7, 7, -3, 2, -5, 1, 0,
    -- filter=135 channel=40
    -1, 6, 6, -1, 2, 1, 0, -6, 0,
    -- filter=135 channel=41
    5, 0, 6, 2, 2, -2, 0, -5, -4,
    -- filter=135 channel=42
    5, -1, 0, 0, 0, 6, 0, 3, 1,
    -- filter=135 channel=43
    4, -5, -6, 7, 6, -2, -6, 5, 5,
    -- filter=135 channel=44
    3, -3, -7, 5, -3, 4, -1, -3, -5,
    -- filter=135 channel=45
    1, -6, -4, 5, 5, -1, 1, 0, -5,
    -- filter=135 channel=46
    -4, -4, 5, -1, -2, -4, 0, 5, 0,
    -- filter=135 channel=47
    0, 0, 1, -6, 3, -2, -6, 3, -5,
    -- filter=135 channel=48
    -2, -5, 2, -4, 0, 0, -5, -7, 2,
    -- filter=135 channel=49
    5, -3, -4, -3, 3, -4, 4, 2, 2,
    -- filter=135 channel=50
    0, -3, 0, 0, 3, 3, 1, 1, -6,
    -- filter=135 channel=51
    -4, -2, 4, 0, -1, 6, -3, 0, 0,
    -- filter=135 channel=52
    -6, 3, 6, 6, -1, -4, 7, 1, 4,
    -- filter=135 channel=53
    -1, 1, 7, -5, 1, -1, 6, -5, -2,
    -- filter=135 channel=54
    1, -4, 4, -7, 3, 6, -1, 3, 5,
    -- filter=135 channel=55
    -5, 5, 7, -6, 0, 4, -6, -6, 0,
    -- filter=135 channel=56
    1, 2, -2, -2, -3, 5, -6, 2, -4,
    -- filter=135 channel=57
    -6, -3, 3, -2, 2, 0, -5, 3, -1,
    -- filter=135 channel=58
    5, -6, 0, 3, -2, 3, 4, -1, 1,
    -- filter=135 channel=59
    -6, 0, -6, 2, -6, 4, 2, 3, 1,
    -- filter=135 channel=60
    3, -2, -3, -1, 1, 1, 6, -1, 3,
    -- filter=135 channel=61
    0, 4, 0, -3, 4, -3, 4, 7, -1,
    -- filter=135 channel=62
    -7, 6, -2, -5, -4, 3, 5, -5, -1,
    -- filter=135 channel=63
    2, -5, -5, 4, -2, -6, -2, 0, -3,
    -- filter=135 channel=64
    0, -5, 2, -5, 3, -3, 1, 2, 1,
    -- filter=135 channel=65
    1, -7, 0, 4, 1, 2, 0, 0, -5,
    -- filter=135 channel=66
    0, 6, -2, 6, -3, -4, 5, 3, -5,
    -- filter=135 channel=67
    1, -5, -7, 0, 2, 6, -1, -3, 4,
    -- filter=135 channel=68
    4, -6, -4, 1, 0, -6, -2, 7, -3,
    -- filter=135 channel=69
    7, 2, -4, -4, 7, -2, -5, 4, 0,
    -- filter=135 channel=70
    -3, -2, -5, 1, -2, 1, 2, -4, 5,
    -- filter=135 channel=71
    -6, -7, 0, 0, -6, -5, 3, 4, -1,
    -- filter=135 channel=72
    -1, 0, -1, -6, -4, 2, -7, 4, 7,
    -- filter=135 channel=73
    -6, -7, 5, 2, 0, 5, 3, 6, 3,
    -- filter=135 channel=74
    0, -5, 4, 1, -1, -6, 6, -6, -1,
    -- filter=135 channel=75
    2, -7, 0, 5, 1, -2, 0, 5, 5,
    -- filter=135 channel=76
    -5, -5, 2, -7, 0, 5, -1, 0, 0,
    -- filter=135 channel=77
    -3, 3, -5, 3, -4, -3, 5, -3, 1,
    -- filter=135 channel=78
    -7, -5, -6, -4, -6, -7, -5, -2, 1,
    -- filter=135 channel=79
    0, 2, -6, 1, 6, -4, 0, 5, 3,
    -- filter=135 channel=80
    0, 1, -6, -7, 5, 5, 0, 5, -1,
    -- filter=135 channel=81
    3, 2, 1, -2, -1, 6, -5, -3, -1,
    -- filter=135 channel=82
    1, -2, 2, 5, 0, 1, 0, 3, -3,
    -- filter=135 channel=83
    4, 0, 0, 3, 3, -3, 1, 2, -1,
    -- filter=135 channel=84
    -6, 7, -1, 0, 4, -6, -3, 6, -4,
    -- filter=135 channel=85
    0, -4, -7, -6, -5, 6, -2, 5, -5,
    -- filter=135 channel=86
    2, 6, -3, 1, -2, 0, -5, -3, -1,
    -- filter=135 channel=87
    -4, -4, 0, 0, 0, 2, 0, 1, 1,
    -- filter=135 channel=88
    -4, 0, 2, -3, 4, -1, 4, 1, -1,
    -- filter=135 channel=89
    2, 0, 3, -1, -3, -7, 3, -3, 4,
    -- filter=135 channel=90
    -6, -7, -6, -5, -4, 6, 0, 1, -3,
    -- filter=135 channel=91
    2, 5, 5, 5, 4, 4, -6, 5, 4,
    -- filter=135 channel=92
    2, 3, -4, 6, 7, -1, 4, -1, 6,
    -- filter=135 channel=93
    -6, -3, -1, 5, 4, -3, 6, -2, 1,
    -- filter=135 channel=94
    -3, 7, 2, 0, 4, -3, -2, 2, 7,
    -- filter=135 channel=95
    0, 4, 3, 4, 4, -1, -2, -4, -6,
    -- filter=135 channel=96
    -2, 2, 0, -7, 4, -3, -1, -1, -5,
    -- filter=135 channel=97
    3, 4, -4, -3, 5, -1, -5, -1, -2,
    -- filter=135 channel=98
    7, 4, 5, 5, -7, -4, 0, -3, -6,
    -- filter=135 channel=99
    -2, 6, 2, 2, 4, 2, 0, -5, 4,
    -- filter=135 channel=100
    4, -6, 2, 2, -5, -4, 4, -6, 0,
    -- filter=135 channel=101
    1, 7, -7, 3, 0, 3, -7, -4, -2,
    -- filter=135 channel=102
    4, -7, 5, 4, 1, -4, 0, -2, -6,
    -- filter=135 channel=103
    5, 0, 2, 7, -3, 6, -4, 5, -6,
    -- filter=135 channel=104
    1, 4, -1, 5, -4, -7, 1, -5, -4,
    -- filter=135 channel=105
    -4, 4, -2, 0, 1, 4, 3, -1, 0,
    -- filter=135 channel=106
    -4, 7, -6, 3, -2, 0, -4, -7, -3,
    -- filter=135 channel=107
    2, 2, -7, 0, -2, 0, 4, -7, 1,
    -- filter=135 channel=108
    2, 5, -1, -3, -4, -1, 5, 1, 4,
    -- filter=135 channel=109
    2, 4, 4, 1, -5, 2, -1, -5, 1,
    -- filter=135 channel=110
    5, -4, 0, 0, -5, -5, -2, -6, 6,
    -- filter=135 channel=111
    5, 3, -2, 4, -6, -2, 3, 2, -3,
    -- filter=135 channel=112
    6, -6, 4, -3, 4, -2, -5, -7, 4,
    -- filter=135 channel=113
    -4, 3, 2, -2, -5, 6, 5, 4, 4,
    -- filter=135 channel=114
    -2, -2, 4, 1, 0, -3, -5, -1, -1,
    -- filter=135 channel=115
    2, -5, -6, -3, 0, -2, 6, -7, 0,
    -- filter=135 channel=116
    0, 4, 2, -3, -2, -3, 0, 1, 5,
    -- filter=135 channel=117
    4, -3, 3, -4, -2, -4, 1, -2, 0,
    -- filter=135 channel=118
    2, -7, -4, 5, 0, 4, 3, 3, 0,
    -- filter=135 channel=119
    0, 3, 3, -7, -2, -6, -2, -2, 4,
    -- filter=135 channel=120
    6, 7, -2, 1, 3, 4, 3, -2, 3,
    -- filter=135 channel=121
    -2, -6, -1, -6, 6, 4, 0, -2, 1,
    -- filter=135 channel=122
    -5, 0, 1, -1, -3, 1, 1, 0, -4,
    -- filter=135 channel=123
    -6, -3, 1, 0, 5, -5, 1, -2, 1,
    -- filter=135 channel=124
    -5, 3, -1, -3, -1, -7, -3, -4, -6,
    -- filter=135 channel=125
    -2, -1, -2, 3, -3, -2, 3, -6, -1,
    -- filter=135 channel=126
    -3, 0, 6, 2, -5, 0, 0, 2, 0,
    -- filter=135 channel=127
    -6, 0, -2, 0, -1, 3, 2, -7, 7,
    -- filter=136 channel=0
    3, -12, -29, 19, 0, -31, 22, 8, -9,
    -- filter=136 channel=1
    4, -10, -14, 18, -4, -17, 17, 18, -1,
    -- filter=136 channel=2
    1, 1, -2, 2, 0, -3, 0, 3, -6,
    -- filter=136 channel=3
    -1, -10, -9, -5, -8, -10, 11, 7, -7,
    -- filter=136 channel=4
    3, -7, -12, -1, 3, -9, 1, 2, -7,
    -- filter=136 channel=5
    -11, -5, -13, -4, -6, -20, 0, -3, 2,
    -- filter=136 channel=6
    -5, -7, -12, -9, 0, 0, -3, -2, -3,
    -- filter=136 channel=7
    0, 3, 3, -5, -3, -7, 3, -2, -4,
    -- filter=136 channel=8
    3, -9, 5, -2, 2, 1, -4, 4, 2,
    -- filter=136 channel=9
    0, 3, 1, 1, 1, 2, -1, -4, 4,
    -- filter=136 channel=10
    -15, -5, 3, -19, -14, 10, -8, -6, 8,
    -- filter=136 channel=11
    -6, -2, 8, -9, 5, 12, -3, 0, 8,
    -- filter=136 channel=12
    0, -13, 4, -3, -17, 0, -5, -2, 11,
    -- filter=136 channel=13
    -6, -9, 9, -12, 0, 5, 9, 2, 3,
    -- filter=136 channel=14
    -5, -1, -1, -4, 6, 2, 2, 2, 6,
    -- filter=136 channel=15
    0, -8, -7, -7, -2, -12, 5, 1, 0,
    -- filter=136 channel=16
    0, -13, -4, -11, -5, 4, -7, -1, 0,
    -- filter=136 channel=17
    2, -5, -2, 0, -4, -5, -6, -1, -3,
    -- filter=136 channel=18
    -8, -12, -11, -9, -7, -9, 5, 3, -3,
    -- filter=136 channel=19
    5, 4, -5, 6, 0, 1, 1, -3, -5,
    -- filter=136 channel=20
    0, 4, 8, -4, 0, 6, -4, 6, 4,
    -- filter=136 channel=21
    3, -3, 17, -2, 9, 28, -1, 0, 10,
    -- filter=136 channel=22
    -1, -4, -11, 4, 2, -11, 4, -4, -4,
    -- filter=136 channel=23
    -6, 2, 1, -2, 4, 3, 5, -4, 7,
    -- filter=136 channel=24
    -2, 6, -6, 0, 0, -2, -2, -4, 5,
    -- filter=136 channel=25
    -4, -5, -10, 0, -4, 2, 12, 3, -7,
    -- filter=136 channel=26
    1, -4, -2, 4, -8, -1, 3, 2, 6,
    -- filter=136 channel=27
    0, -3, -8, 13, 1, -5, 8, 2, -13,
    -- filter=136 channel=28
    5, 7, 5, 5, -1, 2, 2, 4, -2,
    -- filter=136 channel=29
    -7, -4, 0, -7, -1, -2, -3, -1, -6,
    -- filter=136 channel=30
    8, -4, -16, 0, 3, -6, 6, 9, -3,
    -- filter=136 channel=31
    -12, 8, 25, -20, 9, 25, -10, -6, 13,
    -- filter=136 channel=32
    0, -3, -15, 8, -5, -10, 4, 13, -3,
    -- filter=136 channel=33
    7, -1, -9, 7, -6, -17, 13, 7, -2,
    -- filter=136 channel=34
    -1, -6, 1, -13, -11, -16, 2, -5, -2,
    -- filter=136 channel=35
    0, -3, 4, 0, -3, -4, 1, -5, -3,
    -- filter=136 channel=36
    0, 4, 13, -10, -2, 23, -8, -2, 13,
    -- filter=136 channel=37
    5, -5, -18, 15, 0, -18, 21, 18, 4,
    -- filter=136 channel=38
    1, 0, 1, 3, -8, -4, 7, -5, -1,
    -- filter=136 channel=39
    -3, 3, -3, -2, 2, 3, -3, -5, 9,
    -- filter=136 channel=40
    0, 3, 0, 7, 3, 6, 5, 2, 2,
    -- filter=136 channel=41
    1, -12, -2, -4, -11, -2, -1, -4, -6,
    -- filter=136 channel=42
    3, 5, -5, 9, 1, -4, 4, 5, -2,
    -- filter=136 channel=43
    -5, -10, -4, 0, -10, -15, 9, 0, 1,
    -- filter=136 channel=44
    3, -6, 3, 13, 7, 0, 9, 10, -4,
    -- filter=136 channel=45
    11, 9, -5, 13, 3, 2, 11, 4, 3,
    -- filter=136 channel=46
    -8, 0, 2, -2, -6, -8, 0, -5, -1,
    -- filter=136 channel=47
    0, -2, 4, 8, 0, 9, 1, 4, 7,
    -- filter=136 channel=48
    -4, -1, -1, -1, 11, 4, 11, 8, 0,
    -- filter=136 channel=49
    3, 4, -5, -1, 7, -7, 1, 7, -8,
    -- filter=136 channel=50
    -4, 0, 4, 1, 6, 9, 7, 9, -5,
    -- filter=136 channel=51
    7, -5, 2, 1, -4, 4, 1, -2, -3,
    -- filter=136 channel=52
    1, -9, 9, 0, -8, 2, 0, 3, 0,
    -- filter=136 channel=53
    -5, 2, 7, -11, -5, 9, -6, 1, 6,
    -- filter=136 channel=54
    -6, 3, -4, 4, -5, -3, -5, 0, 4,
    -- filter=136 channel=55
    -9, -5, 8, -17, -13, 14, 2, -1, 7,
    -- filter=136 channel=56
    1, -2, 0, -6, -9, -11, 0, 3, 3,
    -- filter=136 channel=57
    4, 3, 0, 0, 4, -3, 5, 3, 0,
    -- filter=136 channel=58
    -14, -11, -4, 1, 2, -2, -1, -3, 4,
    -- filter=136 channel=59
    -3, 0, -5, -7, -4, 3, 6, 4, 0,
    -- filter=136 channel=60
    0, -1, -2, 2, 6, -4, 3, -5, -4,
    -- filter=136 channel=61
    -3, -1, 6, -10, 0, 0, -2, -6, 4,
    -- filter=136 channel=62
    1, -1, 0, -3, 1, 5, 0, 4, 0,
    -- filter=136 channel=63
    -1, -7, 1, -4, 3, -7, 0, -5, 0,
    -- filter=136 channel=64
    0, 0, 2, -7, -4, 11, -8, -6, 0,
    -- filter=136 channel=65
    0, -6, -1, 0, 6, 5, -1, 5, -4,
    -- filter=136 channel=66
    4, -9, 0, 0, -13, 4, -7, 1, -2,
    -- filter=136 channel=67
    0, -2, 0, 1, 1, 5, 4, -4, 3,
    -- filter=136 channel=68
    -1, -1, -3, 9, 9, 11, -3, 8, 9,
    -- filter=136 channel=69
    -1, 4, -3, -2, -4, 7, -4, -1, 1,
    -- filter=136 channel=70
    7, 2, -2, 2, 5, -1, 5, 1, 3,
    -- filter=136 channel=71
    -3, 5, 7, 5, -6, 0, 4, -3, 2,
    -- filter=136 channel=72
    -8, 2, 6, -4, -3, 27, -3, -10, 2,
    -- filter=136 channel=73
    0, -5, -4, 3, 4, 0, 8, 7, 3,
    -- filter=136 channel=74
    -7, -7, 0, 4, 8, 0, 9, 6, 5,
    -- filter=136 channel=75
    -3, -4, -16, 1, -11, -29, 6, 4, -10,
    -- filter=136 channel=76
    8, -2, 7, -8, 4, 11, 7, 9, 3,
    -- filter=136 channel=77
    -5, -4, 1, 6, 6, -5, -6, 6, 2,
    -- filter=136 channel=78
    -10, -10, -1, -5, -5, 3, 4, -7, -3,
    -- filter=136 channel=79
    1, -4, -22, -2, -2, -15, 20, 12, -9,
    -- filter=136 channel=80
    -3, -5, 16, 5, 0, 21, -1, 3, 12,
    -- filter=136 channel=81
    -5, 0, 2, 5, -1, 2, -1, -2, 5,
    -- filter=136 channel=82
    1, -7, -4, 0, 2, 2, 4, 7, 5,
    -- filter=136 channel=83
    2, 3, 4, 7, 0, 12, -1, 3, -2,
    -- filter=136 channel=84
    -1, -3, -2, 7, 0, -12, 9, 5, -1,
    -- filter=136 channel=85
    -5, 3, 5, 0, 2, 6, -3, 0, -2,
    -- filter=136 channel=86
    -1, -10, -3, -2, -5, -8, 0, 1, -6,
    -- filter=136 channel=87
    -8, 1, -2, 1, -4, -7, 0, 1, -4,
    -- filter=136 channel=88
    -6, -5, 10, -8, 10, 17, -16, -14, 14,
    -- filter=136 channel=89
    -1, -11, 2, -6, -9, 10, 0, -4, 3,
    -- filter=136 channel=90
    -6, 4, 12, -10, 0, 18, -3, -7, 4,
    -- filter=136 channel=91
    4, 5, -12, 6, 1, -7, 17, 2, 4,
    -- filter=136 channel=92
    0, 0, -2, -8, -3, -4, -3, -2, 6,
    -- filter=136 channel=93
    2, 0, -4, 12, 5, 0, 0, -1, -9,
    -- filter=136 channel=94
    3, 2, 2, -1, 2, -2, 0, 1, 0,
    -- filter=136 channel=95
    0, 4, -5, -4, 2, -1, 0, -7, 5,
    -- filter=136 channel=96
    5, 6, 1, 3, 7, -5, -1, -3, 0,
    -- filter=136 channel=97
    0, -5, -7, -6, 2, 3, 7, 0, -2,
    -- filter=136 channel=98
    0, -3, -1, -3, -9, 0, 7, -6, 0,
    -- filter=136 channel=99
    -10, -6, 16, -19, -6, 22, -19, -10, 1,
    -- filter=136 channel=100
    -1, -4, -2, -11, -8, -4, -12, -2, 2,
    -- filter=136 channel=101
    5, -8, -5, -5, 0, 1, 5, 7, -6,
    -- filter=136 channel=102
    3, -5, 1, 7, 5, -5, 5, -2, 2,
    -- filter=136 channel=103
    -4, -6, 6, -1, -1, 13, 10, 8, 7,
    -- filter=136 channel=104
    -2, 0, 12, -4, 7, 25, -13, -8, 4,
    -- filter=136 channel=105
    3, 1, -8, -9, -6, -3, -7, -2, 0,
    -- filter=136 channel=106
    -1, 9, 3, 0, 7, -3, -3, 3, 6,
    -- filter=136 channel=107
    -1, -7, -14, 8, -5, -16, 7, 6, -8,
    -- filter=136 channel=108
    3, 0, -10, -10, 4, -7, -8, -4, -5,
    -- filter=136 channel=109
    -9, -14, -2, -6, -4, -4, 5, 4, 2,
    -- filter=136 channel=110
    -4, -6, 4, -8, -1, 15, -12, -7, 2,
    -- filter=136 channel=111
    -7, -8, -5, -7, 4, -7, 0, 1, -2,
    -- filter=136 channel=112
    2, -3, -3, 2, 0, -9, 8, -4, 4,
    -- filter=136 channel=113
    2, -9, -2, 0, -13, 0, 1, -8, 2,
    -- filter=136 channel=114
    -1, -15, -30, 14, -4, -30, 10, 2, -23,
    -- filter=136 channel=115
    2, -6, -3, 0, -7, 3, 0, -5, 3,
    -- filter=136 channel=116
    -8, -2, 5, -8, 1, 8, -3, -5, -1,
    -- filter=136 channel=117
    9, 0, -2, 6, -4, 6, -4, 2, 5,
    -- filter=136 channel=118
    0, -4, 0, 2, -5, -3, -6, -5, -1,
    -- filter=136 channel=119
    0, -3, -4, -10, -12, -7, -14, -11, -3,
    -- filter=136 channel=120
    8, 0, 0, -2, 4, 5, 14, 12, -7,
    -- filter=136 channel=121
    -13, -6, 4, -9, -13, 6, -3, -4, 3,
    -- filter=136 channel=122
    -7, 1, 13, -5, 7, 23, -3, 0, 11,
    -- filter=136 channel=123
    -8, -1, -2, -2, 0, 3, -8, -2, 10,
    -- filter=136 channel=124
    -3, 2, 1, 4, 3, -3, 1, -7, -9,
    -- filter=136 channel=125
    -14, -11, 14, -8, -8, 20, -2, -7, 5,
    -- filter=136 channel=126
    -6, -11, -4, -10, -10, -2, 7, 6, -6,
    -- filter=136 channel=127
    -1, -3, -2, -2, -9, -7, 0, -5, 7,
    -- filter=137 channel=0
    -5, 1, 4, 3, 7, -10, 6, 3, -11,
    -- filter=137 channel=1
    -4, 0, -3, -7, -4, -11, -2, 6, -4,
    -- filter=137 channel=2
    -6, -2, 0, -3, 0, 0, -5, -4, 0,
    -- filter=137 channel=3
    -12, -15, 3, -2, 3, 2, -9, 2, -17,
    -- filter=137 channel=4
    0, 0, -14, 3, -8, -13, 4, -10, -9,
    -- filter=137 channel=5
    3, 2, 6, -8, -1, 0, 7, -5, -1,
    -- filter=137 channel=6
    0, 0, -5, 2, 11, -4, 3, 11, -11,
    -- filter=137 channel=7
    -4, -1, -2, -4, 4, 0, -4, -4, 6,
    -- filter=137 channel=8
    3, 4, 2, -6, 3, 0, 4, 0, -1,
    -- filter=137 channel=9
    -1, -5, -6, 5, -6, -3, -1, 3, -4,
    -- filter=137 channel=10
    -5, -5, 2, -5, 8, 6, -4, 0, -1,
    -- filter=137 channel=11
    -2, 0, 3, 6, 17, -12, 5, 0, -15,
    -- filter=137 channel=12
    0, 1, -1, 5, 11, 5, -1, 3, -5,
    -- filter=137 channel=13
    -2, 7, -1, -12, 20, -2, -4, 9, -2,
    -- filter=137 channel=14
    -4, -7, -6, -2, 0, -4, -4, 2, 3,
    -- filter=137 channel=15
    -10, 5, 0, -5, 17, -8, 7, 16, -9,
    -- filter=137 channel=16
    6, 1, 2, 0, -8, 12, -6, -8, 4,
    -- filter=137 channel=17
    2, -1, 6, -6, 7, 2, -3, -6, -4,
    -- filter=137 channel=18
    -6, 9, 0, -6, 30, -21, 8, 25, -27,
    -- filter=137 channel=19
    -6, -5, -1, 4, 0, 5, 2, 3, 1,
    -- filter=137 channel=20
    -16, 9, -5, -5, 21, -7, 3, 12, -11,
    -- filter=137 channel=21
    11, -5, 6, 5, -3, 11, 0, -5, 16,
    -- filter=137 channel=22
    -6, 1, -1, 4, 6, -1, 3, 7, 2,
    -- filter=137 channel=23
    -6, 14, -11, 0, 15, -10, 2, 6, -9,
    -- filter=137 channel=24
    5, 7, -3, -6, 0, -2, 6, -2, -5,
    -- filter=137 channel=25
    2, 3, -1, -7, 5, -8, 3, 7, -2,
    -- filter=137 channel=26
    1, 3, -2, 2, -5, 9, -1, 1, 6,
    -- filter=137 channel=27
    -8, 19, -8, 2, -1, -12, 4, -2, 1,
    -- filter=137 channel=28
    3, 2, 7, 0, -4, -2, 5, 0, -1,
    -- filter=137 channel=29
    -12, -1, -7, -6, 21, -11, 3, 7, -13,
    -- filter=137 channel=30
    -5, 4, 4, 3, 2, -2, 8, 1, 1,
    -- filter=137 channel=31
    -3, 5, -6, -4, -7, 3, -13, -15, 0,
    -- filter=137 channel=32
    -8, 15, -4, 0, 13, -20, 3, 14, -20,
    -- filter=137 channel=33
    2, -3, 10, -2, 11, -2, 4, 1, -8,
    -- filter=137 channel=34
    -3, 4, 4, -3, 0, 8, 4, 1, 13,
    -- filter=137 channel=35
    6, -4, 4, -7, 7, 0, 0, 5, 4,
    -- filter=137 channel=36
    -1, 0, -9, -6, 1, 4, 0, -6, 10,
    -- filter=137 channel=37
    0, 1, -6, -1, -9, -10, 10, -5, -1,
    -- filter=137 channel=38
    -9, 2, 6, 3, 4, -7, -4, -3, -7,
    -- filter=137 channel=39
    0, 9, 5, -7, 9, -4, 4, 11, -4,
    -- filter=137 channel=40
    3, -1, 0, 5, 5, -4, 0, 4, -3,
    -- filter=137 channel=41
    -4, -7, 11, 2, 17, 12, 5, 31, 10,
    -- filter=137 channel=42
    10, -1, 4, 0, -10, -6, 3, -1, -8,
    -- filter=137 channel=43
    0, 4, 6, -7, 10, -11, -8, 11, -11,
    -- filter=137 channel=44
    3, 3, 2, 6, 0, -5, 0, -9, 6,
    -- filter=137 channel=45
    0, -2, 0, 0, 5, 4, -2, 5, 4,
    -- filter=137 channel=46
    2, -2, 2, -4, 4, 5, 1, 3, 6,
    -- filter=137 channel=47
    6, 2, 4, 0, -12, 3, 5, -14, 15,
    -- filter=137 channel=48
    6, 7, 0, 3, -14, -9, 4, -11, 5,
    -- filter=137 channel=49
    -6, 1, -10, 1, 3, -7, 2, -3, -15,
    -- filter=137 channel=50
    2, 4, -1, 9, -9, -2, -3, -6, -3,
    -- filter=137 channel=51
    1, -4, 7, 0, -2, 6, 0, 4, -3,
    -- filter=137 channel=52
    -3, 0, -4, 0, 6, 6, -10, -1, 1,
    -- filter=137 channel=53
    -12, 10, 4, -7, 10, -1, 4, 3, -1,
    -- filter=137 channel=54
    -2, 0, -6, 3, 4, 1, 3, 6, 1,
    -- filter=137 channel=55
    -6, 13, 0, -9, 14, -4, -5, 16, -18,
    -- filter=137 channel=56
    -7, 6, 1, 7, 6, 1, 7, 8, 10,
    -- filter=137 channel=57
    -1, -5, -3, -4, -2, 4, 2, -6, 6,
    -- filter=137 channel=58
    6, -8, 7, -4, -4, 9, 4, -6, 0,
    -- filter=137 channel=59
    -2, 6, 5, 2, 8, 4, -1, 6, 2,
    -- filter=137 channel=60
    -1, -3, -5, 3, -2, 2, 4, -4, 2,
    -- filter=137 channel=61
    -2, 0, -6, 4, 1, -5, -5, -4, 8,
    -- filter=137 channel=62
    6, 1, 7, 5, 5, -4, -2, 0, -4,
    -- filter=137 channel=63
    1, 2, 0, 1, -6, 7, -2, -2, 0,
    -- filter=137 channel=64
    3, -6, 1, -5, 6, -2, -6, 4, 4,
    -- filter=137 channel=65
    -1, 0, -4, 3, -4, 0, 4, 2, 2,
    -- filter=137 channel=66
    -2, 4, 1, -9, 20, -5, -2, 14, 7,
    -- filter=137 channel=67
    2, -2, -3, -6, -6, 0, 0, 6, -4,
    -- filter=137 channel=68
    -4, -3, -9, -3, 3, -9, -5, -1, -1,
    -- filter=137 channel=69
    0, 7, -3, -5, 8, 4, -2, -1, -4,
    -- filter=137 channel=70
    -4, 9, -12, 9, 6, -9, 9, 0, 0,
    -- filter=137 channel=71
    -6, -3, 3, -3, -7, -1, 0, -6, -2,
    -- filter=137 channel=72
    -4, 0, 8, -3, 2, -6, 6, -5, 9,
    -- filter=137 channel=73
    -1, 3, -7, -4, 9, -17, -1, 3, -5,
    -- filter=137 channel=74
    -6, 13, 1, 9, -1, -4, 0, -1, 0,
    -- filter=137 channel=75
    -5, -10, 8, -11, 2, -9, 4, 1, -7,
    -- filter=137 channel=76
    -15, 4, -1, -8, 25, -14, -6, 14, -5,
    -- filter=137 channel=77
    2, 2, 6, -7, -3, -7, -5, 4, 0,
    -- filter=137 channel=78
    3, -3, 3, 0, -4, -7, 4, -3, 4,
    -- filter=137 channel=79
    -6, 8, -2, -5, 29, -24, 8, 23, -27,
    -- filter=137 channel=80
    0, 4, 0, -7, -9, -7, 4, -2, 4,
    -- filter=137 channel=81
    1, 0, 3, -4, -3, 0, 0, 0, 0,
    -- filter=137 channel=82
    -5, 0, 6, -6, -3, 5, 0, -1, -1,
    -- filter=137 channel=83
    1, -1, -6, 1, -11, 6, 2, 0, -3,
    -- filter=137 channel=84
    -12, 12, -5, -6, 10, -13, 2, 5, -6,
    -- filter=137 channel=85
    3, 3, -5, 3, -2, 5, 1, 5, 2,
    -- filter=137 channel=86
    3, 2, 6, 1, 3, -6, -8, 4, 1,
    -- filter=137 channel=87
    -1, 14, 3, -3, 1, 0, -6, 5, -7,
    -- filter=137 channel=88
    3, 7, -9, -8, -1, 9, -1, -8, 11,
    -- filter=137 channel=89
    -3, 0, 0, -2, 23, -10, -3, 13, -11,
    -- filter=137 channel=90
    4, 8, -4, -2, 2, 10, -2, -15, 9,
    -- filter=137 channel=91
    -4, 8, -2, 0, 9, -17, 7, 1, -12,
    -- filter=137 channel=92
    4, 7, -7, 3, -4, 3, 1, 0, 5,
    -- filter=137 channel=93
    2, -2, -3, 0, -5, -4, 9, -13, 8,
    -- filter=137 channel=94
    -7, 0, 5, -1, -2, -6, 1, -2, 5,
    -- filter=137 channel=95
    6, 2, -4, -2, 3, 2, 5, 5, -3,
    -- filter=137 channel=96
    7, -3, -4, 0, 5, 1, 5, -1, 4,
    -- filter=137 channel=97
    -1, -10, -1, -2, 1, 2, -1, -5, -7,
    -- filter=137 channel=98
    0, 1, 0, 4, 2, -8, 1, 0, -1,
    -- filter=137 channel=99
    -16, 11, -6, -8, 7, -14, 0, 0, 5,
    -- filter=137 channel=100
    4, 2, 0, 4, 0, 6, 0, 2, 7,
    -- filter=137 channel=101
    -11, -2, -7, 1, -9, -10, 6, 1, -6,
    -- filter=137 channel=102
    3, -7, -6, -4, -4, 5, -6, 6, 0,
    -- filter=137 channel=103
    4, 0, 12, -3, -9, 3, -5, -15, 6,
    -- filter=137 channel=104
    -1, -3, -3, 6, -13, 4, -6, -13, 11,
    -- filter=137 channel=105
    -15, 8, 6, -1, 5, -3, 2, 14, -6,
    -- filter=137 channel=106
    -2, 1, 7, -1, 1, -3, 0, 0, 0,
    -- filter=137 channel=107
    -2, 11, -12, -8, 12, -15, 6, 5, -15,
    -- filter=137 channel=108
    5, 4, -1, 2, 2, 2, 0, 12, -4,
    -- filter=137 channel=109
    -13, 8, -9, 7, 5, -7, 14, 3, -3,
    -- filter=137 channel=110
    0, 0, 4, -4, -5, -1, -6, -1, 6,
    -- filter=137 channel=111
    3, 2, -4, -5, 5, 4, 4, 7, 6,
    -- filter=137 channel=112
    2, 12, 0, 3, 2, -1, -5, -3, 5,
    -- filter=137 channel=113
    3, -6, 11, -7, 3, -5, 1, 2, -1,
    -- filter=137 channel=114
    -17, 19, -3, -2, 20, -29, 3, 22, -25,
    -- filter=137 channel=115
    2, -1, 4, -2, 3, -6, -5, 3, 0,
    -- filter=137 channel=116
    -4, 13, 4, 2, 1, -8, 11, 2, -3,
    -- filter=137 channel=117
    -6, -2, -4, 0, 0, -1, 5, 4, 7,
    -- filter=137 channel=118
    0, 2, -3, 5, 0, -4, -4, 2, 6,
    -- filter=137 channel=119
    0, 7, 8, -1, -2, 16, -3, 10, 13,
    -- filter=137 channel=120
    -17, 12, -20, 7, 3, -19, 10, 1, 0,
    -- filter=137 channel=121
    0, 0, 2, 0, 14, -1, 0, 4, -3,
    -- filter=137 channel=122
    8, -9, 17, 0, -13, 18, -10, -16, 31,
    -- filter=137 channel=123
    -2, -3, -6, -3, -1, -3, 2, -3, 4,
    -- filter=137 channel=124
    -1, 6, -4, -7, 0, -11, 2, 6, -6,
    -- filter=137 channel=125
    -4, 8, 3, -6, -4, -4, 4, -4, -3,
    -- filter=137 channel=126
    0, -8, 6, -10, 7, 0, 0, 21, -7,
    -- filter=137 channel=127
    -3, 4, 7, 1, 0, 7, -1, 10, 7,
    -- filter=138 channel=0
    -17, 0, -9, -9, 2, 1, 4, 8, 0,
    -- filter=138 channel=1
    -9, 6, -1, -14, 12, 6, -7, 7, 2,
    -- filter=138 channel=2
    6, 5, -8, 1, 2, 1, 4, 1, 6,
    -- filter=138 channel=3
    1, 2, 2, -10, 6, -10, 3, 0, 1,
    -- filter=138 channel=4
    -2, 0, -2, -5, 1, 7, 0, -5, 6,
    -- filter=138 channel=5
    -3, -3, 5, 8, -1, 6, -1, -2, 6,
    -- filter=138 channel=6
    2, 13, 3, -6, 4, -2, 5, 0, -2,
    -- filter=138 channel=7
    -2, -1, 6, 4, -1, 3, 0, 0, -7,
    -- filter=138 channel=8
    1, -2, -9, 3, -1, 2, -8, 0, 3,
    -- filter=138 channel=9
    5, -8, -5, 1, -1, -11, -4, 1, -5,
    -- filter=138 channel=10
    -1, 2, -3, 2, 9, -1, 0, 4, -6,
    -- filter=138 channel=11
    0, 2, -4, -5, 7, -1, 0, 2, -6,
    -- filter=138 channel=12
    4, 14, 1, 0, 8, -4, -1, 5, 0,
    -- filter=138 channel=13
    2, 10, -12, 3, 15, -4, -2, 5, -5,
    -- filter=138 channel=14
    -2, -5, 2, 2, 7, 0, -4, -3, 0,
    -- filter=138 channel=15
    0, 2, -4, -3, 12, -8, -4, 0, 0,
    -- filter=138 channel=16
    4, 4, -3, 0, 0, -5, 1, 3, 3,
    -- filter=138 channel=17
    -2, -5, 2, -6, 0, -6, 6, 4, -2,
    -- filter=138 channel=18
    -7, 13, -12, -5, 23, -15, -5, 0, -5,
    -- filter=138 channel=19
    -3, -6, 2, 1, 6, 1, 6, -4, -3,
    -- filter=138 channel=20
    8, 8, 3, -4, 0, 4, 1, -9, -4,
    -- filter=138 channel=21
    8, 3, -6, 8, -8, 3, 6, 1, 6,
    -- filter=138 channel=22
    -8, -5, -9, 6, -1, 4, -7, 1, -7,
    -- filter=138 channel=23
    6, -11, -24, 8, -6, -23, -7, 0, -17,
    -- filter=138 channel=24
    5, -1, 0, -1, -2, 6, -6, 6, 0,
    -- filter=138 channel=25
    2, 10, -20, 2, 12, -16, 7, -3, -1,
    -- filter=138 channel=26
    0, -4, 4, -7, 1, 1, -5, -5, 3,
    -- filter=138 channel=27
    6, 0, -38, 19, 0, -17, 3, -1, -4,
    -- filter=138 channel=28
    6, -5, -3, 3, -4, -5, 5, -3, 7,
    -- filter=138 channel=29
    8, 19, 10, 5, -1, -8, -3, -7, 9,
    -- filter=138 channel=30
    0, 1, -15, 6, -7, -9, 5, 5, 7,
    -- filter=138 channel=31
    13, -7, -29, 24, 1, -13, 10, 2, -1,
    -- filter=138 channel=32
    5, 0, -18, 6, 13, -21, 0, -6, -10,
    -- filter=138 channel=33
    0, 1, -18, 0, 14, -19, 3, -1, -3,
    -- filter=138 channel=34
    5, 2, -5, 6, -3, -4, 2, -5, -9,
    -- filter=138 channel=35
    -3, 5, -5, -2, 5, -3, 2, 0, 3,
    -- filter=138 channel=36
    6, 9, 7, -4, -9, 1, -5, 0, 10,
    -- filter=138 channel=37
    -6, -2, -3, -7, -1, 8, 4, -5, 3,
    -- filter=138 channel=38
    4, 3, -4, 5, 2, -8, 8, 5, -8,
    -- filter=138 channel=39
    4, 6, 5, -4, 0, -7, -5, -6, 0,
    -- filter=138 channel=40
    1, 0, -7, 5, 2, -7, 1, 3, 0,
    -- filter=138 channel=41
    9, 16, 18, -3, 27, -1, -7, 12, 4,
    -- filter=138 channel=42
    7, 2, -8, 5, -1, -3, -1, 3, 2,
    -- filter=138 channel=43
    -8, 0, -5, -5, 9, 6, -4, -5, -9,
    -- filter=138 channel=44
    -3, -9, -16, 12, -12, -6, 12, -6, 3,
    -- filter=138 channel=45
    -3, 5, 0, -6, 4, 6, -6, 6, 6,
    -- filter=138 channel=46
    0, 5, 5, 2, 6, 6, 0, -7, 1,
    -- filter=138 channel=47
    -6, -2, -14, 8, 1, -6, 15, -4, 3,
    -- filter=138 channel=48
    9, 7, -19, -1, -6, -13, 6, -5, 7,
    -- filter=138 channel=49
    2, 8, -7, 1, 4, -7, -1, 3, 9,
    -- filter=138 channel=50
    2, -7, -23, 10, -5, -13, -3, -6, -6,
    -- filter=138 channel=51
    1, -1, 2, -2, -2, 4, 4, 0, -5,
    -- filter=138 channel=52
    -6, 5, -4, 6, -3, -1, -11, -10, -1,
    -- filter=138 channel=53
    7, 2, 2, 6, -5, -4, -9, 2, -4,
    -- filter=138 channel=54
    4, -5, -5, -6, -2, 3, 6, 0, -1,
    -- filter=138 channel=55
    6, 0, -12, 0, 5, -20, -12, -5, -2,
    -- filter=138 channel=56
    -2, 8, -9, -4, 0, -1, -8, -2, -6,
    -- filter=138 channel=57
    -3, 0, 1, 3, 4, 3, -2, 2, -3,
    -- filter=138 channel=58
    3, 2, 1, -1, 1, 3, -6, -3, 2,
    -- filter=138 channel=59
    5, -1, -12, 1, 6, -11, 9, 0, -9,
    -- filter=138 channel=60
    2, 1, 5, 0, -4, -3, -4, 5, 3,
    -- filter=138 channel=61
    8, 6, -2, 7, -7, 4, 0, -2, 6,
    -- filter=138 channel=62
    1, 4, -2, -3, 4, -3, 0, -6, -3,
    -- filter=138 channel=63
    -5, 7, -1, 0, 0, 9, -5, -1, 10,
    -- filter=138 channel=64
    0, 8, 5, -4, 0, 6, 0, 2, -2,
    -- filter=138 channel=65
    -4, 2, -6, 0, -4, -5, 5, 5, 3,
    -- filter=138 channel=66
    9, 3, 9, 0, 10, -5, -4, 0, -4,
    -- filter=138 channel=67
    -4, -6, 0, 1, -6, -4, -4, 2, 0,
    -- filter=138 channel=68
    1, -3, 5, 2, -5, -4, 5, 0, 4,
    -- filter=138 channel=69
    4, 2, 5, 0, -1, 5, -5, -4, 2,
    -- filter=138 channel=70
    -3, -15, -16, 10, -14, -10, -6, 0, -15,
    -- filter=138 channel=71
    -2, 1, 3, -6, -6, 5, -4, 1, -2,
    -- filter=138 channel=72
    2, 10, -13, 14, -2, -6, 5, 0, -6,
    -- filter=138 channel=73
    7, 12, -13, -3, 8, -3, -7, -7, 4,
    -- filter=138 channel=74
    6, -13, -14, 8, -9, -11, -8, 1, -5,
    -- filter=138 channel=75
    -3, -10, 4, 0, 18, 0, 8, -1, -9,
    -- filter=138 channel=76
    5, 4, 7, 4, 15, -2, -10, -2, -4,
    -- filter=138 channel=77
    -2, 0, 2, 2, 2, -4, 4, 1, -3,
    -- filter=138 channel=78
    2, -6, 0, 2, -4, 5, -3, 0, 5,
    -- filter=138 channel=79
    2, 3, -24, 0, 16, -14, -5, 2, -15,
    -- filter=138 channel=80
    4, 4, -19, 18, 13, -15, 14, -2, 5,
    -- filter=138 channel=81
    1, 3, 4, -3, 0, -6, 3, 5, 4,
    -- filter=138 channel=82
    2, -8, -2, 0, -6, 1, 5, 0, -5,
    -- filter=138 channel=83
    10, -2, 1, 5, -6, -7, -3, 5, 7,
    -- filter=138 channel=84
    3, 0, -8, -1, 3, -10, 1, 5, 2,
    -- filter=138 channel=85
    -3, 2, 1, 6, 0, 7, 0, 0, -2,
    -- filter=138 channel=86
    3, 2, -3, 6, 2, 4, 7, -1, -2,
    -- filter=138 channel=87
    -1, 9, -3, 5, -4, 0, 0, 4, 0,
    -- filter=138 channel=88
    9, -2, 0, 8, -13, 0, -3, -7, 7,
    -- filter=138 channel=89
    -4, 9, -3, 2, 14, -17, 0, -5, -6,
    -- filter=138 channel=90
    -4, -4, -4, 3, -8, -3, 4, -6, -8,
    -- filter=138 channel=91
    9, -6, -16, 7, -5, -11, -2, 0, 0,
    -- filter=138 channel=92
    3, -6, -9, 0, -7, 0, 5, 5, -1,
    -- filter=138 channel=93
    6, 0, -9, -3, 0, 4, 3, 1, 6,
    -- filter=138 channel=94
    -1, -5, -2, 7, 6, -2, 7, -3, -3,
    -- filter=138 channel=95
    3, 4, 4, -6, 0, -6, -6, 0, 3,
    -- filter=138 channel=96
    4, -2, -6, 2, -3, -7, 0, -3, 3,
    -- filter=138 channel=97
    -4, -11, 2, -2, -6, -3, -6, 3, -7,
    -- filter=138 channel=98
    12, 7, -14, 16, 11, -19, 6, -1, 0,
    -- filter=138 channel=99
    10, -5, -13, 20, -9, -12, 5, -10, -9,
    -- filter=138 channel=100
    -2, -1, -2, 3, -4, 0, -1, -2, 2,
    -- filter=138 channel=101
    4, -3, 1, -10, -3, -2, -4, -4, 11,
    -- filter=138 channel=102
    -3, -6, 1, -3, 6, 3, 0, -4, -2,
    -- filter=138 channel=103
    -6, -5, -16, 7, 0, -2, 16, 2, -7,
    -- filter=138 channel=104
    3, 1, -9, 8, -4, -5, 3, 1, 2,
    -- filter=138 channel=105
    0, 5, 10, -3, 11, 4, -5, -4, 3,
    -- filter=138 channel=106
    2, 0, -1, 2, -1, -4, 4, 0, 0,
    -- filter=138 channel=107
    -3, 11, 0, -1, 7, 0, -1, -2, 4,
    -- filter=138 channel=108
    0, 6, 12, 3, 7, 5, 4, 0, 4,
    -- filter=138 channel=109
    14, 10, -22, 13, 1, -18, -1, 0, -7,
    -- filter=138 channel=110
    -3, -6, -9, 4, 8, 4, 8, 6, -6,
    -- filter=138 channel=111
    3, 9, 5, 6, 3, -3, -7, 5, 2,
    -- filter=138 channel=112
    -1, -7, -14, 11, -7, -4, 0, 3, 0,
    -- filter=138 channel=113
    6, -6, -14, 13, 2, -8, 3, -7, -4,
    -- filter=138 channel=114
    -5, 6, -9, -8, 9, -3, 0, -1, -2,
    -- filter=138 channel=115
    8, -4, 2, -1, 7, 2, 0, -4, -6,
    -- filter=138 channel=116
    8, 11, -10, -1, -1, -8, 4, -6, 8,
    -- filter=138 channel=117
    0, 0, 0, 0, -1, -6, 6, 2, 6,
    -- filter=138 channel=118
    0, 2, 7, -3, 3, -5, -5, 1, 2,
    -- filter=138 channel=119
    0, -1, -2, 8, 0, -10, -2, -4, 2,
    -- filter=138 channel=120
    8, -2, -25, 19, -9, -15, -11, -8, -3,
    -- filter=138 channel=121
    -4, 6, 6, 1, 5, 1, 5, -4, -9,
    -- filter=138 channel=122
    5, 0, -17, 0, -10, 0, 13, 5, -2,
    -- filter=138 channel=123
    -4, 1, -11, 1, 2, -5, 0, 4, -4,
    -- filter=138 channel=124
    -4, 2, 9, -4, 4, 3, 4, 4, -3,
    -- filter=138 channel=125
    11, 7, -11, 13, 0, -6, -3, 6, -7,
    -- filter=138 channel=126
    0, 2, 0, 1, 22, -5, 4, 0, -11,
    -- filter=138 channel=127
    -4, 3, 4, 3, 3, 0, -3, 2, 1,
    -- filter=139 channel=0
    0, -1, -4, 5, 3, 6, 5, 3, 6,
    -- filter=139 channel=1
    -7, 0, -3, 4, 6, 1, -5, 3, 0,
    -- filter=139 channel=2
    -2, 5, 5, -1, -5, -5, -5, 0, 3,
    -- filter=139 channel=3
    -3, 0, 4, -3, -5, -5, -7, -6, -4,
    -- filter=139 channel=4
    -5, 2, 3, -4, -6, 2, 1, -6, 1,
    -- filter=139 channel=5
    0, -5, -6, -7, -5, -6, -3, -3, -6,
    -- filter=139 channel=6
    2, 0, -5, 1, 6, -6, 1, 4, 0,
    -- filter=139 channel=7
    3, 2, -6, 0, -6, 1, 3, 1, 0,
    -- filter=139 channel=8
    0, -2, -6, 2, 0, 1, -1, 0, -4,
    -- filter=139 channel=9
    4, -3, -3, -5, -5, 1, 0, -5, 4,
    -- filter=139 channel=10
    -3, 4, 0, 5, 4, -7, 0, -7, 0,
    -- filter=139 channel=11
    3, -6, -4, 1, 5, -2, -4, 2, 1,
    -- filter=139 channel=12
    2, 0, 4, 6, -4, -2, -5, -5, 3,
    -- filter=139 channel=13
    -7, -6, -6, -5, -4, 6, 0, -4, -4,
    -- filter=139 channel=14
    -7, 5, 0, 2, 0, -1, -4, -3, 1,
    -- filter=139 channel=15
    4, -3, 0, -5, 1, 1, 6, 0, -3,
    -- filter=139 channel=16
    6, 4, 2, 5, -4, -1, -3, 4, -6,
    -- filter=139 channel=17
    5, 3, 6, -2, -5, 2, -1, -4, -5,
    -- filter=139 channel=18
    -7, 0, -4, -5, 2, 6, 0, 0, -1,
    -- filter=139 channel=19
    4, 0, -3, -2, 6, -3, 2, -4, 1,
    -- filter=139 channel=20
    -3, 0, -7, 4, 6, -1, -6, -1, 0,
    -- filter=139 channel=21
    -7, 0, 3, -7, 5, -5, -5, -3, 1,
    -- filter=139 channel=22
    5, -1, 3, 0, 5, 3, -7, 2, 6,
    -- filter=139 channel=23
    -3, 1, 0, 5, 5, 1, 1, 0, 0,
    -- filter=139 channel=24
    3, -3, -4, 2, 2, 3, 1, 0, 1,
    -- filter=139 channel=25
    0, 0, 5, -1, -2, -2, 0, -2, -6,
    -- filter=139 channel=26
    3, -2, -1, 0, -2, 3, 4, 4, 0,
    -- filter=139 channel=27
    7, 4, -3, -6, 2, -2, 1, 3, 5,
    -- filter=139 channel=28
    3, 2, 2, -3, 0, -5, -3, -5, 5,
    -- filter=139 channel=29
    3, -6, -1, -6, 5, 7, 0, 1, 4,
    -- filter=139 channel=30
    -3, -3, -3, 0, 1, 4, 0, -7, -6,
    -- filter=139 channel=31
    3, 3, -1, 5, -3, 0, -2, 6, 0,
    -- filter=139 channel=32
    -5, 2, -6, -1, -6, 3, 5, 6, 1,
    -- filter=139 channel=33
    -5, 4, -3, -2, -6, 3, -6, 1, -5,
    -- filter=139 channel=34
    -3, -3, 0, 0, 4, 0, 6, -6, -7,
    -- filter=139 channel=35
    -3, 7, 5, 5, -4, -7, 0, 5, 0,
    -- filter=139 channel=36
    3, -5, 0, 6, -5, -1, -5, 7, 2,
    -- filter=139 channel=37
    0, -2, 0, 0, -2, 4, -3, -1, -1,
    -- filter=139 channel=38
    -5, 5, -2, -3, 2, -5, -6, -6, 0,
    -- filter=139 channel=39
    6, 1, 4, -5, 7, 0, 6, -5, 0,
    -- filter=139 channel=40
    -4, 2, 5, -6, -3, 4, -1, 0, -1,
    -- filter=139 channel=41
    0, -3, -2, -4, -2, 0, 3, -7, -3,
    -- filter=139 channel=42
    -7, -3, -3, -5, 1, 3, -6, 4, 2,
    -- filter=139 channel=43
    0, 5, -5, -1, 0, 4, -6, -5, 3,
    -- filter=139 channel=44
    5, -3, -3, 2, 6, 0, -1, -4, 0,
    -- filter=139 channel=45
    1, 5, -5, 4, 1, 7, -6, -2, 4,
    -- filter=139 channel=46
    -1, 0, 6, -4, 0, 0, -4, -1, 1,
    -- filter=139 channel=47
    4, 3, -2, -4, -7, -6, 2, 0, -7,
    -- filter=139 channel=48
    3, 1, -1, 6, 1, -2, -3, 0, 3,
    -- filter=139 channel=49
    2, -2, 2, 0, 5, -3, -6, 5, -7,
    -- filter=139 channel=50
    0, -1, 4, 7, 4, 3, -2, -3, 4,
    -- filter=139 channel=51
    0, 5, 1, 5, -4, 3, 0, -6, 3,
    -- filter=139 channel=52
    -5, -6, 0, 6, -3, -7, 1, 3, -2,
    -- filter=139 channel=53
    0, -1, -3, 6, -1, -7, -6, 3, -3,
    -- filter=139 channel=54
    3, 2, 0, 5, 3, -2, -6, 0, 2,
    -- filter=139 channel=55
    -3, -3, 2, -5, -6, -3, -5, -7, 4,
    -- filter=139 channel=56
    -5, 2, 2, -7, -6, -1, 1, -2, 6,
    -- filter=139 channel=57
    -3, -2, 2, 4, 2, 6, -6, 2, 0,
    -- filter=139 channel=58
    -6, -3, -6, 5, 4, -7, -2, -4, -1,
    -- filter=139 channel=59
    -5, 4, 5, 0, 6, 0, -1, 0, 1,
    -- filter=139 channel=60
    5, -6, -5, 0, 4, 5, -1, 0, 7,
    -- filter=139 channel=61
    -1, 5, 0, 1, -3, 5, 5, 0, 3,
    -- filter=139 channel=62
    -3, -6, 1, -5, 3, 4, -6, 7, 0,
    -- filter=139 channel=63
    4, 3, -2, 0, -6, 2, 0, -7, -1,
    -- filter=139 channel=64
    -4, -4, -5, 4, -6, -7, -4, 4, 3,
    -- filter=139 channel=65
    -6, -4, 4, 3, -3, -6, 5, 6, 3,
    -- filter=139 channel=66
    -5, 0, -1, -4, -4, 2, -3, 3, -3,
    -- filter=139 channel=67
    4, 0, 4, -6, 6, -5, -1, 3, 1,
    -- filter=139 channel=68
    0, 0, 4, -4, -6, 7, 4, 2, 3,
    -- filter=139 channel=69
    -3, 1, 6, 4, 2, 4, 4, 4, -3,
    -- filter=139 channel=70
    -6, 0, 6, 0, 1, 2, -6, 4, 6,
    -- filter=139 channel=71
    -3, 0, 0, -3, 1, 7, 4, -2, 0,
    -- filter=139 channel=72
    6, -2, -2, -4, 5, -2, 4, -4, -6,
    -- filter=139 channel=73
    2, 4, -4, 7, 0, -6, -5, 2, -2,
    -- filter=139 channel=74
    -3, -3, -3, 0, -6, -6, 5, -1, 0,
    -- filter=139 channel=75
    5, -6, -1, -1, 0, -2, 5, 6, -4,
    -- filter=139 channel=76
    0, 0, 6, -1, 3, -7, -6, 6, 1,
    -- filter=139 channel=77
    3, 3, 6, -4, 6, -3, 1, -2, -3,
    -- filter=139 channel=78
    6, 2, 7, -3, 6, -7, 1, 5, 1,
    -- filter=139 channel=79
    6, 2, -1, -4, -7, 4, 3, 6, 5,
    -- filter=139 channel=80
    6, 6, -7, 5, -5, -7, -3, -4, -2,
    -- filter=139 channel=81
    4, -7, -3, -5, 0, 5, -4, -2, 6,
    -- filter=139 channel=82
    0, -3, -5, -6, 2, -3, -6, -3, -5,
    -- filter=139 channel=83
    4, -7, 2, 1, -6, 2, 5, 2, 6,
    -- filter=139 channel=84
    0, -7, -7, 3, 0, -7, -1, -1, 3,
    -- filter=139 channel=85
    -7, -7, 4, 4, -6, -2, 3, -2, 3,
    -- filter=139 channel=86
    2, -1, -3, 3, 3, 3, -4, 6, 2,
    -- filter=139 channel=87
    -7, -4, 1, -3, 1, 3, -5, -1, -3,
    -- filter=139 channel=88
    7, 5, 7, -6, -4, 2, -4, -1, -3,
    -- filter=139 channel=89
    5, 1, 4, -5, -7, -2, 4, 3, -6,
    -- filter=139 channel=90
    0, -3, 1, -2, -5, -1, -3, -4, -1,
    -- filter=139 channel=91
    -6, -1, -7, 6, -4, 5, -4, 1, -1,
    -- filter=139 channel=92
    -6, 0, -6, 0, -2, 0, -1, 2, 0,
    -- filter=139 channel=93
    6, 0, -7, 2, 5, -4, -2, -3, 0,
    -- filter=139 channel=94
    5, 3, 1, 3, 6, -7, -2, -4, 4,
    -- filter=139 channel=95
    1, -4, 4, 1, -5, 6, -2, 5, -7,
    -- filter=139 channel=96
    0, 5, 3, -4, 1, 0, 4, -6, 7,
    -- filter=139 channel=97
    -3, -4, 0, -1, 6, 0, 3, 0, 4,
    -- filter=139 channel=98
    -6, -5, -2, -5, 0, 0, 6, -2, -6,
    -- filter=139 channel=99
    -4, 6, -5, -2, -6, 1, -5, -6, 1,
    -- filter=139 channel=100
    0, -1, 0, 0, -5, 7, 1, 0, 1,
    -- filter=139 channel=101
    -2, 1, 4, 3, 3, -3, -3, -6, 6,
    -- filter=139 channel=102
    -3, 2, 4, -4, 6, 2, 0, 5, 1,
    -- filter=139 channel=103
    -5, -7, 0, 4, -1, -2, 6, 5, -1,
    -- filter=139 channel=104
    -6, 6, -4, -3, 6, -4, -1, 3, -6,
    -- filter=139 channel=105
    -4, 4, -2, -3, 6, 4, 4, -1, -4,
    -- filter=139 channel=106
    -1, -3, 0, -6, -4, 0, 0, 6, -4,
    -- filter=139 channel=107
    -5, 3, 6, 6, 0, 1, -5, 4, -4,
    -- filter=139 channel=108
    0, -3, -2, -3, 4, -6, -2, -4, 1,
    -- filter=139 channel=109
    4, 6, 1, -5, -1, 0, 0, 0, 6,
    -- filter=139 channel=110
    -1, 6, 5, 5, 3, -4, -7, -3, -5,
    -- filter=139 channel=111
    -4, -1, -4, 5, -5, 1, 3, 4, 2,
    -- filter=139 channel=112
    -5, -7, -2, -7, -4, 0, 2, 0, -3,
    -- filter=139 channel=113
    2, -5, 0, -1, -4, 6, -6, 2, -2,
    -- filter=139 channel=114
    3, -1, 7, 3, -4, 0, 3, -6, 4,
    -- filter=139 channel=115
    -5, 5, -5, 0, -1, 6, -2, -2, 0,
    -- filter=139 channel=116
    0, 0, 0, -2, 1, 4, 5, 2, 2,
    -- filter=139 channel=117
    -4, 0, -6, 4, -3, -4, 3, -3, 5,
    -- filter=139 channel=118
    -4, 0, 6, 5, 0, 4, -6, -2, -4,
    -- filter=139 channel=119
    7, 3, 4, 4, -1, 0, -6, 2, 3,
    -- filter=139 channel=120
    0, -5, -3, -3, -4, 5, -3, 7, 3,
    -- filter=139 channel=121
    6, -1, -3, 4, -6, 2, 2, -2, 1,
    -- filter=139 channel=122
    -2, -7, 6, 4, -3, 1, 0, 5, 0,
    -- filter=139 channel=123
    -2, 6, 3, 5, -5, -1, 7, -4, -4,
    -- filter=139 channel=124
    -1, 7, 0, 1, 2, -5, -3, 3, -5,
    -- filter=139 channel=125
    3, 6, 0, -7, -3, 0, 2, -3, 6,
    -- filter=139 channel=126
    1, -5, 1, -4, 0, 4, -3, 5, -5,
    -- filter=139 channel=127
    -5, -2, 3, 4, 0, -6, 0, 4, -2,
    -- filter=140 channel=0
    -6, -4, 4, -2, 1, -6, -2, 6, 0,
    -- filter=140 channel=1
    -7, 3, 0, 6, 4, 6, 4, 0, 3,
    -- filter=140 channel=2
    -3, 5, -7, 5, 3, -4, 2, 0, 0,
    -- filter=140 channel=3
    3, 5, 0, 3, 1, -1, -2, 6, -5,
    -- filter=140 channel=4
    3, -5, 4, -7, 7, -3, 5, 5, 0,
    -- filter=140 channel=5
    -1, 6, -6, 0, -1, 4, -2, 1, 4,
    -- filter=140 channel=6
    6, -6, -5, 6, -5, 0, 7, -6, 0,
    -- filter=140 channel=7
    -3, 6, 1, 2, 0, -1, 3, -7, -1,
    -- filter=140 channel=8
    -5, 4, 1, -7, 3, 5, 0, -2, -6,
    -- filter=140 channel=9
    -7, -4, -5, -4, 7, -1, -1, 0, 5,
    -- filter=140 channel=10
    0, 0, 0, 1, 0, -7, 3, 0, 3,
    -- filter=140 channel=11
    -4, 4, -5, 7, -7, 3, 4, 1, 0,
    -- filter=140 channel=12
    0, 3, 2, -4, -5, -5, 7, 7, 0,
    -- filter=140 channel=13
    0, -3, 0, 5, 1, -1, 2, 2, 0,
    -- filter=140 channel=14
    -3, 5, 5, -4, -2, 1, 6, -2, -4,
    -- filter=140 channel=15
    -6, 0, -4, 7, 0, 1, 0, 0, -4,
    -- filter=140 channel=16
    -4, -6, 4, 6, -5, 6, 6, 6, -4,
    -- filter=140 channel=17
    -4, 0, 0, -4, -7, 4, -6, 5, -1,
    -- filter=140 channel=18
    3, 4, -1, 3, 3, -4, -4, -4, 3,
    -- filter=140 channel=19
    1, -1, -5, 4, -7, -6, -5, 5, -1,
    -- filter=140 channel=20
    -2, -1, -2, -4, 5, -6, 2, -1, 5,
    -- filter=140 channel=21
    -4, 0, -7, 6, 6, 3, 5, -4, -5,
    -- filter=140 channel=22
    -6, 0, 2, 0, 6, 1, 2, -6, 7,
    -- filter=140 channel=23
    3, 7, -1, -3, -1, -6, -1, 0, -6,
    -- filter=140 channel=24
    0, 3, 6, 6, -5, -4, -3, -1, -3,
    -- filter=140 channel=25
    0, 0, -4, -1, 3, -3, 5, -6, -5,
    -- filter=140 channel=26
    -1, 0, -6, 1, -3, 0, 4, 1, 3,
    -- filter=140 channel=27
    -8, 1, 0, -7, 6, 4, -1, -2, 8,
    -- filter=140 channel=28
    3, -1, 2, 6, 7, 6, 4, -5, -6,
    -- filter=140 channel=29
    -7, -7, -1, -3, 4, 3, 0, 3, -2,
    -- filter=140 channel=30
    0, -6, -1, 0, 5, 1, 2, 8, 3,
    -- filter=140 channel=31
    0, -2, -7, 2, 6, -1, -6, 1, 1,
    -- filter=140 channel=32
    1, 2, 3, 0, 5, -7, -4, 4, 0,
    -- filter=140 channel=33
    0, 1, 2, -3, -7, -3, -4, -2, -5,
    -- filter=140 channel=34
    6, 0, -7, 0, 0, -6, 6, 3, -4,
    -- filter=140 channel=35
    0, 4, 3, -1, -5, 6, 6, 6, -4,
    -- filter=140 channel=36
    4, 3, 1, -3, 0, 5, -4, -5, 1,
    -- filter=140 channel=37
    6, -4, -1, -2, 0, 0, 7, 0, -4,
    -- filter=140 channel=38
    -4, -3, -1, 5, -3, 0, -2, 3, -2,
    -- filter=140 channel=39
    -6, 1, 0, -6, 5, -1, 1, 0, -2,
    -- filter=140 channel=40
    3, 7, -6, 3, -1, 4, -5, -7, 0,
    -- filter=140 channel=41
    -7, -3, -4, 4, 6, -1, -2, 1, -5,
    -- filter=140 channel=42
    1, -6, 7, 3, 2, -3, 0, 2, 1,
    -- filter=140 channel=43
    -6, -2, -5, -1, 7, -6, -6, -4, -3,
    -- filter=140 channel=44
    -3, 2, -2, 0, -4, -1, -3, -5, 4,
    -- filter=140 channel=45
    6, 1, -2, 0, -6, 4, -2, -3, -6,
    -- filter=140 channel=46
    -1, 0, -6, -2, -7, -4, -2, 7, -3,
    -- filter=140 channel=47
    0, -6, -5, 1, 3, -1, 5, 0, -3,
    -- filter=140 channel=48
    -4, -7, 0, -4, -2, 7, -3, -4, 6,
    -- filter=140 channel=49
    -6, 4, -5, -5, -4, 2, 5, 3, 0,
    -- filter=140 channel=50
    -1, 6, 3, -5, -4, -6, -6, -4, 7,
    -- filter=140 channel=51
    -3, -3, 3, 6, -6, 0, -7, 1, -7,
    -- filter=140 channel=52
    -1, 3, -2, 0, 6, 5, 5, -4, -4,
    -- filter=140 channel=53
    0, -4, 0, 6, 5, -2, -1, 0, 1,
    -- filter=140 channel=54
    -4, -5, 0, -7, 4, 6, -5, 2, -4,
    -- filter=140 channel=55
    -1, 3, -4, 1, -1, 2, -4, -7, 6,
    -- filter=140 channel=56
    0, 6, -4, 0, 0, -1, -3, 2, -4,
    -- filter=140 channel=57
    2, 0, 2, 5, 3, 1, 6, 5, -2,
    -- filter=140 channel=58
    -3, -3, 1, 1, -6, -2, 3, 2, 1,
    -- filter=140 channel=59
    -5, 4, -3, -1, 0, 7, 1, 4, 4,
    -- filter=140 channel=60
    -5, -7, 3, 0, -1, 3, 5, 2, -3,
    -- filter=140 channel=61
    3, 6, 6, -1, -6, 3, -6, 4, -2,
    -- filter=140 channel=62
    3, -1, 6, -1, 7, -3, -1, -7, 5,
    -- filter=140 channel=63
    1, 4, 0, 5, -4, 0, -6, -5, 5,
    -- filter=140 channel=64
    0, 3, 2, 4, -4, 6, -1, 0, -6,
    -- filter=140 channel=65
    -1, 5, 2, -4, -1, -5, -6, 0, -2,
    -- filter=140 channel=66
    1, -4, 4, 4, -6, 3, 5, 5, -3,
    -- filter=140 channel=67
    0, 1, 4, -4, 3, 2, 3, 0, 1,
    -- filter=140 channel=68
    -2, -5, -7, 4, -5, -1, -1, 3, -2,
    -- filter=140 channel=69
    -6, -4, -6, -1, -4, -5, -7, 7, -1,
    -- filter=140 channel=70
    3, 6, -2, -8, -1, 2, 3, 2, -5,
    -- filter=140 channel=71
    -1, 0, 2, -4, 3, 2, -1, 6, -4,
    -- filter=140 channel=72
    5, -3, 6, -3, -5, 5, -5, 4, 2,
    -- filter=140 channel=73
    -8, -2, 0, -7, -3, -1, -5, -3, 4,
    -- filter=140 channel=74
    6, -2, 5, 0, 5, -4, -3, 5, -1,
    -- filter=140 channel=75
    4, 2, -5, -6, 1, 2, -6, -1, -3,
    -- filter=140 channel=76
    4, -4, -5, -1, -5, 6, -5, 4, -5,
    -- filter=140 channel=77
    6, 6, -5, -5, 0, 6, 1, 2, 2,
    -- filter=140 channel=78
    -7, 3, 4, 0, 0, 0, -3, 0, 0,
    -- filter=140 channel=79
    -6, 3, 0, -1, 2, 5, 5, -6, 7,
    -- filter=140 channel=80
    0, 1, 0, 1, 1, 6, -4, -1, -6,
    -- filter=140 channel=81
    0, 7, -5, 4, 2, 3, -1, -3, 5,
    -- filter=140 channel=82
    -4, 5, -7, -6, -6, -6, -3, 4, 0,
    -- filter=140 channel=83
    -3, -2, 4, 4, 4, 0, 4, -2, 6,
    -- filter=140 channel=84
    4, 3, 1, -4, 5, -1, -4, -1, 6,
    -- filter=140 channel=85
    6, -2, 5, -1, -3, -3, -5, 6, -2,
    -- filter=140 channel=86
    6, 5, -2, 7, -3, -1, -2, 6, 2,
    -- filter=140 channel=87
    0, -5, 4, -4, -1, 6, 1, 2, 0,
    -- filter=140 channel=88
    0, 4, 4, 5, 2, 5, 6, 2, 0,
    -- filter=140 channel=89
    3, -2, -4, -1, -4, -5, -4, -5, 3,
    -- filter=140 channel=90
    -5, 2, -3, 4, -4, -3, 1, 4, -5,
    -- filter=140 channel=91
    5, -4, 4, 0, 3, -3, 3, 1, 2,
    -- filter=140 channel=92
    -5, 7, -7, -7, 0, -7, -5, -4, 0,
    -- filter=140 channel=93
    -1, -3, -4, 6, 4, 6, 7, -5, 1,
    -- filter=140 channel=94
    -1, -6, 2, -1, -6, 4, 0, 2, 5,
    -- filter=140 channel=95
    0, 0, 3, -6, -5, 7, 7, 2, 3,
    -- filter=140 channel=96
    6, -5, -6, -3, 5, -5, -6, 0, -5,
    -- filter=140 channel=97
    -1, 7, 5, -6, 2, -3, -2, 1, 1,
    -- filter=140 channel=98
    -4, 0, -2, -4, -5, 5, -4, -2, 5,
    -- filter=140 channel=99
    -3, 1, 0, -7, 7, -3, -6, 7, -6,
    -- filter=140 channel=100
    -3, -2, 2, 3, 0, 4, 3, -6, 1,
    -- filter=140 channel=101
    0, 3, 2, 5, 5, 0, 7, -2, -2,
    -- filter=140 channel=102
    1, 4, 2, 2, 3, 4, 2, -6, -4,
    -- filter=140 channel=103
    -3, -1, -2, 0, 0, -5, -3, 4, 6,
    -- filter=140 channel=104
    0, 2, 4, -7, -1, 0, -3, -5, 2,
    -- filter=140 channel=105
    -3, -6, 5, 2, 7, -5, -6, -4, 6,
    -- filter=140 channel=106
    -3, -6, -5, -6, 2, 3, 0, 2, 6,
    -- filter=140 channel=107
    -4, 7, 0, -1, -2, -5, 2, 0, 1,
    -- filter=140 channel=108
    5, 2, -5, -5, 0, -5, 4, -4, 0,
    -- filter=140 channel=109
    6, 5, 0, 0, -3, 0, 0, 7, -1,
    -- filter=140 channel=110
    5, -6, 0, 0, 5, 2, -2, 0, -2,
    -- filter=140 channel=111
    2, 4, 4, 2, 2, 0, -5, 0, 3,
    -- filter=140 channel=112
    2, -3, -6, 1, 0, 7, -3, 2, -6,
    -- filter=140 channel=113
    -1, 0, -6, 6, -3, 0, -7, -3, 5,
    -- filter=140 channel=114
    1, 2, 0, -5, 1, -2, 2, 6, -6,
    -- filter=140 channel=115
    2, 4, -5, -5, 4, 0, -5, -2, 2,
    -- filter=140 channel=116
    2, 6, 0, -2, 1, -1, -3, -5, -4,
    -- filter=140 channel=117
    1, 3, 0, 1, 3, 0, -2, -5, -6,
    -- filter=140 channel=118
    3, 7, -1, -7, 6, 3, -5, 0, -5,
    -- filter=140 channel=119
    -4, -1, -1, -4, 5, -2, -1, 5, -2,
    -- filter=140 channel=120
    4, 1, -6, -6, -5, 4, -6, 8, 2,
    -- filter=140 channel=121
    -1, 2, 0, 1, 1, 6, -5, -2, -1,
    -- filter=140 channel=122
    -2, -1, -1, -5, -2, -4, -7, -4, -4,
    -- filter=140 channel=123
    -3, -3, 2, -4, -5, 1, -1, 4, 0,
    -- filter=140 channel=124
    -5, 5, -5, 7, 1, -2, 5, 4, -7,
    -- filter=140 channel=125
    0, 2, -4, -4, 1, 0, -1, 0, -3,
    -- filter=140 channel=126
    2, 0, 5, 2, 4, 7, -1, 6, -1,
    -- filter=140 channel=127
    -6, -4, 1, 0, 1, 0, 5, 1, 1,
    -- filter=141 channel=0
    6, -8, 3, -1, -8, 9, 10, -3, 13,
    -- filter=141 channel=1
    -7, 0, 0, -4, -20, 1, 12, -4, 1,
    -- filter=141 channel=2
    -7, 0, 7, 0, -8, 3, 6, -6, 0,
    -- filter=141 channel=3
    3, 0, 0, -10, -2, -4, -3, -4, -3,
    -- filter=141 channel=4
    -4, 3, 0, 8, -11, -3, -2, -9, -13,
    -- filter=141 channel=5
    -5, 1, -5, -3, 9, -3, 12, -1, 0,
    -- filter=141 channel=6
    -1, 1, 5, 3, 3, 5, 1, 8, -1,
    -- filter=141 channel=7
    -5, -4, 0, 7, 3, 1, -2, -4, -1,
    -- filter=141 channel=8
    -3, 0, 0, 0, -2, 6, -11, -3, 1,
    -- filter=141 channel=9
    -5, 8, -5, -4, -6, 10, -2, -8, 0,
    -- filter=141 channel=10
    0, 5, 8, -8, 3, 2, 0, 0, -1,
    -- filter=141 channel=11
    2, -2, -1, -6, 2, 5, 4, -10, -2,
    -- filter=141 channel=12
    2, 4, 4, 4, -5, 15, 4, 8, 1,
    -- filter=141 channel=13
    -8, -11, 1, -7, -19, 15, 4, -9, -1,
    -- filter=141 channel=14
    -5, -1, 5, -4, -1, -2, 1, 3, 3,
    -- filter=141 channel=15
    0, -10, 9, -7, -4, 1, -1, -11, 0,
    -- filter=141 channel=16
    0, 12, -4, -6, 0, 3, 2, 0, -1,
    -- filter=141 channel=17
    2, -3, 0, 2, 0, 5, 2, -3, 2,
    -- filter=141 channel=18
    3, -7, 10, -8, -13, 18, 5, -6, 9,
    -- filter=141 channel=19
    0, 2, 2, 0, -5, 0, -5, 1, -3,
    -- filter=141 channel=20
    0, -3, 7, -5, 4, 0, -2, 0, 9,
    -- filter=141 channel=21
    7, 11, -1, 1, 0, 2, -5, 2, 3,
    -- filter=141 channel=22
    0, 6, 4, -3, -3, 1, 1, 3, 5,
    -- filter=141 channel=23
    -5, 0, 5, -29, 8, 10, -9, -18, 19,
    -- filter=141 channel=24
    0, 6, 5, 1, 5, 5, -4, 5, -1,
    -- filter=141 channel=25
    -4, -6, 4, -1, -18, 19, 13, -6, -2,
    -- filter=141 channel=26
    3, 6, 8, 9, 6, 5, 5, 6, -4,
    -- filter=141 channel=27
    -9, -6, 8, -15, -3, 19, 4, -24, 15,
    -- filter=141 channel=28
    0, 4, -1, 6, -7, -6, -5, 0, 2,
    -- filter=141 channel=29
    3, 4, 0, 0, 4, -1, 2, 4, -3,
    -- filter=141 channel=30
    -7, 0, 7, -5, -7, 11, 0, -2, -3,
    -- filter=141 channel=31
    -10, 8, 7, -19, 10, 12, -9, -16, -2,
    -- filter=141 channel=32
    1, -5, 15, -8, -11, 13, 9, -16, 10,
    -- filter=141 channel=33
    0, -6, 0, -16, -5, 19, 5, -16, 10,
    -- filter=141 channel=34
    13, 17, 5, -3, 18, 11, -3, 11, 22,
    -- filter=141 channel=35
    2, 4, -5, -4, -2, 5, 6, 3, -4,
    -- filter=141 channel=36
    2, 9, -2, -5, 6, -7, -6, -3, -8,
    -- filter=141 channel=37
    -6, -5, 5, -5, -7, 6, 2, -3, -4,
    -- filter=141 channel=38
    3, 0, 7, -9, 1, 1, -4, -6, 2,
    -- filter=141 channel=39
    -3, 1, 0, 6, 5, 1, 3, 5, -4,
    -- filter=141 channel=40
    6, -3, -7, -8, 0, 4, -9, -11, 9,
    -- filter=141 channel=41
    14, 7, 12, 9, -6, 20, 1, 5, -1,
    -- filter=141 channel=42
    3, -10, 8, -3, 0, -4, -3, -4, -6,
    -- filter=141 channel=43
    9, 1, -5, -4, 3, 0, 1, -7, 4,
    -- filter=141 channel=44
    -5, -4, -3, -1, -5, 3, -4, 3, 1,
    -- filter=141 channel=45
    -3, -4, -3, 0, 5, 3, 1, -2, 2,
    -- filter=141 channel=46
    1, 5, -2, -4, 1, 4, 0, -2, -2,
    -- filter=141 channel=47
    4, 0, -3, 1, 6, 9, 6, -5, 4,
    -- filter=141 channel=48
    0, 5, 8, -1, -1, 4, 4, 0, -1,
    -- filter=141 channel=49
    -12, -11, 0, -8, -2, 1, -3, -1, -4,
    -- filter=141 channel=50
    -5, -3, 6, -9, -4, 3, -1, -15, 0,
    -- filter=141 channel=51
    -3, -1, 0, 1, 7, 0, 3, 0, 3,
    -- filter=141 channel=52
    1, 7, -1, -3, 6, 0, 0, -2, 3,
    -- filter=141 channel=53
    7, 4, 5, -2, 1, 1, 8, -8, 8,
    -- filter=141 channel=54
    3, 1, 1, 0, 3, -2, 2, 1, 3,
    -- filter=141 channel=55
    -4, -4, 0, -13, -9, 8, 4, -10, 0,
    -- filter=141 channel=56
    3, 2, 10, -7, 1, -1, -10, -4, 12,
    -- filter=141 channel=57
    5, 2, 1, 9, -2, 0, -4, 8, 3,
    -- filter=141 channel=58
    2, 8, -2, 2, 2, 8, 3, 7, -3,
    -- filter=141 channel=59
    0, -10, 8, 2, -5, 13, 8, 1, 1,
    -- filter=141 channel=60
    -4, -1, -1, 7, 2, -5, -4, 5, 4,
    -- filter=141 channel=61
    2, 2, 6, 4, 0, -1, 3, -5, -4,
    -- filter=141 channel=62
    6, -7, -3, 2, -7, -1, 2, -7, -2,
    -- filter=141 channel=63
    9, 12, 2, 2, 2, 3, 7, 6, 3,
    -- filter=141 channel=64
    1, -5, 2, -1, 4, -1, -4, -6, -4,
    -- filter=141 channel=65
    -2, 6, -4, -4, 4, -1, 4, 3, 2,
    -- filter=141 channel=66
    1, 4, 8, 11, -1, 22, 4, 0, 4,
    -- filter=141 channel=67
    -6, 3, -4, 1, -5, -4, 0, 3, 7,
    -- filter=141 channel=68
    -1, -9, 5, 2, -6, 2, -3, -6, -8,
    -- filter=141 channel=69
    4, 2, 3, 4, -1, 8, 8, 0, 6,
    -- filter=141 channel=70
    -7, 0, 11, -17, 2, 11, -8, -18, 6,
    -- filter=141 channel=71
    -1, 3, -9, -9, -8, -8, -6, -1, -2,
    -- filter=141 channel=72
    0, 0, 9, 0, -9, 7, -7, 0, -7,
    -- filter=141 channel=73
    -5, -2, 0, 0, -7, 3, 8, -2, -4,
    -- filter=141 channel=74
    -5, 2, -2, -13, 12, 14, -3, -13, 6,
    -- filter=141 channel=75
    -2, -4, -4, -3, -14, 4, 8, -8, 1,
    -- filter=141 channel=76
    -1, -2, 3, 5, -3, 0, 3, 2, -5,
    -- filter=141 channel=77
    -5, 6, -6, -6, 6, -6, 2, -3, -4,
    -- filter=141 channel=78
    6, 2, 6, 0, 0, -4, -4, 4, 5,
    -- filter=141 channel=79
    -3, -12, 10, -17, -22, 24, 6, -20, 10,
    -- filter=141 channel=80
    -7, 0, 0, -2, -2, 7, 0, -8, -6,
    -- filter=141 channel=81
    -4, 0, 4, -4, 1, -2, 3, 2, 6,
    -- filter=141 channel=82
    6, 5, 4, -9, 3, -2, 0, -8, 1,
    -- filter=141 channel=83
    2, -5, 3, -1, -9, -7, 7, 4, -2,
    -- filter=141 channel=84
    -7, -1, 9, -9, -5, 9, 2, 1, 3,
    -- filter=141 channel=85
    5, 1, 1, -4, -7, 0, -3, 6, -6,
    -- filter=141 channel=86
    0, 2, 2, -2, -3, 9, -1, 2, 5,
    -- filter=141 channel=87
    -5, 6, 5, -9, 7, 9, 0, -1, 9,
    -- filter=141 channel=88
    4, 12, 4, -10, 14, -4, -1, 3, 2,
    -- filter=141 channel=89
    -8, -10, -1, -14, -15, 9, -7, -17, -8,
    -- filter=141 channel=90
    6, 11, 5, -1, 16, 4, -16, 5, 3,
    -- filter=141 channel=91
    -7, -5, 3, -15, -5, 13, 7, -9, 5,
    -- filter=141 channel=92
    6, -1, 0, 0, 7, 1, -6, 3, 8,
    -- filter=141 channel=93
    -7, 9, 1, 3, -5, 2, 3, 0, -2,
    -- filter=141 channel=94
    4, -7, 3, 1, -7, -2, 5, 0, 4,
    -- filter=141 channel=95
    -4, 3, 3, -7, 4, 2, -5, 0, 0,
    -- filter=141 channel=96
    -8, -3, 3, -1, 0, 2, -2, 3, 2,
    -- filter=141 channel=97
    9, 0, -2, -3, 4, 0, 0, 0, 8,
    -- filter=141 channel=98
    -8, 0, 14, -6, -4, 22, 4, -10, 2,
    -- filter=141 channel=99
    -8, 9, -1, -20, 17, 10, -11, -12, 2,
    -- filter=141 channel=100
    -7, -3, 5, -7, -1, 2, 2, -4, 3,
    -- filter=141 channel=101
    -1, -5, 4, 6, -7, -3, 0, -7, -8,
    -- filter=141 channel=102
    4, 4, 4, -2, -5, -6, 0, 0, -7,
    -- filter=141 channel=103
    6, 0, -8, -9, -4, 1, -2, -11, 9,
    -- filter=141 channel=104
    -2, 6, 0, -3, -6, 4, 3, 2, 5,
    -- filter=141 channel=105
    9, 0, 0, 0, 1, -4, 4, 3, -4,
    -- filter=141 channel=106
    2, -8, -3, -1, -6, 0, -1, 2, 0,
    -- filter=141 channel=107
    1, 1, 8, -13, 5, 0, 1, -9, 13,
    -- filter=141 channel=108
    9, 6, 2, 5, 0, 8, 8, 0, -4,
    -- filter=141 channel=109
    -3, -4, 8, -7, -6, 19, 6, -10, -3,
    -- filter=141 channel=110
    6, 10, 6, -4, 0, 7, -10, 0, 3,
    -- filter=141 channel=111
    8, -6, 6, 1, -5, -4, 5, -5, 0,
    -- filter=141 channel=112
    -6, -1, -3, -11, -1, 10, -2, -5, 8,
    -- filter=141 channel=113
    -2, -2, -3, -5, -6, 0, -5, -10, 8,
    -- filter=141 channel=114
    -13, -9, 15, -5, -17, 13, 7, -12, 9,
    -- filter=141 channel=115
    3, 0, -4, -2, -2, 0, 5, 0, -1,
    -- filter=141 channel=116
    -10, -5, 12, -4, -10, 3, 13, -9, -5,
    -- filter=141 channel=117
    5, -7, 0, -4, -2, 3, -7, -7, -7,
    -- filter=141 channel=118
    -1, 1, 7, -3, 3, 0, 3, -3, -1,
    -- filter=141 channel=119
    5, 13, 1, -13, 21, 11, -2, 12, 19,
    -- filter=141 channel=120
    -1, 12, 14, -21, -1, 13, 0, -14, 11,
    -- filter=141 channel=121
    0, 1, 2, 3, -9, 3, -1, -9, -5,
    -- filter=141 channel=122
    6, 17, -10, -3, 1, 7, -7, -2, 1,
    -- filter=141 channel=123
    6, 8, 3, -7, 15, 8, 2, 5, 11,
    -- filter=141 channel=124
    7, 1, 7, 4, -3, 7, -2, -7, 3,
    -- filter=141 channel=125
    -14, 3, 0, -9, -3, 15, -2, -14, 4,
    -- filter=141 channel=126
    1, -2, 5, -8, -10, 12, 0, 0, 4,
    -- filter=141 channel=127
    -2, 2, 6, -2, -6, 0, 8, 1, -2,
    -- filter=142 channel=0
    1, -5, -4, 2, 4, 0, -6, -4, -1,
    -- filter=142 channel=1
    1, 3, 3, 2, 0, -6, 0, -4, 2,
    -- filter=142 channel=2
    -3, -3, -1, -4, -4, 0, -2, 4, 6,
    -- filter=142 channel=3
    0, 1, 0, -6, 7, -1, 4, 4, 8,
    -- filter=142 channel=4
    -3, 2, 2, 2, -4, 2, 1, -6, 5,
    -- filter=142 channel=5
    -5, -1, 4, 2, 2, 4, 2, -1, 2,
    -- filter=142 channel=6
    0, -1, -2, -5, 0, 5, 7, 0, 0,
    -- filter=142 channel=7
    4, 0, 1, 7, -2, 7, 2, 1, 4,
    -- filter=142 channel=8
    -2, -4, -3, 0, 0, -6, 1, -5, -4,
    -- filter=142 channel=9
    0, -4, 2, 6, 3, 5, 0, 1, 5,
    -- filter=142 channel=10
    0, -1, -6, 2, -2, 0, 5, 6, 0,
    -- filter=142 channel=11
    -4, 0, -6, 0, 0, -6, -6, 1, -1,
    -- filter=142 channel=12
    0, -1, 0, 0, -1, 5, 7, -1, 5,
    -- filter=142 channel=13
    1, 4, -5, -3, -4, -5, -5, -5, 6,
    -- filter=142 channel=14
    -1, 6, 0, 1, 0, 7, 0, 5, -6,
    -- filter=142 channel=15
    1, -2, 0, 6, -2, -3, 2, -2, -6,
    -- filter=142 channel=16
    5, -4, 0, -1, 0, 3, 6, -2, 5,
    -- filter=142 channel=17
    -3, 2, -6, -3, 2, 5, 5, 4, -3,
    -- filter=142 channel=18
    6, -3, -4, -2, 5, 4, 2, 2, 4,
    -- filter=142 channel=19
    -6, 2, 0, 1, 0, 4, 0, -4, -4,
    -- filter=142 channel=20
    -2, 1, 1, 2, -3, -7, 6, 0, -6,
    -- filter=142 channel=21
    6, 2, 1, 2, -1, 5, 6, -4, -2,
    -- filter=142 channel=22
    7, -4, -5, -1, 0, 0, 0, -3, -6,
    -- filter=142 channel=23
    -2, -4, -1, 1, 7, 6, -5, -6, 0,
    -- filter=142 channel=24
    -4, 6, 4, -3, -6, -3, 3, -3, 0,
    -- filter=142 channel=25
    -4, -5, -4, -3, -3, -5, -4, 2, -6,
    -- filter=142 channel=26
    6, -7, -6, 3, 7, -7, -1, 0, -6,
    -- filter=142 channel=27
    -3, -1, 3, 5, -4, -5, 6, -3, 6,
    -- filter=142 channel=28
    -2, -2, -2, -5, -4, 1, -7, -4, -4,
    -- filter=142 channel=29
    0, 6, -2, 3, -7, 3, -4, 3, 5,
    -- filter=142 channel=30
    -3, 1, -2, 7, 1, 7, -3, 0, 4,
    -- filter=142 channel=31
    -3, 0, -5, 3, 2, -2, -7, 3, -6,
    -- filter=142 channel=32
    0, -1, 5, -1, 1, 2, 0, -1, 2,
    -- filter=142 channel=33
    -2, 7, -2, -1, -3, 5, -1, -5, -5,
    -- filter=142 channel=34
    -3, 3, 2, 8, 2, -4, 1, 1, -6,
    -- filter=142 channel=35
    1, 5, 4, -4, 5, -2, -7, -4, -6,
    -- filter=142 channel=36
    0, 5, 1, -6, 0, 1, 1, 5, 0,
    -- filter=142 channel=37
    -6, -3, 7, -3, 0, -6, 6, -5, 5,
    -- filter=142 channel=38
    0, 1, 5, 7, -4, -3, -5, -3, 7,
    -- filter=142 channel=39
    3, -3, -1, 2, -5, -1, -3, 0, 0,
    -- filter=142 channel=40
    0, -1, 5, 4, -1, 7, -1, -4, 5,
    -- filter=142 channel=41
    -2, -5, -3, -3, 6, 4, -4, 0, 0,
    -- filter=142 channel=42
    1, 0, -4, -1, -3, 0, -6, 0, -3,
    -- filter=142 channel=43
    -1, -7, 2, 2, 4, 2, 0, 7, -4,
    -- filter=142 channel=44
    0, 0, 2, 6, 2, 0, 2, -7, 5,
    -- filter=142 channel=45
    3, 0, 0, -3, -6, -3, 5, 0, 4,
    -- filter=142 channel=46
    -4, 3, -1, -7, 7, 3, -3, 6, 0,
    -- filter=142 channel=47
    0, 4, 1, -1, 2, 6, 0, -3, 0,
    -- filter=142 channel=48
    0, -2, 4, -1, -2, -4, 6, 0, 3,
    -- filter=142 channel=49
    6, 0, -2, 4, -2, -2, 1, 2, 4,
    -- filter=142 channel=50
    0, -5, 3, -3, 1, 2, -4, -5, -3,
    -- filter=142 channel=51
    5, -4, 4, 2, -7, 0, 6, 5, 0,
    -- filter=142 channel=52
    -1, -4, -3, 4, -1, -3, -6, -5, -2,
    -- filter=142 channel=53
    -1, 2, -6, 7, 0, -4, 6, 0, 0,
    -- filter=142 channel=54
    -2, 0, 3, 2, 4, 4, -1, 6, 0,
    -- filter=142 channel=55
    1, 5, -6, 6, -3, -3, 0, -2, -2,
    -- filter=142 channel=56
    4, 0, -5, -6, 1, 5, 6, 0, -6,
    -- filter=142 channel=57
    5, 1, -6, -5, 0, -4, 5, -5, -1,
    -- filter=142 channel=58
    3, -5, 6, 0, 1, -1, 4, 1, 0,
    -- filter=142 channel=59
    1, 1, 7, 1, 3, 0, 1, -2, -3,
    -- filter=142 channel=60
    -1, 5, -1, 0, 4, 0, 0, -2, 7,
    -- filter=142 channel=61
    3, 7, -4, 4, 1, 7, -3, 5, -4,
    -- filter=142 channel=62
    0, -5, -5, 5, 2, 1, 0, -6, -3,
    -- filter=142 channel=63
    5, 6, -4, -3, 2, -1, 7, 6, -5,
    -- filter=142 channel=64
    -2, 6, -4, 3, -4, -1, 4, -6, -3,
    -- filter=142 channel=65
    3, 7, 7, 6, 3, 0, -3, 0, -5,
    -- filter=142 channel=66
    4, 7, 7, -2, -7, 1, -1, -1, 3,
    -- filter=142 channel=67
    1, 0, -2, -4, 3, -6, -1, 4, -1,
    -- filter=142 channel=68
    -1, 2, 1, 3, 2, -6, 5, 7, -6,
    -- filter=142 channel=69
    -3, 0, 1, -2, -4, -7, -6, 6, -5,
    -- filter=142 channel=70
    4, 5, 4, 3, -2, -4, -5, -2, -4,
    -- filter=142 channel=71
    0, -2, -6, 5, -3, -6, 4, -4, -3,
    -- filter=142 channel=72
    1, 5, -3, -7, 0, 4, 3, 3, -5,
    -- filter=142 channel=73
    2, 0, -6, -6, 3, 0, 1, -2, -1,
    -- filter=142 channel=74
    9, 4, 6, 5, 4, 0, 5, 5, 0,
    -- filter=142 channel=75
    -7, 8, 1, -1, 3, -4, 8, -4, 4,
    -- filter=142 channel=76
    4, -6, -3, -1, -3, -7, -3, 5, 4,
    -- filter=142 channel=77
    2, -5, 5, 0, 3, 5, -3, -3, -4,
    -- filter=142 channel=78
    -5, -5, 6, -1, -2, -1, 5, -6, -2,
    -- filter=142 channel=79
    -7, -6, 4, -4, 4, 0, 0, -2, 0,
    -- filter=142 channel=80
    -5, -4, -2, 0, 1, 2, 6, -7, 0,
    -- filter=142 channel=81
    2, 6, 2, 0, -6, -4, 0, -2, 1,
    -- filter=142 channel=82
    2, 3, 5, -3, -3, -3, 6, 1, 5,
    -- filter=142 channel=83
    -1, 0, 7, -2, 6, -3, -5, 6, 6,
    -- filter=142 channel=84
    2, -4, -7, 1, 4, 5, -1, 4, 0,
    -- filter=142 channel=85
    4, 1, 0, 4, -2, -3, 7, 0, -6,
    -- filter=142 channel=86
    3, 7, 1, -3, -6, 3, 4, -3, 0,
    -- filter=142 channel=87
    -3, 0, 2, 1, -1, -4, 1, 7, 3,
    -- filter=142 channel=88
    8, -1, 0, 1, -4, 5, -6, -4, -5,
    -- filter=142 channel=89
    -7, 3, 4, 4, 7, 0, 0, -6, -1,
    -- filter=142 channel=90
    2, -4, 7, -2, 0, 4, -3, -5, 7,
    -- filter=142 channel=91
    1, -4, -7, 6, -1, 0, 4, -5, 1,
    -- filter=142 channel=92
    -4, -3, 7, 6, -4, -1, 7, -5, -2,
    -- filter=142 channel=93
    -5, 6, 3, 0, 2, 0, -4, 6, -6,
    -- filter=142 channel=94
    4, 3, -4, -5, 1, 4, -4, 0, -4,
    -- filter=142 channel=95
    -5, 6, -1, -3, 1, -1, 0, -6, 5,
    -- filter=142 channel=96
    -3, -6, 5, -7, -5, -2, -3, -2, -1,
    -- filter=142 channel=97
    1, 0, -3, 4, -3, 4, 2, 4, 6,
    -- filter=142 channel=98
    -2, 7, -3, 2, 0, 0, -2, -6, -7,
    -- filter=142 channel=99
    8, -5, 0, 0, -8, -1, 2, -8, -7,
    -- filter=142 channel=100
    4, 4, 3, -1, 7, -5, 1, 0, 0,
    -- filter=142 channel=101
    0, 1, 2, -1, -2, -4, -4, -7, 4,
    -- filter=142 channel=102
    -6, 6, 4, -1, -1, 4, 1, -4, 1,
    -- filter=142 channel=103
    1, 2, -4, -1, -1, 8, -5, -3, 6,
    -- filter=142 channel=104
    1, -5, 6, -7, -7, -2, 0, -1, -6,
    -- filter=142 channel=105
    0, -4, 3, 1, -5, -7, 7, -2, -1,
    -- filter=142 channel=106
    6, -3, -7, 7, 6, 6, -5, 1, -5,
    -- filter=142 channel=107
    6, 5, 0, 7, -7, -5, -7, 0, -1,
    -- filter=142 channel=108
    2, -2, 5, 0, 7, 1, 1, -5, 0,
    -- filter=142 channel=109
    -6, 1, -3, 6, 0, 2, -5, -8, 3,
    -- filter=142 channel=110
    0, 5, 0, -1, -6, 7, 0, -6, -1,
    -- filter=142 channel=111
    0, 7, 3, 0, -4, 1, -1, 7, -7,
    -- filter=142 channel=112
    -2, -5, 0, 2, -3, -2, 0, -3, 5,
    -- filter=142 channel=113
    0, -2, 2, -2, 6, -6, 1, 6, -3,
    -- filter=142 channel=114
    0, -4, -8, 0, -6, 0, 1, -1, -2,
    -- filter=142 channel=115
    3, -3, -1, 3, 0, -6, 2, 0, -5,
    -- filter=142 channel=116
    -3, 0, 1, 3, 0, 1, -7, -3, 6,
    -- filter=142 channel=117
    2, 7, 3, -5, 2, 5, -7, 1, -3,
    -- filter=142 channel=118
    -6, 4, 5, 0, -5, -5, 1, -2, 1,
    -- filter=142 channel=119
    1, 0, -6, 0, 2, 5, 2, -5, 7,
    -- filter=142 channel=120
    -3, -4, -3, 7, 2, -3, 2, 0, 2,
    -- filter=142 channel=121
    -5, 0, -2, -3, -5, 5, 1, -7, 1,
    -- filter=142 channel=122
    2, 2, 8, -6, 3, 0, -3, -7, -5,
    -- filter=142 channel=123
    -4, 1, -6, 3, -4, 3, 5, 2, -1,
    -- filter=142 channel=124
    0, 2, 0, 7, 3, 1, 5, 3, 7,
    -- filter=142 channel=125
    -1, -5, 5, 0, -4, -4, 5, 1, -7,
    -- filter=142 channel=126
    -3, -2, -1, -6, 4, -5, 2, 1, -5,
    -- filter=142 channel=127
    -6, 0, 4, -5, 2, -5, 0, 1, 2,
    -- filter=143 channel=0
    -3, -4, 2, 1, 5, 0, -5, 3, 5,
    -- filter=143 channel=1
    -8, 4, -2, -1, -2, -5, -9, -7, 3,
    -- filter=143 channel=2
    0, -3, 0, 0, 6, 0, 0, 2, 2,
    -- filter=143 channel=3
    -7, -2, 2, 1, -1, 0, 1, 1, 4,
    -- filter=143 channel=4
    3, 6, 1, 5, 1, 1, -3, 3, 0,
    -- filter=143 channel=5
    1, -3, 4, -3, 2, -2, 4, 3, 4,
    -- filter=143 channel=6
    -1, 1, -6, 6, -4, 2, 0, -6, -6,
    -- filter=143 channel=7
    -4, 4, -5, -2, 0, -1, -7, 7, -6,
    -- filter=143 channel=8
    -1, 5, -5, -7, 0, -3, -2, 2, 5,
    -- filter=143 channel=9
    -1, 6, 6, 3, -1, 4, -5, 2, -3,
    -- filter=143 channel=10
    0, 6, 1, 3, 1, 2, -3, -2, -3,
    -- filter=143 channel=11
    -3, -5, -5, -5, 1, -4, 4, -2, 0,
    -- filter=143 channel=12
    -8, 1, 7, -5, 4, 7, 4, -7, 8,
    -- filter=143 channel=13
    -6, 4, -1, -3, 0, 2, -5, -8, 6,
    -- filter=143 channel=14
    -4, 0, -5, -6, 2, 0, 5, 1, 0,
    -- filter=143 channel=15
    1, -6, -1, -2, -8, -5, 0, 0, 5,
    -- filter=143 channel=16
    -1, -5, 0, 2, 3, -4, -2, 2, 8,
    -- filter=143 channel=17
    -1, -4, -1, -7, 6, 5, -1, 4, 2,
    -- filter=143 channel=18
    -5, -8, 3, -9, -5, 0, -10, 0, 0,
    -- filter=143 channel=19
    -5, -1, -6, -6, -5, 0, 3, -1, -2,
    -- filter=143 channel=20
    6, -2, 3, 7, 5, -7, -5, 8, -1,
    -- filter=143 channel=21
    -5, 0, -5, -4, -2, 6, 3, 5, 0,
    -- filter=143 channel=22
    -2, 0, -1, 3, -3, -2, 2, 4, 7,
    -- filter=143 channel=23
    -2, -1, 0, -7, 2, 4, -10, -3, 1,
    -- filter=143 channel=24
    6, 0, -4, -1, -3, -3, -6, -6, -4,
    -- filter=143 channel=25
    -7, 1, 8, -6, -5, 6, -3, -6, 0,
    -- filter=143 channel=26
    -6, 0, -1, 0, -5, 4, 8, -6, 0,
    -- filter=143 channel=27
    -3, -4, 3, 0, -4, 6, -8, -7, 1,
    -- filter=143 channel=28
    -5, 0, 0, 2, 5, 0, 2, 0, -4,
    -- filter=143 channel=29
    -5, 0, -6, 6, -1, 4, -1, 3, -5,
    -- filter=143 channel=30
    -5, 0, -4, -7, 4, -1, 1, -8, 2,
    -- filter=143 channel=31
    -2, -6, 0, 1, -6, 3, -4, -5, -1,
    -- filter=143 channel=32
    1, 2, 4, -8, -3, -4, -4, -7, 5,
    -- filter=143 channel=33
    -9, 4, 6, -4, 0, 8, 1, 5, 0,
    -- filter=143 channel=34
    -4, 2, 0, -2, 7, 5, 2, 4, 0,
    -- filter=143 channel=35
    3, -2, -3, 6, -5, 0, 7, -5, -1,
    -- filter=143 channel=36
    -2, 7, 2, 1, 0, -4, 7, -1, 4,
    -- filter=143 channel=37
    -4, -2, 5, -8, 3, 9, 0, 0, -4,
    -- filter=143 channel=38
    -1, -6, 2, 0, 1, 7, 4, -6, 6,
    -- filter=143 channel=39
    -2, 4, 7, 6, 3, -1, -6, -2, -3,
    -- filter=143 channel=40
    -5, -5, 3, 7, -6, 8, 0, 2, 7,
    -- filter=143 channel=41
    0, -1, 0, 2, 4, 5, 1, -4, -3,
    -- filter=143 channel=42
    3, 2, -1, 3, 3, -1, -7, -2, -2,
    -- filter=143 channel=43
    -5, 0, -2, -6, -1, 3, 4, 0, 4,
    -- filter=143 channel=44
    0, 2, -6, 2, 1, 1, -6, -4, -5,
    -- filter=143 channel=45
    -4, 0, -4, 6, 7, 3, -3, -6, 3,
    -- filter=143 channel=46
    -3, 4, -1, -6, 7, 0, -6, -4, -7,
    -- filter=143 channel=47
    2, 4, -1, -4, 6, 0, -9, -8, 6,
    -- filter=143 channel=48
    -2, -1, 5, 1, 1, -1, -1, 2, -3,
    -- filter=143 channel=49
    1, -7, -1, 5, 0, -7, -6, -3, 3,
    -- filter=143 channel=50
    -8, 2, 6, -6, 5, -7, 3, -2, 5,
    -- filter=143 channel=51
    1, 0, -1, -1, 4, 0, 3, 6, -7,
    -- filter=143 channel=52
    -4, 2, -1, 0, 2, 2, -4, 2, 4,
    -- filter=143 channel=53
    5, 4, 3, -4, -3, 0, -5, 6, 0,
    -- filter=143 channel=54
    -4, 4, -3, -3, 0, 2, -4, -1, 1,
    -- filter=143 channel=55
    -4, -4, 7, 0, -9, 0, -6, 5, 7,
    -- filter=143 channel=56
    0, 6, -4, -6, 6, -2, -4, 8, 6,
    -- filter=143 channel=57
    -7, -6, 3, 0, -6, 1, -4, -5, 5,
    -- filter=143 channel=58
    2, -3, 2, -4, 6, 1, -1, -1, -6,
    -- filter=143 channel=59
    3, -4, 2, 0, 0, 0, 4, 0, -2,
    -- filter=143 channel=60
    -6, 3, -3, 3, 1, 1, 4, -2, -3,
    -- filter=143 channel=61
    -2, 3, 1, 3, -4, 7, -4, 5, 5,
    -- filter=143 channel=62
    -6, 5, 2, 6, 0, -5, 5, 3, -6,
    -- filter=143 channel=63
    3, -2, 6, -6, 4, 2, 4, -6, 0,
    -- filter=143 channel=64
    5, -5, -4, 5, 7, 2, 7, 0, 3,
    -- filter=143 channel=65
    4, -1, 6, 2, 5, -1, 3, 1, 5,
    -- filter=143 channel=66
    5, -6, 0, 0, -7, 6, -8, 2, 6,
    -- filter=143 channel=67
    4, 2, -4, 0, -4, 0, 5, -4, 0,
    -- filter=143 channel=68
    -3, -5, 7, 0, -3, 0, -2, -4, -3,
    -- filter=143 channel=69
    0, 5, -5, -4, 0, 3, 2, -6, 2,
    -- filter=143 channel=70
    4, -1, 9, 2, 3, 4, 1, 1, 6,
    -- filter=143 channel=71
    -5, 7, 4, 7, 0, 0, -4, 3, 6,
    -- filter=143 channel=72
    2, -7, 2, -6, 4, 4, 3, -5, -2,
    -- filter=143 channel=73
    5, 5, 4, -6, -4, 6, -3, -7, 7,
    -- filter=143 channel=74
    -6, 5, 3, 3, 6, 8, -5, -5, 0,
    -- filter=143 channel=75
    -6, -7, 4, -5, -8, 2, -6, 4, 8,
    -- filter=143 channel=76
    3, 2, -2, -3, -4, 0, 3, -1, -1,
    -- filter=143 channel=77
    6, 5, -4, -5, 6, -6, 3, 4, 0,
    -- filter=143 channel=78
    4, 5, 2, 2, -1, 0, 0, 6, 3,
    -- filter=143 channel=79
    -7, -3, 6, -7, -2, 2, -13, -10, 1,
    -- filter=143 channel=80
    -9, -6, -5, -2, 0, 6, 0, 2, 1,
    -- filter=143 channel=81
    -5, 1, -6, -1, 1, -4, 0, -6, 6,
    -- filter=143 channel=82
    -6, 1, 1, -3, 1, 0, 5, 3, -3,
    -- filter=143 channel=83
    4, 5, 0, 2, -3, 5, -4, 0, -3,
    -- filter=143 channel=84
    -3, -5, -4, -6, 0, 1, 3, -3, 1,
    -- filter=143 channel=85
    -1, -3, 7, -3, -1, -4, -5, 4, 0,
    -- filter=143 channel=86
    6, -4, 9, 3, 3, 0, -2, -1, 1,
    -- filter=143 channel=87
    -2, 3, 0, -2, 0, -4, -3, 0, 6,
    -- filter=143 channel=88
    -4, 7, 4, -4, -4, -6, 1, 9, 7,
    -- filter=143 channel=89
    3, 2, -3, -2, -5, -5, -3, 4, 6,
    -- filter=143 channel=90
    -5, 8, 6, 0, 3, 4, -5, 8, 8,
    -- filter=143 channel=91
    1, -5, -1, 0, 2, 5, 2, -6, 1,
    -- filter=143 channel=92
    2, -3, -6, -2, -4, 6, 0, 3, 0,
    -- filter=143 channel=93
    2, 0, -6, 6, -5, 0, -3, -8, 6,
    -- filter=143 channel=94
    5, -1, 0, 6, -6, -3, 2, -5, 5,
    -- filter=143 channel=95
    -1, 2, -5, -5, 0, -2, 0, -1, -4,
    -- filter=143 channel=96
    0, 4, -6, -4, -3, 3, 1, 1, 5,
    -- filter=143 channel=97
    -4, -1, 6, -4, 4, 7, -3, 5, 0,
    -- filter=143 channel=98
    -6, -4, 1, -7, -1, -3, 4, -3, -5,
    -- filter=143 channel=99
    0, -1, 3, -4, -3, -1, -1, -3, -1,
    -- filter=143 channel=100
    0, -3, 2, 3, 3, 3, -3, -7, 3,
    -- filter=143 channel=101
    -5, 7, 0, -3, 2, 1, -3, 4, -6,
    -- filter=143 channel=102
    -6, -2, 6, 0, 7, -4, -1, 1, -1,
    -- filter=143 channel=103
    -6, 0, -2, 4, -6, 6, -3, 4, 5,
    -- filter=143 channel=104
    4, -5, 3, 0, 0, 0, -6, -4, 1,
    -- filter=143 channel=105
    7, 3, 0, -6, 3, -3, 5, 1, -3,
    -- filter=143 channel=106
    -5, -1, 3, 7, 3, 6, -1, -7, -1,
    -- filter=143 channel=107
    -5, 7, 8, -1, 4, 6, -6, -3, 3,
    -- filter=143 channel=108
    0, -5, 2, 2, 4, -1, 0, -6, 5,
    -- filter=143 channel=109
    -9, 1, 3, -2, -3, 1, -10, -8, -1,
    -- filter=143 channel=110
    -6, 1, 5, 3, -1, 5, -1, -5, 3,
    -- filter=143 channel=111
    -5, -6, -3, -5, 6, 3, -5, -3, -6,
    -- filter=143 channel=112
    0, 0, -1, 0, 0, 6, -5, 0, 0,
    -- filter=143 channel=113
    -7, 0, -1, 5, 6, -6, -3, 1, 7,
    -- filter=143 channel=114
    -5, -7, 1, -4, -8, 1, 0, -8, 8,
    -- filter=143 channel=115
    -2, -4, 7, 4, -3, -4, -6, 3, -5,
    -- filter=143 channel=116
    -2, 1, 0, -6, -5, -6, -8, -1, 1,
    -- filter=143 channel=117
    0, 0, -5, -5, 4, 2, -4, -7, 4,
    -- filter=143 channel=118
    3, -5, 5, 1, 5, 2, -5, -2, 1,
    -- filter=143 channel=119
    0, 0, 6, -4, 7, 0, -7, 0, 3,
    -- filter=143 channel=120
    -3, 9, 0, 3, -5, -5, 3, 0, 0,
    -- filter=143 channel=121
    2, -2, -3, 0, -2, 0, 3, -4, 4,
    -- filter=143 channel=122
    4, 3, -5, 3, 0, -3, 3, 4, 0,
    -- filter=143 channel=123
    -6, 6, 5, 4, 1, 4, 3, -2, 2,
    -- filter=143 channel=124
    -1, -3, 1, 0, 7, -5, -4, -4, 6,
    -- filter=143 channel=125
    3, -8, -1, -8, -6, -5, 0, -4, -2,
    -- filter=143 channel=126
    5, 0, 6, 5, -7, 0, -6, 0, -2,
    -- filter=143 channel=127
    6, -5, 3, -6, 1, 3, -4, 1, -6,
    -- filter=144 channel=0
    2, 5, 4, 0, -2, -5, 1, -11, 1,
    -- filter=144 channel=1
    6, -2, 0, -3, 3, 5, 0, 0, -2,
    -- filter=144 channel=2
    -1, -5, -6, 3, 1, -4, 3, 7, 5,
    -- filter=144 channel=3
    -7, 4, 5, 4, 3, 8, 2, -4, -3,
    -- filter=144 channel=4
    -6, 2, 0, 0, -2, -10, 12, 5, 5,
    -- filter=144 channel=5
    10, 3, 9, 2, -4, 6, -7, 0, 3,
    -- filter=144 channel=6
    -7, -7, 4, -5, 1, 6, -3, 8, 1,
    -- filter=144 channel=7
    -5, -4, 7, 0, 0, -1, -6, 3, -5,
    -- filter=144 channel=8
    -6, 4, 3, -3, -7, 2, 0, -8, -6,
    -- filter=144 channel=9
    -2, 2, -6, 2, -3, 2, 0, 4, -1,
    -- filter=144 channel=10
    6, 2, -1, -5, -4, 0, 0, 7, 1,
    -- filter=144 channel=11
    2, -3, -8, 6, -3, -1, 0, 11, 4,
    -- filter=144 channel=12
    0, -2, 0, -6, -7, -3, -7, -8, 3,
    -- filter=144 channel=13
    -3, 0, 0, -5, 2, -6, 8, 6, -4,
    -- filter=144 channel=14
    2, 7, 0, 5, -6, -2, -1, -1, 3,
    -- filter=144 channel=15
    -1, 0, -5, 7, 0, 0, 13, 8, -6,
    -- filter=144 channel=16
    -3, -3, 4, 0, 1, -1, 0, -2, 5,
    -- filter=144 channel=17
    5, 0, -4, 1, 0, 7, -2, -3, 0,
    -- filter=144 channel=18
    -6, -11, 1, 7, -1, -4, 13, 7, -6,
    -- filter=144 channel=19
    -4, 2, -6, -5, -2, 6, 7, 2, 2,
    -- filter=144 channel=20
    -1, -7, -7, -5, -4, 4, 19, 8, 10,
    -- filter=144 channel=21
    1, 8, -3, 6, 7, 5, 0, -1, -1,
    -- filter=144 channel=22
    3, -2, 4, -4, 2, -5, 4, 0, -5,
    -- filter=144 channel=23
    -6, -10, 4, -1, -14, 0, 16, -3, -8,
    -- filter=144 channel=24
    0, -3, 0, -5, 3, 5, 1, -6, -1,
    -- filter=144 channel=25
    1, -2, 1, 5, -9, -10, 10, 2, 1,
    -- filter=144 channel=26
    3, 3, 4, 6, 2, -3, -2, 4, 4,
    -- filter=144 channel=27
    0, -9, 1, 1, -2, -9, 10, -1, -9,
    -- filter=144 channel=28
    1, 3, 4, 5, -7, -6, 3, 2, 4,
    -- filter=144 channel=29
    -3, 0, -5, -2, 1, -5, 10, 5, 4,
    -- filter=144 channel=30
    -1, 7, 5, 0, 0, -2, -2, 3, -6,
    -- filter=144 channel=31
    -1, 9, -4, 3, 4, -3, 7, 4, 2,
    -- filter=144 channel=32
    4, -8, -3, -1, -3, -1, 8, -3, -6,
    -- filter=144 channel=33
    4, -5, -4, -7, -3, 1, 10, -7, -5,
    -- filter=144 channel=34
    -1, 0, -3, -11, -10, -1, 0, -6, -6,
    -- filter=144 channel=35
    -3, 6, -1, -6, -4, 3, -3, 6, 6,
    -- filter=144 channel=36
    0, -3, 3, 8, -4, -2, 9, 7, 10,
    -- filter=144 channel=37
    9, 7, 10, 6, -6, 6, -11, -12, 2,
    -- filter=144 channel=38
    0, 5, -4, -7, -6, -7, 5, -6, -1,
    -- filter=144 channel=39
    -8, 2, -6, 1, -4, -2, 8, 0, 3,
    -- filter=144 channel=40
    -5, -2, -2, 0, 6, 0, 1, -1, -4,
    -- filter=144 channel=41
    4, -9, -5, 7, -2, -3, -5, -3, -4,
    -- filter=144 channel=42
    -2, -3, 2, -1, 6, 4, 5, -6, -6,
    -- filter=144 channel=43
    3, -5, 9, -3, -7, -4, 6, 7, 1,
    -- filter=144 channel=44
    3, 7, 2, 0, -6, -6, 0, -4, 2,
    -- filter=144 channel=45
    -6, 5, -3, -6, 7, 2, -1, 0, -1,
    -- filter=144 channel=46
    1, 0, -5, -6, -4, 0, -2, 0, 2,
    -- filter=144 channel=47
    9, 10, 12, -4, 3, 7, -9, -4, 0,
    -- filter=144 channel=48
    10, 5, -3, 0, -4, 2, -3, -2, 0,
    -- filter=144 channel=49
    -8, 2, -7, 1, -3, -6, 11, -1, -6,
    -- filter=144 channel=50
    -3, 2, 0, -3, -4, -3, 9, 2, 0,
    -- filter=144 channel=51
    2, -4, 1, -4, 7, 0, 4, -6, -5,
    -- filter=144 channel=52
    -7, 2, 4, -3, 0, 1, 0, 3, -8,
    -- filter=144 channel=53
    3, 1, -6, 3, -1, 1, 9, 8, -5,
    -- filter=144 channel=54
    -1, -4, -3, 0, 6, 0, 1, 1, -2,
    -- filter=144 channel=55
    3, -14, 4, -2, -6, -6, 13, 13, -1,
    -- filter=144 channel=56
    6, -4, 5, 4, -6, 1, 0, -4, 0,
    -- filter=144 channel=57
    -2, -3, -4, 9, 0, -3, 3, 7, -1,
    -- filter=144 channel=58
    0, 2, 3, -5, -3, 1, -3, -3, -7,
    -- filter=144 channel=59
    -5, 5, 0, -3, -6, -4, -1, -1, 5,
    -- filter=144 channel=60
    2, -4, 0, 0, 3, 0, 5, -2, -2,
    -- filter=144 channel=61
    -4, -3, 1, 3, -7, 6, 5, 3, 2,
    -- filter=144 channel=62
    -5, 0, 5, -2, 4, 6, 0, -5, 1,
    -- filter=144 channel=63
    -4, 6, -3, 2, 3, -5, 4, -3, 1,
    -- filter=144 channel=64
    2, -5, 5, 2, 3, 1, 8, -1, -3,
    -- filter=144 channel=65
    -2, -4, 0, 7, 4, 0, -3, 6, 0,
    -- filter=144 channel=66
    0, -2, 0, -5, 2, 2, 2, 0, 1,
    -- filter=144 channel=67
    5, -4, -5, -4, -6, -2, 7, -4, -4,
    -- filter=144 channel=68
    2, -3, -7, 5, -4, -6, 3, 2, -1,
    -- filter=144 channel=69
    -4, 3, 2, -4, 1, 7, -6, 0, -6,
    -- filter=144 channel=70
    -9, 0, 0, -9, -10, -2, 7, -8, 1,
    -- filter=144 channel=71
    6, -4, -4, 5, 4, -2, 4, 5, -7,
    -- filter=144 channel=72
    -5, -2, -5, -6, -8, -6, 0, 2, -1,
    -- filter=144 channel=73
    -1, -10, -6, 1, -5, -2, 10, 5, -3,
    -- filter=144 channel=74
    -8, 6, -5, -2, 0, -6, -2, -5, -7,
    -- filter=144 channel=75
    -2, 9, -1, 1, -8, -1, 3, -4, -1,
    -- filter=144 channel=76
    -5, -2, -5, 9, -4, -4, 9, 13, 7,
    -- filter=144 channel=77
    -4, 6, 2, 7, 4, 4, 1, 0, 6,
    -- filter=144 channel=78
    3, 4, 4, 4, 4, 7, 0, -1, -4,
    -- filter=144 channel=79
    -7, -11, -2, 0, -13, -7, 11, 0, 0,
    -- filter=144 channel=80
    0, -7, 7, 4, 2, -8, 9, 3, -3,
    -- filter=144 channel=81
    -2, -2, -6, 1, 0, -2, -4, -3, -2,
    -- filter=144 channel=82
    -7, 4, -5, -1, 4, 7, 6, 0, 0,
    -- filter=144 channel=83
    1, 4, -8, 3, 6, 3, -5, 5, -6,
    -- filter=144 channel=84
    3, -5, -4, -3, 3, -2, 0, 5, 0,
    -- filter=144 channel=85
    1, 0, 2, -7, 6, -3, 1, 0, 0,
    -- filter=144 channel=86
    -7, 4, 0, -9, -6, -5, -6, -5, 6,
    -- filter=144 channel=87
    -1, -7, 0, -1, 1, 2, 7, 3, 6,
    -- filter=144 channel=88
    5, -1, -1, -5, 0, 0, -4, -4, 4,
    -- filter=144 channel=89
    0, 1, 3, 0, 0, -8, 10, 10, 0,
    -- filter=144 channel=90
    6, 0, 6, -5, 2, 4, 6, -4, 4,
    -- filter=144 channel=91
    -4, -8, -8, 7, -8, -4, 8, 8, -2,
    -- filter=144 channel=92
    -1, -6, -1, 5, 3, -6, 3, -1, 0,
    -- filter=144 channel=93
    8, 3, 2, -4, -1, 6, 0, -5, -6,
    -- filter=144 channel=94
    6, -1, 4, -3, -2, -7, -5, -4, -7,
    -- filter=144 channel=95
    -1, -2, 3, -6, 4, -3, 0, 7, 0,
    -- filter=144 channel=96
    7, 0, -7, -1, -4, 5, -4, 6, 5,
    -- filter=144 channel=97
    -7, 3, 0, -6, -7, -4, 1, -4, -3,
    -- filter=144 channel=98
    -5, -6, -2, 0, -6, -6, 0, -3, 1,
    -- filter=144 channel=99
    0, -2, -3, -1, -9, 0, 7, 8, -8,
    -- filter=144 channel=100
    3, -3, -5, 0, 0, -7, 5, 2, 1,
    -- filter=144 channel=101
    -5, 3, -6, 1, 0, 4, 4, 4, 10,
    -- filter=144 channel=102
    -1, -7, -6, -6, -7, -2, -3, -5, -3,
    -- filter=144 channel=103
    9, 0, 0, -5, 3, 2, -3, -8, -8,
    -- filter=144 channel=104
    1, -3, 0, -3, 3, 1, 7, 0, -6,
    -- filter=144 channel=105
    -2, 2, 4, 6, 5, 3, 10, 9, 3,
    -- filter=144 channel=106
    -6, -8, 3, 0, 2, -5, 6, -2, 4,
    -- filter=144 channel=107
    -7, -5, 4, 2, 1, 1, -1, -2, 0,
    -- filter=144 channel=108
    6, -5, 0, 3, -6, -5, 4, 2, 7,
    -- filter=144 channel=109
    0, -12, 4, 5, -5, -12, 7, 5, -2,
    -- filter=144 channel=110
    -2, -6, -2, -9, -5, -1, 8, 6, -6,
    -- filter=144 channel=111
    0, 5, -4, 1, 5, -4, 4, -2, -6,
    -- filter=144 channel=112
    3, -1, 2, -4, 2, 4, 3, -1, 2,
    -- filter=144 channel=113
    1, 2, -3, -4, 2, 0, 1, -5, -1,
    -- filter=144 channel=114
    -6, -11, 0, 3, -12, -5, 5, -2, 2,
    -- filter=144 channel=115
    -6, 0, -1, 0, -4, 0, -2, 6, 3,
    -- filter=144 channel=116
    6, 0, 4, -1, 5, -12, 7, 2, -2,
    -- filter=144 channel=117
    -3, -6, -5, 2, 2, 0, -2, 3, -1,
    -- filter=144 channel=118
    -4, 6, 0, -4, 5, 0, 6, 2, 4,
    -- filter=144 channel=119
    0, -3, -7, -7, -4, 0, 3, -10, -7,
    -- filter=144 channel=120
    -11, -9, 3, 3, -12, -16, 13, 0, -10,
    -- filter=144 channel=121
    0, -8, 6, 0, 0, 0, -3, -2, -5,
    -- filter=144 channel=122
    11, 11, 5, 1, -3, 1, -1, -7, 1,
    -- filter=144 channel=123
    -6, -2, -3, -7, 0, 2, 2, 0, -5,
    -- filter=144 channel=124
    -6, -9, 2, 1, 4, 1, 6, 0, 8,
    -- filter=144 channel=125
    -5, -7, 6, -3, 0, -11, 10, 2, 1,
    -- filter=144 channel=126
    -1, 4, 2, -2, -8, -2, 9, 9, 0,
    -- filter=144 channel=127
    -6, 6, -6, -4, -2, 2, 2, 2, -2,
    -- filter=145 channel=0
    7, -11, -8, 4, -10, -9, 6, -1, 0,
    -- filter=145 channel=1
    6, 8, 0, -3, 2, 0, -2, 4, 10,
    -- filter=145 channel=2
    5, -5, 6, 5, -4, -4, -4, -6, 5,
    -- filter=145 channel=3
    2, -14, -5, -4, -14, -4, 8, 2, -3,
    -- filter=145 channel=4
    0, 2, -5, -10, -9, -12, 7, -11, -8,
    -- filter=145 channel=5
    -14, -10, 0, -1, -5, -11, -5, 0, 2,
    -- filter=145 channel=6
    5, -10, 1, -1, -3, -10, 2, -15, -7,
    -- filter=145 channel=7
    0, 4, -5, -4, 6, 7, -4, -1, -6,
    -- filter=145 channel=8
    5, -1, 7, -2, -3, -7, -1, -3, 0,
    -- filter=145 channel=9
    0, -3, 3, 0, 3, -1, -10, -6, 0,
    -- filter=145 channel=10
    -9, -10, -8, -7, 0, 4, 2, 5, -5,
    -- filter=145 channel=11
    -9, -15, 0, -2, -13, -3, 4, -2, 0,
    -- filter=145 channel=12
    2, -8, 13, -2, -6, 0, 1, -6, 1,
    -- filter=145 channel=13
    8, -10, 7, -3, 0, 3, 12, 3, 0,
    -- filter=145 channel=14
    0, 7, -1, -5, 0, -5, -2, 5, -4,
    -- filter=145 channel=15
    -3, -11, -11, 0, -16, -7, 9, -2, 1,
    -- filter=145 channel=16
    -10, -10, 6, -5, -7, 5, -7, -1, 8,
    -- filter=145 channel=17
    4, -6, 1, -4, 3, 6, -1, 0, -6,
    -- filter=145 channel=18
    7, -6, -6, -3, -19, -11, 0, -6, -3,
    -- filter=145 channel=19
    5, 0, 0, -5, 1, 0, -4, 4, -6,
    -- filter=145 channel=20
    -2, -15, -17, -3, -27, -10, -3, -16, -4,
    -- filter=145 channel=21
    -7, 0, 2, 2, 6, 10, -11, 0, 10,
    -- filter=145 channel=22
    0, -2, -9, -2, -8, -10, 6, 4, 0,
    -- filter=145 channel=23
    1, -6, -1, -4, -10, -10, 18, 3, 4,
    -- filter=145 channel=24
    -2, -4, -6, -4, -6, 4, 4, 4, 1,
    -- filter=145 channel=25
    4, -9, 8, -7, 3, 10, -5, 3, 15,
    -- filter=145 channel=26
    -6, 1, -7, 1, -1, -2, -8, -12, 0,
    -- filter=145 channel=27
    7, 0, 2, 3, 7, 14, -3, 9, 15,
    -- filter=145 channel=28
    3, -3, 4, 7, -6, 0, -3, 0, 1,
    -- filter=145 channel=29
    -10, -7, -13, 5, -9, -13, 0, -4, -4,
    -- filter=145 channel=30
    6, -3, 3, 2, 6, 0, -2, 7, -5,
    -- filter=145 channel=31
    -6, 2, 4, 1, 23, 6, -6, 7, 9,
    -- filter=145 channel=32
    8, 0, -9, -6, -11, -3, 3, -10, -2,
    -- filter=145 channel=33
    0, -4, -5, -2, 5, -4, 0, -1, 11,
    -- filter=145 channel=34
    1, -9, 0, -4, -8, -14, -1, -8, 9,
    -- filter=145 channel=35
    -3, 4, -2, 4, -2, -3, -5, -6, 4,
    -- filter=145 channel=36
    5, -7, 7, 7, 0, -5, 2, 1, -5,
    -- filter=145 channel=37
    0, 16, 15, -1, 13, 3, 3, -2, 9,
    -- filter=145 channel=38
    -1, -6, -2, -10, 5, -2, 1, -1, 8,
    -- filter=145 channel=39
    0, -5, 1, -2, -12, -14, -4, -5, -12,
    -- filter=145 channel=40
    1, -4, -3, -1, -4, -5, 6, 2, -1,
    -- filter=145 channel=41
    3, -9, 8, -8, -33, -2, -1, -20, -1,
    -- filter=145 channel=42
    8, 5, 0, -7, 8, 2, 0, 3, -4,
    -- filter=145 channel=43
    8, -15, -20, -10, -19, -12, 2, 4, -7,
    -- filter=145 channel=44
    -5, -1, 15, -1, 9, 13, 1, 10, 4,
    -- filter=145 channel=45
    3, 4, -2, 7, 5, 5, -2, 2, 4,
    -- filter=145 channel=46
    1, 0, 2, 6, 3, -1, 0, 2, 2,
    -- filter=145 channel=47
    -20, -5, 11, -3, 9, 19, -14, 13, 6,
    -- filter=145 channel=48
    5, 5, 14, -1, 22, 9, 0, 9, 9,
    -- filter=145 channel=49
    8, 0, 0, 0, -12, -13, 7, -2, -7,
    -- filter=145 channel=50
    5, 10, -5, 1, 5, 2, 3, 3, 2,
    -- filter=145 channel=51
    -2, -4, 5, 5, -5, -4, 7, 2, -6,
    -- filter=145 channel=52
    2, -4, 3, 7, -6, 0, 0, -9, 0,
    -- filter=145 channel=53
    3, -5, 1, -4, -9, 1, -4, -7, -9,
    -- filter=145 channel=54
    0, 4, 4, -6, -5, 2, 0, -5, -4,
    -- filter=145 channel=55
    -2, -6, -7, 7, -4, -9, 11, 0, 0,
    -- filter=145 channel=56
    5, 2, 2, -6, -15, 1, 3, 0, 5,
    -- filter=145 channel=57
    -6, 0, 5, -8, -11, 0, 1, -3, -5,
    -- filter=145 channel=58
    -7, -3, -6, -3, -14, -14, 0, 2, 0,
    -- filter=145 channel=59
    -10, -7, 10, -8, 16, 14, -8, 8, 4,
    -- filter=145 channel=60
    -4, -6, 1, -3, -5, -7, 6, 1, -2,
    -- filter=145 channel=61
    -6, -9, 2, 1, -1, 2, -1, 1, -2,
    -- filter=145 channel=62
    -6, -1, -3, 0, -7, -7, 7, 0, -4,
    -- filter=145 channel=63
    -12, -4, 0, -4, -10, -9, -11, -13, -4,
    -- filter=145 channel=64
    -9, -1, -3, 4, -9, 0, -1, -6, -1,
    -- filter=145 channel=65
    6, 3, 5, -6, 3, 5, 0, 2, 3,
    -- filter=145 channel=66
    -12, -6, 4, -3, -22, -2, -6, -10, 8,
    -- filter=145 channel=67
    0, 0, 4, 0, -8, 1, 6, -8, 5,
    -- filter=145 channel=68
    3, -5, -7, 0, 3, -6, 2, 4, -8,
    -- filter=145 channel=69
    -2, -5, 6, -5, -3, -6, -5, -11, 0,
    -- filter=145 channel=70
    9, 2, 9, 0, 10, 7, 11, 10, 14,
    -- filter=145 channel=71
    2, -4, -1, 6, 7, 4, 5, 2, 2,
    -- filter=145 channel=72
    0, 2, -1, 5, 18, 1, 2, 9, -1,
    -- filter=145 channel=73
    -3, -1, 5, -5, 0, -3, -2, 3, 3,
    -- filter=145 channel=74
    -4, 2, 14, 4, 0, 4, -2, -4, 9,
    -- filter=145 channel=75
    7, -3, 5, -2, -8, 7, -2, 2, 16,
    -- filter=145 channel=76
    -2, -7, -14, 0, -7, -5, 0, -11, -9,
    -- filter=145 channel=77
    -6, -3, -2, -2, -4, -2, 3, 6, 7,
    -- filter=145 channel=78
    -6, -1, -7, 3, -10, -1, -5, -3, -1,
    -- filter=145 channel=79
    16, -1, -5, -9, -18, -13, 15, -5, 10,
    -- filter=145 channel=80
    -8, -7, 3, -9, 14, 16, -9, 7, 13,
    -- filter=145 channel=81
    2, -3, -5, 6, 3, -1, 6, -4, 1,
    -- filter=145 channel=82
    -3, -4, 0, 0, -5, 5, 5, -6, -3,
    -- filter=145 channel=83
    -8, 2, 3, 0, 3, 8, -4, -3, 0,
    -- filter=145 channel=84
    0, -4, 4, -4, -12, 0, 0, -6, 3,
    -- filter=145 channel=85
    3, -6, 0, 4, -4, 0, 6, 4, 2,
    -- filter=145 channel=86
    -2, -14, 7, -7, -9, 2, 2, -12, -2,
    -- filter=145 channel=87
    2, -8, -1, -2, -18, -13, -5, -17, 1,
    -- filter=145 channel=88
    -7, -10, 7, -1, 2, -8, 7, 0, -3,
    -- filter=145 channel=89
    -2, -6, 0, 0, 3, 5, 0, 2, 5,
    -- filter=145 channel=90
    -7, -15, 4, 7, 1, -6, 6, 1, 2,
    -- filter=145 channel=91
    3, 0, 1, 2, -4, 0, 13, -2, 5,
    -- filter=145 channel=92
    -5, 2, -3, 0, -9, -7, -8, 1, 5,
    -- filter=145 channel=93
    -8, -2, 1, -8, 13, 11, -8, -4, 7,
    -- filter=145 channel=94
    -5, 5, 7, -5, -2, 2, 0, 6, -5,
    -- filter=145 channel=95
    -7, 5, -2, 1, -3, -4, 0, -1, -5,
    -- filter=145 channel=96
    -7, -6, -1, 2, 7, -2, -5, -5, 4,
    -- filter=145 channel=97
    0, -7, -4, 2, 0, 4, 7, 8, -2,
    -- filter=145 channel=98
    -5, -11, 5, -16, 0, 2, -10, -3, 11,
    -- filter=145 channel=99
    -3, -13, 0, 3, 0, -7, 7, -2, 0,
    -- filter=145 channel=100
    -9, -4, -10, 3, -7, -11, -3, -3, -9,
    -- filter=145 channel=101
    8, 1, -9, -7, -12, -13, 5, -8, -9,
    -- filter=145 channel=102
    5, 4, 1, 1, 5, 5, -3, 1, 6,
    -- filter=145 channel=103
    -9, -13, 2, 2, 9, 8, -21, 13, 15,
    -- filter=145 channel=104
    -9, 1, 4, 0, 19, 19, -13, -4, 8,
    -- filter=145 channel=105
    -6, -14, -8, -8, -2, -7, 0, -5, -7,
    -- filter=145 channel=106
    0, -5, 2, 2, -1, -4, -2, -3, -2,
    -- filter=145 channel=107
    -2, -10, -7, 0, -22, -10, 8, -18, -11,
    -- filter=145 channel=108
    -9, -12, -6, 2, -7, -4, -9, -8, -7,
    -- filter=145 channel=109
    -6, -11, 2, -4, 1, 11, -1, -1, 4,
    -- filter=145 channel=110
    -9, -15, -2, 3, 4, -4, -9, -3, -7,
    -- filter=145 channel=111
    -6, -8, -7, 2, -6, -1, -5, -8, 6,
    -- filter=145 channel=112
    0, -1, 0, -2, 9, 7, -8, 9, 0,
    -- filter=145 channel=113
    3, 0, 6, -6, 7, 10, -5, 9, 12,
    -- filter=145 channel=114
    9, -16, -9, -5, -29, -19, 7, -18, -19,
    -- filter=145 channel=115
    4, -7, 1, 3, 3, -2, -2, -7, -7,
    -- filter=145 channel=116
    1, 0, 0, -4, -4, 6, 2, 2, 2,
    -- filter=145 channel=117
    9, -3, -2, 0, 0, 1, 9, 9, 7,
    -- filter=145 channel=118
    -4, 6, 7, -3, -3, 4, -4, -6, 5,
    -- filter=145 channel=119
    -3, -5, 7, -2, -20, -4, -6, -10, 0,
    -- filter=145 channel=120
    -3, 3, 11, -4, -3, -1, 9, 5, -5,
    -- filter=145 channel=121
    -8, -2, -1, 0, -3, -2, 5, -2, 2,
    -- filter=145 channel=122
    -10, -10, 4, -1, 28, 27, -17, 0, 18,
    -- filter=145 channel=123
    0, -7, 7, -5, 1, -5, -5, 0, 6,
    -- filter=145 channel=124
    -6, 1, -7, 1, -11, 0, -3, -6, -13,
    -- filter=145 channel=125
    -6, -11, 2, -4, 16, 9, -2, 4, 0,
    -- filter=145 channel=126
    -3, -7, -3, 2, -11, 2, -3, 3, -3,
    -- filter=145 channel=127
    -8, -6, -5, -4, -1, 0, 5, 1, 1,
    -- filter=146 channel=0
    -8, 0, -3, 0, -1, 4, 0, 10, -4,
    -- filter=146 channel=1
    4, 1, 0, -7, 13, 10, 7, 12, 7,
    -- filter=146 channel=2
    -4, 5, -5, -5, 3, -8, 6, 1, -3,
    -- filter=146 channel=3
    0, -4, 7, -6, 1, -6, 1, 13, 7,
    -- filter=146 channel=4
    3, 8, 0, -2, 0, -4, -4, -2, -3,
    -- filter=146 channel=5
    -7, -3, 12, 0, 5, 4, 4, 0, 2,
    -- filter=146 channel=6
    -2, -8, -6, 1, -11, 2, -9, -1, -7,
    -- filter=146 channel=7
    5, 3, 3, 0, 5, 7, -6, 2, 6,
    -- filter=146 channel=8
    -3, 3, 4, -1, 2, -7, 1, 5, -2,
    -- filter=146 channel=9
    -1, 5, 0, 5, 5, 0, -5, -8, -8,
    -- filter=146 channel=10
    -6, -4, -1, 6, -6, -2, 3, -2, -11,
    -- filter=146 channel=11
    -9, -3, -7, -8, -6, -8, 1, 1, -15,
    -- filter=146 channel=12
    5, 8, 1, -6, 5, -5, -3, 11, 6,
    -- filter=146 channel=13
    -1, -4, -3, 7, -2, 0, 6, -4, -3,
    -- filter=146 channel=14
    -7, -2, -3, 2, -4, -2, -6, 1, 0,
    -- filter=146 channel=15
    -15, -5, -19, -6, -6, -10, 5, -5, -14,
    -- filter=146 channel=16
    -1, 8, 6, 0, 9, 0, 3, 4, 2,
    -- filter=146 channel=17
    -3, -2, -3, 2, -4, 5, -5, 2, -5,
    -- filter=146 channel=18
    -10, -11, -22, -10, -7, -19, 10, -8, -18,
    -- filter=146 channel=19
    -1, -1, 2, 3, 7, -4, -5, -1, 6,
    -- filter=146 channel=20
    -9, -16, -10, 2, -11, -8, -4, -10, -20,
    -- filter=146 channel=21
    7, 5, 5, 1, 9, 0, -11, 0, 2,
    -- filter=146 channel=22
    3, 0, -5, -2, 1, -6, 1, 1, -7,
    -- filter=146 channel=23
    -6, -23, -13, 3, -7, -12, 5, -6, -16,
    -- filter=146 channel=24
    0, 0, -2, 6, 6, 5, -5, -2, 1,
    -- filter=146 channel=25
    6, 13, -3, 12, 4, -5, 9, 2, -6,
    -- filter=146 channel=26
    7, 0, -2, 1, 5, 6, -8, -4, 2,
    -- filter=146 channel=27
    11, -1, -14, 11, -5, -10, 7, 0, -19,
    -- filter=146 channel=28
    -5, -4, -2, 1, 1, -3, -1, -7, -5,
    -- filter=146 channel=29
    -4, -7, -10, -2, -4, -3, -3, -7, -15,
    -- filter=146 channel=30
    7, 0, 4, 6, -5, -8, 7, 5, -2,
    -- filter=146 channel=31
    -5, -5, -6, -3, -4, -22, -6, -12, -14,
    -- filter=146 channel=32
    -5, -9, -14, 4, 1, -3, 3, -7, -13,
    -- filter=146 channel=33
    -7, -5, -6, 5, -2, -12, 4, -4, -3,
    -- filter=146 channel=34
    2, -1, -2, -1, -6, 1, 1, -5, 11,
    -- filter=146 channel=35
    1, 6, -2, 0, 2, 0, 0, 4, -3,
    -- filter=146 channel=36
    -6, 3, 0, -11, -8, -5, -2, -9, -11,
    -- filter=146 channel=37
    6, 11, 12, -4, 7, -2, -7, 2, 2,
    -- filter=146 channel=38
    1, 2, -9, -2, -6, -9, -2, 3, -3,
    -- filter=146 channel=39
    1, -7, -4, -3, 0, -2, -3, -10, -6,
    -- filter=146 channel=40
    0, -9, -11, 0, -5, -10, 5, 1, -13,
    -- filter=146 channel=41
    7, 18, 9, 7, 3, 11, 13, 8, 17,
    -- filter=146 channel=42
    -3, 7, -6, -2, 9, 1, -5, 4, 0,
    -- filter=146 channel=43
    -12, -13, 0, -8, -10, -12, -2, 1, 6,
    -- filter=146 channel=44
    0, 9, 10, 0, 1, 1, 0, 7, -6,
    -- filter=146 channel=45
    -3, -9, -3, 0, -6, -3, -8, -8, -7,
    -- filter=146 channel=46
    5, 5, 3, -4, 3, 7, -1, 0, 2,
    -- filter=146 channel=47
    10, 5, 6, 11, 19, 3, 4, 0, -1,
    -- filter=146 channel=48
    6, 10, 0, 6, 11, -6, 0, 2, 0,
    -- filter=146 channel=49
    -7, 2, -6, -4, -11, 0, 3, -7, -1,
    -- filter=146 channel=50
    2, -3, -8, 0, 3, -4, -4, -6, -3,
    -- filter=146 channel=51
    4, -2, -4, 0, 2, 6, 4, -4, 0,
    -- filter=146 channel=52
    4, -3, -3, -6, -3, 0, 0, -3, 6,
    -- filter=146 channel=53
    1, -4, -1, -8, 0, -2, 0, -5, -12,
    -- filter=146 channel=54
    0, 1, -6, -7, 1, 4, -1, -3, 7,
    -- filter=146 channel=55
    -13, -20, -26, 0, -13, -14, -3, -17, -13,
    -- filter=146 channel=56
    9, 1, 0, 8, -6, -5, -4, -1, 1,
    -- filter=146 channel=57
    5, 0, 5, 0, 5, -4, 8, 5, -3,
    -- filter=146 channel=58
    -10, -4, 9, 2, 5, 5, -10, -3, 6,
    -- filter=146 channel=59
    9, 1, -2, 14, 0, -4, 6, -5, -9,
    -- filter=146 channel=60
    -4, 5, -2, 0, 1, -7, -4, 4, -1,
    -- filter=146 channel=61
    -4, -4, 4, 0, -3, 1, 2, 1, 2,
    -- filter=146 channel=62
    -5, -7, 7, -5, -6, 0, 6, -1, -2,
    -- filter=146 channel=63
    -5, -3, 7, -9, 6, 0, 0, 3, -3,
    -- filter=146 channel=64
    1, -9, 0, -9, -5, 2, 2, -11, -2,
    -- filter=146 channel=65
    1, 2, -1, -3, -6, -5, 4, -3, -5,
    -- filter=146 channel=66
    -4, 11, 8, -6, 8, 0, 7, 2, 5,
    -- filter=146 channel=67
    6, 0, 6, 3, 4, -6, 2, 0, -3,
    -- filter=146 channel=68
    2, -2, 0, 3, 4, -3, -5, -7, 4,
    -- filter=146 channel=69
    -2, 3, 4, 5, -2, 0, -1, 7, 6,
    -- filter=146 channel=70
    -1, -5, -16, 2, -2, -8, 3, -8, -6,
    -- filter=146 channel=71
    0, 1, -5, 4, -6, -5, 0, -2, 3,
    -- filter=146 channel=72
    3, 4, -10, 4, -3, -8, -2, -5, -21,
    -- filter=146 channel=73
    0, -1, -2, 7, 3, -8, -1, -2, -6,
    -- filter=146 channel=74
    1, -12, -7, -1, -3, -11, -5, -9, 3,
    -- filter=146 channel=75
    -10, 9, 4, -7, 6, 9, 1, 17, 8,
    -- filter=146 channel=76
    -15, -16, -17, -6, -18, -4, -6, -7, -12,
    -- filter=146 channel=77
    5, -3, 7, 0, -5, -2, -1, -2, 1,
    -- filter=146 channel=78
    -1, 2, -4, -3, -1, 0, 1, -6, 5,
    -- filter=146 channel=79
    -11, -10, -20, 0, 0, -20, 10, -3, -16,
    -- filter=146 channel=80
    6, 4, -5, 10, 8, -2, 4, -5, -12,
    -- filter=146 channel=81
    5, 1, -5, -6, -3, 3, 0, 1, 1,
    -- filter=146 channel=82
    -7, -4, 6, 3, 1, -4, -6, 3, 4,
    -- filter=146 channel=83
    -1, 7, 0, 4, 1, -6, 4, 2, -4,
    -- filter=146 channel=84
    -2, 0, -5, 2, 0, -3, 4, 2, -4,
    -- filter=146 channel=85
    -2, 0, -1, 1, 7, 0, -3, 7, 2,
    -- filter=146 channel=86
    0, -9, -3, 3, 0, 1, -7, 0, 0,
    -- filter=146 channel=87
    1, -4, -8, -9, -9, -1, -1, 1, -3,
    -- filter=146 channel=88
    -5, -5, 4, -8, -14, -4, -2, -16, -10,
    -- filter=146 channel=89
    4, 1, -16, 0, -2, -2, 3, -1, -13,
    -- filter=146 channel=90
    -9, 0, 4, -1, -2, 3, -3, -5, -1,
    -- filter=146 channel=91
    5, -8, -13, 3, -2, -13, 2, -5, -16,
    -- filter=146 channel=92
    6, 5, 6, 4, -8, -3, 2, -3, -1,
    -- filter=146 channel=93
    3, 12, 11, 0, 9, 8, -4, 3, 8,
    -- filter=146 channel=94
    -5, -2, 6, 1, -6, 4, 0, 1, 1,
    -- filter=146 channel=95
    -1, 6, -5, -5, 5, 6, 1, 0, -7,
    -- filter=146 channel=96
    2, 4, -4, -3, 2, -2, 0, -2, -4,
    -- filter=146 channel=97
    1, 5, 2, 0, -1, -8, -3, 0, 6,
    -- filter=146 channel=98
    9, 0, -11, 10, 6, -2, 15, 6, -16,
    -- filter=146 channel=99
    2, -12, -16, 1, -18, -12, -3, -14, -12,
    -- filter=146 channel=100
    2, -2, 2, 7, 2, 7, 3, -3, 6,
    -- filter=146 channel=101
    5, 5, -5, -6, -7, 0, 1, 9, -1,
    -- filter=146 channel=102
    0, 0, -5, -7, -5, -5, 4, 2, -6,
    -- filter=146 channel=103
    -3, 10, 7, 15, 14, 1, 0, 3, 4,
    -- filter=146 channel=104
    4, -3, -8, 4, -2, -6, -3, -8, -15,
    -- filter=146 channel=105
    -8, -6, 0, 4, 0, 0, -2, -8, -3,
    -- filter=146 channel=106
    -6, -6, -9, 0, 0, -8, -6, -5, -6,
    -- filter=146 channel=107
    -7, -14, -13, -13, -13, -3, 0, -13, -11,
    -- filter=146 channel=108
    -4, 1, 8, 2, 8, 10, 9, -1, 8,
    -- filter=146 channel=109
    5, 1, -8, 16, -1, -6, 12, 2, -9,
    -- filter=146 channel=110
    -11, -8, -8, -3, -5, -3, -1, -10, -6,
    -- filter=146 channel=111
    5, -4, -1, -1, 0, -5, 6, 1, 8,
    -- filter=146 channel=112
    1, -13, 4, 2, -10, 2, 9, 1, -2,
    -- filter=146 channel=113
    -2, -7, -3, 9, 1, -8, 1, -3, -5,
    -- filter=146 channel=114
    -3, -18, -11, -2, -7, -22, 7, 1, -14,
    -- filter=146 channel=115
    -3, -4, 1, -3, 0, 4, 1, 2, 3,
    -- filter=146 channel=116
    2, 7, -4, 9, -7, -6, 0, 1, -12,
    -- filter=146 channel=117
    -6, -3, 1, 5, -5, 0, 1, -2, -5,
    -- filter=146 channel=118
    2, -6, -5, 4, -2, -1, -2, -5, 0,
    -- filter=146 channel=119
    11, -5, -2, -1, -1, 1, 10, -4, 11,
    -- filter=146 channel=120
    6, -15, -8, 7, -14, -17, 0, -9, -6,
    -- filter=146 channel=121
    -3, 10, 8, 2, 8, 6, 9, 9, -5,
    -- filter=146 channel=122
    13, 21, 15, 12, 11, 4, 5, -2, 8,
    -- filter=146 channel=123
    2, -1, 0, 1, 3, 2, 8, -1, -4,
    -- filter=146 channel=124
    2, -1, -10, -6, -1, -8, -6, -9, -9,
    -- filter=146 channel=125
    7, -2, -6, 6, -6, -4, -3, -3, -20,
    -- filter=146 channel=126
    -6, 10, -10, -2, 6, 0, 4, 13, -7,
    -- filter=146 channel=127
    5, -4, -2, -4, -4, 6, -4, 1, -5,
    -- filter=147 channel=0
    0, 4, 5, 4, 4, -14, 3, -8, -7,
    -- filter=147 channel=1
    1, 2, 2, 11, 12, -18, 4, -4, -30,
    -- filter=147 channel=2
    2, 0, -4, 6, -2, 0, 3, 0, 2,
    -- filter=147 channel=3
    -3, -7, -2, -4, -9, -10, -7, -3, 0,
    -- filter=147 channel=4
    -10, -6, 3, -10, -11, 2, -1, -6, 4,
    -- filter=147 channel=5
    6, 25, 12, 6, 11, -13, 9, 5, -16,
    -- filter=147 channel=6
    -1, 4, -4, 0, 4, 2, 7, -2, -1,
    -- filter=147 channel=7
    5, 3, -6, -6, -2, -6, 0, 0, 4,
    -- filter=147 channel=8
    0, 5, -7, 0, 2, 1, -7, -3, 6,
    -- filter=147 channel=9
    10, 5, 7, 0, -2, -1, 10, 5, 0,
    -- filter=147 channel=10
    -2, -5, -1, -8, -9, -5, 4, 0, 0,
    -- filter=147 channel=11
    3, -6, -1, -9, -9, 8, -1, -1, 24,
    -- filter=147 channel=12
    -2, -8, 7, 0, -6, -2, 0, -6, -2,
    -- filter=147 channel=13
    -3, -20, -1, -12, -3, 6, -4, 2, 12,
    -- filter=147 channel=14
    -6, 6, -3, 3, -4, 5, -4, -7, 0,
    -- filter=147 channel=15
    6, -13, 6, -13, -6, 4, -2, 5, 22,
    -- filter=147 channel=16
    0, 13, -5, 0, 3, 0, 2, 7, -13,
    -- filter=147 channel=17
    -3, 6, 2, -3, -6, -3, 5, -3, 3,
    -- filter=147 channel=18
    6, -16, 0, -9, -3, 12, 10, 5, 14,
    -- filter=147 channel=19
    -3, -5, -4, -4, -2, -7, -5, 7, 1,
    -- filter=147 channel=20
    3, -8, 3, -12, -9, 20, -6, -6, 28,
    -- filter=147 channel=21
    11, 10, -3, 1, 15, -5, -4, -3, -10,
    -- filter=147 channel=22
    0, 3, -10, 0, 3, -6, 5, 3, 2,
    -- filter=147 channel=23
    -8, -18, -3, -21, -14, 19, 4, 0, 23,
    -- filter=147 channel=24
    2, -3, 6, -5, 0, -5, -2, 2, 1,
    -- filter=147 channel=25
    -2, -3, 2, 0, -7, 1, 2, -10, -4,
    -- filter=147 channel=26
    0, 12, -2, 11, 15, 7, 11, 13, -11,
    -- filter=147 channel=27
    -7, -1, 2, -3, 2, 1, 12, -1, 7,
    -- filter=147 channel=28
    0, -2, 0, 4, 3, 2, 5, 0, -2,
    -- filter=147 channel=29
    6, -7, 15, -8, 0, 18, 9, 0, 18,
    -- filter=147 channel=30
    7, 12, 5, 2, 7, -6, 7, -6, -7,
    -- filter=147 channel=31
    -5, 1, -1, 2, 13, 9, 0, 10, 10,
    -- filter=147 channel=32
    4, -14, -7, -10, -1, 11, -4, -6, 11,
    -- filter=147 channel=33
    4, -1, -4, 4, -3, -6, 6, 0, 0,
    -- filter=147 channel=34
    -7, -9, -12, -14, -10, -7, -4, -10, 1,
    -- filter=147 channel=35
    -4, 2, 0, 3, 3, -2, -6, -6, -5,
    -- filter=147 channel=36
    -7, -6, -5, -3, -4, 7, -8, -8, 6,
    -- filter=147 channel=37
    -3, 8, -1, 0, 10, -10, -7, 0, -28,
    -- filter=147 channel=38
    -2, -6, 3, 0, 0, 0, 0, 0, 4,
    -- filter=147 channel=39
    6, -3, -1, -7, 2, 6, 6, 0, 6,
    -- filter=147 channel=40
    6, 2, 2, -3, 1, 9, 0, -1, 13,
    -- filter=147 channel=41
    -1, -14, -19, -16, -14, -18, -8, -14, -16,
    -- filter=147 channel=42
    4, 2, 8, 8, 10, -3, 7, -2, 2,
    -- filter=147 channel=43
    -1, -13, 2, -4, -6, -7, -9, -8, 1,
    -- filter=147 channel=44
    1, 7, 4, 9, 6, -14, -7, -5, -18,
    -- filter=147 channel=45
    -4, 10, -4, -3, -1, 4, 1, -4, 0,
    -- filter=147 channel=46
    -1, 4, 0, 0, 0, -9, 0, -6, 1,
    -- filter=147 channel=47
    1, 5, 0, 17, 13, -7, -2, -4, -16,
    -- filter=147 channel=48
    -2, -3, -8, 15, 10, 0, 3, -4, -6,
    -- filter=147 channel=49
    0, -5, 10, -1, -3, 8, 0, 4, 14,
    -- filter=147 channel=50
    0, 2, 0, -3, -1, 8, 7, 6, 3,
    -- filter=147 channel=51
    -2, -6, 6, -6, -3, -2, 1, -6, -5,
    -- filter=147 channel=52
    2, -10, 3, -1, -13, -5, -13, -8, 9,
    -- filter=147 channel=53
    -2, 3, 7, -1, -10, 9, 5, -2, 9,
    -- filter=147 channel=54
    -6, -5, 3, 1, 5, 2, -1, 0, 0,
    -- filter=147 channel=55
    3, -22, 1, -4, -5, 10, 9, -4, 27,
    -- filter=147 channel=56
    -4, -5, -4, -1, -3, -8, 0, 4, -4,
    -- filter=147 channel=57
    -8, -6, -10, -7, 0, -4, 6, -6, -8,
    -- filter=147 channel=58
    7, 11, -1, 12, 10, 5, 7, -5, -3,
    -- filter=147 channel=59
    3, 4, -6, 8, 3, -1, 11, -4, -9,
    -- filter=147 channel=60
    0, -1, 4, -1, 1, -6, 2, -5, -4,
    -- filter=147 channel=61
    -3, -2, 5, -3, 0, -4, -8, -7, 0,
    -- filter=147 channel=62
    0, 4, 6, -7, 0, -5, -5, 3, 2,
    -- filter=147 channel=63
    2, 7, 3, 1, 7, -6, 0, -1, -8,
    -- filter=147 channel=64
    -5, -5, -6, -9, -5, -4, -6, 7, -5,
    -- filter=147 channel=65
    -5, -6, -5, 3, 6, 7, -5, 7, -7,
    -- filter=147 channel=66
    -6, -13, -7, -10, -14, -8, -12, -16, -2,
    -- filter=147 channel=67
    0, -2, -2, -1, -1, 2, 6, -4, -6,
    -- filter=147 channel=68
    4, -4, 7, 1, -5, 1, 2, 5, -4,
    -- filter=147 channel=69
    -4, -2, 2, 6, 0, -4, -1, -2, -6,
    -- filter=147 channel=70
    -12, -11, 0, -4, -3, 0, -6, -3, 13,
    -- filter=147 channel=71
    -1, 0, -9, -7, 0, -10, 1, -1, 3,
    -- filter=147 channel=72
    3, -5, 0, -2, -4, 4, 6, 7, 2,
    -- filter=147 channel=73
    -6, 0, 3, -3, -4, 2, 8, 4, 15,
    -- filter=147 channel=74
    -8, -7, -10, -2, 2, -4, -6, 4, 10,
    -- filter=147 channel=75
    4, 8, -6, 3, -1, -13, 2, -6, -21,
    -- filter=147 channel=76
    9, -9, -1, -4, -13, 7, -1, 6, 23,
    -- filter=147 channel=77
    -6, 3, 0, 7, -7, 0, -1, 4, -3,
    -- filter=147 channel=78
    -5, 1, 6, -5, 7, -4, 6, 2, 5,
    -- filter=147 channel=79
    3, -20, 1, -4, -14, 15, 6, -2, 18,
    -- filter=147 channel=80
    10, 3, -2, 3, 13, -5, 7, 6, -9,
    -- filter=147 channel=81
    -1, 2, 1, -4, 0, -7, -4, 3, 1,
    -- filter=147 channel=82
    3, -6, 5, -5, 0, -4, 2, 4, 3,
    -- filter=147 channel=83
    -2, 2, -5, 5, 9, -2, 11, 6, 1,
    -- filter=147 channel=84
    -2, -5, 0, -7, 3, 2, -2, -1, 9,
    -- filter=147 channel=85
    4, -2, 0, 0, -4, 3, -3, 3, -3,
    -- filter=147 channel=86
    1, -3, 2, -5, -1, 5, 0, -4, 5,
    -- filter=147 channel=87
    -4, -5, 0, -4, -11, 0, -5, -3, 5,
    -- filter=147 channel=88
    -5, -6, -5, -1, 7, -2, 1, -5, 1,
    -- filter=147 channel=89
    2, -7, 1, 0, -14, 11, 2, -3, 18,
    -- filter=147 channel=90
    -4, -2, 0, -6, -4, -8, -6, -3, 4,
    -- filter=147 channel=91
    -10, -12, 7, -6, -9, 13, 0, 0, 9,
    -- filter=147 channel=92
    -7, -1, -1, 2, -8, 1, 0, -4, 0,
    -- filter=147 channel=93
    -1, 16, 10, 14, 18, -9, 6, -9, -25,
    -- filter=147 channel=94
    0, -7, 2, 6, 6, -1, 0, 7, 1,
    -- filter=147 channel=95
    4, 3, 1, 0, -6, 7, 6, -3, 0,
    -- filter=147 channel=96
    6, -5, 4, -5, -1, 7, 6, -1, -3,
    -- filter=147 channel=97
    0, 2, -9, 0, -5, 0, 1, -6, -5,
    -- filter=147 channel=98
    -7, 0, -9, 1, -1, 5, 5, 0, -2,
    -- filter=147 channel=99
    -7, -9, -6, -6, -8, 4, -3, 0, 17,
    -- filter=147 channel=100
    -3, 0, -1, 2, -8, 1, -8, 0, -1,
    -- filter=147 channel=101
    -8, -3, 0, 2, -8, -6, 0, -2, 4,
    -- filter=147 channel=102
    0, 5, 0, 7, -1, 2, 7, -5, -3,
    -- filter=147 channel=103
    0, 11, -3, 15, 14, -20, -4, -2, -22,
    -- filter=147 channel=104
    -2, 0, 0, 12, 1, 2, -1, 9, -3,
    -- filter=147 channel=105
    3, -6, 4, 1, -3, 8, 3, 0, 8,
    -- filter=147 channel=106
    -6, -8, 2, -2, 0, 7, 7, 2, 5,
    -- filter=147 channel=107
    -4, -10, 6, -3, -7, 15, -6, 0, 16,
    -- filter=147 channel=108
    0, 9, -4, 5, 1, -7, -1, -2, 0,
    -- filter=147 channel=109
    -7, 0, -6, 7, -2, 5, 2, 5, 9,
    -- filter=147 channel=110
    -3, 0, -2, -7, 3, 9, -10, 7, 1,
    -- filter=147 channel=111
    7, 4, 2, 5, 1, 3, -5, 3, -3,
    -- filter=147 channel=112
    1, -7, 0, 0, 0, -4, 0, 4, -6,
    -- filter=147 channel=113
    -1, -14, -1, -1, -9, -2, -5, 0, 6,
    -- filter=147 channel=114
    8, -4, 3, -2, 0, 8, 10, -9, 1,
    -- filter=147 channel=115
    0, 5, 4, 0, 6, -7, 3, -1, 4,
    -- filter=147 channel=116
    -1, -6, 0, 8, 3, 5, 10, -6, 5,
    -- filter=147 channel=117
    1, 0, -7, 6, -3, -6, -7, 5, 2,
    -- filter=147 channel=118
    -1, -5, -3, 1, -5, 0, -4, -4, -1,
    -- filter=147 channel=119
    -15, -5, -14, -3, -2, -6, -5, 0, 0,
    -- filter=147 channel=120
    -3, 0, 1, -1, 9, 17, 4, -2, 24,
    -- filter=147 channel=121
    -2, -12, -5, -7, 0, 0, 5, -3, 4,
    -- filter=147 channel=122
    1, 18, -1, 21, 13, -19, -3, -2, -31,
    -- filter=147 channel=123
    -2, 2, 0, 2, 0, -8, 0, 1, -8,
    -- filter=147 channel=124
    -4, -4, 3, -3, 0, 11, 8, 3, 6,
    -- filter=147 channel=125
    0, -1, 6, -3, 6, 0, 3, 5, 3,
    -- filter=147 channel=126
    11, -9, 0, 0, -4, -5, 5, 2, 0,
    -- filter=147 channel=127
    -4, 0, 2, 3, 2, 3, -6, 4, -2,
    -- filter=148 channel=0
    2, 2, -4, 10, 13, -30, 12, 23, -25,
    -- filter=148 channel=1
    -2, 6, -17, -2, 13, -27, 11, 7, -14,
    -- filter=148 channel=2
    2, -4, 2, 4, -5, -2, -7, -2, 5,
    -- filter=148 channel=3
    -6, 4, 8, -17, 2, 5, -8, 1, -8,
    -- filter=148 channel=4
    -4, -1, -2, -16, 0, -3, -11, 7, -1,
    -- filter=148 channel=5
    3, 1, -9, 11, 9, -9, 21, 1, -9,
    -- filter=148 channel=6
    -4, 6, 3, 0, 5, 6, -5, -2, -2,
    -- filter=148 channel=7
    -4, 6, 0, 0, 0, -1, -3, 1, -1,
    -- filter=148 channel=8
    -7, 5, -1, 5, 1, -2, 0, -1, -1,
    -- filter=148 channel=9
    11, -1, -1, 13, -1, -3, 11, -10, -6,
    -- filter=148 channel=10
    8, -4, -4, 8, -7, -2, 12, -10, -10,
    -- filter=148 channel=11
    -5, 9, 6, 2, 1, 16, -8, 0, 8,
    -- filter=148 channel=12
    0, 0, -9, 0, 7, -6, -3, -3, 3,
    -- filter=148 channel=13
    4, -7, -4, 9, -3, -17, 10, 5, -1,
    -- filter=148 channel=14
    0, 2, -4, 0, -4, 4, -5, 0, -1,
    -- filter=148 channel=15
    -5, -8, -2, 3, 3, -4, 9, -5, 1,
    -- filter=148 channel=16
    5, 1, -1, 14, -10, -14, 1, 1, -7,
    -- filter=148 channel=17
    6, -2, 4, -1, 6, 5, 1, 5, 4,
    -- filter=148 channel=18
    5, -2, -2, 12, 1, -13, 17, 7, -4,
    -- filter=148 channel=19
    1, -3, -5, 1, 6, 1, 0, 0, -5,
    -- filter=148 channel=20
    -6, 8, 14, -8, 0, 14, -2, -2, 18,
    -- filter=148 channel=21
    10, -12, -7, 6, -17, -19, 4, -10, -12,
    -- filter=148 channel=22
    -7, 0, -6, 5, -1, -3, 4, 6, -11,
    -- filter=148 channel=23
    -14, -9, 16, 3, -26, -4, 6, -7, 4,
    -- filter=148 channel=24
    0, -7, -5, -2, -5, 1, 3, 7, 6,
    -- filter=148 channel=25
    19, -3, -5, 16, -11, -19, 24, 0, -6,
    -- filter=148 channel=26
    6, 4, -8, 12, -3, -3, -4, 1, -4,
    -- filter=148 channel=27
    3, -10, -4, 20, -18, -33, 26, -13, -26,
    -- filter=148 channel=28
    -2, -7, -6, 7, 3, 2, -4, -2, 0,
    -- filter=148 channel=29
    -9, 4, 5, -10, 13, 12, 1, 0, 5,
    -- filter=148 channel=30
    11, 4, 0, 11, 0, -13, 11, 0, -5,
    -- filter=148 channel=31
    1, -5, 12, 21, -33, -16, 22, -21, 2,
    -- filter=148 channel=32
    9, 0, -1, 10, 0, -20, 12, 2, -11,
    -- filter=148 channel=33
    0, 1, -7, 15, -2, -22, 8, 0, -23,
    -- filter=148 channel=34
    0, 3, -8, 7, 0, -10, 9, 6, -9,
    -- filter=148 channel=35
    5, 4, 4, 0, 5, 1, 2, -1, 0,
    -- filter=148 channel=36
    0, -6, 4, -6, -12, 7, -8, -2, 0,
    -- filter=148 channel=37
    6, -2, -9, 8, 10, -25, 4, 11, -17,
    -- filter=148 channel=38
    3, 2, 5, 12, -4, -9, 18, -8, 0,
    -- filter=148 channel=39
    0, 7, 5, -10, 1, 10, -8, 3, 6,
    -- filter=148 channel=40
    -9, -3, 1, -11, 5, 1, -6, 1, -2,
    -- filter=148 channel=41
    14, -3, -15, 31, 30, -23, 24, 29, -13,
    -- filter=148 channel=42
    9, 4, 1, 5, 11, -4, 6, 4, 1,
    -- filter=148 channel=43
    -12, -2, 11, -11, 12, -1, 4, 8, 2,
    -- filter=148 channel=44
    13, -6, -3, 6, -11, -18, 5, -1, -11,
    -- filter=148 channel=45
    0, -2, 0, 3, -1, 7, 3, -2, -6,
    -- filter=148 channel=46
    -1, 1, 1, 9, 8, -9, 1, 4, 0,
    -- filter=148 channel=47
    18, 5, 0, 20, -10, -19, 12, -1, -14,
    -- filter=148 channel=48
    14, -9, -3, 19, -10, -28, 22, -3, -3,
    -- filter=148 channel=49
    -7, 0, 1, -4, 6, -8, 0, 9, -9,
    -- filter=148 channel=50
    7, -1, 2, 13, -9, -4, 7, -12, -8,
    -- filter=148 channel=51
    -4, -3, 0, 1, -3, 6, -2, 0, 2,
    -- filter=148 channel=52
    -9, -8, -3, 0, -13, 6, -6, -9, -5,
    -- filter=148 channel=53
    -7, 0, 7, -1, 0, 0, -5, 5, -2,
    -- filter=148 channel=54
    0, -6, -7, -5, 4, -3, 3, -5, 0,
    -- filter=148 channel=55
    -2, -9, 4, -1, -11, 0, 5, -5, 4,
    -- filter=148 channel=56
    0, -2, -11, 1, 4, -2, 8, -5, -5,
    -- filter=148 channel=57
    4, -1, -6, 3, -2, 0, 5, 7, -4,
    -- filter=148 channel=58
    8, -3, 0, 8, 13, -11, 1, 19, -11,
    -- filter=148 channel=59
    8, -7, -9, 16, -10, -22, 24, 6, -13,
    -- filter=148 channel=60
    -3, 1, -1, 0, 6, 0, -3, 3, -6,
    -- filter=148 channel=61
    4, 3, 2, 2, 0, 4, -5, -6, 6,
    -- filter=148 channel=62
    -4, -2, -4, -7, -3, 0, 0, -5, 1,
    -- filter=148 channel=63
    -1, -5, -3, 3, 13, -6, 11, 1, 0,
    -- filter=148 channel=64
    1, 1, 5, 0, 0, 4, -8, -2, 0,
    -- filter=148 channel=65
    -1, -6, -1, 7, -2, 0, 6, 7, 2,
    -- filter=148 channel=66
    -3, -5, -11, 7, 6, -12, 1, 5, -3,
    -- filter=148 channel=67
    -5, 6, -5, -6, -2, 6, 5, 4, -3,
    -- filter=148 channel=68
    4, -6, -2, -8, -2, 4, -1, 3, 0,
    -- filter=148 channel=69
    -2, 3, 3, 4, 4, -1, 4, -4, -8,
    -- filter=148 channel=70
    -2, -7, 2, 5, -8, -3, 1, -4, -11,
    -- filter=148 channel=71
    -10, -1, 0, -4, 2, 7, -1, -3, 0,
    -- filter=148 channel=72
    10, -2, 11, 16, -11, -13, 8, -12, -2,
    -- filter=148 channel=73
    4, 0, -1, 0, -8, -4, 4, 4, -3,
    -- filter=148 channel=74
    3, -12, -3, 5, -11, -16, 7, -11, -10,
    -- filter=148 channel=75
    5, 7, -1, 15, 18, -18, 18, 17, -23,
    -- filter=148 channel=76
    -3, 3, 4, -1, -2, 16, -13, -7, 10,
    -- filter=148 channel=77
    -5, -4, -8, 5, 4, -7, 7, 0, -5,
    -- filter=148 channel=78
    -1, 0, 4, 5, -3, -9, 8, 0, -9,
    -- filter=148 channel=79
    -2, -7, -11, 15, 0, -25, 19, 11, -16,
    -- filter=148 channel=80
    13, -13, 6, 19, -21, -16, 33, 2, -1,
    -- filter=148 channel=81
    3, -2, -4, -6, 0, 1, -2, -5, 0,
    -- filter=148 channel=82
    -1, 5, 0, -4, -1, 3, 2, 1, -7,
    -- filter=148 channel=83
    5, 2, -6, 3, -5, 2, 8, -3, 0,
    -- filter=148 channel=84
    5, 0, -8, 6, -4, -8, 0, 0, 0,
    -- filter=148 channel=85
    -4, -5, 6, 3, -2, 3, -3, -7, 6,
    -- filter=148 channel=86
    8, -5, -13, 7, -2, -16, 1, 5, -10,
    -- filter=148 channel=87
    3, 4, 5, 2, -7, 9, 3, 0, 1,
    -- filter=148 channel=88
    -8, -5, -1, -5, -12, 6, -6, -18, 0,
    -- filter=148 channel=89
    12, -5, 9, 10, -7, -14, 7, 0, -6,
    -- filter=148 channel=90
    -2, -10, 0, 0, -12, 9, -1, -9, 5,
    -- filter=148 channel=91
    1, -11, 1, 1, -18, -13, 0, 5, -3,
    -- filter=148 channel=92
    -2, -4, -2, -1, -5, -4, 8, 5, -3,
    -- filter=148 channel=93
    10, 3, -6, 9, 0, -17, 8, 6, -8,
    -- filter=148 channel=94
    -2, -5, 0, -6, -4, -1, -6, 4, -6,
    -- filter=148 channel=95
    6, 3, -2, 7, -2, -5, 7, 0, 1,
    -- filter=148 channel=96
    9, 2, -4, 7, -2, -6, 2, 4, 0,
    -- filter=148 channel=97
    1, 0, 3, 2, 5, 6, -10, -4, -8,
    -- filter=148 channel=98
    14, -5, -4, 25, 4, -22, 30, 4, -6,
    -- filter=148 channel=99
    0, -12, 11, 9, -25, -2, 17, -11, 0,
    -- filter=148 channel=100
    10, 9, 5, 1, 9, 5, 3, 7, -6,
    -- filter=148 channel=101
    0, -6, -6, -8, -6, 0, -2, -2, 8,
    -- filter=148 channel=102
    6, 4, 2, 1, 1, -6, 4, -7, -3,
    -- filter=148 channel=103
    6, -3, -1, 14, -8, -9, 22, -5, -11,
    -- filter=148 channel=104
    13, -5, 1, 19, -19, -17, 20, -12, -12,
    -- filter=148 channel=105
    -8, 11, 14, -11, 0, 5, 0, -1, 14,
    -- filter=148 channel=106
    -2, 0, -2, -7, 6, -3, -9, 3, 9,
    -- filter=148 channel=107
    -5, 1, 7, -8, 2, 6, -12, -4, 4,
    -- filter=148 channel=108
    13, -2, -5, 6, 9, -3, 1, 0, -4,
    -- filter=148 channel=109
    14, -4, -11, 27, -14, -20, 24, -7, -20,
    -- filter=148 channel=110
    2, 0, 8, 3, -11, 1, 0, -6, 2,
    -- filter=148 channel=111
    9, -9, -4, 0, -4, -10, 3, -2, -5,
    -- filter=148 channel=112
    0, -6, 0, 14, -17, -15, 10, -2, -19,
    -- filter=148 channel=113
    0, -10, 2, 6, -8, -10, 10, -1, -11,
    -- filter=148 channel=114
    -1, 6, -16, 7, 5, -34, 12, 15, -17,
    -- filter=148 channel=115
    7, -4, -5, -6, -1, 5, -6, 1, -7,
    -- filter=148 channel=116
    13, -2, -3, 5, -15, -16, 21, -1, -1,
    -- filter=148 channel=117
    -3, -3, 3, 5, 3, 3, 4, -7, 0,
    -- filter=148 channel=118
    -1, 5, -8, 5, 1, -1, 6, 2, 2,
    -- filter=148 channel=119
    -1, 1, -3, 13, -2, -7, 11, 7, -2,
    -- filter=148 channel=120
    3, -10, -4, 16, -26, -11, 0, -17, -16,
    -- filter=148 channel=121
    -1, 0, -6, 1, 0, -3, 12, 3, -8,
    -- filter=148 channel=122
    17, 0, -9, 15, -19, -26, 14, -12, -16,
    -- filter=148 channel=123
    0, 5, 5, 0, 4, 0, 0, 1, -2,
    -- filter=148 channel=124
    -4, -2, 0, -6, 2, 13, 2, 6, 4,
    -- filter=148 channel=125
    16, -7, -4, 19, -18, -13, 25, -7, -15,
    -- filter=148 channel=126
    0, 4, 2, 10, 0, -11, 5, 2, -11,
    -- filter=148 channel=127
    0, -3, -5, 8, 0, 3, -2, 8, -1,
    -- filter=149 channel=0
    3, 0, 9, -2, 6, -9, -2, 7, -8,
    -- filter=149 channel=1
    0, -3, 6, 0, 12, 1, -4, -1, -10,
    -- filter=149 channel=2
    1, 0, 2, -2, 1, 2, 0, 0, 7,
    -- filter=149 channel=3
    -4, -10, -4, 7, -4, -4, -14, 0, 0,
    -- filter=149 channel=4
    2, -8, -5, 0, 7, -2, 4, -11, 5,
    -- filter=149 channel=5
    0, 0, -3, 7, 3, 1, -5, 5, -9,
    -- filter=149 channel=6
    -2, 6, -5, 0, 4, -3, 7, 6, -7,
    -- filter=149 channel=7
    0, 3, 2, -5, 0, -4, 6, 2, -1,
    -- filter=149 channel=8
    0, 4, -5, -1, 0, -1, 3, 5, 1,
    -- filter=149 channel=9
    -3, -5, -2, 6, 0, -4, -5, -4, 1,
    -- filter=149 channel=10
    0, -1, -1, 0, 0, 2, -4, 7, -5,
    -- filter=149 channel=11
    -1, 1, 5, -3, 3, -2, 11, -7, 0,
    -- filter=149 channel=12
    3, 3, 6, 0, 2, 8, 3, 9, -6,
    -- filter=149 channel=13
    -7, -5, 3, 0, 5, 2, -7, 16, -3,
    -- filter=149 channel=14
    3, -4, 0, 4, 0, 4, 0, 3, -5,
    -- filter=149 channel=15
    -3, -4, 8, 2, 3, -2, -4, 12, -11,
    -- filter=149 channel=16
    -1, 5, 1, 7, 6, 2, 4, 6, 2,
    -- filter=149 channel=17
    2, 2, -4, 3, 7, 1, 1, 3, 4,
    -- filter=149 channel=18
    -5, -5, 4, -8, 6, -4, 3, 15, -11,
    -- filter=149 channel=19
    -1, -1, 5, 0, 3, 6, -5, 2, -3,
    -- filter=149 channel=20
    1, 0, -3, 1, -6, -1, 7, 6, -10,
    -- filter=149 channel=21
    0, 6, 1, -3, 8, -3, 7, 0, -11,
    -- filter=149 channel=22
    -4, 9, 3, -4, 3, -1, 3, -4, -7,
    -- filter=149 channel=23
    -2, -2, 2, -2, 6, -13, -4, 5, 2,
    -- filter=149 channel=24
    -2, -6, 0, -4, 2, 0, 7, -6, 7,
    -- filter=149 channel=25
    -2, 4, 3, -10, 10, -9, -7, 13, -16,
    -- filter=149 channel=26
    1, 3, 1, 1, 0, 0, 4, -4, -3,
    -- filter=149 channel=27
    -10, 6, 6, 0, 9, -4, 6, 7, -4,
    -- filter=149 channel=28
    0, 5, 0, 4, 5, -6, 1, 0, -1,
    -- filter=149 channel=29
    -9, -7, 6, 3, -3, -6, 2, 9, -9,
    -- filter=149 channel=30
    0, 2, -2, 0, 2, -5, -2, 6, -3,
    -- filter=149 channel=31
    -13, 0, 4, -7, 5, -10, 1, 2, -5,
    -- filter=149 channel=32
    -6, 4, 7, -2, 17, -8, -5, 14, -8,
    -- filter=149 channel=33
    -4, -1, 16, -1, 7, -8, -5, 6, -16,
    -- filter=149 channel=34
    -7, -3, 4, 2, 2, 1, 0, -1, 11,
    -- filter=149 channel=35
    3, -7, -2, -2, 3, 2, -1, 3, 2,
    -- filter=149 channel=36
    -7, -5, -4, -1, 9, 2, 9, 8, -1,
    -- filter=149 channel=37
    -6, 2, 0, 0, 7, 0, 4, -4, -11,
    -- filter=149 channel=38
    -8, 0, 10, 0, 1, 1, 0, 6, -5,
    -- filter=149 channel=39
    -3, 0, 2, 0, -3, -3, 6, 4, 2,
    -- filter=149 channel=40
    -4, 1, -5, -5, -2, 3, 0, 4, 2,
    -- filter=149 channel=41
    16, -10, 0, 6, 5, 4, -5, 25, 0,
    -- filter=149 channel=42
    -3, -2, 6, 1, 0, 0, 4, -6, 4,
    -- filter=149 channel=43
    4, -5, 3, 0, -4, 5, -7, -5, -9,
    -- filter=149 channel=44
    1, 0, 7, -7, 13, -2, 0, 0, -6,
    -- filter=149 channel=45
    -7, 0, -2, 3, 2, 0, 4, -3, -6,
    -- filter=149 channel=46
    0, 7, 2, -4, 0, 7, 5, -7, 3,
    -- filter=149 channel=47
    -2, 0, -3, -5, 12, -2, -4, 14, -14,
    -- filter=149 channel=48
    -5, 7, 1, -3, 6, -13, 3, -3, -8,
    -- filter=149 channel=49
    -9, 3, -8, -7, 3, 0, 8, -5, -5,
    -- filter=149 channel=50
    -9, 4, 0, 2, 7, -11, 5, -8, -5,
    -- filter=149 channel=51
    6, 3, -2, 4, 6, 3, 4, -2, 0,
    -- filter=149 channel=52
    -2, -4, 5, 3, 12, -7, 0, -2, -3,
    -- filter=149 channel=53
    -5, 4, 2, -7, -5, 2, 7, 4, 3,
    -- filter=149 channel=54
    0, -5, 0, -7, 5, -5, 5, 6, -3,
    -- filter=149 channel=55
    -5, -7, 5, -1, 8, -9, 3, 17, -4,
    -- filter=149 channel=56
    -6, 9, -7, 1, 10, -4, -2, 4, 0,
    -- filter=149 channel=57
    2, -3, -3, -1, 5, -5, 4, 7, -6,
    -- filter=149 channel=58
    -1, 0, -2, -1, -1, -3, 9, -3, 0,
    -- filter=149 channel=59
    -4, -4, 7, -11, 14, 1, 3, 15, -12,
    -- filter=149 channel=60
    -5, -4, -2, -6, 4, 3, 0, 5, 7,
    -- filter=149 channel=61
    -6, 1, 2, 0, 10, -6, 5, 2, -2,
    -- filter=149 channel=62
    0, 0, 3, 1, -4, -1, -4, 5, -5,
    -- filter=149 channel=63
    -4, 0, -4, 3, 4, 0, -2, -1, 4,
    -- filter=149 channel=64
    0, 0, 1, 2, 0, 2, 0, -3, 3,
    -- filter=149 channel=65
    -3, -6, -6, 3, 5, 3, 3, 7, -3,
    -- filter=149 channel=66
    9, -7, -1, 0, 11, 1, 0, 20, 3,
    -- filter=149 channel=67
    3, 6, -3, -1, 5, 6, 4, 4, -4,
    -- filter=149 channel=68
    -6, 5, -5, -3, -2, 3, 0, 3, 4,
    -- filter=149 channel=69
    0, -2, -2, 0, -4, -3, -7, 3, -2,
    -- filter=149 channel=70
    -8, -1, 4, -1, 0, 1, 5, 0, 0,
    -- filter=149 channel=71
    1, -4, -5, -6, 4, -3, -8, 3, -5,
    -- filter=149 channel=72
    -7, -2, 9, -4, -1, -13, -2, 6, -14,
    -- filter=149 channel=73
    -12, 0, 2, 2, 11, -8, 10, -2, -3,
    -- filter=149 channel=74
    -2, 0, -1, 1, 3, -11, 0, 3, 5,
    -- filter=149 channel=75
    2, 5, 4, -3, 2, -1, 0, 6, -8,
    -- filter=149 channel=76
    -6, 1, -2, -6, 0, 4, 0, 11, -6,
    -- filter=149 channel=77
    -7, 6, 0, 4, 3, 1, 2, 3, -5,
    -- filter=149 channel=78
    -2, 6, 0, 7, 3, 1, 9, -5, -5,
    -- filter=149 channel=79
    -7, 6, 10, -9, 6, -3, -3, 20, -17,
    -- filter=149 channel=80
    -3, 5, 4, -7, 6, -4, -1, 7, -10,
    -- filter=149 channel=81
    2, 0, 0, 5, 3, -1, 6, 6, 6,
    -- filter=149 channel=82
    -2, 3, -6, 0, 4, -3, -3, 6, -2,
    -- filter=149 channel=83
    -7, -4, -1, 0, -6, 2, 7, -1, 0,
    -- filter=149 channel=84
    -7, -1, -4, 1, 16, -5, 0, 0, -5,
    -- filter=149 channel=85
    0, 2, -5, 4, -4, 2, 7, -6, -2,
    -- filter=149 channel=86
    -7, 0, 0, -1, 5, 4, 2, -1, -7,
    -- filter=149 channel=87
    5, -1, -4, 1, 0, -5, 10, 0, 3,
    -- filter=149 channel=88
    0, 0, 0, 6, 4, -10, -2, 0, 2,
    -- filter=149 channel=89
    -4, -5, 3, -12, 10, -7, -5, 11, -3,
    -- filter=149 channel=90
    -3, 5, -9, 1, 0, -2, 6, 5, 5,
    -- filter=149 channel=91
    -12, 6, -4, -3, 7, -13, 0, 0, 1,
    -- filter=149 channel=92
    -2, -3, -2, 0, -7, -4, 2, -7, 3,
    -- filter=149 channel=93
    -2, 7, -4, -7, 9, 0, -3, 4, -3,
    -- filter=149 channel=94
    -2, 3, -1, 7, 1, -7, 6, -4, -5,
    -- filter=149 channel=95
    -5, 6, -4, 3, 2, -2, 4, 1, -6,
    -- filter=149 channel=96
    2, 2, 2, -7, -5, -2, -6, 5, -6,
    -- filter=149 channel=97
    3, -10, 5, -3, -1, 5, -8, -6, -3,
    -- filter=149 channel=98
    -10, 3, 5, -8, 17, -13, -7, 12, -13,
    -- filter=149 channel=99
    -6, 1, 6, -7, 3, -6, 12, 6, -6,
    -- filter=149 channel=100
    2, 0, -3, 8, 2, 7, 4, -2, 5,
    -- filter=149 channel=101
    2, -5, -5, 9, 6, -8, -7, -8, 3,
    -- filter=149 channel=102
    3, -4, -6, 3, -1, 3, 5, 1, -5,
    -- filter=149 channel=103
    -6, 1, -3, -3, 5, -12, -8, 2, -9,
    -- filter=149 channel=104
    -10, 1, 0, 3, 0, -8, 8, 0, -15,
    -- filter=149 channel=105
    -2, -4, 4, -4, -1, -1, 9, -3, -4,
    -- filter=149 channel=106
    -4, -2, -5, 4, -7, -1, 4, -5, -1,
    -- filter=149 channel=107
    -7, -5, -5, 0, 7, -10, 5, 0, 4,
    -- filter=149 channel=108
    8, 3, 2, 4, -1, 4, -4, -2, -4,
    -- filter=149 channel=109
    -2, 0, 1, -9, 10, -14, 4, 12, -10,
    -- filter=149 channel=110
    -7, 4, 7, 3, 4, -3, 0, 9, -2,
    -- filter=149 channel=111
    -1, 5, 0, 1, -1, 8, 4, 8, 0,
    -- filter=149 channel=112
    -10, -1, -4, 0, -2, -6, -2, 0, -7,
    -- filter=149 channel=113
    -7, 4, 3, -5, 2, -7, -10, 10, -2,
    -- filter=149 channel=114
    -11, 0, -2, -7, 10, -9, 0, 14, -15,
    -- filter=149 channel=115
    -4, 7, -6, 2, -3, 3, 5, 0, 0,
    -- filter=149 channel=116
    -11, -1, 0, 0, 11, -6, -3, 5, -8,
    -- filter=149 channel=117
    5, 0, 4, -4, 8, 4, -7, -3, 1,
    -- filter=149 channel=118
    -7, 5, 6, -2, 7, 3, -3, 4, -1,
    -- filter=149 channel=119
    1, 10, -3, 8, 2, 1, 12, 6, 4,
    -- filter=149 channel=120
    -16, 0, 6, -3, 15, -18, 17, -10, -9,
    -- filter=149 channel=121
    3, -2, -1, 1, -2, 9, -3, 13, -2,
    -- filter=149 channel=122
    5, 8, -1, -4, 17, -12, -2, 10, -7,
    -- filter=149 channel=123
    1, 6, -4, 7, 2, -3, 5, 0, 5,
    -- filter=149 channel=124
    5, -2, 0, -3, -5, -8, 2, 0, 0,
    -- filter=149 channel=125
    -13, -3, 4, -5, 13, -10, 8, 4, -5,
    -- filter=149 channel=126
    8, -11, -1, -4, 10, -2, 0, 9, -2,
    -- filter=149 channel=127
    0, -2, 0, 0, -5, 2, 5, 11, 0,
    -- filter=150 channel=0
    -4, 8, 15, -10, -6, 10, -12, -17, 3,
    -- filter=150 channel=1
    -3, 10, 4, -8, -7, 7, 0, -10, -5,
    -- filter=150 channel=2
    -5, 0, -4, 0, -8, -1, 0, -1, 0,
    -- filter=150 channel=3
    3, 4, 6, 10, 14, -3, -1, 9, 11,
    -- filter=150 channel=4
    -2, 1, 5, -2, -12, 5, 5, 5, -5,
    -- filter=150 channel=5
    6, 0, 12, 0, 1, 4, -9, -8, 8,
    -- filter=150 channel=6
    2, -2, 0, 4, 6, -2, 0, 3, 8,
    -- filter=150 channel=7
    1, 0, 0, 0, 5, 0, -4, -2, 3,
    -- filter=150 channel=8
    -2, 2, -4, -2, 2, -1, 0, 0, -5,
    -- filter=150 channel=9
    3, 0, -3, -5, 1, 7, -4, -9, -2,
    -- filter=150 channel=10
    4, -5, -2, -2, 7, -1, 8, -7, 0,
    -- filter=150 channel=11
    1, 0, -4, -5, 5, 2, 5, -3, 12,
    -- filter=150 channel=12
    0, -7, -5, 0, -2, 4, -3, -5, 3,
    -- filter=150 channel=13
    2, 0, -8, -3, -2, 7, 10, -11, -6,
    -- filter=150 channel=14
    -2, -6, 0, 0, 5, 4, 3, 2, -1,
    -- filter=150 channel=15
    8, 4, -3, 2, 11, 6, -10, -14, 9,
    -- filter=150 channel=16
    4, 0, -4, -8, 6, -1, -1, -12, -3,
    -- filter=150 channel=17
    1, 7, -7, 5, -1, -1, -5, 0, -3,
    -- filter=150 channel=18
    -1, -2, 6, 0, -3, 18, -1, -19, -7,
    -- filter=150 channel=19
    4, 0, -6, 7, 0, 3, 7, -3, 7,
    -- filter=150 channel=20
    -9, -3, -5, -1, 14, -2, 1, 10, 16,
    -- filter=150 channel=21
    6, -3, 5, 5, 0, -2, -1, 1, -7,
    -- filter=150 channel=22
    2, 3, 6, -11, 3, 5, -14, 2, 0,
    -- filter=150 channel=23
    3, -5, -11, -9, 29, 11, -14, -12, 15,
    -- filter=150 channel=24
    -5, 0, -6, 3, 3, 0, 4, -1, 0,
    -- filter=150 channel=25
    3, 8, 5, -11, -4, 15, 7, -21, -8,
    -- filter=150 channel=26
    1, 0, 7, 2, -1, 10, -1, 7, -1,
    -- filter=150 channel=27
    8, 16, 10, -13, 6, 16, -16, -23, 0,
    -- filter=150 channel=28
    -3, -2, 6, 6, 5, -5, -4, -3, 0,
    -- filter=150 channel=29
    1, -1, -4, 6, -3, 8, 10, 4, 14,
    -- filter=150 channel=30
    -3, 0, 11, -3, 4, 6, 1, -18, -9,
    -- filter=150 channel=31
    0, -4, 3, -3, 5, 9, -11, -16, -3,
    -- filter=150 channel=32
    5, 10, -2, -4, 2, 14, -9, -17, 0,
    -- filter=150 channel=33
    9, 2, 3, -8, 13, 12, -5, -18, 7,
    -- filter=150 channel=34
    -1, -6, -7, -1, 10, 4, -9, 13, 18,
    -- filter=150 channel=35
    3, 5, -6, 0, 0, 5, 3, 3, 4,
    -- filter=150 channel=36
    -4, -3, 1, 3, -4, -4, 6, -8, -13,
    -- filter=150 channel=37
    -3, 3, 7, 0, -9, 6, -1, -12, -2,
    -- filter=150 channel=38
    1, -3, 1, 0, 9, 11, 1, 1, 2,
    -- filter=150 channel=39
    -7, 0, -8, -6, 3, -6, 1, 1, 7,
    -- filter=150 channel=40
    5, 0, -13, -4, 0, -6, -1, -1, 6,
    -- filter=150 channel=41
    -8, -8, 3, 3, -9, 5, 20, 3, 0,
    -- filter=150 channel=42
    -4, 6, 6, -6, -4, 4, 4, -5, 2,
    -- filter=150 channel=43
    1, 5, 6, 3, 13, -2, 2, -2, 17,
    -- filter=150 channel=44
    5, 2, 13, -11, -7, 11, 0, -10, -9,
    -- filter=150 channel=45
    -4, -1, 7, -9, -6, 2, 3, -2, -5,
    -- filter=150 channel=46
    3, 8, -6, 8, -4, -5, 3, 0, -5,
    -- filter=150 channel=47
    -2, 9, 8, -3, 0, 7, 2, -11, 0,
    -- filter=150 channel=48
    5, 5, 12, -5, -1, 11, 11, -15, -16,
    -- filter=150 channel=49
    -5, 3, 6, -4, -8, 1, 2, -12, -5,
    -- filter=150 channel=50
    11, 10, 6, -11, 9, 4, -10, -18, -7,
    -- filter=150 channel=51
    4, 0, -7, -6, 5, 6, 2, -4, 5,
    -- filter=150 channel=52
    -3, 0, -10, 0, 3, 5, -2, -3, 10,
    -- filter=150 channel=53
    0, -2, 2, 5, 8, 0, 7, 6, -1,
    -- filter=150 channel=54
    2, 0, 2, -6, -2, 5, 2, 6, -4,
    -- filter=150 channel=55
    -2, 1, -2, -6, 4, 11, 0, -10, 5,
    -- filter=150 channel=56
    0, -8, -7, -1, 4, 2, 2, -2, -1,
    -- filter=150 channel=57
    -5, 4, 5, -3, 3, 0, 5, 2, -7,
    -- filter=150 channel=58
    2, -4, 9, -6, 6, 4, -6, 1, 7,
    -- filter=150 channel=59
    -1, 6, 4, -5, -12, 7, 1, -8, 0,
    -- filter=150 channel=60
    1, -4, 1, 6, 6, -2, 0, 0, 7,
    -- filter=150 channel=61
    -3, -7, 0, 0, 2, -7, 8, 1, 3,
    -- filter=150 channel=62
    -5, 1, 5, -5, 5, 2, 0, 6, 0,
    -- filter=150 channel=63
    3, -4, 8, 6, 0, -2, -3, 3, -2,
    -- filter=150 channel=64
    -4, 2, -3, 6, 5, -1, -2, 3, 1,
    -- filter=150 channel=65
    1, 2, -6, 3, 6, -6, -5, 4, 4,
    -- filter=150 channel=66
    1, -1, -11, -1, 0, -2, 6, -6, -1,
    -- filter=150 channel=67
    -6, 3, 2, 5, 5, -1, -4, -5, -5,
    -- filter=150 channel=68
    -6, -8, 4, -1, 2, -4, 7, 0, 0,
    -- filter=150 channel=69
    6, 0, -1, 3, 0, 7, 7, 5, 8,
    -- filter=150 channel=70
    9, 4, 0, -12, 3, 12, -8, -12, 4,
    -- filter=150 channel=71
    0, -1, 0, 1, 3, 1, -6, 6, -2,
    -- filter=150 channel=72
    2, 0, -1, 3, -5, 2, 9, -16, -5,
    -- filter=150 channel=73
    3, 3, -4, 3, -2, 6, 3, -16, 0,
    -- filter=150 channel=74
    -3, 7, -2, -7, 9, 5, -2, -2, 1,
    -- filter=150 channel=75
    10, 6, 11, -7, 1, 0, -3, -21, -2,
    -- filter=150 channel=76
    -8, -10, -17, 4, 1, -5, 7, -2, 11,
    -- filter=150 channel=77
    -7, -4, 2, 5, -3, -7, 3, -4, 6,
    -- filter=150 channel=78
    -6, -1, 3, 1, -3, 4, -4, 1, 4,
    -- filter=150 channel=79
    -1, 3, 1, -12, 5, 19, -1, -27, 4,
    -- filter=150 channel=80
    1, 0, 13, -2, -2, 13, 13, -16, -9,
    -- filter=150 channel=81
    0, 0, -2, -2, 7, -6, -1, 5, 1,
    -- filter=150 channel=82
    -2, 2, 0, -4, 1, 6, 0, 8, -2,
    -- filter=150 channel=83
    0, 3, 2, 0, 1, 6, -2, -4, -11,
    -- filter=150 channel=84
    -8, -2, -3, -1, 1, 4, -3, -15, -8,
    -- filter=150 channel=85
    -1, 1, -2, -1, 0, 3, 6, 5, 0,
    -- filter=150 channel=86
    -7, 4, 0, -7, -4, 0, 2, 0, 12,
    -- filter=150 channel=87
    -10, 0, -15, -2, 7, -7, 3, 1, 0,
    -- filter=150 channel=88
    -5, 0, -7, -4, -9, -7, -1, -5, -13,
    -- filter=150 channel=89
    0, 2, -1, 5, -2, 1, 11, -18, -3,
    -- filter=150 channel=90
    -6, -15, -9, -4, 2, -10, -1, 5, 1,
    -- filter=150 channel=91
    -2, 0, -4, -12, 2, 6, 0, -24, 0,
    -- filter=150 channel=92
    -4, -5, 0, 3, 12, 4, -1, -1, 11,
    -- filter=150 channel=93
    -2, 8, 7, -8, -11, 14, -4, -15, -15,
    -- filter=150 channel=94
    2, 6, 3, -5, 0, 6, 3, -4, 3,
    -- filter=150 channel=95
    0, 3, 1, -1, -2, -8, -7, 0, 0,
    -- filter=150 channel=96
    0, 8, 5, 1, -3, -3, 8, -1, -5,
    -- filter=150 channel=97
    -1, 8, 1, 4, 7, -3, -9, -1, 11,
    -- filter=150 channel=98
    10, 14, 16, -2, 3, 13, 3, -9, -7,
    -- filter=150 channel=99
    0, -9, -13, -10, 12, 0, -12, -10, 5,
    -- filter=150 channel=100
    -5, -2, -2, 5, 3, 0, -3, 0, 3,
    -- filter=150 channel=101
    -6, 1, -2, -4, -4, 0, -1, -7, -10,
    -- filter=150 channel=102
    -7, -5, 2, -6, -1, -2, 6, -3, 4,
    -- filter=150 channel=103
    7, 0, 10, 5, -5, 7, 0, -12, 4,
    -- filter=150 channel=104
    10, 5, 9, -9, -3, 2, 0, -13, -12,
    -- filter=150 channel=105
    -2, -8, -8, 3, 8, 0, 5, 5, 3,
    -- filter=150 channel=106
    3, -10, -10, -2, 3, -6, -4, 6, 1,
    -- filter=150 channel=107
    1, -8, -8, -9, 0, 7, -12, -2, 8,
    -- filter=150 channel=108
    -4, -4, -1, 5, 1, 1, 7, 1, 0,
    -- filter=150 channel=109
    2, 12, 6, -12, 5, 22, -2, -25, -3,
    -- filter=150 channel=110
    7, 2, -2, -4, 7, 0, 1, -7, 7,
    -- filter=150 channel=111
    -2, 1, -2, 4, -7, 2, 5, -1, 5,
    -- filter=150 channel=112
    9, 9, 7, -2, 12, 10, -13, -4, 1,
    -- filter=150 channel=113
    0, 7, 5, -7, 9, 0, -9, -5, 9,
    -- filter=150 channel=114
    -6, 4, 2, -13, 0, 24, -1, -24, 7,
    -- filter=150 channel=115
    -3, -4, 5, -5, 7, 0, -5, 1, 2,
    -- filter=150 channel=116
    1, 9, 2, -4, -5, 18, 5, -18, -13,
    -- filter=150 channel=117
    4, 3, -4, -2, -9, -7, 8, -7, 0,
    -- filter=150 channel=118
    6, 6, -7, -2, -5, 1, -3, 0, 5,
    -- filter=150 channel=119
    -5, 2, 4, 0, 6, 1, -7, 14, 3,
    -- filter=150 channel=120
    -7, 2, -4, -14, 15, 6, -8, -18, 4,
    -- filter=150 channel=121
    6, 0, -4, -1, 5, 1, -2, -3, 1,
    -- filter=150 channel=122
    -2, -3, 4, 0, -15, -6, 2, -14, -9,
    -- filter=150 channel=123
    4, -1, -3, 2, 14, 0, -5, 3, 0,
    -- filter=150 channel=124
    -1, -9, 3, 0, 1, 6, -6, 0, 11,
    -- filter=150 channel=125
    -1, 10, -2, 0, 0, 9, 6, -21, -10,
    -- filter=150 channel=126
    8, -5, 4, 3, -1, 8, 4, -5, 1,
    -- filter=150 channel=127
    -3, -7, -6, 7, 1, -3, 4, 0, -3,
    -- filter=151 channel=0
    7, 4, 16, -13, -13, 0, -11, -37, -20,
    -- filter=151 channel=1
    7, 14, 19, -9, -26, -12, -26, -37, -12,
    -- filter=151 channel=2
    2, -1, 4, -8, -2, 2, -10, -10, -8,
    -- filter=151 channel=3
    8, 2, -2, -10, -4, 5, -9, 4, -3,
    -- filter=151 channel=4
    -12, -5, 3, -18, -13, -5, -15, -12, -17,
    -- filter=151 channel=5
    4, 10, 13, -6, -12, 8, -16, -19, -5,
    -- filter=151 channel=6
    -1, -13, -10, 7, 7, -3, -1, 12, 3,
    -- filter=151 channel=7
    0, 0, -6, 6, -1, 2, -4, 0, 3,
    -- filter=151 channel=8
    1, -1, -4, 0, 0, 0, -3, -6, -6,
    -- filter=151 channel=9
    -5, 3, 3, -2, -6, 11, 3, 0, -7,
    -- filter=151 channel=10
    12, -2, 5, -3, 3, 11, 3, 3, 2,
    -- filter=151 channel=11
    -3, -19, -20, 0, 14, -7, 6, 12, 1,
    -- filter=151 channel=12
    2, -3, 8, -5, 0, 3, -6, 5, 6,
    -- filter=151 channel=13
    -5, -6, 0, -2, -1, 7, -6, 0, -4,
    -- filter=151 channel=14
    -3, 1, -1, 7, -6, -5, -1, 3, 4,
    -- filter=151 channel=15
    -5, 2, -13, 4, 14, -1, 1, 3, 12,
    -- filter=151 channel=16
    0, 8, 10, -5, -11, 6, -10, -8, -4,
    -- filter=151 channel=17
    -2, -1, 0, 4, -4, -3, 7, -6, -1,
    -- filter=151 channel=18
    5, -4, -3, 13, 5, -1, 0, -10, -6,
    -- filter=151 channel=19
    6, 2, 6, 6, -2, -2, -3, 6, -2,
    -- filter=151 channel=20
    -14, -20, -36, 4, 14, -8, 5, 36, 22,
    -- filter=151 channel=21
    3, 1, 17, -5, -10, 6, -9, -7, 3,
    -- filter=151 channel=22
    7, 8, -1, -1, 0, 8, -7, -8, -2,
    -- filter=151 channel=23
    2, -11, 2, 7, 10, 14, 3, 17, 0,
    -- filter=151 channel=24
    -6, -3, -1, 0, 0, -7, 4, -2, 7,
    -- filter=151 channel=25
    -1, 14, 20, 1, -10, 11, -10, -19, -11,
    -- filter=151 channel=26
    3, 10, 9, -10, 3, -2, 0, -4, -5,
    -- filter=151 channel=27
    9, 3, 26, -9, 7, 15, -15, -24, -10,
    -- filter=151 channel=28
    -2, -7, -4, -7, -2, 2, 7, 0, 4,
    -- filter=151 channel=29
    -10, -20, -23, 1, 9, 2, 8, 25, 13,
    -- filter=151 channel=30
    -1, 4, 14, -2, -5, 11, -7, -18, -8,
    -- filter=151 channel=31
    8, 14, 24, -13, 5, 10, -5, -2, 0,
    -- filter=151 channel=32
    6, -4, 2, -1, 3, 11, -1, -10, 1,
    -- filter=151 channel=33
    6, 14, 15, -9, 9, 15, -15, -8, -1,
    -- filter=151 channel=34
    -7, -2, 8, 1, 8, 4, 0, -3, 7,
    -- filter=151 channel=35
    -1, 4, -1, 7, 1, 2, -4, 6, -7,
    -- filter=151 channel=36
    -1, -2, -1, 0, -3, -11, 7, 9, -1,
    -- filter=151 channel=37
    3, 0, 16, -13, -21, -10, -28, -40, -14,
    -- filter=151 channel=38
    0, 1, 11, -7, 6, 15, 0, -2, 5,
    -- filter=151 channel=39
    -6, -17, -12, 6, -1, 4, 8, 9, 7,
    -- filter=151 channel=40
    -9, -1, -4, 0, 8, 7, 8, 6, -2,
    -- filter=151 channel=41
    0, 5, -2, 6, 4, -3, -1, 4, -6,
    -- filter=151 channel=42
    7, -3, 1, -8, -1, -1, 3, -2, -3,
    -- filter=151 channel=43
    5, 1, -2, 2, 1, 2, 5, 0, 4,
    -- filter=151 channel=44
    2, 9, 24, -14, -17, 4, -6, -26, -13,
    -- filter=151 channel=45
    -7, -2, 2, 4, -3, -2, 2, 5, 3,
    -- filter=151 channel=46
    7, -3, 0, -5, -3, 1, -9, 0, 0,
    -- filter=151 channel=47
    2, 6, 26, -13, -19, 7, -12, -25, -7,
    -- filter=151 channel=48
    1, 11, 18, -6, -4, 0, -15, -22, -7,
    -- filter=151 channel=49
    -10, -8, 2, -5, 3, 1, -3, -1, -5,
    -- filter=151 channel=50
    4, 10, 14, 3, 5, 5, -1, -6, -3,
    -- filter=151 channel=51
    -7, 1, 5, 5, -3, 5, -2, 0, 2,
    -- filter=151 channel=52
    -1, -13, 3, -6, -3, 2, 5, 4, 7,
    -- filter=151 channel=53
    -3, -11, -14, 7, 0, 6, -3, 14, 0,
    -- filter=151 channel=54
    6, 0, 4, -1, 0, -6, -6, -3, -4,
    -- filter=151 channel=55
    -1, -17, -25, 11, 12, -2, 2, 22, 11,
    -- filter=151 channel=56
    -2, -5, 0, 2, -6, 4, 4, -3, 2,
    -- filter=151 channel=57
    0, -4, 6, -6, -1, -6, 0, 3, -3,
    -- filter=151 channel=58
    0, -1, 1, -10, 0, 4, -8, -13, -8,
    -- filter=151 channel=59
    12, 14, 19, -9, 0, 5, -7, -9, -14,
    -- filter=151 channel=60
    4, -7, 4, 2, 0, 6, -3, 4, 0,
    -- filter=151 channel=61
    2, 1, -1, -9, 5, 0, 5, -2, 4,
    -- filter=151 channel=62
    -1, 4, 1, 7, 5, 0, -5, -1, 3,
    -- filter=151 channel=63
    4, 8, 12, 3, -9, -2, 5, -2, -7,
    -- filter=151 channel=64
    -3, 0, -14, 0, 0, 4, 6, 9, 6,
    -- filter=151 channel=65
    0, 7, -2, 5, -2, 6, 0, 0, 5,
    -- filter=151 channel=66
    0, -7, 0, -6, -7, 5, -5, 0, -5,
    -- filter=151 channel=67
    2, -2, 0, 4, 4, 7, -5, 4, 5,
    -- filter=151 channel=68
    0, 0, -3, -4, 1, 1, -7, -2, -7,
    -- filter=151 channel=69
    -4, -2, 4, -3, -3, -6, 0, -4, 6,
    -- filter=151 channel=70
    11, 4, 6, -2, 1, 7, -2, -14, -3,
    -- filter=151 channel=71
    -2, -2, 0, 4, 9, 9, -9, 3, -2,
    -- filter=151 channel=72
    2, 0, 7, -7, -5, 4, 8, 4, -6,
    -- filter=151 channel=73
    -5, -6, -7, -2, -1, 2, 0, -8, 0,
    -- filter=151 channel=74
    4, 5, 14, 0, 1, 9, -9, -13, -4,
    -- filter=151 channel=75
    13, 9, 17, -8, -11, -3, -23, -33, -15,
    -- filter=151 channel=76
    -19, -21, -37, 13, 10, -1, 15, 18, 19,
    -- filter=151 channel=77
    4, -5, 0, 2, 4, 3, -2, 7, 7,
    -- filter=151 channel=78
    -3, -2, 13, 4, 4, 9, 1, 4, 4,
    -- filter=151 channel=79
    10, 0, 2, 7, -2, 9, -8, -4, -4,
    -- filter=151 channel=80
    14, 17, 20, 1, -3, 4, 3, -8, -13,
    -- filter=151 channel=81
    0, 0, -2, -5, -3, -2, -6, 1, -4,
    -- filter=151 channel=82
    4, -2, -4, 1, 7, 7, 4, 3, 0,
    -- filter=151 channel=83
    9, 10, 15, -3, -8, -5, 1, -9, -9,
    -- filter=151 channel=84
    0, -7, -10, -5, -3, -6, -5, -6, -1,
    -- filter=151 channel=85
    -2, -1, -3, 0, 2, -5, 4, 0, 3,
    -- filter=151 channel=86
    1, 0, 11, -12, -10, 0, -3, -7, -7,
    -- filter=151 channel=87
    -4, -18, -19, 1, 3, 0, 2, 13, 12,
    -- filter=151 channel=88
    -2, -4, -6, -2, -1, -8, 9, 3, 7,
    -- filter=151 channel=89
    8, -9, 0, 6, -3, 6, 5, 5, -3,
    -- filter=151 channel=90
    2, -3, 0, -6, 0, 7, 2, -2, 7,
    -- filter=151 channel=91
    -4, -6, -1, -8, -1, 2, -3, -3, -15,
    -- filter=151 channel=92
    -3, -2, -3, 0, 3, 6, 4, -5, 1,
    -- filter=151 channel=93
    0, 11, 33, -5, -10, -7, -12, -25, -18,
    -- filter=151 channel=94
    2, 1, -6, 0, 3, -1, -2, 3, 3,
    -- filter=151 channel=95
    -2, -4, -3, 0, -3, 4, -3, 0, -3,
    -- filter=151 channel=96
    3, 2, 7, 1, 5, 2, -3, -4, -1,
    -- filter=151 channel=97
    3, -1, 1, -4, 6, 9, -4, -10, -8,
    -- filter=151 channel=98
    6, 17, 16, -9, -1, 7, -1, -11, -2,
    -- filter=151 channel=99
    -6, -8, 6, 0, 12, 7, 6, 2, 0,
    -- filter=151 channel=100
    2, 0, -3, 9, 1, 1, -3, -2, 1,
    -- filter=151 channel=101
    0, -3, 3, -13, -11, -4, -13, -5, -4,
    -- filter=151 channel=102
    -4, 0, 0, 0, 1, 2, -5, 0, 0,
    -- filter=151 channel=103
    10, 0, 24, -7, -19, 11, -11, -25, -15,
    -- filter=151 channel=104
    10, 7, 11, -8, -8, 1, 5, -6, -2,
    -- filter=151 channel=105
    -7, -15, -21, 0, 10, -4, 14, 13, 4,
    -- filter=151 channel=106
    -5, -2, -15, 6, 2, 0, 3, 6, 3,
    -- filter=151 channel=107
    -9, -16, -5, 8, 3, 4, 0, 2, 3,
    -- filter=151 channel=108
    -8, -5, 1, 2, -2, -8, 0, 4, 2,
    -- filter=151 channel=109
    7, 6, 16, -6, 0, 6, -16, -6, -10,
    -- filter=151 channel=110
    6, -6, -3, 5, 3, 0, 4, 6, -1,
    -- filter=151 channel=111
    0, 1, 2, 6, -7, 3, 0, 5, 3,
    -- filter=151 channel=112
    7, 14, 9, -5, -5, 2, -13, -18, -2,
    -- filter=151 channel=113
    4, 2, 9, 2, -3, 14, 2, -10, 2,
    -- filter=151 channel=114
    2, -5, 7, 5, -1, 0, -8, -25, -3,
    -- filter=151 channel=115
    0, 3, 1, 3, -1, 4, -7, -4, -1,
    -- filter=151 channel=116
    0, 0, 2, -3, 3, 2, 2, -3, -13,
    -- filter=151 channel=117
    4, -2, -1, -4, 0, 4, -4, -1, 1,
    -- filter=151 channel=118
    -2, -5, 0, 4, 0, 1, 0, 0, -2,
    -- filter=151 channel=119
    -2, -3, 10, 3, 5, 1, -1, 0, -4,
    -- filter=151 channel=120
    -4, 1, 1, 4, 11, 0, -4, 2, 0,
    -- filter=151 channel=121
    4, -2, -2, 0, -5, -6, -6, -5, 0,
    -- filter=151 channel=122
    -4, 11, 33, -20, -21, 5, -21, -30, -18,
    -- filter=151 channel=123
    -3, -1, 3, 0, 0, -1, -4, -8, 0,
    -- filter=151 channel=124
    -11, -6, -8, 10, 1, 4, 2, 13, 2,
    -- filter=151 channel=125
    6, 7, 7, -7, -2, 11, 1, -10, -2,
    -- filter=151 channel=126
    6, -2, 1, -4, 2, 7, 8, 3, -7,
    -- filter=151 channel=127
    -2, 4, -2, 0, 3, -3, -1, -4, -7,
    -- filter=152 channel=0
    15, 10, -14, 10, 2, -12, 10, -4, -12,
    -- filter=152 channel=1
    10, 6, -10, -1, -2, -6, 0, 4, -7,
    -- filter=152 channel=2
    1, 1, -6, -7, -3, 5, 3, -2, 8,
    -- filter=152 channel=3
    14, 4, 5, -1, 2, 5, -7, -3, -8,
    -- filter=152 channel=4
    0, 3, -5, -3, -2, 7, 1, 6, 6,
    -- filter=152 channel=5
    19, 6, -11, 9, 9, -18, 14, -1, -17,
    -- filter=152 channel=6
    -4, 4, -7, 3, 6, 7, -1, -4, 7,
    -- filter=152 channel=7
    5, -6, -7, -3, -3, -4, -7, 1, 7,
    -- filter=152 channel=8
    -8, 2, 4, 4, -4, 10, 0, 4, -1,
    -- filter=152 channel=9
    0, 7, 1, 0, 0, -11, 3, 3, 3,
    -- filter=152 channel=10
    10, 11, 5, 1, 0, -6, 2, 6, -2,
    -- filter=152 channel=11
    1, -1, 0, 1, 4, 5, -3, 7, 1,
    -- filter=152 channel=12
    4, 9, 4, -3, 7, 1, 3, 9, 0,
    -- filter=152 channel=13
    1, 7, 10, 1, 15, 0, 0, 1, -4,
    -- filter=152 channel=14
    4, -1, 7, 1, -6, 2, 5, 3, -2,
    -- filter=152 channel=15
    -5, 0, 2, 0, 10, -5, 3, -4, 0,
    -- filter=152 channel=16
    -3, 10, -5, 1, 7, -12, -6, -6, -1,
    -- filter=152 channel=17
    7, 4, 2, -6, 5, 2, 3, 5, -3,
    -- filter=152 channel=18
    4, 6, -12, 0, 12, -1, -2, -6, 1,
    -- filter=152 channel=19
    1, 0, -5, -2, -3, 4, 0, -2, 6,
    -- filter=152 channel=20
    -3, 0, -7, 6, 24, 0, 6, 12, 1,
    -- filter=152 channel=21
    -4, 11, 0, 4, 5, -11, 8, 5, -5,
    -- filter=152 channel=22
    3, 4, 4, 7, -4, 1, -2, 1, 3,
    -- filter=152 channel=23
    3, -6, -12, -3, 5, -12, -8, -9, 4,
    -- filter=152 channel=24
    -2, 1, 1, 4, 0, -1, 3, 0, -6,
    -- filter=152 channel=25
    0, 9, -14, -3, 9, -11, 2, 5, -6,
    -- filter=152 channel=26
    8, 6, 0, 12, 9, 0, 11, -6, -4,
    -- filter=152 channel=27
    3, 8, -26, -10, 0, -30, -11, -4, -5,
    -- filter=152 channel=28
    -3, -3, 6, 1, -6, -1, 6, 7, 6,
    -- filter=152 channel=29
    2, -4, -13, 14, 19, 2, 5, 9, 2,
    -- filter=152 channel=30
    14, 10, 0, 1, 2, -10, -1, -5, -8,
    -- filter=152 channel=31
    8, 0, -17, -10, -5, -19, -5, -2, -5,
    -- filter=152 channel=32
    2, 5, -14, 0, 14, -6, -8, 2, -7,
    -- filter=152 channel=33
    12, 8, -8, 2, -3, -10, 1, -2, -6,
    -- filter=152 channel=34
    2, 9, 13, -5, -1, 15, 1, 3, 2,
    -- filter=152 channel=35
    5, 3, -2, 5, -4, 2, 4, 2, 0,
    -- filter=152 channel=36
    -1, 9, 9, 8, 14, 10, -1, 0, 7,
    -- filter=152 channel=37
    13, 16, -13, 6, 10, -10, -2, -4, -11,
    -- filter=152 channel=38
    1, 3, 3, 5, 3, -10, -2, -1, 2,
    -- filter=152 channel=39
    -3, -3, 4, 9, 11, -2, 0, 4, 0,
    -- filter=152 channel=40
    2, -5, 0, 6, 6, 8, -5, 2, 7,
    -- filter=152 channel=41
    -2, 8, 22, -8, 11, 19, -2, -4, 9,
    -- filter=152 channel=42
    7, 5, -8, 1, -8, -1, -4, -7, -3,
    -- filter=152 channel=43
    6, -2, 6, 5, 1, 5, 4, -7, 3,
    -- filter=152 channel=44
    11, 10, -14, -4, -1, -18, 7, -5, -3,
    -- filter=152 channel=45
    7, 1, -7, 3, 2, 1, 0, -6, -6,
    -- filter=152 channel=46
    -6, -6, 4, 5, 3, 11, 1, -3, 0,
    -- filter=152 channel=47
    3, 9, -7, -3, -3, -18, 8, -4, -15,
    -- filter=152 channel=48
    -2, 4, -11, -6, 3, -18, -3, -10, 0,
    -- filter=152 channel=49
    -9, -2, -11, 2, -2, 0, -5, -3, -3,
    -- filter=152 channel=50
    2, -2, -10, -2, 1, -12, 1, -3, -2,
    -- filter=152 channel=51
    -5, -5, 0, 4, -3, 0, -4, -5, 4,
    -- filter=152 channel=52
    -3, -3, 0, 0, 1, 6, 2, -2, 0,
    -- filter=152 channel=53
    -5, -6, 3, -2, 0, -5, 1, 4, 0,
    -- filter=152 channel=54
    -3, 0, -2, 5, 2, 3, 0, 2, 0,
    -- filter=152 channel=55
    3, -2, -4, -1, 20, -2, -1, 3, -7,
    -- filter=152 channel=56
    0, 0, 0, 0, 4, 1, 1, 7, 7,
    -- filter=152 channel=57
    -6, -4, 6, 0, -2, 1, -4, -1, 8,
    -- filter=152 channel=58
    12, 9, 0, 8, 0, 0, 2, 5, 0,
    -- filter=152 channel=59
    1, 9, -9, -3, 1, -18, -3, -3, -10,
    -- filter=152 channel=60
    -1, -3, -6, 6, -6, 6, -3, 2, 4,
    -- filter=152 channel=61
    6, 9, 9, 7, 1, 9, -3, 7, 0,
    -- filter=152 channel=62
    3, -6, -5, 7, 6, -2, -2, -7, 0,
    -- filter=152 channel=63
    5, 2, 9, 1, 9, 0, 6, 9, -9,
    -- filter=152 channel=64
    3, 5, 10, 2, 4, 9, 2, -1, 9,
    -- filter=152 channel=65
    0, -2, 0, 3, 3, -5, 1, 2, -5,
    -- filter=152 channel=66
    -1, 13, 6, 0, 15, 5, -6, 7, 5,
    -- filter=152 channel=67
    5, 4, 7, 4, 0, 0, -2, 4, -2,
    -- filter=152 channel=68
    -2, 1, 5, -1, 5, -1, -6, -6, -1,
    -- filter=152 channel=69
    0, 1, 5, 7, 11, -1, 0, 8, -7,
    -- filter=152 channel=70
    5, 5, -7, -3, -3, -5, -5, -2, 5,
    -- filter=152 channel=71
    5, -4, 0, 0, -7, -7, 2, -5, 1,
    -- filter=152 channel=72
    0, 11, -15, -6, 6, -18, -5, -1, -11,
    -- filter=152 channel=73
    -6, -1, -5, 1, 1, -3, -8, 4, 7,
    -- filter=152 channel=74
    4, -2, -7, -1, 3, -5, 2, -4, 9,
    -- filter=152 channel=75
    18, 10, 5, 9, 7, -19, 10, -8, -14,
    -- filter=152 channel=76
    -6, -1, 10, 3, 21, 14, 2, 3, 1,
    -- filter=152 channel=77
    6, 6, 5, -6, 2, -4, -1, 6, 3,
    -- filter=152 channel=78
    -1, 3, 7, 7, 1, 0, 9, 0, 3,
    -- filter=152 channel=79
    11, 3, -3, 0, 13, -16, -9, -2, -13,
    -- filter=152 channel=80
    10, 5, -8, -10, 1, -25, 3, -3, -17,
    -- filter=152 channel=81
    1, -6, -4, -5, 0, 4, -6, 7, 1,
    -- filter=152 channel=82
    0, 0, -6, 3, -6, 4, -4, -5, -1,
    -- filter=152 channel=83
    2, -3, -8, 1, -2, -6, 5, 4, -8,
    -- filter=152 channel=84
    3, 4, -7, 0, 9, -1, -4, -3, 8,
    -- filter=152 channel=85
    -5, 6, 0, -5, -2, -6, -4, -2, -5,
    -- filter=152 channel=86
    0, 11, 5, 2, 16, 7, 2, 0, 0,
    -- filter=152 channel=87
    3, 0, 2, 7, 4, 15, 0, -1, 7,
    -- filter=152 channel=88
    -6, 7, 3, 5, 9, 10, 0, 0, 8,
    -- filter=152 channel=89
    -1, 0, -8, -14, 10, -13, -11, 4, -7,
    -- filter=152 channel=90
    -2, 10, 0, 3, 10, 4, 1, 11, 4,
    -- filter=152 channel=91
    -1, 0, -11, -11, -2, -14, -12, -2, -4,
    -- filter=152 channel=92
    -4, -5, -4, 0, -6, 4, -6, -2, 7,
    -- filter=152 channel=93
    6, 11, -7, -2, 8, -20, 7, -1, -4,
    -- filter=152 channel=94
    0, 5, -4, -5, 6, -2, -2, 3, 7,
    -- filter=152 channel=95
    2, 2, -2, -1, -1, 4, 0, -5, 0,
    -- filter=152 channel=96
    6, 0, 4, -3, -7, -1, -6, 3, -8,
    -- filter=152 channel=97
    8, -3, 1, 7, 6, 4, -1, 3, 1,
    -- filter=152 channel=98
    -1, 11, -11, -5, 3, -16, -3, 0, -12,
    -- filter=152 channel=99
    -4, 3, -10, -10, 2, -15, -6, 8, 7,
    -- filter=152 channel=100
    -2, 0, 10, 3, 5, 9, 5, 6, -1,
    -- filter=152 channel=101
    -4, 9, -5, 0, -7, 0, 1, 8, 12,
    -- filter=152 channel=102
    -4, -4, 6, -4, -7, 5, 0, -4, 4,
    -- filter=152 channel=103
    8, 12, -14, -1, 4, -26, -1, 1, -11,
    -- filter=152 channel=104
    0, 7, -11, -4, -7, -15, 2, 3, 1,
    -- filter=152 channel=105
    -1, -2, 1, 6, 10, 4, 0, -3, 2,
    -- filter=152 channel=106
    -6, -3, 2, 3, 10, 2, -3, -5, 3,
    -- filter=152 channel=107
    1, 0, -10, 11, 8, 0, 5, -5, -1,
    -- filter=152 channel=108
    -1, -2, 7, 4, -2, 3, 6, 0, 1,
    -- filter=152 channel=109
    4, -4, -20, -7, 1, -11, 2, 0, 2,
    -- filter=152 channel=110
    5, 8, -1, 4, 7, -7, 2, 2, -5,
    -- filter=152 channel=111
    5, 2, 7, 0, 6, 0, -4, 3, -3,
    -- filter=152 channel=112
    -6, 3, -12, -4, -1, -13, -7, 5, -7,
    -- filter=152 channel=113
    9, 5, 3, -8, 0, -4, -10, 3, -8,
    -- filter=152 channel=114
    3, 1, -21, 4, 7, -13, 5, -10, -8,
    -- filter=152 channel=115
    -5, 0, 5, -2, 2, 3, -1, 1, -1,
    -- filter=152 channel=116
    -1, 8, -5, -8, -2, -6, -8, -6, 0,
    -- filter=152 channel=117
    -2, 0, -2, -3, 6, -1, 2, 3, 2,
    -- filter=152 channel=118
    2, 6, 3, -5, 4, -1, -7, -2, -6,
    -- filter=152 channel=119
    3, -2, 1, 7, -2, 7, -2, 10, 4,
    -- filter=152 channel=120
    -1, -4, -12, -7, 8, -9, -15, -1, -5,
    -- filter=152 channel=121
    2, 11, 11, 2, 9, 2, -5, 5, 6,
    -- filter=152 channel=122
    -2, 16, -7, 4, -6, -12, -3, -2, -8,
    -- filter=152 channel=123
    7, 4, 3, 0, -2, 3, -1, 1, 1,
    -- filter=152 channel=124
    -4, -5, -3, 10, 5, 7, 2, -4, 3,
    -- filter=152 channel=125
    -4, 2, -9, -7, -3, -18, -8, 0, -7,
    -- filter=152 channel=126
    6, 8, 3, -3, 5, 1, 1, 4, 0,
    -- filter=152 channel=127
    2, 5, 6, 2, 3, 8, 1, 2, -1,
    -- filter=153 channel=0
    2, -3, -8, 3, -4, -19, 1, -12, -13,
    -- filter=153 channel=1
    -4, -2, -14, -4, -11, -17, 0, 0, -3,
    -- filter=153 channel=2
    -3, 4, 5, -5, -3, 0, 10, -1, -3,
    -- filter=153 channel=3
    8, 4, 3, -7, -1, 0, -3, -12, -1,
    -- filter=153 channel=4
    -1, -4, -2, -4, -8, 0, 7, 14, -2,
    -- filter=153 channel=5
    3, 5, -3, 1, 2, -11, 4, 4, -6,
    -- filter=153 channel=6
    -7, 2, 0, -5, 6, 5, -4, 1, -5,
    -- filter=153 channel=7
    -4, -5, 4, -2, 3, 6, 0, -2, -4,
    -- filter=153 channel=8
    -2, -5, 1, 7, -9, -4, 5, -5, 4,
    -- filter=153 channel=9
    -7, 3, 3, -7, 4, -1, 0, 5, -1,
    -- filter=153 channel=10
    -1, 4, 1, -2, 0, 4, 0, 4, -2,
    -- filter=153 channel=11
    6, 3, 6, -4, 13, 13, 4, 1, 4,
    -- filter=153 channel=12
    5, -7, -4, 3, 4, -2, 7, 1, 1,
    -- filter=153 channel=13
    0, 2, -3, 1, -7, -10, 4, -10, -9,
    -- filter=153 channel=14
    -1, -6, 1, -6, -4, 0, 3, -5, 7,
    -- filter=153 channel=15
    1, -4, -1, -5, -6, 4, -3, -10, 3,
    -- filter=153 channel=16
    4, 8, 4, 3, 0, -1, 0, 3, 2,
    -- filter=153 channel=17
    -4, 2, 1, 4, 0, -2, 1, 5, -2,
    -- filter=153 channel=18
    -1, -9, 1, -9, -3, -7, -1, -12, -9,
    -- filter=153 channel=19
    4, -4, 2, -6, 4, 3, 1, 2, 5,
    -- filter=153 channel=20
    0, 8, 22, 10, 13, 25, 7, 8, 9,
    -- filter=153 channel=21
    2, 7, 1, 10, 13, 6, 3, 10, 8,
    -- filter=153 channel=22
    5, -8, -11, -8, -9, -10, -8, 0, -7,
    -- filter=153 channel=23
    3, 0, 8, -1, -13, 5, 4, -6, 2,
    -- filter=153 channel=24
    3, 5, 4, -1, -6, 3, 1, 3, -6,
    -- filter=153 channel=25
    5, -12, -3, 0, -7, -10, -3, 0, -8,
    -- filter=153 channel=26
    -3, 5, -4, 8, 4, 8, 0, 9, 9,
    -- filter=153 channel=27
    -2, -4, -16, -2, -12, -8, -4, -13, -17,
    -- filter=153 channel=28
    -1, 5, 2, 0, 5, 2, 1, 3, 2,
    -- filter=153 channel=29
    5, 11, 16, 0, 4, 16, 0, 8, 7,
    -- filter=153 channel=30
    -9, 4, 0, -1, -8, -7, -5, 0, -11,
    -- filter=153 channel=31
    6, 12, 8, 9, 6, 7, 1, 6, -3,
    -- filter=153 channel=32
    -3, -12, -2, -9, -10, -3, -2, -4, -6,
    -- filter=153 channel=33
    7, -4, -8, 0, -6, -16, -2, -8, -16,
    -- filter=153 channel=34
    -2, -5, 0, -1, 3, -4, -7, -2, -6,
    -- filter=153 channel=35
    0, 0, -6, 2, -1, 7, 6, 3, -1,
    -- filter=153 channel=36
    5, 4, 6, 4, 10, 2, 14, 16, 16,
    -- filter=153 channel=37
    0, -8, -7, 0, -5, -14, -2, -9, -5,
    -- filter=153 channel=38
    -3, 0, -3, -1, -3, -4, -3, 0, -4,
    -- filter=153 channel=39
    5, -2, 12, 6, 12, 2, 2, 7, 8,
    -- filter=153 channel=40
    3, -2, 7, 7, 2, 12, -5, 3, 7,
    -- filter=153 channel=41
    3, -2, 8, 9, 7, -14, 23, 5, -5,
    -- filter=153 channel=42
    -4, -7, -1, -2, -3, -2, -1, 1, 0,
    -- filter=153 channel=43
    0, 6, 0, 2, -7, 1, 0, 0, -3,
    -- filter=153 channel=44
    -8, -4, -12, 0, -6, -15, -3, 2, -7,
    -- filter=153 channel=45
    4, 7, -4, 5, -6, 7, 2, 2, -4,
    -- filter=153 channel=46
    7, 1, -1, 0, 2, -8, -4, 6, 5,
    -- filter=153 channel=47
    -5, -1, -5, -8, 1, -2, -9, 0, -7,
    -- filter=153 channel=48
    1, -9, -4, -5, -4, -7, 2, 0, 1,
    -- filter=153 channel=49
    -1, -6, -1, 0, -5, -9, -4, 0, 5,
    -- filter=153 channel=50
    -4, -11, -11, 5, -12, -7, 0, -2, -9,
    -- filter=153 channel=51
    0, -6, 6, 0, 0, 7, 4, -5, -1,
    -- filter=153 channel=52
    6, 4, -3, -3, -5, 5, 6, 2, 7,
    -- filter=153 channel=53
    3, 1, 0, -1, 4, 5, -5, -4, 4,
    -- filter=153 channel=54
    -4, -5, -5, -7, 1, 2, 5, 7, -2,
    -- filter=153 channel=55
    6, -1, 10, -1, 4, 11, 2, 1, -3,
    -- filter=153 channel=56
    0, 1, 0, 7, -3, -9, 3, -2, -6,
    -- filter=153 channel=57
    2, 0, 6, -2, -3, -8, 6, 4, 6,
    -- filter=153 channel=58
    1, -3, 4, -1, -1, -9, -1, 6, 4,
    -- filter=153 channel=59
    5, -2, -6, -2, 2, -4, 5, -6, 2,
    -- filter=153 channel=60
    1, -3, -1, -2, -5, 3, 5, -3, 0,
    -- filter=153 channel=61
    6, 0, 2, 2, -1, 2, 7, 4, 9,
    -- filter=153 channel=62
    0, -3, 7, 4, -2, 5, -5, -6, 0,
    -- filter=153 channel=63
    8, -3, 0, 2, -2, 3, 8, 7, 6,
    -- filter=153 channel=64
    7, 2, 10, 1, -1, 9, 5, 7, 4,
    -- filter=153 channel=65
    0, 5, 0, -4, -3, 5, -5, -3, -4,
    -- filter=153 channel=66
    5, -7, -3, 8, 5, -1, 12, 7, 3,
    -- filter=153 channel=67
    0, 9, 0, 8, 9, 4, -3, 1, 4,
    -- filter=153 channel=68
    6, 0, -2, 0, 0, 1, 3, 6, 8,
    -- filter=153 channel=69
    6, 3, 5, 7, 4, -5, 0, -5, 0,
    -- filter=153 channel=70
    4, -15, -12, 0, -19, -4, -9, -6, -11,
    -- filter=153 channel=71
    5, 7, -1, 1, 7, -3, -4, 2, -7,
    -- filter=153 channel=72
    3, 7, 1, 10, 5, 0, 9, -1, 7,
    -- filter=153 channel=73
    2, -4, -2, 0, 0, 3, 3, 0, -1,
    -- filter=153 channel=74
    2, -9, -1, 6, -13, 2, 7, -9, -8,
    -- filter=153 channel=75
    2, 0, 1, 1, -10, -14, -8, -3, -5,
    -- filter=153 channel=76
    8, 3, 17, 7, 16, 20, 5, 0, 10,
    -- filter=153 channel=77
    5, -6, -3, 0, 3, 4, 4, -1, 6,
    -- filter=153 channel=78
    2, 6, -3, -7, 1, -5, 1, 4, 0,
    -- filter=153 channel=79
    -3, -16, 0, -5, -19, -19, 2, -5, -8,
    -- filter=153 channel=80
    8, -2, -3, -5, -1, -3, 5, 7, 1,
    -- filter=153 channel=81
    -3, 2, 3, -3, 2, -1, 4, 6, -5,
    -- filter=153 channel=82
    -1, 3, 2, -2, 5, 5, 5, -5, -6,
    -- filter=153 channel=83
    -2, 4, -2, -3, -3, -3, 4, 11, -4,
    -- filter=153 channel=84
    0, -7, -8, -6, -12, 4, 5, 6, 7,
    -- filter=153 channel=85
    7, 6, 0, -6, 2, 0, 0, 4, -3,
    -- filter=153 channel=86
    -3, -9, -3, 5, -10, -9, 6, -1, -3,
    -- filter=153 channel=87
    -1, 6, 3, 9, 9, 12, 0, 0, 1,
    -- filter=153 channel=88
    -1, 1, 14, 2, 3, 13, 6, 9, 13,
    -- filter=153 channel=89
    7, -7, -3, -5, -5, 0, -1, 0, -2,
    -- filter=153 channel=90
    12, 12, 5, -2, 11, 13, 8, 4, 9,
    -- filter=153 channel=91
    -8, -9, -8, 4, -18, -12, 2, 5, 0,
    -- filter=153 channel=92
    6, -5, 1, 7, 0, 4, -6, -6, -8,
    -- filter=153 channel=93
    -7, 1, -4, -5, -12, -7, 6, 6, -7,
    -- filter=153 channel=94
    6, 6, 5, -3, -7, -6, 2, -5, 5,
    -- filter=153 channel=95
    0, 6, -2, -5, -7, 4, 6, 4, -1,
    -- filter=153 channel=96
    0, 5, -5, -7, 4, -5, -5, 0, -5,
    -- filter=153 channel=97
    0, -3, 6, 3, -1, 0, 0, -3, -7,
    -- filter=153 channel=98
    0, 4, -7, -4, -14, -8, 5, -10, -7,
    -- filter=153 channel=99
    10, 0, 0, 8, 7, 14, 0, 0, 8,
    -- filter=153 channel=100
    0, 4, 0, -1, 8, -4, 1, 7, -2,
    -- filter=153 channel=101
    -2, -6, 1, 2, 5, -4, -1, 10, 7,
    -- filter=153 channel=102
    3, -7, -4, -5, 0, -5, -1, -4, 7,
    -- filter=153 channel=103
    0, 4, -2, 2, -9, -12, -6, -1, -6,
    -- filter=153 channel=104
    1, 4, 6, -1, 9, 4, 8, 7, -2,
    -- filter=153 channel=105
    4, 12, 4, 4, 11, 15, -3, 8, 13,
    -- filter=153 channel=106
    -1, 2, 3, 10, 10, 0, -2, 7, 10,
    -- filter=153 channel=107
    -2, 4, 3, -4, -5, 6, -5, -6, 0,
    -- filter=153 channel=108
    -3, 1, 7, 5, 8, 4, -1, 0, 0,
    -- filter=153 channel=109
    1, -13, -9, -3, -19, -13, 5, 2, -10,
    -- filter=153 channel=110
    1, 1, -1, 6, 9, 1, -5, 0, 9,
    -- filter=153 channel=111
    7, 7, 0, 3, 0, 4, 7, 8, 4,
    -- filter=153 channel=112
    -7, -7, -8, 1, -12, -9, -1, -5, -9,
    -- filter=153 channel=113
    -3, -4, -3, 4, -8, -7, 2, -8, -4,
    -- filter=153 channel=114
    -4, -16, -16, -9, -24, -18, 1, -9, -14,
    -- filter=153 channel=115
    -1, 3, 1, -2, -2, 0, -2, 3, 4,
    -- filter=153 channel=116
    4, 0, -9, -2, -6, -6, 11, 9, 5,
    -- filter=153 channel=117
    -5, 5, 5, -6, -6, -6, 6, 0, 0,
    -- filter=153 channel=118
    6, 2, -2, 6, 6, 0, -5, 4, 7,
    -- filter=153 channel=119
    0, 0, -4, 0, 0, 1, -4, 4, -4,
    -- filter=153 channel=120
    0, -2, -9, -5, -15, 4, 1, -8, -2,
    -- filter=153 channel=121
    -1, -4, 4, 0, 7, 4, 1, 0, -9,
    -- filter=153 channel=122
    2, 4, -2, -1, 0, -3, -2, 0, 0,
    -- filter=153 channel=123
    -2, 4, -7, 6, 0, -1, 6, 5, -6,
    -- filter=153 channel=124
    -4, 3, 10, 7, -1, 1, -5, 3, -1,
    -- filter=153 channel=125
    8, -6, -4, 0, 3, -1, 9, 3, 7,
    -- filter=153 channel=126
    9, 0, -4, 1, 6, -2, 4, -1, -9,
    -- filter=153 channel=127
    -1, 7, 2, 0, 0, -7, 6, -4, 4,
    -- filter=154 channel=0
    2, -22, -37, 17, -21, -40, 25, 0, -19,
    -- filter=154 channel=1
    7, -19, -35, 3, -16, -45, 13, -2, -26,
    -- filter=154 channel=2
    3, 3, 6, 0, -3, 4, 7, -3, -4,
    -- filter=154 channel=3
    0, -8, -1, -4, -2, -14, -4, 0, -3,
    -- filter=154 channel=4
    5, 1, -6, -7, -14, -14, 6, 6, 0,
    -- filter=154 channel=5
    2, -7, -20, 8, -18, -13, 2, 5, -15,
    -- filter=154 channel=6
    -2, 5, -1, -4, -7, -6, 6, 1, -4,
    -- filter=154 channel=7
    0, 6, -3, -1, -3, 4, 1, -4, 6,
    -- filter=154 channel=8
    0, -13, 0, -5, -9, 2, -1, -7, -8,
    -- filter=154 channel=9
    2, 2, 1, 2, 3, 2, 5, 6, 2,
    -- filter=154 channel=10
    0, 7, 5, -4, 3, 4, -5, 0, 1,
    -- filter=154 channel=11
    0, 5, 13, -6, 8, 22, -8, 0, 13,
    -- filter=154 channel=12
    2, -10, 2, -5, 1, -7, -10, 0, -6,
    -- filter=154 channel=13
    -2, -6, -5, -6, -1, 0, -13, -1, -7,
    -- filter=154 channel=14
    7, -5, -3, 1, -6, -6, -4, 0, 4,
    -- filter=154 channel=15
    -2, -4, -7, 3, -4, 1, 8, -2, 5,
    -- filter=154 channel=16
    -2, -8, -14, -2, -6, -1, -7, -2, -11,
    -- filter=154 channel=17
    -5, -6, 5, -5, 0, 6, 6, 3, -3,
    -- filter=154 channel=18
    1, -5, -9, 2, -10, -19, 6, -1, -6,
    -- filter=154 channel=19
    -4, 2, 5, 6, 3, -1, -5, 0, 0,
    -- filter=154 channel=20
    2, 9, 20, 6, -1, 19, -13, 0, 14,
    -- filter=154 channel=21
    -3, 9, -2, 4, 7, -1, 4, 13, 1,
    -- filter=154 channel=22
    5, -7, -3, -2, -4, -14, 1, -6, -3,
    -- filter=154 channel=23
    -3, -15, 7, 5, -9, 6, 0, -6, 0,
    -- filter=154 channel=24
    -2, 6, 0, -7, -5, 0, 0, 2, -6,
    -- filter=154 channel=25
    9, -3, -12, 7, -3, -13, 4, 5, -3,
    -- filter=154 channel=26
    3, -2, -5, -3, 0, 2, 4, -2, -3,
    -- filter=154 channel=27
    16, -7, -8, 17, -2, -8, 17, 0, -16,
    -- filter=154 channel=28
    5, -6, 3, -1, 6, 4, -1, 3, -6,
    -- filter=154 channel=29
    1, 7, 17, -1, 10, 18, 3, -6, 11,
    -- filter=154 channel=30
    12, -11, -9, 8, -10, -4, 14, 1, -14,
    -- filter=154 channel=31
    0, 11, 0, 15, 14, 16, 2, 4, 9,
    -- filter=154 channel=32
    5, -4, -12, 1, -8, -10, 3, 2, -2,
    -- filter=154 channel=33
    6, 1, -20, 12, 0, -7, 7, 5, -10,
    -- filter=154 channel=34
    -5, -13, 1, -5, -27, -5, 1, -20, -9,
    -- filter=154 channel=35
    7, -7, 6, 2, -7, 4, -6, 7, -3,
    -- filter=154 channel=36
    -9, 8, 12, -6, 12, 10, -10, 2, 6,
    -- filter=154 channel=37
    6, -14, -27, 14, -26, -29, 18, -1, -12,
    -- filter=154 channel=38
    7, 0, -4, -2, 1, 7, 0, 2, -7,
    -- filter=154 channel=39
    7, 6, 8, 8, -1, 7, -3, -6, 6,
    -- filter=154 channel=40
    -8, 1, -2, 6, 0, 7, -8, 0, 0,
    -- filter=154 channel=41
    -9, -16, -5, -1, -14, -24, 0, -10, -8,
    -- filter=154 channel=42
    1, -5, -10, 3, -3, -1, 10, 1, 0,
    -- filter=154 channel=43
    -5, -9, -8, 3, -8, -8, 5, 0, -6,
    -- filter=154 channel=44
    10, 0, -19, 8, -6, -8, 12, 7, -2,
    -- filter=154 channel=45
    9, 1, 4, 6, -1, -6, 9, -2, -2,
    -- filter=154 channel=46
    -2, -4, -1, -8, 1, -11, 4, -10, -6,
    -- filter=154 channel=47
    5, 0, -7, 5, 2, -17, -4, 1, -10,
    -- filter=154 channel=48
    7, 6, -14, 15, -3, -2, 10, 4, -4,
    -- filter=154 channel=49
    14, 5, -5, 3, 2, 4, 4, 7, 0,
    -- filter=154 channel=50
    12, -2, -2, 3, 9, 10, 10, 9, 7,
    -- filter=154 channel=51
    -7, 4, 4, -3, 0, 3, 0, 7, 3,
    -- filter=154 channel=52
    -8, -7, -1, -5, -12, 0, -8, -7, -6,
    -- filter=154 channel=53
    0, 3, 13, 4, 0, 13, -3, -1, 7,
    -- filter=154 channel=54
    -2, 6, 6, -5, -3, 2, 0, 4, 4,
    -- filter=154 channel=55
    0, 6, 4, -2, 0, 20, -12, -8, 1,
    -- filter=154 channel=56
    -11, -3, -6, -4, -11, -8, -10, -9, -6,
    -- filter=154 channel=57
    4, 1, 3, 4, -8, -5, 0, -10, -5,
    -- filter=154 channel=58
    0, 1, -14, -2, -8, -5, 8, -3, -13,
    -- filter=154 channel=59
    -1, 7, -1, 0, 2, -3, -2, 8, -6,
    -- filter=154 channel=60
    -4, 2, 1, -4, 5, -4, -1, 1, -4,
    -- filter=154 channel=61
    -9, -9, 6, -12, -4, 6, -8, 0, 0,
    -- filter=154 channel=62
    3, -6, -4, -6, -1, -2, -4, -3, 3,
    -- filter=154 channel=63
    7, -5, -2, 3, 0, -3, -1, 4, -4,
    -- filter=154 channel=64
    -3, 4, 0, -10, 5, 0, 1, -3, 2,
    -- filter=154 channel=65
    1, 3, -5, -6, 0, -1, 0, -4, 3,
    -- filter=154 channel=66
    -1, -2, 4, -3, -9, -15, -10, -6, 3,
    -- filter=154 channel=67
    5, 1, 2, 2, -5, -5, 5, 5, 4,
    -- filter=154 channel=68
    2, -2, 0, 7, 2, 8, -5, -4, -2,
    -- filter=154 channel=69
    -2, -5, -1, 5, -4, 0, 4, 2, 1,
    -- filter=154 channel=70
    2, -12, -9, 4, -12, -10, 1, -11, -10,
    -- filter=154 channel=71
    4, -4, 3, 5, 0, -7, 4, 5, 1,
    -- filter=154 channel=72
    7, 5, 7, 5, 20, 8, 2, 9, -1,
    -- filter=154 channel=73
    5, 5, 1, 4, -4, 11, -1, -6, -8,
    -- filter=154 channel=74
    2, -11, 0, -3, -6, -1, 5, -7, -1,
    -- filter=154 channel=75
    -7, -21, -30, 8, -25, -32, 9, 1, -20,
    -- filter=154 channel=76
    -4, 4, 20, -8, 3, 9, -13, -2, 12,
    -- filter=154 channel=77
    3, 7, 2, 0, 2, 6, 2, 2, 0,
    -- filter=154 channel=78
    6, -2, -7, 4, -8, 0, 9, 0, 4,
    -- filter=154 channel=79
    10, -7, -20, 11, -9, -18, 9, -9, -19,
    -- filter=154 channel=80
    10, 4, 3, 8, 20, 0, 1, 11, 3,
    -- filter=154 channel=81
    4, 5, 7, 4, 2, 6, -2, 7, 0,
    -- filter=154 channel=82
    -3, -5, -8, 1, -4, 2, -5, 7, 5,
    -- filter=154 channel=83
    2, -2, -2, 8, 7, 4, 5, 9, -5,
    -- filter=154 channel=84
    5, 0, -6, 5, -7, 2, 8, -13, 0,
    -- filter=154 channel=85
    5, 3, 0, 5, -5, 4, 6, 1, 2,
    -- filter=154 channel=86
    -5, -14, 0, -1, -13, -16, -1, -1, -9,
    -- filter=154 channel=87
    2, -13, 13, -1, -3, 3, -14, -4, 6,
    -- filter=154 channel=88
    -5, -2, 18, 0, 5, 20, -2, -5, 10,
    -- filter=154 channel=89
    5, 3, 1, 5, 13, 9, 0, 5, 0,
    -- filter=154 channel=90
    -8, -3, 11, -13, -4, 13, -9, -14, -2,
    -- filter=154 channel=91
    7, -2, 5, 10, 5, 9, 3, 6, -5,
    -- filter=154 channel=92
    -9, -9, 0, -2, -6, -4, 2, -9, -4,
    -- filter=154 channel=93
    3, -2, -16, 10, -11, -25, 7, 5, -9,
    -- filter=154 channel=94
    0, 6, -3, 2, 2, 0, -2, -4, 5,
    -- filter=154 channel=95
    3, -4, 1, -1, -8, -8, -2, -3, 1,
    -- filter=154 channel=96
    9, -2, -3, -2, 7, -5, 8, -3, 4,
    -- filter=154 channel=97
    -3, 1, -10, 6, 1, -10, 2, -6, 2,
    -- filter=154 channel=98
    9, 4, -9, 14, 9, -2, 5, 5, -11,
    -- filter=154 channel=99
    -5, 0, 20, 0, 3, 32, -16, 0, 10,
    -- filter=154 channel=100
    1, 2, 3, 5, 0, 5, 0, -2, -3,
    -- filter=154 channel=101
    5, 0, -3, -11, 2, -7, -5, -5, 3,
    -- filter=154 channel=102
    -4, -4, 6, -3, 3, -1, -4, 0, 1,
    -- filter=154 channel=103
    1, 1, -17, 15, 0, -14, 6, 9, -5,
    -- filter=154 channel=104
    4, 6, 2, 1, 21, 2, -1, 9, 1,
    -- filter=154 channel=105
    5, 4, 0, 0, -6, 0, -1, 2, 11,
    -- filter=154 channel=106
    0, -1, 1, 1, -3, 7, -7, -4, 11,
    -- filter=154 channel=107
    5, -8, -10, 0, -16, -9, -5, -11, -3,
    -- filter=154 channel=108
    -7, -8, 1, -6, -12, -13, -1, -1, -6,
    -- filter=154 channel=109
    0, -11, -3, 3, -4, 5, 10, 7, -5,
    -- filter=154 channel=110
    0, 3, 0, 0, 9, 7, -4, -1, 2,
    -- filter=154 channel=111
    6, 0, -3, -5, -4, 0, -2, 1, 0,
    -- filter=154 channel=112
    0, -5, -5, 1, -5, -7, 9, -7, -2,
    -- filter=154 channel=113
    5, -7, -11, -2, 5, 1, 6, 0, -6,
    -- filter=154 channel=114
    18, -11, -22, 18, -25, -34, 19, -10, -30,
    -- filter=154 channel=115
    -2, -1, -1, -1, 6, 1, -5, 5, 2,
    -- filter=154 channel=116
    4, 9, 2, 10, 17, 8, 3, 1, -1,
    -- filter=154 channel=117
    -5, -1, 6, -4, 1, 1, -1, 6, -1,
    -- filter=154 channel=118
    3, 3, -1, -5, -2, 6, -5, 7, 3,
    -- filter=154 channel=119
    -4, -14, -6, -2, -14, -9, -1, -13, 0,
    -- filter=154 channel=120
    13, -4, 14, 2, -1, 16, 13, 2, 0,
    -- filter=154 channel=121
    -7, -4, -3, 0, 0, -9, -12, -12, 2,
    -- filter=154 channel=122
    2, 0, -13, 8, 13, -5, 1, -3, -4,
    -- filter=154 channel=123
    -11, -5, 2, -1, -1, -3, 0, -8, -6,
    -- filter=154 channel=124
    -3, 1, 7, 3, 3, 4, -2, 1, -2,
    -- filter=154 channel=125
    0, 1, 9, -4, 19, 9, -2, 10, 3,
    -- filter=154 channel=126
    -6, 0, -7, 7, -1, -1, 5, 0, 5,
    -- filter=154 channel=127
    3, -3, 0, 3, 2, -4, -6, 4, 4,
    -- filter=155 channel=0
    -4, -10, -12, -4, -7, -2, 4, 3, -4,
    -- filter=155 channel=1
    -1, -3, 2, 1, -3, -6, 6, 1, 6,
    -- filter=155 channel=2
    0, 2, 0, -6, 7, 4, -2, 7, 12,
    -- filter=155 channel=3
    -7, -18, -2, -6, -10, 0, -10, -1, 2,
    -- filter=155 channel=4
    -15, -8, -5, -10, 0, 4, -3, 3, 9,
    -- filter=155 channel=5
    -2, -6, 1, -6, -13, -7, 11, 3, 1,
    -- filter=155 channel=6
    2, -6, -1, 0, -1, -3, -6, 4, 5,
    -- filter=155 channel=7
    4, 2, -5, 3, -6, 4, 0, -4, 0,
    -- filter=155 channel=8
    -11, 1, -4, -2, 2, 2, -6, 6, -1,
    -- filter=155 channel=9
    -4, -4, 1, 7, 1, -2, 0, 3, 10,
    -- filter=155 channel=10
    -7, -4, -5, -4, -4, -7, 0, -2, -9,
    -- filter=155 channel=11
    0, 6, 6, 1, 0, 9, -7, -4, 0,
    -- filter=155 channel=12
    -4, 1, -4, -2, 4, -8, 2, -5, -5,
    -- filter=155 channel=13
    -5, -15, -9, -10, 0, -1, 3, -5, 10,
    -- filter=155 channel=14
    -1, 4, -6, 6, 6, 1, -3, 3, 1,
    -- filter=155 channel=15
    -9, -10, -14, 0, -5, -6, 6, 4, 7,
    -- filter=155 channel=16
    5, -6, 8, 4, -5, 2, -6, -3, -10,
    -- filter=155 channel=17
    3, -7, -5, 0, 0, 3, -5, -2, 2,
    -- filter=155 channel=18
    -9, -5, -18, -3, 4, 2, 2, 2, 21,
    -- filter=155 channel=19
    -2, 2, -2, -6, -2, 7, 0, 5, 0,
    -- filter=155 channel=20
    7, 6, -2, -2, 2, 8, 3, 0, 12,
    -- filter=155 channel=21
    -3, 0, 4, -1, -2, 2, 9, 8, -4,
    -- filter=155 channel=22
    -5, -5, -5, 1, -2, 3, -2, -5, 5,
    -- filter=155 channel=23
    3, -15, -19, 8, 0, 0, 0, 7, 11,
    -- filter=155 channel=24
    -5, 4, 4, 5, 5, -6, 6, 2, 1,
    -- filter=155 channel=25
    -8, -2, -5, -6, 0, -6, -3, 7, 13,
    -- filter=155 channel=26
    5, 2, 10, 4, 7, 7, -4, 6, 4,
    -- filter=155 channel=27
    -3, -11, -16, 3, 1, -6, 5, 16, 16,
    -- filter=155 channel=28
    6, -1, 0, 3, -4, -5, 4, 5, -3,
    -- filter=155 channel=29
    8, 2, -3, 7, 5, 2, 0, 0, 14,
    -- filter=155 channel=30
    4, -13, -1, 3, 1, 0, -2, 4, 15,
    -- filter=155 channel=31
    0, -3, -1, 6, -2, -10, 6, 11, 3,
    -- filter=155 channel=32
    0, -6, -9, 1, -2, 4, 3, 0, 14,
    -- filter=155 channel=33
    -12, -13, -7, 3, 0, -10, -5, -1, 8,
    -- filter=155 channel=34
    -4, 1, -2, -4, -7, -1, 5, 4, -7,
    -- filter=155 channel=35
    1, 0, -5, -7, 1, -6, 0, -7, -6,
    -- filter=155 channel=36
    7, 2, 0, 2, -1, 9, -3, 3, -3,
    -- filter=155 channel=37
    0, -15, -4, 1, -11, -1, 7, 0, 5,
    -- filter=155 channel=38
    1, -12, 0, 6, -4, 1, 0, 5, 3,
    -- filter=155 channel=39
    7, 0, -3, -2, 0, 4, 6, 3, 4,
    -- filter=155 channel=40
    -4, 6, -1, 3, -5, 5, 2, -2, 5,
    -- filter=155 channel=41
    5, 5, -16, 3, 10, -13, -2, -16, -14,
    -- filter=155 channel=42
    4, 0, 2, 7, -6, -5, 6, -2, 4,
    -- filter=155 channel=43
    0, -8, 0, -1, -5, -7, -7, -1, -3,
    -- filter=155 channel=44
    4, -2, 4, -3, -8, 0, -1, 5, -2,
    -- filter=155 channel=45
    -2, 6, 4, -3, -3, 7, -5, -2, 2,
    -- filter=155 channel=46
    2, -2, -6, 5, 3, 5, 1, -6, -6,
    -- filter=155 channel=47
    -2, -7, 5, -9, 0, 5, -3, 2, 0,
    -- filter=155 channel=48
    -9, 5, 4, 0, 10, 0, 10, 15, 16,
    -- filter=155 channel=49
    2, -6, -5, 6, 0, 5, 4, 0, 9,
    -- filter=155 channel=50
    6, 0, -5, 4, 3, 5, 2, 12, 3,
    -- filter=155 channel=51
    3, 0, 0, -2, 3, -5, 4, 1, -1,
    -- filter=155 channel=52
    -5, 0, -4, 2, -1, 0, -5, 0, 8,
    -- filter=155 channel=53
    -4, -5, 2, 4, -2, -1, 1, -1, -1,
    -- filter=155 channel=54
    -6, 5, -5, -6, 4, 0, -3, 7, 2,
    -- filter=155 channel=55
    -9, -15, -6, -1, 2, 0, -6, -4, 12,
    -- filter=155 channel=56
    -9, -4, -6, 5, -7, -2, -3, 0, 2,
    -- filter=155 channel=57
    4, 0, -1, 0, 6, -2, -5, -2, 5,
    -- filter=155 channel=58
    -7, -9, -8, -1, -6, 0, -4, 1, 1,
    -- filter=155 channel=59
    -8, 0, 1, 1, 11, 6, -5, 9, 2,
    -- filter=155 channel=60
    4, 0, -2, -4, 6, 0, -5, 1, 3,
    -- filter=155 channel=61
    -4, -4, 5, 5, 0, 6, 2, -4, 4,
    -- filter=155 channel=62
    -5, 4, 2, -3, -1, 4, 6, -5, -6,
    -- filter=155 channel=63
    -3, -2, 0, -4, 0, -5, 3, 0, -8,
    -- filter=155 channel=64
    2, -2, 7, -2, 1, 1, -7, -4, -7,
    -- filter=155 channel=65
    -2, -1, -6, 6, -4, 3, -5, -7, -3,
    -- filter=155 channel=66
    -2, -11, -6, -9, -1, 0, -1, -11, -1,
    -- filter=155 channel=67
    -3, -4, -6, 1, 2, -8, -1, 3, -1,
    -- filter=155 channel=68
    -2, 8, 6, 4, 0, 3, 4, -1, 3,
    -- filter=155 channel=69
    0, 5, -4, -7, 5, 3, 2, 3, 2,
    -- filter=155 channel=70
    0, -10, -4, 4, 4, 0, 0, 0, 4,
    -- filter=155 channel=71
    5, -5, -6, -4, -3, -2, -1, -3, -7,
    -- filter=155 channel=72
    -3, -2, -10, 0, 8, -7, 0, 11, 5,
    -- filter=155 channel=73
    2, -3, -5, -1, 2, 9, 4, 0, 17,
    -- filter=155 channel=74
    -4, -2, -6, 3, 4, -1, 10, 2, 9,
    -- filter=155 channel=75
    -11, -20, -8, -11, -11, -10, 0, 5, -3,
    -- filter=155 channel=76
    1, 1, 10, 3, 1, 4, 6, 0, 7,
    -- filter=155 channel=77
    1, 2, -6, -4, 0, 4, 0, -3, -1,
    -- filter=155 channel=78
    -6, -4, -2, -6, 0, -6, 1, -5, 2,
    -- filter=155 channel=79
    -2, -16, -19, 0, -7, -8, 0, 6, 16,
    -- filter=155 channel=80
    3, -5, 5, -1, 2, 0, -3, 9, 8,
    -- filter=155 channel=81
    7, 5, -5, 0, 3, -6, 1, -7, -1,
    -- filter=155 channel=82
    4, -7, -3, 5, -1, 1, 4, 5, -7,
    -- filter=155 channel=83
    -7, 4, -3, -3, 2, -1, 6, 12, 6,
    -- filter=155 channel=84
    -7, 0, -6, -2, 5, 3, -3, 6, 9,
    -- filter=155 channel=85
    2, -4, -7, -6, -6, -1, -4, -4, -3,
    -- filter=155 channel=86
    4, -11, 7, -3, -1, -7, 5, 4, 1,
    -- filter=155 channel=87
    -1, -4, 2, 0, -6, -5, -2, -3, 6,
    -- filter=155 channel=88
    4, 12, 3, 5, 3, 2, 8, 7, -5,
    -- filter=155 channel=89
    -9, -17, -6, 2, 3, -12, 5, 2, 0,
    -- filter=155 channel=90
    4, -1, -1, -1, 0, 7, 1, 3, -2,
    -- filter=155 channel=91
    -2, -11, -12, 6, 1, 6, -1, 14, 19,
    -- filter=155 channel=92
    -9, -7, -9, 2, -9, -8, 0, 5, -6,
    -- filter=155 channel=93
    -10, -6, -5, -3, -6, -7, 9, 10, 5,
    -- filter=155 channel=94
    3, 3, 1, -5, 0, 6, -2, 7, 2,
    -- filter=155 channel=95
    -3, 3, 3, 1, -5, 0, -4, -7, -4,
    -- filter=155 channel=96
    0, 0, -7, -1, 3, 6, -4, 7, -3,
    -- filter=155 channel=97
    -8, -4, -10, -1, -4, 1, -6, 3, -8,
    -- filter=155 channel=98
    1, -7, -13, -2, -2, 0, -6, 2, 7,
    -- filter=155 channel=99
    -4, -12, -3, 1, 1, -7, 0, 12, 0,
    -- filter=155 channel=100
    4, 0, -5, -3, 5, -2, 1, 3, 1,
    -- filter=155 channel=101
    -6, -8, -6, 1, 0, 6, 0, 5, 2,
    -- filter=155 channel=102
    -2, -4, 0, 7, 0, 3, -5, 5, 4,
    -- filter=155 channel=103
    -5, -6, -7, -5, -2, 0, 6, 9, -7,
    -- filter=155 channel=104
    -1, -4, 3, 4, 4, -4, 0, 11, 4,
    -- filter=155 channel=105
    3, 1, 0, 3, -9, 6, -6, -4, -5,
    -- filter=155 channel=106
    -1, 4, -5, 0, 0, 0, 3, -7, -1,
    -- filter=155 channel=107
    -1, -3, 0, 4, -6, 8, -3, -4, 7,
    -- filter=155 channel=108
    -8, 0, 1, -3, -5, 4, -1, -4, -9,
    -- filter=155 channel=109
    -7, -12, -2, 3, 9, 3, 8, 13, 23,
    -- filter=155 channel=110
    -2, 0, -11, -3, -10, -2, 2, 1, 1,
    -- filter=155 channel=111
    -1, -1, -6, -7, 0, 0, 5, 3, 3,
    -- filter=155 channel=112
    3, -4, -5, 7, -1, 4, -4, 0, 10,
    -- filter=155 channel=113
    -2, -8, -7, -2, -7, -14, 5, 6, 0,
    -- filter=155 channel=114
    -6, -15, -16, 5, -6, -2, -5, 5, 25,
    -- filter=155 channel=115
    4, -2, -4, 0, -4, 0, 5, 3, -1,
    -- filter=155 channel=116
    3, -4, -6, 3, 3, 8, 5, 0, 7,
    -- filter=155 channel=117
    -2, 5, -2, 7, 2, -1, 5, 2, 3,
    -- filter=155 channel=118
    1, -1, -6, 0, 0, -3, 6, -2, -4,
    -- filter=155 channel=119
    0, -2, -7, 8, 0, -5, 4, 2, -8,
    -- filter=155 channel=120
    1, -11, -2, 10, 1, -4, 5, 12, 15,
    -- filter=155 channel=121
    0, -6, 1, 3, -2, -6, 0, -4, -2,
    -- filter=155 channel=122
    4, -2, 13, 1, 5, 0, 5, 6, -2,
    -- filter=155 channel=123
    -4, -10, -6, -4, -7, 4, -5, -1, -5,
    -- filter=155 channel=124
    -1, 1, -1, 6, 2, -3, 6, -8, 1,
    -- filter=155 channel=125
    4, -12, -9, 4, 10, 6, -5, 18, 18,
    -- filter=155 channel=126
    -9, -8, -9, -11, -3, -3, 0, -4, -7,
    -- filter=155 channel=127
    -4, -2, 0, 2, -2, -4, -3, 2, -7,
    -- filter=156 channel=0
    13, 1, -8, 12, -1, -16, 12, -5, -10,
    -- filter=156 channel=1
    6, 13, -3, 11, 8, 0, 9, 1, -8,
    -- filter=156 channel=2
    5, -3, 6, -1, 5, -8, -9, 0, 5,
    -- filter=156 channel=3
    -6, 3, -3, 15, -6, -18, 3, -7, -13,
    -- filter=156 channel=4
    5, 1, 0, 11, 0, -11, 0, 0, -11,
    -- filter=156 channel=5
    4, -10, -5, 3, -17, -12, -2, -8, -13,
    -- filter=156 channel=6
    -8, -7, 2, 3, -3, -9, -9, -5, -8,
    -- filter=156 channel=7
    4, 5, -2, 0, -1, -2, 5, 0, 3,
    -- filter=156 channel=8
    -2, 0, 8, -3, 2, 10, -1, 5, 4,
    -- filter=156 channel=9
    7, 0, -2, 0, -5, -7, -6, -8, 2,
    -- filter=156 channel=10
    -4, -7, 0, 0, -3, 2, -2, -11, 5,
    -- filter=156 channel=11
    0, -6, -12, 7, -2, -3, -6, -3, -11,
    -- filter=156 channel=12
    -3, -2, 9, 1, 8, 9, 0, -2, 6,
    -- filter=156 channel=13
    -5, 7, 1, 0, 9, -4, -2, 2, 0,
    -- filter=156 channel=14
    4, -7, 5, -4, 5, 7, -1, -2, -7,
    -- filter=156 channel=15
    -6, 4, -6, 3, 8, -2, 8, 0, 1,
    -- filter=156 channel=16
    1, -8, 12, -2, -12, 11, -6, -12, 11,
    -- filter=156 channel=17
    -3, 4, -5, -3, 6, -3, -4, -7, 0,
    -- filter=156 channel=18
    -4, 9, 0, 15, 12, -3, -9, -2, -7,
    -- filter=156 channel=19
    0, 4, 5, 0, -7, 6, 6, 3, 0,
    -- filter=156 channel=20
    2, 2, -6, 8, 6, -2, -2, 4, -13,
    -- filter=156 channel=21
    2, -14, 5, -12, -17, 6, -5, -6, 6,
    -- filter=156 channel=22
    4, 0, 4, 1, -3, 6, 8, 3, 0,
    -- filter=156 channel=23
    -3, 7, 6, 3, 0, 16, -1, -2, 1,
    -- filter=156 channel=24
    0, 4, -5, 0, 1, -4, -5, -4, 0,
    -- filter=156 channel=25
    -3, 6, 5, -5, 2, -2, -12, 2, -4,
    -- filter=156 channel=26
    0, -11, 5, 0, -17, 1, 0, -14, -1,
    -- filter=156 channel=27
    -1, -5, 11, 18, -1, 11, 0, 0, 2,
    -- filter=156 channel=28
    -1, -4, 0, 6, 2, 0, 7, -6, 3,
    -- filter=156 channel=29
    -6, -2, -15, 0, 0, -14, -1, -5, -16,
    -- filter=156 channel=30
    9, 6, 0, 15, -1, -7, 10, 1, -1,
    -- filter=156 channel=31
    -2, -15, 10, -14, -16, 19, -7, 0, 18,
    -- filter=156 channel=32
    -5, 2, -4, 8, 9, -1, -6, -4, -14,
    -- filter=156 channel=33
    0, 11, 3, 11, -1, -10, -3, 0, 0,
    -- filter=156 channel=34
    -10, 0, 18, -2, 1, 19, -6, -6, 16,
    -- filter=156 channel=35
    0, 0, 6, 4, -1, 4, 2, 2, -4,
    -- filter=156 channel=36
    -7, -10, 11, -9, -2, 13, -5, 6, 4,
    -- filter=156 channel=37
    19, 4, -3, 5, -4, 6, 14, 3, 4,
    -- filter=156 channel=38
    -2, 3, 2, 2, -3, -8, 5, -11, -5,
    -- filter=156 channel=39
    -7, 2, -11, 10, -2, -2, -2, 3, -13,
    -- filter=156 channel=40
    4, 11, -3, 10, 4, 7, 10, 12, 6,
    -- filter=156 channel=41
    -12, -8, 6, -12, -2, -3, -15, -15, 3,
    -- filter=156 channel=42
    8, 5, -8, 9, -6, -6, 11, -3, 0,
    -- filter=156 channel=43
    0, 6, -12, 5, 0, -5, 1, -8, -8,
    -- filter=156 channel=44
    11, 0, 6, -3, -9, 13, 9, 1, 13,
    -- filter=156 channel=45
    2, 10, 1, 13, -1, 4, 4, 2, -7,
    -- filter=156 channel=46
    0, 5, 9, 2, 3, 5, -5, -7, 3,
    -- filter=156 channel=47
    11, -8, 3, 3, -16, 0, -4, -11, 6,
    -- filter=156 channel=48
    0, 2, 10, 8, -8, 11, -7, 2, 7,
    -- filter=156 channel=49
    6, 3, -2, 8, 0, -5, 3, 3, -13,
    -- filter=156 channel=50
    -3, 0, 15, 1, 0, 6, 12, 7, 7,
    -- filter=156 channel=51
    -2, 4, -2, -5, -7, 0, -1, 0, 6,
    -- filter=156 channel=52
    -2, -1, 6, -9, -5, 16, 4, 4, 5,
    -- filter=156 channel=53
    -6, -8, 0, 6, 5, -4, -7, 2, -7,
    -- filter=156 channel=54
    -4, 6, 0, 0, 6, 5, 4, -4, -1,
    -- filter=156 channel=55
    -14, 4, -5, -3, -1, 0, -8, -6, 2,
    -- filter=156 channel=56
    -1, -3, 3, -1, -2, 15, 2, 3, 13,
    -- filter=156 channel=57
    -1, 5, 0, 0, -5, 2, 3, 1, 0,
    -- filter=156 channel=58
    -7, -7, -2, 3, -10, -8, -6, -6, -14,
    -- filter=156 channel=59
    1, -1, 0, 1, -8, 5, -1, -2, 13,
    -- filter=156 channel=60
    -1, -5, 6, -4, -5, 1, -1, -1, -4,
    -- filter=156 channel=61
    -5, 1, -6, -8, 3, 4, -5, -2, -2,
    -- filter=156 channel=62
    0, -5, 5, 1, -4, -5, -7, 4, -4,
    -- filter=156 channel=63
    0, -7, -9, -9, -9, -3, -12, -14, -9,
    -- filter=156 channel=64
    -6, 3, 2, 0, -2, 4, 0, 1, 9,
    -- filter=156 channel=65
    7, -4, 5, 0, 2, -1, 5, -1, -4,
    -- filter=156 channel=66
    -12, -2, 9, -13, -3, 2, -6, 0, 0,
    -- filter=156 channel=67
    -3, 5, -1, -7, 2, 11, 3, -8, 0,
    -- filter=156 channel=68
    8, 7, 0, 0, 3, -4, -7, 1, 6,
    -- filter=156 channel=69
    0, 0, 5, -5, 6, -2, -8, 1, 3,
    -- filter=156 channel=70
    1, 11, 20, 15, 17, 17, 6, 12, 13,
    -- filter=156 channel=71
    -1, 7, -2, 1, 6, 0, 0, 7, 5,
    -- filter=156 channel=72
    -6, -3, 10, -6, -14, 2, -7, -13, 13,
    -- filter=156 channel=73
    -11, 2, -4, 0, 2, 5, -11, 0, -3,
    -- filter=156 channel=74
    -3, -3, 10, -7, -2, 25, -5, 7, 15,
    -- filter=156 channel=75
    0, 6, -4, 11, -6, -11, 1, -2, -9,
    -- filter=156 channel=76
    -6, 5, -3, 10, 8, -9, 4, 11, -3,
    -- filter=156 channel=77
    -3, -4, 4, 6, -4, 5, -6, -1, 2,
    -- filter=156 channel=78
    1, 0, 1, 5, -11, 2, 2, -12, -5,
    -- filter=156 channel=79
    1, 5, -6, 26, 20, -8, 2, 6, -11,
    -- filter=156 channel=80
    -6, -6, 5, 1, -19, 0, -9, -5, 16,
    -- filter=156 channel=81
    0, 0, -6, 1, 1, 5, 5, -2, 4,
    -- filter=156 channel=82
    -5, 4, -4, -2, -1, 4, -1, -1, -3,
    -- filter=156 channel=83
    6, -6, 2, 4, -1, -4, 1, -8, 5,
    -- filter=156 channel=84
    -5, 0, 1, 8, 4, 0, 0, -8, 3,
    -- filter=156 channel=85
    0, -3, -4, -4, 5, 3, 5, -1, -6,
    -- filter=156 channel=86
    6, -4, -4, 3, 0, 2, 0, -5, -3,
    -- filter=156 channel=87
    0, -9, -3, -6, 6, 9, -8, -7, 0,
    -- filter=156 channel=88
    -5, -9, 12, -4, -16, 6, -5, 4, 16,
    -- filter=156 channel=89
    -11, -2, 5, 7, -5, 5, -9, 0, 0,
    -- filter=156 channel=90
    -2, -11, 9, -7, -10, 21, -1, 0, 12,
    -- filter=156 channel=91
    0, -1, 5, 16, 10, 9, -9, 2, 0,
    -- filter=156 channel=92
    3, 7, 13, -5, -1, 14, -4, -5, 1,
    -- filter=156 channel=93
    13, 2, 0, 0, -10, 0, -6, -7, 3,
    -- filter=156 channel=94
    2, 0, 2, -6, 0, 1, -4, 1, 0,
    -- filter=156 channel=95
    1, 2, 3, -3, 3, -8, -6, 0, 3,
    -- filter=156 channel=96
    1, 6, -5, 1, 3, -6, 5, 2, -5,
    -- filter=156 channel=97
    -5, 3, 2, 1, 4, 2, 5, 3, 4,
    -- filter=156 channel=98
    0, -6, -3, 3, -4, -1, -5, -6, -6,
    -- filter=156 channel=99
    -12, -18, 0, -20, -23, 10, -18, -16, 15,
    -- filter=156 channel=100
    -5, -2, 1, -7, -4, 7, -1, -2, 6,
    -- filter=156 channel=101
    -5, -9, 0, 3, 3, -12, 0, -9, -2,
    -- filter=156 channel=102
    -5, -5, 4, 0, -2, -5, 5, 0, -2,
    -- filter=156 channel=103
    6, -6, -3, -4, -18, 10, -5, 0, 6,
    -- filter=156 channel=104
    -1, -10, -3, -3, -13, 9, -2, -7, 16,
    -- filter=156 channel=105
    -5, -1, -12, -3, 3, -5, -1, 3, -13,
    -- filter=156 channel=106
    -6, 7, 2, 1, -4, 7, 0, 0, 6,
    -- filter=156 channel=107
    6, 8, 0, 16, 1, -4, 8, -2, 0,
    -- filter=156 channel=108
    0, 0, -2, -3, 3, -12, -6, -7, -2,
    -- filter=156 channel=109
    -7, -5, 0, -7, -7, 0, -17, -10, 11,
    -- filter=156 channel=110
    -4, -3, 0, -1, -5, -5, -11, -2, 0,
    -- filter=156 channel=111
    0, -4, 3, -2, -5, -4, -6, 2, -4,
    -- filter=156 channel=112
    4, -2, 6, 0, -6, 13, -2, 0, 9,
    -- filter=156 channel=113
    -5, 6, 9, 7, -12, 8, 0, -3, 5,
    -- filter=156 channel=114
    4, 7, -8, 17, 9, -18, -6, -2, -12,
    -- filter=156 channel=115
    -8, 4, 1, -6, 4, -8, 0, -2, -5,
    -- filter=156 channel=116
    -14, -2, -6, -8, -13, 3, -10, -11, 0,
    -- filter=156 channel=117
    4, 0, -5, 0, -3, -3, 3, 6, -5,
    -- filter=156 channel=118
    1, -5, 4, 1, -7, -7, 5, -2, 4,
    -- filter=156 channel=119
    -5, -10, 16, -20, 4, 36, -11, -3, 20,
    -- filter=156 channel=120
    -2, -10, 3, 8, -11, 14, -10, -5, 9,
    -- filter=156 channel=121
    -11, -6, 11, -4, -7, -1, -1, 0, 0,
    -- filter=156 channel=122
    11, -10, 23, -3, -28, 24, 6, -11, 25,
    -- filter=156 channel=123
    -8, 2, 6, -4, -4, 16, -3, 1, 11,
    -- filter=156 channel=124
    0, -5, -6, 5, 4, 2, 2, -4, -6,
    -- filter=156 channel=125
    -4, -8, 5, -5, -11, 12, -17, -5, 14,
    -- filter=156 channel=126
    -14, -5, -5, 5, -7, -6, 0, -4, -9,
    -- filter=156 channel=127
    -11, -5, -2, -9, -3, -4, -1, -1, 0,
    -- filter=157 channel=0
    5, 4, 11, 0, -5, 0, -11, 3, -9,
    -- filter=157 channel=1
    13, 2, 2, -10, 5, -11, -10, 5, 1,
    -- filter=157 channel=2
    -8, -5, 2, 5, -1, -5, 8, 3, 1,
    -- filter=157 channel=3
    13, 2, 1, -2, 6, -2, 1, 7, 2,
    -- filter=157 channel=4
    -4, 9, -4, 17, 11, -4, 14, -13, 1,
    -- filter=157 channel=5
    11, 5, 6, -8, 0, -1, 0, 7, -4,
    -- filter=157 channel=6
    0, 0, 4, 6, 3, -5, 0, 0, -1,
    -- filter=157 channel=7
    -1, 6, 0, -4, -6, 0, 5, -2, -2,
    -- filter=157 channel=8
    0, 10, -4, 13, -3, 3, 7, -4, 4,
    -- filter=157 channel=9
    -8, -8, 7, 0, -1, 6, 7, -1, 2,
    -- filter=157 channel=10
    -8, -8, -4, -2, 0, 0, 3, 14, 3,
    -- filter=157 channel=11
    -5, 0, 5, 6, 9, -1, 4, -6, 0,
    -- filter=157 channel=12
    7, -3, -1, -8, 7, -5, -3, -1, -7,
    -- filter=157 channel=13
    4, -6, -1, -6, 3, 2, 1, 12, -10,
    -- filter=157 channel=14
    6, -4, -7, -4, 6, 6, -1, 7, 4,
    -- filter=157 channel=15
    -5, 2, 0, -7, -3, -1, 5, 0, -4,
    -- filter=157 channel=16
    1, 6, 2, -2, -8, 0, -3, 4, -1,
    -- filter=157 channel=17
    5, 0, -1, 5, -4, -4, -3, 2, 7,
    -- filter=157 channel=18
    -10, 2, 2, -19, 7, 2, 1, 2, -10,
    -- filter=157 channel=19
    -2, 1, 1, 7, -4, -1, 6, 3, 4,
    -- filter=157 channel=20
    -9, 11, -1, -2, 11, -8, -3, 3, 0,
    -- filter=157 channel=21
    -7, -9, -4, -2, -3, -1, 2, 9, 0,
    -- filter=157 channel=22
    6, 10, 6, 2, 5, -6, -2, -3, 1,
    -- filter=157 channel=23
    -8, 5, -4, -14, 8, -8, 5, 2, 1,
    -- filter=157 channel=24
    -1, 3, 1, -6, -3, -6, -5, -3, 6,
    -- filter=157 channel=25
    -7, 5, -8, -20, 6, -3, 5, 10, -4,
    -- filter=157 channel=26
    -3, -5, 1, 4, 5, -1, 0, 0, -4,
    -- filter=157 channel=27
    -16, 7, 1, -5, 11, -8, 16, 0, -2,
    -- filter=157 channel=28
    0, -6, -3, -3, -7, -7, -6, 1, 1,
    -- filter=157 channel=29
    0, 6, -1, 4, 11, -5, 2, -3, -4,
    -- filter=157 channel=30
    -8, 9, 8, -9, -1, 0, 0, -3, -2,
    -- filter=157 channel=31
    -17, 0, 1, -15, -2, 4, 9, 1, 12,
    -- filter=157 channel=32
    -12, 8, -4, -21, 11, -10, -2, -1, -1,
    -- filter=157 channel=33
    -7, 3, 6, -20, 1, 0, -4, 13, 1,
    -- filter=157 channel=34
    -5, 14, -7, 6, 4, -4, 3, -1, -6,
    -- filter=157 channel=35
    1, 2, 4, 6, -7, 2, -4, 0, -4,
    -- filter=157 channel=36
    -8, -3, 2, 8, -1, 2, 12, -4, 6,
    -- filter=157 channel=37
    5, 7, -4, -6, -2, -9, 4, -1, -7,
    -- filter=157 channel=38
    3, 4, 1, -7, 5, 0, 4, 2, -2,
    -- filter=157 channel=39
    -2, 8, 0, -7, 1, 1, 6, 3, -7,
    -- filter=157 channel=40
    -5, 7, -4, 1, 0, 0, 1, 6, -5,
    -- filter=157 channel=41
    0, 1, -1, -8, 8, 1, -14, 11, 0,
    -- filter=157 channel=42
    -1, 0, 0, 1, -2, -6, 4, 0, 6,
    -- filter=157 channel=43
    7, -2, -4, -12, -2, 2, -2, 0, 4,
    -- filter=157 channel=44
    -3, 10, -8, 0, -2, -4, 5, 1, 3,
    -- filter=157 channel=45
    -1, 1, -6, 8, 7, -5, -6, 6, -5,
    -- filter=157 channel=46
    8, 0, -4, 0, 1, -4, -5, 0, 5,
    -- filter=157 channel=47
    0, 2, 0, -15, 0, -1, 0, 6, 3,
    -- filter=157 channel=48
    -4, -5, 3, -13, 5, -2, 19, 6, 5,
    -- filter=157 channel=49
    0, 10, -8, 0, 4, -8, 8, 0, -11,
    -- filter=157 channel=50
    -14, 4, -3, -9, 0, 6, 4, -7, 3,
    -- filter=157 channel=51
    3, 3, -2, -3, -5, -2, -1, 1, -2,
    -- filter=157 channel=52
    -11, 3, -6, 0, 0, 1, 8, -5, -8,
    -- filter=157 channel=53
    -4, 7, -4, 3, 0, 1, 6, -1, -6,
    -- filter=157 channel=54
    -3, -5, 2, -6, -6, -6, 0, -5, -6,
    -- filter=157 channel=55
    -11, 0, 5, -3, 0, 5, 12, 0, -3,
    -- filter=157 channel=56
    0, 5, -1, 0, -5, 3, -1, -4, -2,
    -- filter=157 channel=57
    0, 5, 3, 2, -4, -3, 4, 0, -6,
    -- filter=157 channel=58
    0, 6, 6, -2, 3, 0, -1, -5, 3,
    -- filter=157 channel=59
    -13, -7, -1, -14, 2, 0, 12, 11, 3,
    -- filter=157 channel=60
    -5, 5, -6, 5, 3, 5, 0, -1, 0,
    -- filter=157 channel=61
    -1, -2, -5, -6, -1, -2, -3, 3, 6,
    -- filter=157 channel=62
    -2, -4, -5, -4, 0, 4, 1, 5, -3,
    -- filter=157 channel=63
    9, -3, 2, -1, 0, -7, -6, 6, 4,
    -- filter=157 channel=64
    -2, -5, -3, 0, 3, 0, 1, 2, 1,
    -- filter=157 channel=65
    -7, -3, 5, -4, -2, -3, -1, 0, 1,
    -- filter=157 channel=66
    3, 0, -2, 0, 3, -1, 4, 3, -1,
    -- filter=157 channel=67
    7, 0, 3, 4, 6, 0, 2, -5, 4,
    -- filter=157 channel=68
    1, 0, 6, 2, 0, -2, 6, -5, 6,
    -- filter=157 channel=69
    0, 0, -5, 0, 1, -3, -3, 1, -3,
    -- filter=157 channel=70
    -13, 4, 0, 0, 4, -4, 10, -5, 0,
    -- filter=157 channel=71
    7, -3, 0, -5, 0, -7, -8, -2, 3,
    -- filter=157 channel=72
    -9, -10, 5, -9, 1, -3, 6, 8, 0,
    -- filter=157 channel=73
    -17, 3, 1, -2, 9, 5, 9, 1, 0,
    -- filter=157 channel=74
    -7, 15, -10, 8, 5, -5, 6, -8, -5,
    -- filter=157 channel=75
    11, 0, 10, -3, 0, -9, -12, 13, -6,
    -- filter=157 channel=76
    1, 2, -5, 1, 8, -4, -2, 6, -5,
    -- filter=157 channel=77
    7, 0, 2, 5, -1, -1, 6, 0, -5,
    -- filter=157 channel=78
    -6, 2, 0, -6, 3, 0, -5, 0, -1,
    -- filter=157 channel=79
    -3, 6, 9, -24, 0, -9, 8, 1, -11,
    -- filter=157 channel=80
    -15, -3, -2, -23, 7, 0, 9, 18, 0,
    -- filter=157 channel=81
    6, -3, 1, 0, 1, 4, -6, 5, -5,
    -- filter=157 channel=82
    -6, 5, -7, 0, 0, -7, -4, -2, 4,
    -- filter=157 channel=83
    -9, 1, -3, -3, 2, 5, 3, -4, 0,
    -- filter=157 channel=84
    -13, 0, 4, -4, 4, -2, 3, -4, 0,
    -- filter=157 channel=85
    1, 7, -7, 6, -2, -4, 2, -3, -2,
    -- filter=157 channel=86
    5, 3, 2, -1, 0, -7, -1, -5, -7,
    -- filter=157 channel=87
    -1, 13, -3, 5, 1, 5, 5, 0, 0,
    -- filter=157 channel=88
    -8, 1, 0, -3, 10, 4, 2, 5, -2,
    -- filter=157 channel=89
    -9, -8, 1, -21, 13, 3, 16, 9, 0,
    -- filter=157 channel=90
    -2, 0, -6, -1, -3, -3, -1, 2, 10,
    -- filter=157 channel=91
    -10, 1, -2, 4, 13, 0, 15, -1, -11,
    -- filter=157 channel=92
    4, -1, -3, -2, -4, -6, -6, -3, -5,
    -- filter=157 channel=93
    2, 6, 0, -11, 5, 2, 1, -1, 0,
    -- filter=157 channel=94
    5, 2, -4, -1, 5, 2, -1, 4, -4,
    -- filter=157 channel=95
    6, -4, 0, -2, 6, 5, 7, 8, 4,
    -- filter=157 channel=96
    -3, -2, -3, -7, 6, 4, 2, -3, -1,
    -- filter=157 channel=97
    7, -1, 4, -2, -2, 2, -8, 1, 2,
    -- filter=157 channel=98
    -10, 4, 1, -14, -1, 3, 15, 5, -7,
    -- filter=157 channel=99
    -15, 14, -1, -5, 4, 0, 13, 5, 4,
    -- filter=157 channel=100
    5, 4, -1, 5, -4, 6, -4, 0, -4,
    -- filter=157 channel=101
    -6, 5, -1, 5, 3, 6, 14, -2, 0,
    -- filter=157 channel=102
    -6, -6, 1, -1, 0, 4, -3, -5, 2,
    -- filter=157 channel=103
    -3, -6, -7, -12, -11, -5, -7, 2, 4,
    -- filter=157 channel=104
    -11, -2, -7, -7, -4, -3, 15, 0, 5,
    -- filter=157 channel=105
    0, 6, 1, 0, 4, 1, 2, 6, 1,
    -- filter=157 channel=106
    5, -3, 1, -4, -6, -1, 1, 5, -2,
    -- filter=157 channel=107
    -1, 12, -8, 3, 12, 4, 6, -10, -4,
    -- filter=157 channel=108
    5, -4, 6, -2, 0, 2, -6, -3, 4,
    -- filter=157 channel=109
    -16, 5, -3, -11, 4, -1, 10, 4, -8,
    -- filter=157 channel=110
    -5, 6, 4, -2, -6, -2, 0, 7, 0,
    -- filter=157 channel=111
    -4, 1, 0, 5, 1, 3, -3, -3, -4,
    -- filter=157 channel=112
    -1, 0, 2, 5, -1, -4, 8, -3, 2,
    -- filter=157 channel=113
    0, -9, 0, -5, 1, 0, 0, 11, -1,
    -- filter=157 channel=114
    -10, 14, 0, -15, 6, -12, 9, -5, -5,
    -- filter=157 channel=115
    1, 5, -4, -3, -3, -7, -4, 2, 2,
    -- filter=157 channel=116
    -14, 2, -4, -10, 11, -1, 20, 0, 5,
    -- filter=157 channel=117
    3, 7, 5, -4, 4, 6, 4, 8, -4,
    -- filter=157 channel=118
    2, 0, 5, -3, -1, -5, 0, 4, -4,
    -- filter=157 channel=119
    0, 7, -4, 6, -3, 0, 6, 2, -5,
    -- filter=157 channel=120
    -20, 16, -10, 4, 19, -4, 24, -12, -13,
    -- filter=157 channel=121
    1, -5, -6, -9, -3, -7, -1, 8, -6,
    -- filter=157 channel=122
    -5, -3, -9, -9, -9, -8, 7, 9, 2,
    -- filter=157 channel=123
    0, -3, 3, 0, 6, -3, -2, -4, -3,
    -- filter=157 channel=124
    6, -3, -3, -1, 6, -4, -6, 0, -4,
    -- filter=157 channel=125
    -19, -4, -6, -14, 12, -1, 16, 11, 4,
    -- filter=157 channel=126
    -3, 3, 7, -15, 2, 0, -6, 16, -7,
    -- filter=157 channel=127
    -4, -3, -7, -9, 0, -6, -2, 0, 0,
    -- filter=158 channel=0
    -3, 9, 0, -5, 24, -5, -7, 21, -7,
    -- filter=158 channel=1
    -1, 2, -2, -10, 22, 2, -11, 17, -6,
    -- filter=158 channel=2
    -2, 3, 2, 7, -2, -4, 7, 4, -1,
    -- filter=158 channel=3
    5, 2, 1, -5, 4, 6, 5, 0, 0,
    -- filter=158 channel=4
    -3, -5, -4, -5, 0, 9, -8, 7, 9,
    -- filter=158 channel=5
    -8, 0, 3, -9, 18, -7, -3, 6, -8,
    -- filter=158 channel=6
    -8, 1, -5, 7, 0, -2, -2, 3, 0,
    -- filter=158 channel=7
    -2, -4, 0, -4, 0, -1, 3, 6, 4,
    -- filter=158 channel=8
    0, 0, 7, 1, 2, -1, 8, 4, -1,
    -- filter=158 channel=9
    -5, 0, 4, 0, 0, -8, -1, 5, 0,
    -- filter=158 channel=10
    -5, 0, 1, -5, -6, -8, 5, 4, 2,
    -- filter=158 channel=11
    -1, -5, -6, 6, 3, -6, 6, 0, -2,
    -- filter=158 channel=12
    2, 2, 7, 0, 3, 6, 7, 6, 9,
    -- filter=158 channel=13
    0, 0, 8, 2, -3, 0, 0, -6, -2,
    -- filter=158 channel=14
    1, 7, -2, -4, -2, 5, 0, -5, -6,
    -- filter=158 channel=15
    3, 2, -9, -1, 3, -6, 0, 4, -5,
    -- filter=158 channel=16
    3, -2, 0, -2, -4, -1, -5, -1, 2,
    -- filter=158 channel=17
    1, -1, 0, 1, 6, 6, 4, -6, -3,
    -- filter=158 channel=18
    -8, -6, -10, 0, 0, -12, 2, 2, -7,
    -- filter=158 channel=19
    -4, -2, 1, 2, 3, 6, -5, 0, 1,
    -- filter=158 channel=20
    2, 1, 1, 8, -3, -7, 10, 0, 2,
    -- filter=158 channel=21
    3, -5, 15, -3, -1, -4, -1, 0, -1,
    -- filter=158 channel=22
    -3, 2, -5, 6, 9, 0, 4, 2, 0,
    -- filter=158 channel=23
    0, -11, 10, 3, -11, 0, 0, -2, 1,
    -- filter=158 channel=24
    2, -4, -1, 6, -1, -5, 1, 0, 5,
    -- filter=158 channel=25
    -1, 3, 0, 1, 7, -3, -7, -3, 1,
    -- filter=158 channel=26
    -1, -1, 0, -8, 0, -2, -8, 7, 6,
    -- filter=158 channel=27
    -3, -13, -6, 0, -4, 1, 4, 2, -9,
    -- filter=158 channel=28
    4, -3, 4, 0, 4, 0, 3, -2, -3,
    -- filter=158 channel=29
    0, -5, -5, 3, 2, 2, -6, -6, -1,
    -- filter=158 channel=30
    5, 5, 6, -1, 4, -5, -1, 0, 1,
    -- filter=158 channel=31
    2, -13, 16, -4, -17, 6, 7, -10, 3,
    -- filter=158 channel=32
    0, -2, -9, 1, -1, -1, -4, 3, 0,
    -- filter=158 channel=33
    5, 3, -2, 3, -4, -5, -4, 3, -3,
    -- filter=158 channel=34
    5, 0, 0, 7, 2, -1, 7, -3, -1,
    -- filter=158 channel=35
    0, -7, -3, -1, -4, -5, 0, -1, 2,
    -- filter=158 channel=36
    0, 3, -2, 6, -5, 0, 5, -11, 7,
    -- filter=158 channel=37
    -5, 1, -1, -1, 17, 6, -9, 17, 0,
    -- filter=158 channel=38
    0, 0, 5, 4, -4, -9, -1, -5, 4,
    -- filter=158 channel=39
    4, 3, -8, -4, -9, 0, 0, 3, -6,
    -- filter=158 channel=40
    11, 0, 3, 5, -2, -3, 7, 3, -4,
    -- filter=158 channel=41
    0, 4, -3, -4, 0, 7, 4, 6, -1,
    -- filter=158 channel=42
    -8, 1, 1, -10, 5, -1, -1, 4, -3,
    -- filter=158 channel=43
    5, 1, 0, 0, 5, -4, 0, -3, 6,
    -- filter=158 channel=44
    -7, -2, 7, 3, 9, 2, 0, 0, -3,
    -- filter=158 channel=45
    3, 5, 2, 3, 8, -3, -1, 8, -3,
    -- filter=158 channel=46
    5, -5, 5, 7, 0, -8, -5, 5, -5,
    -- filter=158 channel=47
    -6, 6, 7, -8, -5, 7, -8, 4, -6,
    -- filter=158 channel=48
    3, -3, 5, -8, -4, -1, 1, -2, 4,
    -- filter=158 channel=49
    -6, -3, -3, 5, -4, 4, 2, -2, 0,
    -- filter=158 channel=50
    -1, -2, -3, 4, -6, 4, -6, 0, 2,
    -- filter=158 channel=51
    0, 6, 0, -6, 3, 7, 0, 2, -7,
    -- filter=158 channel=52
    0, -8, -4, 9, -7, 6, 0, 0, 0,
    -- filter=158 channel=53
    7, -5, -2, 7, -2, 5, 0, 2, -2,
    -- filter=158 channel=54
    -4, 0, 1, 7, 7, 5, 7, -7, 0,
    -- filter=158 channel=55
    -1, -12, 3, -1, -1, -3, 0, -2, -5,
    -- filter=158 channel=56
    -4, -5, 3, 8, 2, -2, 3, -1, 0,
    -- filter=158 channel=57
    -4, 0, -5, 4, -6, 3, -5, 0, -6,
    -- filter=158 channel=58
    -9, 5, -1, -8, 7, -4, 1, 10, 7,
    -- filter=158 channel=59
    2, 3, -3, -4, 4, 3, -8, -3, 0,
    -- filter=158 channel=60
    -1, 6, 2, 6, 7, -2, -5, 3, -5,
    -- filter=158 channel=61
    2, -2, 5, -1, -2, -4, -5, 2, 4,
    -- filter=158 channel=62
    3, -2, -6, -2, 3, 7, -5, -6, 6,
    -- filter=158 channel=63
    -10, 6, -2, -9, 3, 0, -6, 2, 0,
    -- filter=158 channel=64
    -3, 2, 3, -6, -7, -6, -1, 0, 0,
    -- filter=158 channel=65
    -2, 0, 3, -6, 0, 3, 5, 1, -7,
    -- filter=158 channel=66
    -1, 2, -3, -4, -2, 5, -1, -1, 7,
    -- filter=158 channel=67
    2, 5, 0, 6, -1, 1, 6, 0, -5,
    -- filter=158 channel=68
    0, -8, 0, -2, 2, 0, 4, -7, -4,
    -- filter=158 channel=69
    -1, 4, 4, 0, -6, 2, 2, 0, -1,
    -- filter=158 channel=70
    -2, 1, 2, -4, 4, -2, 8, 0, 4,
    -- filter=158 channel=71
    -5, -3, -2, -1, -1, -3, 4, 7, -5,
    -- filter=158 channel=72
    4, 1, 2, -7, -4, 1, 1, -9, -5,
    -- filter=158 channel=73
    0, -4, 2, 4, -9, 3, 0, -5, 4,
    -- filter=158 channel=74
    1, -10, 0, 6, 0, -4, 3, -1, 4,
    -- filter=158 channel=75
    -3, 5, 4, -5, 15, 6, -1, 19, -4,
    -- filter=158 channel=76
    1, -4, 0, -3, 1, -2, 1, -2, 1,
    -- filter=158 channel=77
    -7, 5, 6, 7, -3, 0, 0, 5, 4,
    -- filter=158 channel=78
    2, -6, -4, 2, -7, 5, -1, 0, -7,
    -- filter=158 channel=79
    7, -2, -3, -2, -1, -3, 3, 6, 4,
    -- filter=158 channel=80
    5, -4, 13, -10, 0, 0, -5, -8, 1,
    -- filter=158 channel=81
    1, -5, -3, 7, -5, 4, 6, 4, -2,
    -- filter=158 channel=82
    1, 0, 2, 6, 1, 1, 7, 8, -6,
    -- filter=158 channel=83
    6, 3, -2, -6, -4, -1, -7, -2, 0,
    -- filter=158 channel=84
    4, 2, -8, 6, 4, 7, -1, 0, 3,
    -- filter=158 channel=85
    0, -3, -6, -3, 5, 1, 3, -2, -2,
    -- filter=158 channel=86
    -4, -4, 9, 1, 5, -3, -4, 0, 3,
    -- filter=158 channel=87
    6, -4, 4, 8, -3, -3, 8, -3, 1,
    -- filter=158 channel=88
    7, 3, -2, 1, -7, -2, -2, -10, -2,
    -- filter=158 channel=89
    0, 1, 9, -2, -10, -4, -3, -5, 5,
    -- filter=158 channel=90
    7, 0, 13, 7, -1, 2, 8, -10, 8,
    -- filter=158 channel=91
    0, 0, -3, 6, -9, -6, 0, -6, 5,
    -- filter=158 channel=92
    6, 6, 6, 1, -7, 2, 0, 4, 2,
    -- filter=158 channel=93
    3, 3, 9, -17, 12, 9, 0, 10, 7,
    -- filter=158 channel=94
    -2, -6, -3, -1, 4, -7, -5, 1, 0,
    -- filter=158 channel=95
    -5, -2, -1, 3, 2, -3, -7, -4, 3,
    -- filter=158 channel=96
    -3, -5, 0, -2, -6, 6, -2, 0, 5,
    -- filter=158 channel=97
    2, 0, 3, -8, -2, 6, 4, 3, 0,
    -- filter=158 channel=98
    4, -5, 10, -4, -5, -2, -2, 1, 0,
    -- filter=158 channel=99
    5, -14, 1, 1, -8, 0, 9, -10, 4,
    -- filter=158 channel=100
    -3, 2, -7, -2, 2, 1, -1, 8, 2,
    -- filter=158 channel=101
    -2, -3, 4, 2, 6, -1, -2, -6, -3,
    -- filter=158 channel=102
    -4, 3, 0, -4, -1, -1, -4, 1, 4,
    -- filter=158 channel=103
    -1, -3, 6, -11, -4, -7, -7, 7, -5,
    -- filter=158 channel=104
    3, -3, 3, -5, -11, -2, -1, -9, -1,
    -- filter=158 channel=105
    4, -3, 4, 1, 0, -5, 7, -6, 0,
    -- filter=158 channel=106
    -5, -2, -5, -6, -3, -4, 3, 0, -1,
    -- filter=158 channel=107
    0, -5, -1, 7, -1, 1, 9, 5, -5,
    -- filter=158 channel=108
    2, -3, 3, 0, 8, 0, 0, 9, 4,
    -- filter=158 channel=109
    -3, -1, 1, 4, -1, -4, 7, -7, 2,
    -- filter=158 channel=110
    -4, -7, 9, 3, 0, 5, 6, -8, -5,
    -- filter=158 channel=111
    -1, 2, -3, 2, 7, -3, 0, 5, 4,
    -- filter=158 channel=112
    -2, 0, -4, -6, -10, 2, -2, -3, -7,
    -- filter=158 channel=113
    5, -4, 11, 5, -4, 0, -2, 0, 1,
    -- filter=158 channel=114
    -10, 4, -3, 2, 10, -10, -1, 0, -3,
    -- filter=158 channel=115
    1, -5, -4, 6, -6, 3, 2, -5, -5,
    -- filter=158 channel=116
    0, 2, -6, -2, -9, -3, -8, -2, -4,
    -- filter=158 channel=117
    8, -6, 0, 5, 1, -2, 7, 0, 6,
    -- filter=158 channel=118
    2, 0, -7, 0, -2, -6, -5, -1, 2,
    -- filter=158 channel=119
    7, 1, -6, 6, 8, 5, 3, 5, 3,
    -- filter=158 channel=120
    6, -8, 1, 5, -3, -4, 8, -8, -5,
    -- filter=158 channel=121
    4, -7, 2, -7, -1, 4, 0, -2, -2,
    -- filter=158 channel=122
    -2, -1, 19, -2, 0, 1, 0, -7, 2,
    -- filter=158 channel=123
    1, 6, 0, 3, -3, 7, -4, -1, -3,
    -- filter=158 channel=124
    6, 3, -1, -1, -9, 0, 2, 1, 2,
    -- filter=158 channel=125
    7, -8, -3, -3, -13, -5, 7, -4, -2,
    -- filter=158 channel=126
    5, 5, 4, -6, 3, 5, 2, 9, -5,
    -- filter=158 channel=127
    -3, 0, -4, 2, 5, -3, -4, 7, 1,
    -- filter=159 channel=0
    2, -3, -5, -4, -6, -5, -1, -12, -12,
    -- filter=159 channel=1
    2, -1, -11, 2, -7, -14, 0, -5, -3,
    -- filter=159 channel=2
    0, 0, -5, 3, -1, -7, 0, -1, 5,
    -- filter=159 channel=3
    2, -1, 6, -11, -5, -1, -1, -7, 0,
    -- filter=159 channel=4
    3, 5, -3, -7, -6, -5, 2, -8, -1,
    -- filter=159 channel=5
    -1, 0, -7, -6, -1, -2, -3, -1, 3,
    -- filter=159 channel=6
    -5, 7, -6, -6, -8, 3, 1, -4, 0,
    -- filter=159 channel=7
    -6, -3, 2, -3, 2, 4, 6, 2, -2,
    -- filter=159 channel=8
    -7, -9, 4, -2, -1, -7, -6, -2, 2,
    -- filter=159 channel=9
    -2, 7, 1, 4, -2, -2, -1, -4, -1,
    -- filter=159 channel=10
    0, 10, -1, 1, 9, -3, -3, 4, -1,
    -- filter=159 channel=11
    0, 9, 7, 9, -1, 7, 0, 6, -9,
    -- filter=159 channel=12
    -6, 4, 0, 0, 0, 4, -8, -7, -5,
    -- filter=159 channel=13
    4, 10, 8, -3, 0, 4, -9, -1, -9,
    -- filter=159 channel=14
    -3, -1, 1, 3, 2, -4, -4, 2, -5,
    -- filter=159 channel=15
    11, 14, 1, -4, -2, 0, -2, -2, -4,
    -- filter=159 channel=16
    -3, -5, 5, -3, 1, -2, -4, 3, -1,
    -- filter=159 channel=17
    -2, 4, -4, 6, -6, 0, 2, -5, 0,
    -- filter=159 channel=18
    13, 9, 2, -4, -8, 1, -3, -5, -9,
    -- filter=159 channel=19
    2, -6, -6, 2, 1, 0, -5, -1, 3,
    -- filter=159 channel=20
    11, 6, 10, 5, 5, 0, 1, 3, 0,
    -- filter=159 channel=21
    6, -4, -3, -3, 4, 2, 1, 4, 8,
    -- filter=159 channel=22
    6, -5, 4, 5, -10, 1, -2, 2, -11,
    -- filter=159 channel=23
    8, 21, 11, 8, -3, -2, 0, -3, -17,
    -- filter=159 channel=24
    -2, 5, 5, -4, 4, 1, 4, -1, 5,
    -- filter=159 channel=25
    2, 0, 3, -8, 2, -1, -5, 1, 0,
    -- filter=159 channel=26
    -2, -8, 1, 7, 5, 0, 5, 3, 4,
    -- filter=159 channel=27
    5, 10, 0, -4, -3, -8, -9, -6, -16,
    -- filter=159 channel=28
    -5, -5, 1, -7, 3, 6, 0, 6, -3,
    -- filter=159 channel=29
    5, 13, 10, -2, 9, -2, -4, 5, -11,
    -- filter=159 channel=30
    3, -5, -1, 4, 0, 1, 3, -3, -10,
    -- filter=159 channel=31
    11, 15, 6, 0, 14, 0, 5, 14, -8,
    -- filter=159 channel=32
    -2, 13, 4, -9, -7, 0, -8, -12, -5,
    -- filter=159 channel=33
    9, 1, 2, -4, -3, 4, -9, 3, -13,
    -- filter=159 channel=34
    3, -8, -7, -8, -12, -5, -4, -12, -1,
    -- filter=159 channel=35
    -3, -3, -1, 6, 1, 3, 0, 1, -2,
    -- filter=159 channel=36
    1, 8, 2, 6, 2, -5, 8, 0, 7,
    -- filter=159 channel=37
    4, -11, -1, -5, -11, -8, 4, -9, -5,
    -- filter=159 channel=38
    9, 9, 4, -4, -1, 6, -7, 4, 2,
    -- filter=159 channel=39
    -4, 11, 1, 8, 5, -3, 0, -3, -6,
    -- filter=159 channel=40
    -2, 0, 10, 0, 11, 9, 6, -4, -4,
    -- filter=159 channel=41
    -7, -7, 3, -7, -5, -1, -11, -9, 8,
    -- filter=159 channel=42
    8, -6, 0, -4, -7, -2, 5, -5, 0,
    -- filter=159 channel=43
    1, 2, 1, -3, 0, 4, -2, 2, -2,
    -- filter=159 channel=44
    -5, -7, -2, -5, -10, -9, -3, -8, -3,
    -- filter=159 channel=45
    8, 7, 6, -1, 0, 0, 3, 8, -4,
    -- filter=159 channel=46
    -7, -4, -8, -7, -6, 4, -5, 1, -5,
    -- filter=159 channel=47
    6, -7, 5, -8, -7, 2, -3, -2, -4,
    -- filter=159 channel=48
    -6, 1, -8, -4, -6, -12, 2, -3, -12,
    -- filter=159 channel=49
    4, 0, -4, 0, 2, -10, -5, -1, -1,
    -- filter=159 channel=50
    5, 10, 8, 1, 4, -5, -2, 1, -10,
    -- filter=159 channel=51
    5, 0, -5, -5, 3, 1, 1, -3, -3,
    -- filter=159 channel=52
    -6, 0, -5, 0, -9, 0, -5, 4, 0,
    -- filter=159 channel=53
    1, 3, 8, 8, -3, 2, -6, 4, 1,
    -- filter=159 channel=54
    0, 0, -2, 0, -4, 0, 5, 6, 2,
    -- filter=159 channel=55
    2, 17, 12, 7, 4, 2, 3, 5, -13,
    -- filter=159 channel=56
    -3, -2, 2, 4, -4, -5, -8, -3, 4,
    -- filter=159 channel=57
    5, 3, 0, 1, 0, -3, 1, 0, -2,
    -- filter=159 channel=58
    2, 4, -8, 0, 0, 1, -5, -1, -2,
    -- filter=159 channel=59
    2, 7, 0, 0, 9, 1, 0, -5, -8,
    -- filter=159 channel=60
    -7, 0, -6, -6, 2, 2, 2, 3, 0,
    -- filter=159 channel=61
    -6, 6, -1, 0, 1, 1, 0, 1, -1,
    -- filter=159 channel=62
    1, 1, 0, -3, 7, -4, 2, -5, -4,
    -- filter=159 channel=63
    5, 3, -5, -2, 5, -7, 8, -2, -1,
    -- filter=159 channel=64
    -3, -3, 0, -4, 7, 0, 0, 8, 5,
    -- filter=159 channel=65
    -2, -7, 1, -6, -4, -2, 7, -3, 3,
    -- filter=159 channel=66
    1, 2, -3, -1, 6, 6, -5, -2, -1,
    -- filter=159 channel=67
    -6, -3, 1, 6, -3, -5, 5, 4, 4,
    -- filter=159 channel=68
    -3, 7, 4, -2, -5, 0, 9, 2, 5,
    -- filter=159 channel=69
    4, 3, 6, 0, 5, -1, -3, 3, 7,
    -- filter=159 channel=70
    10, 11, -3, 4, -10, 0, -7, -6, -17,
    -- filter=159 channel=71
    11, 11, 2, -6, 3, 6, -3, 8, 1,
    -- filter=159 channel=72
    3, 2, 2, 10, 3, 2, 6, 3, -3,
    -- filter=159 channel=73
    -5, -3, 1, -3, -2, -5, 0, -9, -6,
    -- filter=159 channel=74
    6, -4, -7, 4, 1, -5, 1, -6, -9,
    -- filter=159 channel=75
    -2, -5, -3, -3, -13, -6, 0, -6, -3,
    -- filter=159 channel=76
    0, 5, 15, 5, 1, 12, 3, 8, -2,
    -- filter=159 channel=77
    -1, -1, -5, -5, -1, -5, -2, 7, -4,
    -- filter=159 channel=78
    -2, 0, 5, 6, 6, -1, 4, 4, 0,
    -- filter=159 channel=79
    0, 11, 12, 0, -8, 2, -3, -12, -7,
    -- filter=159 channel=80
    5, 1, 8, 2, 9, 1, -2, 10, 0,
    -- filter=159 channel=81
    3, -1, -1, 1, -3, -5, 0, -6, 6,
    -- filter=159 channel=82
    2, -2, -4, 4, -5, -2, -2, 4, 2,
    -- filter=159 channel=83
    -3, -1, 0, 0, 7, -1, 6, 7, 0,
    -- filter=159 channel=84
    -4, -2, -1, -3, -6, -6, 0, 1, 0,
    -- filter=159 channel=85
    3, -1, 1, -3, -7, -4, -6, 5, -7,
    -- filter=159 channel=86
    1, -3, -7, -10, -2, -6, -1, -10, -4,
    -- filter=159 channel=87
    1, 6, 9, -2, 4, 0, -4, -6, -8,
    -- filter=159 channel=88
    -4, 7, -4, 6, 7, 0, -1, 1, -3,
    -- filter=159 channel=89
    3, 16, 11, -1, 9, -1, 2, -2, 1,
    -- filter=159 channel=90
    -5, 0, 7, 5, 0, 7, 0, -1, 7,
    -- filter=159 channel=91
    6, 0, 2, 0, -6, -10, -4, -1, -13,
    -- filter=159 channel=92
    3, 6, 5, 5, 5, -1, -6, -7, -10,
    -- filter=159 channel=93
    -2, -6, -4, -10, -13, -4, 1, -5, -7,
    -- filter=159 channel=94
    0, 2, 2, 5, 3, 1, -2, -6, 3,
    -- filter=159 channel=95
    2, -7, -4, 4, -3, 4, -1, 3, -2,
    -- filter=159 channel=96
    -6, 4, -4, -5, 3, -1, 3, 4, 0,
    -- filter=159 channel=97
    3, 12, -1, 2, -3, -4, 2, 7, -1,
    -- filter=159 channel=98
    6, 8, -3, -9, 3, -7, -1, -3, -13,
    -- filter=159 channel=99
    5, 13, 0, 1, 6, 0, -4, -4, -15,
    -- filter=159 channel=100
    1, 0, -7, 0, 0, 3, 4, -6, 1,
    -- filter=159 channel=101
    -6, -5, 4, 3, 0, 0, 0, -2, 3,
    -- filter=159 channel=102
    -6, 5, -5, -3, 1, -5, -6, 6, -4,
    -- filter=159 channel=103
    4, 3, 8, 3, -1, 3, -2, 1, -6,
    -- filter=159 channel=104
    8, 7, -2, 1, 5, 0, 0, 6, 1,
    -- filter=159 channel=105
    4, 1, 3, 3, 1, 9, 5, 6, 2,
    -- filter=159 channel=106
    0, -1, 3, 0, 6, 9, 1, -5, 2,
    -- filter=159 channel=107
    9, 5, -5, 0, 0, -6, 5, 2, -12,
    -- filter=159 channel=108
    -7, -7, 0, 3, -6, 0, -7, -4, 8,
    -- filter=159 channel=109
    2, -2, 8, 1, -9, -1, -9, -12, -17,
    -- filter=159 channel=110
    7, 5, 2, 3, 6, 3, 0, 3, 0,
    -- filter=159 channel=111
    -4, 2, -2, -4, 1, -2, 2, -3, 5,
    -- filter=159 channel=112
    0, 4, -7, -1, -6, -4, -4, -6, -11,
    -- filter=159 channel=113
    10, 10, 10, -3, 3, 8, 5, -6, 2,
    -- filter=159 channel=114
    2, -5, -5, -7, -5, -14, 4, -17, -22,
    -- filter=159 channel=115
    -6, -6, -4, 4, 3, -2, 1, 0, -7,
    -- filter=159 channel=116
    8, 8, 5, -2, -1, -12, 0, -8, -11,
    -- filter=159 channel=117
    3, 7, -1, -4, 3, 3, -4, 5, 0,
    -- filter=159 channel=118
    -3, 3, 1, -2, 4, -2, -3, -4, 7,
    -- filter=159 channel=119
    -7, -4, -1, -6, -9, -11, -2, -4, -2,
    -- filter=159 channel=120
    -2, 15, -1, 8, 3, -10, -5, 0, -15,
    -- filter=159 channel=121
    4, -6, 7, -5, 1, -6, 4, 5, -5,
    -- filter=159 channel=122
    -1, -10, -3, 2, -7, -1, 3, 5, 4,
    -- filter=159 channel=123
    -2, 0, 1, 4, 1, -1, -8, -4, 2,
    -- filter=159 channel=124
    -4, 1, 5, 0, -3, 0, 6, -5, -5,
    -- filter=159 channel=125
    -3, 7, -1, -5, 9, -10, -7, 8, 1,
    -- filter=159 channel=126
    0, -2, 12, -7, 0, 4, 0, 1, -5,
    -- filter=159 channel=127
    3, -7, -5, 4, -1, 7, -5, 4, 6,
    -- filter=160 channel=0
    3, -7, 1, -1, 0, 0, 0, 2, -5,
    -- filter=160 channel=1
    9, 5, -8, 4, -4, 1, -1, -9, -9,
    -- filter=160 channel=2
    -3, 2, -1, 1, -1, -2, -2, -2, 1,
    -- filter=160 channel=3
    1, 0, -4, -10, 0, 4, -9, -2, -1,
    -- filter=160 channel=4
    -8, -6, 2, -6, -4, -6, -11, -2, 0,
    -- filter=160 channel=5
    -1, 8, 8, -5, 15, 2, -7, 11, 3,
    -- filter=160 channel=6
    -6, 1, -2, 5, 1, 3, 0, -8, -5,
    -- filter=160 channel=7
    -1, -1, -4, 3, -3, -5, 0, 0, -1,
    -- filter=160 channel=8
    -2, 0, 2, -1, 4, -6, -7, 5, -1,
    -- filter=160 channel=9
    5, -6, -1, 6, -2, -1, 0, -7, 3,
    -- filter=160 channel=10
    0, -9, 0, 10, 1, 5, 11, -6, 8,
    -- filter=160 channel=11
    3, 3, 11, -3, 3, 9, -9, 6, 6,
    -- filter=160 channel=12
    11, -4, 5, 7, -4, -3, -2, 0, 1,
    -- filter=160 channel=13
    11, -3, -1, 9, -10, -2, 10, -4, -1,
    -- filter=160 channel=14
    -5, 0, 0, -4, -7, 0, -3, -6, 0,
    -- filter=160 channel=15
    -1, -11, 2, 3, -7, 6, 1, -11, 8,
    -- filter=160 channel=16
    -5, -4, -10, 5, 0, -3, -7, 8, -5,
    -- filter=160 channel=17
    -1, 4, -7, 2, 0, -7, 0, -6, -4,
    -- filter=160 channel=18
    16, -16, -1, 18, -15, 8, 10, -13, 2,
    -- filter=160 channel=19
    3, -1, 0, -4, 4, 2, -1, -5, -5,
    -- filter=160 channel=20
    -6, -8, 2, -10, -3, 6, -4, 2, 1,
    -- filter=160 channel=21
    2, 7, 1, -3, 10, -5, 4, 7, -9,
    -- filter=160 channel=22
    -4, -9, 0, 0, -7, 5, -2, -7, -5,
    -- filter=160 channel=23
    -3, -7, 0, 0, -11, 2, 1, -6, 13,
    -- filter=160 channel=24
    3, -4, -5, 0, 6, 4, 0, -2, 0,
    -- filter=160 channel=25
    18, -8, -6, 16, -7, -2, 0, -6, 1,
    -- filter=160 channel=26
    -10, -1, -6, -2, 11, -5, -9, 5, 0,
    -- filter=160 channel=27
    10, -14, 3, 8, -11, 11, 4, -11, 2,
    -- filter=160 channel=28
    5, -1, -2, -3, -1, -4, 2, 0, 4,
    -- filter=160 channel=29
    -5, -5, 14, -8, 3, 9, -2, -2, 10,
    -- filter=160 channel=30
    0, -5, -1, -4, 1, -1, -7, -2, 1,
    -- filter=160 channel=31
    -7, 0, 6, -5, 0, 6, 5, 3, 1,
    -- filter=160 channel=32
    5, -11, 9, 13, -12, 4, 3, -12, 9,
    -- filter=160 channel=33
    -2, -2, -1, 4, -3, 9, 10, -12, -1,
    -- filter=160 channel=34
    -3, 10, 6, 4, 13, -4, 3, -2, 0,
    -- filter=160 channel=35
    4, 4, 4, 6, 5, -6, -2, 5, 2,
    -- filter=160 channel=36
    -11, 3, 5, 0, -6, -4, -8, -6, 1,
    -- filter=160 channel=37
    -4, 5, -3, -4, 13, 1, -7, -8, -3,
    -- filter=160 channel=38
    4, 1, 7, 1, -4, 7, 0, -3, -5,
    -- filter=160 channel=39
    1, 2, 0, 0, 3, 0, -2, 6, -3,
    -- filter=160 channel=40
    -5, -4, 0, -1, 0, -3, -5, 0, -1,
    -- filter=160 channel=41
    14, -8, -14, 15, -11, -13, 19, -9, -5,
    -- filter=160 channel=42
    -1, 0, 0, -8, 6, 1, -2, -2, 3,
    -- filter=160 channel=43
    -5, -10, 0, -2, -9, -3, -9, 1, -6,
    -- filter=160 channel=44
    -6, 3, 7, 3, 12, 8, -2, 1, 2,
    -- filter=160 channel=45
    0, -3, 7, -6, -5, 6, -2, 4, 4,
    -- filter=160 channel=46
    2, 4, -6, -1, -5, 2, 5, -2, 0,
    -- filter=160 channel=47
    -4, 0, 1, -3, 9, -5, -6, 10, -8,
    -- filter=160 channel=48
    -4, -2, -6, -2, 5, 7, 4, -8, 1,
    -- filter=160 channel=49
    -6, 0, 1, 4, -5, 6, 1, 0, 0,
    -- filter=160 channel=50
    0, -2, 1, 8, -2, -4, -4, -8, 0,
    -- filter=160 channel=51
    -4, 5, 5, -4, 5, 3, 4, 4, 6,
    -- filter=160 channel=52
    5, -6, 8, -3, 1, -1, -2, -7, 6,
    -- filter=160 channel=53
    0, -5, 9, -3, 4, 3, 0, -1, 10,
    -- filter=160 channel=54
    2, -6, -2, 2, 6, 2, 6, -2, -6,
    -- filter=160 channel=55
    4, -8, 6, 5, -14, 2, 10, -3, 10,
    -- filter=160 channel=56
    -7, 10, 0, -5, 6, 5, -4, 0, -8,
    -- filter=160 channel=57
    2, 1, 4, 8, 1, -4, 3, -1, -6,
    -- filter=160 channel=58
    -9, 0, -5, -3, 6, 2, 0, 3, 1,
    -- filter=160 channel=59
    2, 0, 0, 5, -1, 7, 3, -9, 0,
    -- filter=160 channel=60
    0, 3, 5, 3, -3, 1, -1, 0, -1,
    -- filter=160 channel=61
    4, -3, -5, -7, 0, 0, 1, 5, -5,
    -- filter=160 channel=62
    2, 6, -3, -4, 1, 3, 5, 0, 2,
    -- filter=160 channel=63
    -1, 3, -1, -6, 2, -4, 2, 2, -4,
    -- filter=160 channel=64
    -10, 4, 2, -3, 4, -3, 0, 6, 0,
    -- filter=160 channel=65
    5, -4, 2, 0, 6, 4, 4, 0, 0,
    -- filter=160 channel=66
    5, -9, -2, 8, -1, -6, 5, -5, 0,
    -- filter=160 channel=67
    0, -4, 4, 2, 6, 3, 6, 6, -4,
    -- filter=160 channel=68
    4, -7, -2, 5, 0, 4, 5, 3, -8,
    -- filter=160 channel=69
    3, 5, 1, -3, 0, 3, 4, 5, 6,
    -- filter=160 channel=70
    0, -12, 1, 0, 0, 6, -1, -3, -5,
    -- filter=160 channel=71
    -3, -8, -8, 2, -7, 3, 5, -8, -3,
    -- filter=160 channel=72
    4, -9, -5, 10, -8, 2, 7, -1, 2,
    -- filter=160 channel=73
    11, -5, 11, 9, -11, -2, -2, -1, -2,
    -- filter=160 channel=74
    -1, -7, 1, 1, 3, -7, -7, -6, -5,
    -- filter=160 channel=75
    -6, -1, 0, 4, 12, 11, -2, 0, 1,
    -- filter=160 channel=76
    0, -7, 6, 0, -3, 3, 4, -6, 9,
    -- filter=160 channel=77
    2, -4, -1, -6, 1, -2, -6, 4, -5,
    -- filter=160 channel=78
    -9, 3, 0, -6, 9, -1, -9, 9, -6,
    -- filter=160 channel=79
    12, -16, -4, 17, -17, 6, 2, -9, -4,
    -- filter=160 channel=80
    7, -8, 3, 13, -3, 6, 2, -4, 1,
    -- filter=160 channel=81
    0, -1, 6, 3, -3, 0, 6, 2, 5,
    -- filter=160 channel=82
    -3, 6, 3, -7, 7, -2, -7, 7, 2,
    -- filter=160 channel=83
    1, -4, 3, 5, -3, -7, -4, 5, -1,
    -- filter=160 channel=84
    5, -1, 4, 10, -6, 4, 0, -8, -4,
    -- filter=160 channel=85
    0, -5, 0, -4, 5, 1, -5, 0, 3,
    -- filter=160 channel=86
    6, 2, -3, 8, 7, 5, 1, 3, 2,
    -- filter=160 channel=87
    -7, -2, 3, 0, 1, -4, -5, 0, 6,
    -- filter=160 channel=88
    -7, -2, 4, -5, -4, -7, -6, 7, 2,
    -- filter=160 channel=89
    14, -16, 3, 8, -8, 10, 4, -2, -5,
    -- filter=160 channel=90
    -16, -6, -6, -10, 7, -3, -8, -1, -8,
    -- filter=160 channel=91
    -2, -9, 6, 6, -10, 8, -1, -15, -1,
    -- filter=160 channel=92
    0, 3, 1, -5, 4, 4, 5, 8, 6,
    -- filter=160 channel=93
    -3, 2, 2, -9, 5, 3, 3, 0, 1,
    -- filter=160 channel=94
    -6, -6, 0, -6, 3, 0, 7, 1, 0,
    -- filter=160 channel=95
    4, 0, 2, 4, -6, -3, 5, -1, 0,
    -- filter=160 channel=96
    7, -8, -1, -5, -4, 0, 6, -5, -2,
    -- filter=160 channel=97
    1, 2, -2, -1, 1, 2, -2, 1, 3,
    -- filter=160 channel=98
    14, -10, -2, 14, 0, -1, 7, -5, 2,
    -- filter=160 channel=99
    -7, 2, 12, 5, 6, 6, -1, 6, 6,
    -- filter=160 channel=100
    5, 1, -1, -2, -1, -5, 3, -1, -5,
    -- filter=160 channel=101
    -8, -9, 1, -4, -3, -2, -8, -1, -1,
    -- filter=160 channel=102
    -5, 3, 6, 7, 3, -3, 0, -3, -4,
    -- filter=160 channel=103
    1, 5, 0, -2, 13, 0, 1, 4, 0,
    -- filter=160 channel=104
    -4, 5, -7, 6, 1, -1, 0, 3, 3,
    -- filter=160 channel=105
    -6, 2, 0, 3, -3, -3, -3, 4, -1,
    -- filter=160 channel=106
    6, 0, 1, -1, 0, 4, -5, 7, -1,
    -- filter=160 channel=107
    0, 2, 6, -3, -12, -3, -6, -8, -3,
    -- filter=160 channel=108
    -3, -6, 0, 0, 5, -8, 0, -1, 5,
    -- filter=160 channel=109
    16, -14, 6, 9, -3, 3, -2, -4, 2,
    -- filter=160 channel=110
    -6, -7, -1, 0, 0, 8, -7, 2, 2,
    -- filter=160 channel=111
    8, 5, -7, -4, -5, -6, 6, 6, -4,
    -- filter=160 channel=112
    -3, -6, 0, 6, 4, 3, 4, -8, 6,
    -- filter=160 channel=113
    1, -9, -2, 4, -4, -3, 2, -2, -1,
    -- filter=160 channel=114
    11, -13, 2, 12, -2, 4, -4, -8, -8,
    -- filter=160 channel=115
    3, 6, 4, 1, 6, 3, 0, -2, 0,
    -- filter=160 channel=116
    1, -6, 8, 4, -9, 0, 7, -11, -4,
    -- filter=160 channel=117
    5, 0, 1, 1, -2, 6, -5, -5, -7,
    -- filter=160 channel=118
    6, 0, 0, 2, 6, -6, -5, 0, -4,
    -- filter=160 channel=119
    -2, 4, -4, 0, 1, -7, 0, 8, 0,
    -- filter=160 channel=120
    -4, -12, 14, -5, 0, 3, -6, -4, 8,
    -- filter=160 channel=121
    5, 0, -10, -1, 0, 5, 10, -7, 0,
    -- filter=160 channel=122
    -5, 14, -10, -10, 9, 1, -5, 4, -4,
    -- filter=160 channel=123
    5, -4, -1, 0, 4, 2, -7, 6, 1,
    -- filter=160 channel=124
    -3, -2, 1, -1, 3, -2, -4, 2, 5,
    -- filter=160 channel=125
    5, -10, -4, -2, 2, 10, 5, -9, -5,
    -- filter=160 channel=126
    14, -11, 0, 13, 0, 0, 6, 0, -7,
    -- filter=160 channel=127
    -1, -3, -1, 0, 5, 1, 2, -3, 4,
    -- filter=161 channel=0
    12, 9, 2, 11, 3, -14, -1, 2, -6,
    -- filter=161 channel=1
    13, 0, 5, 11, 5, -14, 4, -6, -14,
    -- filter=161 channel=2
    6, 6, -5, 0, 2, -3, -8, 4, 5,
    -- filter=161 channel=3
    -9, -4, 0, -7, 3, -5, 2, 7, 1,
    -- filter=161 channel=4
    -4, -9, -2, 4, 5, 3, 0, 5, 10,
    -- filter=161 channel=5
    0, -1, 0, 11, 0, -4, 0, 5, -11,
    -- filter=161 channel=6
    3, 3, -7, 0, -3, 7, 3, 0, -1,
    -- filter=161 channel=7
    0, 6, 0, 2, -4, 5, 0, 4, 0,
    -- filter=161 channel=8
    -3, -6, -9, -7, -4, -3, -7, 7, -5,
    -- filter=161 channel=9
    -5, 7, 0, 1, -5, 5, 0, 3, 4,
    -- filter=161 channel=10
    -7, -2, 1, 1, -5, -6, -2, -6, -3,
    -- filter=161 channel=11
    1, -4, -1, -1, -3, 8, -7, -2, 9,
    -- filter=161 channel=12
    2, 4, 4, 3, -2, 2, 3, 1, -6,
    -- filter=161 channel=13
    -9, 0, 2, -4, 0, -3, 0, 1, 0,
    -- filter=161 channel=14
    -1, 0, 4, 6, 1, -5, -6, -4, 4,
    -- filter=161 channel=15
    -1, -1, 2, -7, -8, -4, -5, 7, 13,
    -- filter=161 channel=16
    1, -7, -3, 0, -7, 1, -1, 0, -3,
    -- filter=161 channel=17
    -6, -6, 6, -7, -3, -3, 0, 5, -4,
    -- filter=161 channel=18
    1, 6, -2, -2, 5, 1, -8, 4, 12,
    -- filter=161 channel=19
    -2, -2, -5, -7, -6, 6, -5, 0, 0,
    -- filter=161 channel=20
    0, -6, 0, -14, -2, 7, -2, 1, 20,
    -- filter=161 channel=21
    0, -1, -6, -5, -3, -4, 2, 0, -3,
    -- filter=161 channel=22
    6, 1, 0, 2, 5, -10, 4, -5, -3,
    -- filter=161 channel=23
    -1, 1, -12, -7, -6, -7, 5, 13, 2,
    -- filter=161 channel=24
    0, -3, -5, 4, 5, -6, 7, 4, 5,
    -- filter=161 channel=25
    7, -2, -1, -3, 3, -13, 0, -3, 7,
    -- filter=161 channel=26
    5, -7, 2, -5, 5, 6, -3, -3, 2,
    -- filter=161 channel=27
    0, 0, -8, 3, 0, -17, 2, 10, 8,
    -- filter=161 channel=28
    3, -3, 4, -6, 7, 4, -6, -5, 2,
    -- filter=161 channel=29
    -3, 4, 5, -3, 0, 14, -1, 2, 22,
    -- filter=161 channel=30
    3, 6, -6, 8, 8, -4, 2, 5, 3,
    -- filter=161 channel=31
    -1, 0, 0, -7, 3, -3, -3, 4, 6,
    -- filter=161 channel=32
    -3, -1, -4, 2, 5, -5, -6, -3, 11,
    -- filter=161 channel=33
    -4, 5, -1, 2, -5, -2, 4, 2, -8,
    -- filter=161 channel=34
    -6, 0, -7, 6, 1, -17, 6, 8, -14,
    -- filter=161 channel=35
    -2, 4, -6, 4, -6, 2, -2, -3, -5,
    -- filter=161 channel=36
    -2, 3, 0, 4, 3, 8, -3, 0, 5,
    -- filter=161 channel=37
    1, 1, 3, 12, -4, -4, 1, 0, -11,
    -- filter=161 channel=38
    -4, -6, 6, 7, -3, -9, 0, -3, 1,
    -- filter=161 channel=39
    0, -2, 1, -5, 2, -2, 1, -1, 10,
    -- filter=161 channel=40
    -3, -9, -8, -7, -8, 0, 2, -7, 0,
    -- filter=161 channel=41
    2, 0, 1, -4, 7, -9, 4, 2, -13,
    -- filter=161 channel=42
    1, -6, 2, 0, -4, 0, -3, 6, 3,
    -- filter=161 channel=43
    0, 0, -1, 3, 1, 3, 2, 6, 0,
    -- filter=161 channel=44
    -2, 5, -5, 2, -3, -5, 5, 7, 0,
    -- filter=161 channel=45
    3, 0, -6, 2, -5, -4, -6, 2, -6,
    -- filter=161 channel=46
    -7, -5, 3, 6, -5, 1, 1, 5, 1,
    -- filter=161 channel=47
    7, -6, -3, 8, -2, -9, 4, 0, -9,
    -- filter=161 channel=48
    6, -1, -2, 4, 1, -7, -1, -1, -1,
    -- filter=161 channel=49
    0, 7, 0, 0, -3, 1, -7, 6, 4,
    -- filter=161 channel=50
    -1, -5, -6, -1, -6, 0, -8, 2, 10,
    -- filter=161 channel=51
    4, 6, 0, -5, 2, 0, 5, -2, 4,
    -- filter=161 channel=52
    -5, -2, -12, -1, -7, -2, -5, 2, 4,
    -- filter=161 channel=53
    -2, 4, -4, -8, 5, 3, 4, -5, 4,
    -- filter=161 channel=54
    3, 3, -6, 7, -2, 6, -2, -4, 0,
    -- filter=161 channel=55
    -6, 0, -8, -3, 3, -6, -7, -1, 18,
    -- filter=161 channel=56
    2, 0, 3, 1, -6, -5, 0, -7, 1,
    -- filter=161 channel=57
    0, 2, -3, -4, 5, 6, 1, -4, -5,
    -- filter=161 channel=58
    7, 7, -2, 4, 2, 0, 0, 2, -10,
    -- filter=161 channel=59
    0, -3, 3, -2, 1, -7, 5, 5, -1,
    -- filter=161 channel=60
    -1, 4, 7, 5, -1, -5, 3, 2, -3,
    -- filter=161 channel=61
    2, -3, 1, -2, -4, -2, 3, -6, -6,
    -- filter=161 channel=62
    1, 5, -3, 4, -7, 3, -5, 4, -6,
    -- filter=161 channel=63
    8, -1, 4, 4, -3, -3, -6, 0, -2,
    -- filter=161 channel=64
    -5, 3, 6, -6, 3, -3, -4, 7, 0,
    -- filter=161 channel=65
    4, -5, -3, 0, 6, -5, 0, 4, -1,
    -- filter=161 channel=66
    -1, 1, -8, -3, -1, -5, 7, -4, -10,
    -- filter=161 channel=67
    -5, 0, 5, 5, 1, -6, -5, 7, 1,
    -- filter=161 channel=68
    1, -8, -5, -2, 0, 5, 3, -5, 0,
    -- filter=161 channel=69
    -6, 3, 2, 4, 0, 0, 0, 0, -6,
    -- filter=161 channel=70
    0, -10, -2, -1, -7, -11, -2, 9, 1,
    -- filter=161 channel=71
    -6, -1, 0, -6, -4, -2, -1, -8, -5,
    -- filter=161 channel=72
    -1, -1, -6, 4, 3, 2, -7, 5, 7,
    -- filter=161 channel=73
    -6, 2, -6, 1, 4, 0, -3, -4, 16,
    -- filter=161 channel=74
    4, -3, -9, 6, 0, -2, 6, 5, -5,
    -- filter=161 channel=75
    9, 1, 10, 7, 6, -6, 0, 4, -9,
    -- filter=161 channel=76
    -8, -3, 0, -14, -1, 1, -8, -8, 15,
    -- filter=161 channel=77
    0, 0, 5, -6, 1, -3, -5, -2, 0,
    -- filter=161 channel=78
    4, 3, -1, -3, 4, -8, 6, -4, -8,
    -- filter=161 channel=79
    -9, 5, 1, -1, 3, -7, -1, 9, 7,
    -- filter=161 channel=80
    2, 2, 3, -3, 4, 0, -1, -6, 8,
    -- filter=161 channel=81
    6, 5, -2, 3, 0, -4, -4, -5, -6,
    -- filter=161 channel=82
    1, 5, -4, -4, 6, -5, -2, 2, 4,
    -- filter=161 channel=83
    3, -6, -2, 0, 5, 0, 1, 3, 3,
    -- filter=161 channel=84
    0, -2, 0, -3, 7, 0, -3, 1, 3,
    -- filter=161 channel=85
    5, 0, 0, 0, 3, 3, 4, -4, -6,
    -- filter=161 channel=86
    10, 2, 5, -3, 0, -10, 0, 3, 0,
    -- filter=161 channel=87
    6, 1, 2, -1, 6, 2, -7, 1, 5,
    -- filter=161 channel=88
    0, 3, -5, -6, 0, 4, 3, 2, -5,
    -- filter=161 channel=89
    -12, -1, 4, -7, -3, -5, 4, -4, 10,
    -- filter=161 channel=90
    -9, -4, -11, 4, -2, -5, -5, -4, -9,
    -- filter=161 channel=91
    -5, 5, 0, -5, 0, -5, 2, -1, 12,
    -- filter=161 channel=92
    -5, 0, 0, -6, -8, -9, -6, 0, -9,
    -- filter=161 channel=93
    2, 0, 6, 9, -5, -10, 3, 3, -4,
    -- filter=161 channel=94
    -7, -3, 2, 0, 6, 2, 2, -1, 0,
    -- filter=161 channel=95
    0, 4, -2, -4, -6, -1, -5, -7, -4,
    -- filter=161 channel=96
    0, -4, 4, -3, 1, 0, 5, -2, 7,
    -- filter=161 channel=97
    0, -7, 1, 2, 0, -2, 0, 0, -6,
    -- filter=161 channel=98
    5, -3, -3, 3, 3, -11, -5, -1, 11,
    -- filter=161 channel=99
    -6, 0, -10, -8, 5, 1, 4, 0, 8,
    -- filter=161 channel=100
    7, 2, 4, 0, -4, 3, 1, 1, -10,
    -- filter=161 channel=101
    -6, 2, -1, -1, 2, 3, -5, 7, 2,
    -- filter=161 channel=102
    1, 3, 6, -3, 0, -1, -4, 7, 6,
    -- filter=161 channel=103
    1, 3, 6, 5, -6, -1, 7, 4, -6,
    -- filter=161 channel=104
    -3, 5, 0, -2, -3, 2, -6, 1, 10,
    -- filter=161 channel=105
    -8, -1, 1, 2, -7, 8, 1, -1, 0,
    -- filter=161 channel=106
    -3, -5, 5, -2, 3, 4, -5, 0, 2,
    -- filter=161 channel=107
    -3, 3, -6, 1, -6, -3, -9, 4, 10,
    -- filter=161 channel=108
    5, 8, 0, 5, -5, 0, 4, -4, 3,
    -- filter=161 channel=109
    -3, 4, -11, -3, -3, -10, 0, 5, 14,
    -- filter=161 channel=110
    5, -3, -6, 0, 3, 4, -4, 1, 3,
    -- filter=161 channel=111
    -6, 3, 5, -3, 0, 6, 2, 6, 1,
    -- filter=161 channel=112
    -2, -3, 0, -2, -5, -4, -2, 6, 2,
    -- filter=161 channel=113
    0, 1, -7, 3, -6, -4, 5, 0, -5,
    -- filter=161 channel=114
    -1, 11, 2, -4, 0, 1, -2, 10, 4,
    -- filter=161 channel=115
    -6, -5, 0, 5, -5, -7, -6, -2, -4,
    -- filter=161 channel=116
    -1, 4, -5, -5, 7, 1, 0, -5, 12,
    -- filter=161 channel=117
    -3, -8, 0, -3, 6, 3, 1, 6, -5,
    -- filter=161 channel=118
    4, 0, 2, 2, -5, 4, 4, 0, -1,
    -- filter=161 channel=119
    -2, 5, -8, 7, -5, -14, -3, -6, -12,
    -- filter=161 channel=120
    1, 7, -13, -3, -3, -6, -6, 8, 20,
    -- filter=161 channel=121
    4, -2, 0, -6, -2, -2, -1, 0, -4,
    -- filter=161 channel=122
    -5, -4, -1, -2, -7, -3, -8, -2, -16,
    -- filter=161 channel=123
    -8, -5, 0, 2, -1, 0, -6, 3, -11,
    -- filter=161 channel=124
    4, -4, 1, -8, -7, 3, 3, 2, 10,
    -- filter=161 channel=125
    1, -4, -9, -2, 5, -1, -4, 8, 14,
    -- filter=161 channel=126
    1, 4, 4, 0, 5, -5, 5, -1, 5,
    -- filter=161 channel=127
    -2, 6, 2, -6, -1, -6, -4, 0, 0,
    -- filter=162 channel=0
    4, -5, 10, 2, 2, 10, -4, -1, -5,
    -- filter=162 channel=1
    -2, 3, 8, -1, 4, 2, -6, 1, -3,
    -- filter=162 channel=2
    0, -2, -6, -1, -6, -1, -7, 6, 4,
    -- filter=162 channel=3
    -6, 1, -5, -11, -4, -2, -9, -7, 0,
    -- filter=162 channel=4
    -4, -15, 0, -3, -14, 0, -4, 0, -15,
    -- filter=162 channel=5
    -10, 0, 9, -10, 1, 13, -10, 1, 5,
    -- filter=162 channel=6
    3, 4, -5, 6, -6, 0, 2, -3, -5,
    -- filter=162 channel=7
    -6, -3, 7, 3, -7, 4, -4, 7, -3,
    -- filter=162 channel=8
    -4, 0, -4, 11, -2, 3, 0, -2, -7,
    -- filter=162 channel=9
    1, 2, 2, -5, -3, -2, -7, -5, -9,
    -- filter=162 channel=10
    -2, 4, 0, 3, 1, 3, 3, 3, 3,
    -- filter=162 channel=11
    -6, 1, -1, 5, -6, -6, -4, -9, 0,
    -- filter=162 channel=12
    12, 7, 4, 14, -5, 6, 12, 8, 10,
    -- filter=162 channel=13
    14, 1, 2, 5, 1, -2, 0, 0, -2,
    -- filter=162 channel=14
    6, -2, 1, -4, 2, -5, -4, -1, -2,
    -- filter=162 channel=15
    2, -8, 3, 3, -16, -11, 9, -3, -4,
    -- filter=162 channel=16
    -13, 2, 1, -3, 5, 17, -7, 2, 1,
    -- filter=162 channel=17
    -1, -5, 0, 6, -5, -5, 3, 0, 7,
    -- filter=162 channel=18
    14, 2, -4, 17, 0, -13, 4, -1, -14,
    -- filter=162 channel=19
    2, 2, -4, 2, 5, 3, -4, 2, -7,
    -- filter=162 channel=20
    4, -15, -6, 12, -10, -7, 6, -13, -8,
    -- filter=162 channel=21
    -8, 3, 5, -4, 0, 12, -5, 0, 8,
    -- filter=162 channel=22
    2, 5, -5, 5, 0, -5, 5, 0, -6,
    -- filter=162 channel=23
    2, -9, -7, 9, -25, 1, 13, -17, 4,
    -- filter=162 channel=24
    -3, 3, 3, 1, -3, 3, -1, -2, 0,
    -- filter=162 channel=25
    0, -1, -2, 7, 0, 2, 2, 2, -8,
    -- filter=162 channel=26
    -8, 1, -1, -13, -4, 11, -8, 3, 9,
    -- filter=162 channel=27
    -4, -6, -1, 18, -26, -9, 7, -9, -7,
    -- filter=162 channel=28
    -4, 0, -7, 2, -4, 0, 7, -1, -2,
    -- filter=162 channel=29
    0, -2, 3, 3, -9, -9, 3, -11, -1,
    -- filter=162 channel=30
    -9, -7, -2, -8, -6, -4, -6, -1, -4,
    -- filter=162 channel=31
    -10, 3, -14, 3, -10, 1, -3, -8, 6,
    -- filter=162 channel=32
    -2, -10, 4, 9, -19, 2, 5, 1, -9,
    -- filter=162 channel=33
    3, -2, 0, 3, -17, 2, 3, -5, -12,
    -- filter=162 channel=34
    8, 11, -1, 29, 9, 4, 12, 3, 3,
    -- filter=162 channel=35
    4, 7, 6, 4, -5, 1, 0, -2, 6,
    -- filter=162 channel=36
    2, -7, -7, 7, 5, 8, 1, 10, 4,
    -- filter=162 channel=37
    -3, 0, 13, -3, -9, 5, -4, -6, 6,
    -- filter=162 channel=38
    -3, -3, -7, 6, -7, 4, 4, -2, -4,
    -- filter=162 channel=39
    6, -8, 1, 1, -10, -4, 4, -1, 0,
    -- filter=162 channel=40
    1, 2, -5, -5, -9, -8, 2, -3, 3,
    -- filter=162 channel=41
    13, 11, 18, 14, 33, 5, 20, 19, 1,
    -- filter=162 channel=42
    -4, -5, 1, -10, -6, 6, 3, -10, -3,
    -- filter=162 channel=43
    7, 1, 6, -4, -9, -4, 11, 0, -12,
    -- filter=162 channel=44
    -9, 1, -8, -12, -7, 0, -9, -10, -2,
    -- filter=162 channel=45
    0, -6, 0, -3, -11, 6, 1, 3, -7,
    -- filter=162 channel=46
    9, 9, 5, -1, 1, -10, -2, 2, -3,
    -- filter=162 channel=47
    -7, 1, 1, -10, -2, 5, -12, -4, 11,
    -- filter=162 channel=48
    -13, 2, -7, -8, -1, -1, -3, -7, -3,
    -- filter=162 channel=49
    2, -13, -3, 1, -14, -7, 8, -1, -12,
    -- filter=162 channel=50
    2, 0, -7, -1, -15, -2, 2, -5, 0,
    -- filter=162 channel=51
    -1, -3, 0, -3, -2, 0, -2, -2, 5,
    -- filter=162 channel=52
    5, -6, -8, 16, 1, 4, 5, 5, -5,
    -- filter=162 channel=53
    1, 0, 4, -2, -7, 5, 9, -6, 5,
    -- filter=162 channel=54
    2, -5, -1, 5, 0, 0, -5, -6, 5,
    -- filter=162 channel=55
    12, 0, 2, 15, -5, -5, 13, -10, -4,
    -- filter=162 channel=56
    -1, 9, 3, 13, 5, -6, 10, 1, 5,
    -- filter=162 channel=57
    4, 5, 5, 0, 6, 3, 8, 5, 7,
    -- filter=162 channel=58
    0, 7, 4, -2, 6, 1, -6, 0, -3,
    -- filter=162 channel=59
    0, 6, -5, -3, 9, 4, 1, 2, 3,
    -- filter=162 channel=60
    -7, -7, 0, 6, -3, -3, -2, 4, -5,
    -- filter=162 channel=61
    0, 0, -2, 10, 3, 1, 3, 0, 1,
    -- filter=162 channel=62
    2, -6, -2, -1, -2, -1, 0, 6, 6,
    -- filter=162 channel=63
    2, 6, 10, -3, 2, 6, 0, 1, 6,
    -- filter=162 channel=64
    7, 0, -7, 4, 4, -1, -3, 1, -6,
    -- filter=162 channel=65
    3, -3, 2, -5, -4, 2, -2, 3, -4,
    -- filter=162 channel=66
    16, 4, 4, 17, 6, 7, 6, 13, 9,
    -- filter=162 channel=67
    -2, -3, -1, 1, 7, -8, 1, 6, -1,
    -- filter=162 channel=68
    -1, 2, 0, -1, -1, -8, 3, -4, 2,
    -- filter=162 channel=69
    7, -5, 8, 5, -6, 0, -1, -2, 4,
    -- filter=162 channel=70
    6, -1, -3, 15, -18, -1, 13, -15, -3,
    -- filter=162 channel=71
    -8, 1, 4, 0, 2, 7, -8, -6, 3,
    -- filter=162 channel=72
    -5, 2, 2, 0, 0, 1, -2, -1, -2,
    -- filter=162 channel=73
    2, -6, -3, 14, -14, -2, 8, -4, -8,
    -- filter=162 channel=74
    -5, -4, -10, 14, -3, 7, 4, 1, -7,
    -- filter=162 channel=75
    1, 4, 13, -9, -4, 12, -6, 8, 7,
    -- filter=162 channel=76
    9, -7, 1, 15, -11, -9, 3, -1, -8,
    -- filter=162 channel=77
    7, -6, -2, -4, -6, -6, -5, 5, 6,
    -- filter=162 channel=78
    -6, 4, -1, 1, 4, -2, -1, -6, 7,
    -- filter=162 channel=79
    6, 0, -2, 19, -14, -5, 18, 1, -13,
    -- filter=162 channel=80
    0, 0, 0, -13, -5, 1, -2, 0, 5,
    -- filter=162 channel=81
    1, -4, 1, 4, -5, -6, 2, -1, 2,
    -- filter=162 channel=82
    -7, -3, 1, -7, 1, -1, 0, -4, -2,
    -- filter=162 channel=83
    -3, -3, 1, 2, 0, -1, -8, 0, -2,
    -- filter=162 channel=84
    4, -6, 3, 12, -5, -3, 9, -1, -8,
    -- filter=162 channel=85
    -2, 1, 2, -6, 3, 5, -1, 0, 0,
    -- filter=162 channel=86
    4, 5, -2, 19, 0, 9, 7, -1, 0,
    -- filter=162 channel=87
    8, 7, 4, 17, -7, 1, 6, -5, -7,
    -- filter=162 channel=88
    -3, 5, 0, -3, 6, 2, 6, 3, 4,
    -- filter=162 channel=89
    5, -7, 7, 6, -10, -1, 9, -3, 0,
    -- filter=162 channel=90
    -4, 6, 2, 4, -3, 0, 3, 4, -1,
    -- filter=162 channel=91
    8, -15, 0, 11, -22, -4, 10, -13, -11,
    -- filter=162 channel=92
    -3, 5, 2, 1, 1, -4, -1, -1, -5,
    -- filter=162 channel=93
    -12, 4, -1, -15, 4, 6, -1, 0, 9,
    -- filter=162 channel=94
    -1, -4, 2, 6, 4, 0, 0, 7, -6,
    -- filter=162 channel=95
    -1, 7, 3, -7, 0, 6, -6, -8, 3,
    -- filter=162 channel=96
    2, -3, -5, 1, 4, 1, -3, 0, -7,
    -- filter=162 channel=97
    5, 0, -1, -10, -9, -6, -3, -3, -8,
    -- filter=162 channel=98
    2, -5, 1, -6, -10, -4, 0, -2, -9,
    -- filter=162 channel=99
    -5, 1, -13, 9, -14, 10, 8, 0, 4,
    -- filter=162 channel=100
    7, 10, 7, 3, 4, -7, 4, 3, 3,
    -- filter=162 channel=101
    -5, -1, -10, -3, -5, 0, 2, -1, -5,
    -- filter=162 channel=102
    -1, -3, -1, -4, -4, -6, 0, -7, -1,
    -- filter=162 channel=103
    -6, 2, 0, -21, 3, 10, -11, -8, 0,
    -- filter=162 channel=104
    -2, 4, 0, -10, 7, 4, -5, 7, -1,
    -- filter=162 channel=105
    -2, -3, 8, 6, -1, -2, -2, -11, 0,
    -- filter=162 channel=106
    6, -5, 1, 7, 3, -6, -4, 6, -8,
    -- filter=162 channel=107
    8, 2, 6, 14, -18, 1, 7, -11, -10,
    -- filter=162 channel=108
    5, 4, 8, 7, 11, -3, 3, 11, -4,
    -- filter=162 channel=109
    4, 1, -7, 13, -3, -7, 8, -9, -4,
    -- filter=162 channel=110
    5, 5, 6, 2, -6, 14, 7, 7, 9,
    -- filter=162 channel=111
    5, -4, -5, 4, 0, -7, 7, 0, 3,
    -- filter=162 channel=112
    -1, 0, 0, 6, -17, 4, 1, -5, -2,
    -- filter=162 channel=113
    0, -1, 0, 1, -8, 5, 7, -10, -6,
    -- filter=162 channel=114
    4, -10, -5, 20, -8, -5, 7, -2, -13,
    -- filter=162 channel=115
    8, 4, -1, 0, -3, 5, -4, 7, 3,
    -- filter=162 channel=116
    5, -12, 0, 2, -7, -2, 4, 5, -1,
    -- filter=162 channel=117
    4, 0, 5, 4, -2, 7, 4, 7, 5,
    -- filter=162 channel=118
    -2, 1, -6, -5, -2, 3, 0, -2, 2,
    -- filter=162 channel=119
    3, 11, -13, 28, 15, -9, 18, 17, -9,
    -- filter=162 channel=120
    -10, -14, -17, 12, -31, -8, 5, -18, -2,
    -- filter=162 channel=121
    0, -4, 8, 0, 10, 0, 7, 10, 6,
    -- filter=162 channel=122
    -14, 8, 3, -16, 1, 24, -19, 0, 19,
    -- filter=162 channel=123
    0, 4, -2, 6, 9, 2, 4, 4, 5,
    -- filter=162 channel=124
    8, 0, 1, 7, -10, 5, -3, 1, -6,
    -- filter=162 channel=125
    3, -3, 4, 2, 2, 7, -1, -6, 3,
    -- filter=162 channel=126
    7, 6, 7, 0, 8, -12, 3, 5, -5,
    -- filter=162 channel=127
    7, 0, 5, -3, 3, 3, 0, 6, 2,
    -- filter=163 channel=0
    0, -4, 6, -6, 1, -2, 8, 5, -1,
    -- filter=163 channel=1
    -5, -7, 3, -5, -4, -6, 0, -7, -2,
    -- filter=163 channel=2
    -6, 4, 1, -7, 0, -2, -6, -4, 1,
    -- filter=163 channel=3
    0, 1, 4, -4, 4, -2, 3, 5, 1,
    -- filter=163 channel=4
    0, 7, 6, -5, 0, -1, 3, 0, 6,
    -- filter=163 channel=5
    -1, 4, -3, 3, -5, 5, -4, -1, -2,
    -- filter=163 channel=6
    2, 7, 6, -2, -6, 1, -2, 6, -6,
    -- filter=163 channel=7
    -5, -1, -3, -7, -5, 7, 0, -5, -4,
    -- filter=163 channel=8
    0, -4, 3, -3, 0, -6, -6, 0, 1,
    -- filter=163 channel=9
    3, -6, -2, 3, 0, -7, -2, -1, 1,
    -- filter=163 channel=10
    -2, 5, -2, 0, -5, 0, -3, 5, 4,
    -- filter=163 channel=11
    2, 6, 3, -2, -1, 0, -2, 6, 2,
    -- filter=163 channel=12
    3, -2, 3, 6, -4, 0, -2, -2, -1,
    -- filter=163 channel=13
    6, 0, 6, 4, -5, 2, -7, -7, -3,
    -- filter=163 channel=14
    0, -3, 4, -4, 6, -4, 0, 6, -4,
    -- filter=163 channel=15
    1, -3, 0, -6, 3, 0, -4, -4, 1,
    -- filter=163 channel=16
    5, 7, -2, 7, -2, -4, 0, -4, -5,
    -- filter=163 channel=17
    -6, 0, 0, 3, 0, 4, -2, 1, -1,
    -- filter=163 channel=18
    -4, 1, 0, 6, -7, 0, 1, 2, -4,
    -- filter=163 channel=19
    6, 2, 1, -1, 4, -3, 0, -3, -2,
    -- filter=163 channel=20
    -5, 0, 1, 5, 2, -6, 2, 1, 7,
    -- filter=163 channel=21
    -2, 6, -3, -1, 5, 0, -5, -7, 0,
    -- filter=163 channel=22
    1, -2, 8, 4, -6, 5, 1, -5, 7,
    -- filter=163 channel=23
    -5, 7, 0, -6, -2, -5, 4, -1, -1,
    -- filter=163 channel=24
    -2, -6, 0, 0, 4, 6, -7, -2, -4,
    -- filter=163 channel=25
    -6, 0, -5, 6, -7, -3, 6, 0, -6,
    -- filter=163 channel=26
    4, -6, 0, -2, 3, 0, -5, -2, 4,
    -- filter=163 channel=27
    -9, 0, 1, -8, 3, 1, 5, 1, -3,
    -- filter=163 channel=28
    -2, 7, -1, -3, -3, 1, 6, -3, 4,
    -- filter=163 channel=29
    5, 6, -3, 6, 4, 0, -5, -1, -6,
    -- filter=163 channel=30
    5, -7, 0, 4, 6, 1, 0, 1, 2,
    -- filter=163 channel=31
    -5, -3, -1, -6, -7, -1, -5, 0, 2,
    -- filter=163 channel=32
    5, -7, -3, 0, -3, -6, 2, -3, 1,
    -- filter=163 channel=33
    -5, -5, 6, 0, 2, 2, -2, 4, -5,
    -- filter=163 channel=34
    4, -2, 7, 0, 2, 5, 4, -7, 2,
    -- filter=163 channel=35
    7, -3, -6, -6, -4, 2, 1, -1, 4,
    -- filter=163 channel=36
    -2, 5, 7, 0, -7, 1, 1, -3, -6,
    -- filter=163 channel=37
    -6, -3, 2, 6, -4, -3, 0, 3, -2,
    -- filter=163 channel=38
    0, -7, 5, -5, 6, 6, 4, -5, 0,
    -- filter=163 channel=39
    0, 5, -6, 5, -3, 1, 2, 2, 0,
    -- filter=163 channel=40
    -4, -2, 4, 5, -6, 0, -3, 2, -5,
    -- filter=163 channel=41
    3, 0, -2, 3, 3, 6, 6, -6, -7,
    -- filter=163 channel=42
    -5, 4, 2, 3, 5, 7, -2, -6, -5,
    -- filter=163 channel=43
    5, 0, -2, 0, 6, -3, 1, 5, 0,
    -- filter=163 channel=44
    -5, 6, 4, 5, 3, -3, -4, -6, -6,
    -- filter=163 channel=45
    -6, 0, 7, -3, -7, 4, 0, 0, 4,
    -- filter=163 channel=46
    3, 1, 7, 0, -5, 3, 6, 0, 5,
    -- filter=163 channel=47
    6, 6, -3, 2, 1, 6, 0, -6, 7,
    -- filter=163 channel=48
    -3, -5, 7, -2, 4, 6, 5, -3, 6,
    -- filter=163 channel=49
    6, 5, -6, 0, 6, 0, 4, 4, 0,
    -- filter=163 channel=50
    -6, -7, -1, -6, -3, 3, -8, -4, 0,
    -- filter=163 channel=51
    -4, 7, -3, 1, -2, 3, 4, -5, 4,
    -- filter=163 channel=52
    5, 7, -5, 0, 3, 6, -6, -1, -3,
    -- filter=163 channel=53
    5, 4, -1, 0, 0, -2, -3, 6, 0,
    -- filter=163 channel=54
    -2, -2, -6, 5, 6, -6, -4, 2, 1,
    -- filter=163 channel=55
    4, 2, -4, 1, -4, -2, 3, -3, -8,
    -- filter=163 channel=56
    -5, -3, 8, -5, -4, 6, 0, 6, -6,
    -- filter=163 channel=57
    7, -5, -3, 6, -5, 2, 0, 1, 0,
    -- filter=163 channel=58
    0, -3, -4, 0, 6, -6, -1, -7, 3,
    -- filter=163 channel=59
    0, 6, 2, 5, -4, 0, -1, 4, 0,
    -- filter=163 channel=60
    1, 4, -5, -6, 0, 2, 2, 0, 0,
    -- filter=163 channel=61
    -7, 0, 2, 6, -4, -2, -1, 1, -2,
    -- filter=163 channel=62
    0, -5, 4, 7, -4, -5, -4, -4, 1,
    -- filter=163 channel=63
    7, 4, 6, -6, 0, 3, -2, -6, 7,
    -- filter=163 channel=64
    -4, 1, -1, 0, -3, -5, 2, -6, -5,
    -- filter=163 channel=65
    -4, -7, 2, -3, 5, 0, 0, 2, 3,
    -- filter=163 channel=66
    -6, -6, -2, 1, -2, 5, -7, -5, -2,
    -- filter=163 channel=67
    -3, 7, -2, -3, -7, 4, 6, 0, -2,
    -- filter=163 channel=68
    4, 3, -6, 7, -7, -5, -6, -2, 5,
    -- filter=163 channel=69
    6, 4, -4, -4, 4, -1, 7, 5, -2,
    -- filter=163 channel=70
    -1, 1, -4, 1, -6, 0, -1, -4, -1,
    -- filter=163 channel=71
    -6, 3, -5, 2, 4, -5, 3, -5, 1,
    -- filter=163 channel=72
    0, -7, 5, -4, -6, -5, 5, -6, 2,
    -- filter=163 channel=73
    6, -6, -3, -2, -1, 0, 2, 6, 5,
    -- filter=163 channel=74
    -3, -1, -5, 5, 1, -3, -2, -2, -4,
    -- filter=163 channel=75
    -6, 3, 5, 0, -2, 2, -4, 6, -4,
    -- filter=163 channel=76
    -3, 6, -7, 0, 1, 6, -3, 0, 6,
    -- filter=163 channel=77
    7, 5, -1, -4, -2, -5, -6, -1, -3,
    -- filter=163 channel=78
    3, 5, 2, -5, 0, 6, -4, -3, 0,
    -- filter=163 channel=79
    1, -2, -1, -4, -4, -8, 6, -8, 6,
    -- filter=163 channel=80
    1, -7, -3, 0, 1, -2, -6, 4, -6,
    -- filter=163 channel=81
    5, 1, -2, -6, -3, -4, -2, -7, 5,
    -- filter=163 channel=82
    -5, 5, -1, -3, -4, 1, 2, 0, 5,
    -- filter=163 channel=83
    6, -2, 5, -3, 0, 0, 1, -5, 0,
    -- filter=163 channel=84
    3, -2, -5, -5, 3, -7, -3, -6, 6,
    -- filter=163 channel=85
    4, -1, 2, 1, -2, 2, -1, 4, 1,
    -- filter=163 channel=86
    -2, -3, -5, -4, -6, -3, 2, 0, 6,
    -- filter=163 channel=87
    1, 1, 7, 2, 3, -6, 4, -3, 5,
    -- filter=163 channel=88
    0, 0, 3, -1, -3, 1, 3, 4, 5,
    -- filter=163 channel=89
    -1, 4, -7, 5, 5, -5, -8, -7, 3,
    -- filter=163 channel=90
    6, 0, 1, 6, -4, -6, -3, -2, 0,
    -- filter=163 channel=91
    3, 0, 0, 2, 3, 0, -7, 5, 5,
    -- filter=163 channel=92
    4, 4, 1, -2, -3, 0, 6, 5, -6,
    -- filter=163 channel=93
    -1, -4, 4, 5, -5, -1, -2, 0, -3,
    -- filter=163 channel=94
    0, -4, 4, 1, 4, 6, -6, 2, -4,
    -- filter=163 channel=95
    -4, 3, 0, -7, -7, 7, 6, -5, 0,
    -- filter=163 channel=96
    -1, 2, 3, -2, -2, 1, 6, 0, 0,
    -- filter=163 channel=97
    2, 0, 1, -7, 2, 3, -6, -6, -7,
    -- filter=163 channel=98
    -6, 2, 3, 1, -5, -1, -7, 0, -7,
    -- filter=163 channel=99
    -5, 3, -5, -8, 2, 6, 2, 1, -1,
    -- filter=163 channel=100
    6, 5, -4, 0, -4, -2, 3, -1, 3,
    -- filter=163 channel=101
    6, -4, 2, 5, 5, 1, -6, -2, 2,
    -- filter=163 channel=102
    5, 4, 3, 6, 0, -3, -5, 5, 0,
    -- filter=163 channel=103
    5, -3, -1, 0, -4, 5, -7, -4, 5,
    -- filter=163 channel=104
    2, 0, 4, -6, 5, 1, -2, 3, 1,
    -- filter=163 channel=105
    3, 2, -4, 3, 0, -4, -6, 7, -5,
    -- filter=163 channel=106
    4, -4, 5, -4, 0, -7, 2, 3, 0,
    -- filter=163 channel=107
    0, -3, 4, 2, 2, 3, 7, 3, 7,
    -- filter=163 channel=108
    -5, -5, -6, -6, 3, -1, -3, -1, -5,
    -- filter=163 channel=109
    -9, 5, 6, 0, -2, -1, -1, 4, 1,
    -- filter=163 channel=110
    -1, 0, -1, -3, -2, 0, 6, 0, 7,
    -- filter=163 channel=111
    -7, -4, -4, -4, -7, 0, -6, 5, -1,
    -- filter=163 channel=112
    1, -1, 3, 5, 6, 4, -6, 6, 1,
    -- filter=163 channel=113
    -6, 5, 6, 3, -5, 5, -7, 6, 5,
    -- filter=163 channel=114
    -1, -1, -3, 4, -7, -6, 0, -3, -5,
    -- filter=163 channel=115
    -5, 3, 5, 6, -3, 1, 4, -2, 6,
    -- filter=163 channel=116
    0, -4, -2, -7, -8, 3, 3, -6, 0,
    -- filter=163 channel=117
    2, 4, -4, -2, 0, -3, 0, -1, 4,
    -- filter=163 channel=118
    -6, 7, -3, 0, 3, 2, 4, -3, -6,
    -- filter=163 channel=119
    5, -3, 5, 0, 0, 1, 1, -7, 6,
    -- filter=163 channel=120
    0, -5, 6, -3, 1, -4, -1, -7, 7,
    -- filter=163 channel=121
    6, 2, -5, 5, -2, 6, -6, 1, 3,
    -- filter=163 channel=122
    -5, -3, -2, -3, 0, -1, -3, -4, 1,
    -- filter=163 channel=123
    -2, 0, 1, -2, -7, 5, 5, 4, 0,
    -- filter=163 channel=124
    -4, 1, 3, -3, 0, 7, 2, 0, 5,
    -- filter=163 channel=125
    -5, -6, 2, 6, 3, 4, -4, -7, 0,
    -- filter=163 channel=126
    -2, 6, 0, -2, -2, 2, -7, 0, 4,
    -- filter=163 channel=127
    0, -2, 5, 5, -3, 0, 2, 3, -7,
    -- filter=164 channel=0
    6, 1, -4, -1, 0, 1, 4, 2, -6,
    -- filter=164 channel=1
    2, -2, 4, -3, -7, -1, 1, 7, 5,
    -- filter=164 channel=2
    -7, 2, -4, -1, 6, 8, 6, 1, -4,
    -- filter=164 channel=3
    -1, 6, 5, 0, -1, -1, -9, -5, 1,
    -- filter=164 channel=4
    -2, 0, -2, 0, 9, 13, 12, 1, 8,
    -- filter=164 channel=5
    -5, -8, 0, 6, -10, 2, 0, -7, -3,
    -- filter=164 channel=6
    -4, -2, -1, -5, -9, -3, -4, 2, 1,
    -- filter=164 channel=7
    -1, -5, 1, 0, 1, -6, 7, 6, -3,
    -- filter=164 channel=8
    -4, -4, -7, -4, -2, 9, 2, -4, -1,
    -- filter=164 channel=9
    -11, 0, 0, -4, 0, -2, 5, 9, 1,
    -- filter=164 channel=10
    0, -4, -10, 0, -5, -10, -8, 0, 0,
    -- filter=164 channel=11
    -5, -10, -12, -5, -4, -6, -5, 0, -4,
    -- filter=164 channel=12
    -6, -4, 2, -5, -2, 8, -8, -4, 4,
    -- filter=164 channel=13
    -3, -11, -2, -9, 0, -7, -2, 2, 9,
    -- filter=164 channel=14
    -1, 3, 4, 2, -4, 1, -5, 0, 3,
    -- filter=164 channel=15
    -2, -8, -12, -7, -10, -9, -6, 0, -3,
    -- filter=164 channel=16
    -7, -2, 0, 5, 3, -1, 5, 7, 3,
    -- filter=164 channel=17
    1, 3, 6, -4, 3, 0, 3, -7, -2,
    -- filter=164 channel=18
    -3, -12, -17, -10, -4, 0, -5, -1, 8,
    -- filter=164 channel=19
    7, -3, 0, 7, 3, 2, 3, -5, 7,
    -- filter=164 channel=20
    2, -12, -9, -13, -10, -9, -13, -3, -9,
    -- filter=164 channel=21
    -6, -9, 0, -1, 7, -6, -1, 15, 9,
    -- filter=164 channel=22
    3, -5, -7, -6, -4, -1, 0, -8, 5,
    -- filter=164 channel=23
    -1, -16, -10, -19, -14, -5, 3, 8, 7,
    -- filter=164 channel=24
    4, -3, 4, 0, 3, 3, 6, 3, 4,
    -- filter=164 channel=25
    -10, -15, -9, -7, -6, -2, 1, 10, 11,
    -- filter=164 channel=26
    -8, 3, -3, 1, 0, 5, 0, 7, 0,
    -- filter=164 channel=27
    -11, -5, -3, -13, 2, -3, 7, 12, 18,
    -- filter=164 channel=28
    3, -2, 0, 4, -1, 3, -3, 2, -4,
    -- filter=164 channel=29
    -1, -7, 0, -7, -3, -7, -9, 0, 2,
    -- filter=164 channel=30
    2, -2, 4, -2, -4, -7, 3, 6, 0,
    -- filter=164 channel=31
    -5, -14, -7, -6, 0, -7, 4, 19, 16,
    -- filter=164 channel=32
    -1, -15, -13, -14, -5, -11, 0, 10, -1,
    -- filter=164 channel=33
    -2, -3, -8, -13, -2, 0, 0, 8, 1,
    -- filter=164 channel=34
    -10, 3, 3, -6, -6, -8, 8, -6, 6,
    -- filter=164 channel=35
    5, -5, 6, -4, -6, 0, 7, -3, 0,
    -- filter=164 channel=36
    0, -2, 5, -5, 3, 5, 0, 4, 7,
    -- filter=164 channel=37
    -1, -1, 10, 2, -3, 11, 13, 12, -1,
    -- filter=164 channel=38
    1, -7, -2, -8, -3, -10, -5, 7, 8,
    -- filter=164 channel=39
    1, 0, 0, -6, -8, 0, -4, -7, 3,
    -- filter=164 channel=40
    -1, -1, -5, -7, -3, -5, -7, -4, 3,
    -- filter=164 channel=41
    -2, -1, -12, -6, -5, 3, 1, 1, 4,
    -- filter=164 channel=42
    -8, 1, -3, -3, -5, 4, 2, 5, 0,
    -- filter=164 channel=43
    -4, 0, -8, -8, -7, -6, 0, 1, 0,
    -- filter=164 channel=44
    -7, -7, 1, 0, 3, 6, 3, 14, 15,
    -- filter=164 channel=45
    1, 4, 4, 2, -5, -3, -1, 2, 0,
    -- filter=164 channel=46
    6, -6, 3, -3, -3, 1, -7, 4, -5,
    -- filter=164 channel=47
    1, -7, 4, -1, -7, 4, 8, 5, 12,
    -- filter=164 channel=48
    -10, 1, -5, -10, 1, 0, 5, 16, 8,
    -- filter=164 channel=49
    -5, 2, -12, -10, 1, 0, -6, 4, 4,
    -- filter=164 channel=50
    0, -2, 2, -4, 0, 0, 0, 12, 5,
    -- filter=164 channel=51
    1, -2, -6, -3, 0, 0, -2, -2, 1,
    -- filter=164 channel=52
    -5, -2, -2, 1, 1, -4, 0, -5, 0,
    -- filter=164 channel=53
    -1, -9, -8, -2, 1, -3, 1, -5, -7,
    -- filter=164 channel=54
    6, 0, 0, 0, 2, 0, 4, 0, 2,
    -- filter=164 channel=55
    -8, -14, -12, -18, -2, 0, -6, 3, 1,
    -- filter=164 channel=56
    1, -1, -4, -4, -8, -2, -3, -4, 11,
    -- filter=164 channel=57
    1, 4, -6, -2, 0, -4, -6, 0, -3,
    -- filter=164 channel=58
    0, 7, 3, 3, 1, -5, 3, -4, -5,
    -- filter=164 channel=59
    -10, -9, -3, -7, 4, -7, 1, 16, 9,
    -- filter=164 channel=60
    -3, -5, 6, 4, 4, -5, 3, 6, -3,
    -- filter=164 channel=61
    1, -8, -6, 4, 2, 0, -2, -3, 7,
    -- filter=164 channel=62
    6, -7, 0, 7, 4, -5, 6, 0, 4,
    -- filter=164 channel=63
    -2, -3, 0, -1, -8, -4, 0, -8, -4,
    -- filter=164 channel=64
    -8, -6, 5, -2, 1, -7, 6, -4, 5,
    -- filter=164 channel=65
    0, 2, -7, -5, -2, -2, 6, -4, -6,
    -- filter=164 channel=66
    6, -5, 5, -10, -7, 4, -7, 0, 0,
    -- filter=164 channel=67
    -5, -5, 2, 0, 2, -3, 7, -3, 5,
    -- filter=164 channel=68
    4, -3, 0, -7, 2, 1, 0, 7, -4,
    -- filter=164 channel=69
    1, -8, -7, 5, -2, 1, 1, 2, 0,
    -- filter=164 channel=70
    4, -9, 4, -6, -3, 0, 2, 11, 5,
    -- filter=164 channel=71
    8, 7, -5, 7, 6, -1, -2, -5, 5,
    -- filter=164 channel=72
    -8, -4, 0, -5, 1, -1, 10, 15, 6,
    -- filter=164 channel=73
    -9, -5, -11, -3, 5, -1, 5, -3, 1,
    -- filter=164 channel=74
    -5, -9, 5, 3, 8, 2, 8, 7, 5,
    -- filter=164 channel=75
    3, -3, -3, 2, -17, -2, 6, -4, -2,
    -- filter=164 channel=76
    -5, -8, 0, -10, 0, -12, -8, -6, -6,
    -- filter=164 channel=77
    0, -2, -4, -3, -4, 6, 2, -3, -5,
    -- filter=164 channel=78
    -1, -3, 2, 5, -3, -5, 2, 0, 3,
    -- filter=164 channel=79
    3, -10, -6, -22, -20, -12, -12, 9, 13,
    -- filter=164 channel=80
    -13, -5, 0, -14, 1, 0, 9, 13, 15,
    -- filter=164 channel=81
    -5, -1, -6, 2, 6, 0, -3, -6, -6,
    -- filter=164 channel=82
    3, 2, -4, 2, 5, -4, -5, 5, 4,
    -- filter=164 channel=83
    -7, 5, -4, 7, 9, 0, 10, -1, 9,
    -- filter=164 channel=84
    -6, -8, 1, -8, -7, -6, -6, -3, 0,
    -- filter=164 channel=85
    3, 5, -2, 3, 7, 0, 0, -1, -2,
    -- filter=164 channel=86
    -7, -10, -1, -9, 3, -4, 6, -5, -2,
    -- filter=164 channel=87
    0, -10, -9, -9, -9, -3, -3, 1, 3,
    -- filter=164 channel=88
    -8, -5, 3, -3, 2, 2, 5, 11, 0,
    -- filter=164 channel=89
    -9, -8, -7, -11, -5, -4, -2, 12, 5,
    -- filter=164 channel=90
    -3, 5, 7, 3, 2, -1, 0, 9, 8,
    -- filter=164 channel=91
    -9, -4, -10, -8, 5, 7, 11, 2, 8,
    -- filter=164 channel=92
    -6, -2, 5, -7, 1, 1, -2, 0, -3,
    -- filter=164 channel=93
    -6, -6, 0, 8, 7, 10, 9, 10, 12,
    -- filter=164 channel=94
    0, -1, 0, 2, 0, -1, -7, 2, -2,
    -- filter=164 channel=95
    -5, 0, -3, 5, 0, 0, 6, -6, 1,
    -- filter=164 channel=96
    2, 4, -5, -5, 6, -2, 6, -3, -3,
    -- filter=164 channel=97
    5, -1, -7, 4, -4, 0, -1, 3, -5,
    -- filter=164 channel=98
    -2, -5, -1, -17, -4, 2, 0, 6, 14,
    -- filter=164 channel=99
    -4, -18, -5, -12, -6, -4, 4, 16, 7,
    -- filter=164 channel=100
    -4, 2, -1, -4, -5, -5, -6, -2, 8,
    -- filter=164 channel=101
    -6, -1, 0, -3, 2, 0, 7, 4, 10,
    -- filter=164 channel=102
    -5, -7, 4, -3, -1, 5, 5, -2, 1,
    -- filter=164 channel=103
    -7, 0, 4, 2, -10, -4, 0, 13, 2,
    -- filter=164 channel=104
    -9, -4, 0, -1, 0, -4, 3, 16, 8,
    -- filter=164 channel=105
    1, -2, -4, 3, 4, -5, -8, -6, -6,
    -- filter=164 channel=106
    3, 0, 1, 2, 5, -8, -5, 0, -5,
    -- filter=164 channel=107
    -7, -3, 0, 0, -9, 0, -3, 1, 2,
    -- filter=164 channel=108
    5, -1, -7, -8, 2, -3, -2, 3, 1,
    -- filter=164 channel=109
    -10, -17, -6, -10, -5, -5, 7, 8, 5,
    -- filter=164 channel=110
    -1, -9, -3, -7, -10, -10, -4, 0, 7,
    -- filter=164 channel=111
    -2, 5, 5, 0, 4, -2, -8, -2, 5,
    -- filter=164 channel=112
    -9, -5, -6, -2, -6, 3, 1, 10, 5,
    -- filter=164 channel=113
    5, -3, 4, -2, -3, -7, 5, -2, 8,
    -- filter=164 channel=114
    -7, -18, -7, -13, -2, -1, -6, 4, -4,
    -- filter=164 channel=115
    0, -4, 6, -4, -2, -6, -4, -6, -4,
    -- filter=164 channel=116
    -5, -7, -9, -6, 2, 7, 3, 5, 13,
    -- filter=164 channel=117
    -3, 4, -4, 0, 1, -1, -6, 6, 8,
    -- filter=164 channel=118
    1, 0, -1, -1, 2, 3, 5, 5, 5,
    -- filter=164 channel=119
    -9, 1, -1, 4, 1, 0, 0, 6, 13,
    -- filter=164 channel=120
    -3, -18, -5, -15, -8, 7, 8, 4, 11,
    -- filter=164 channel=121
    1, -3, -3, 0, -5, 3, 3, -4, 8,
    -- filter=164 channel=122
    -6, -8, 9, 5, 2, 8, 20, 22, 18,
    -- filter=164 channel=123
    5, 3, -4, -2, 4, 3, 2, 4, 2,
    -- filter=164 channel=124
    4, -2, -4, 4, -3, -6, 4, -7, 2,
    -- filter=164 channel=125
    -5, -3, -10, -14, 3, 8, 2, 13, 17,
    -- filter=164 channel=126
    0, -2, 1, -6, -7, -12, -2, 2, 3,
    -- filter=164 channel=127
    -2, -1, 0, -7, 2, 0, 4, 5, 6,
    -- filter=165 channel=0
    9, 1, 5, 7, -3, 0, 1, 5, 0,
    -- filter=165 channel=1
    -7, -4, 6, -2, -10, -7, 6, 3, -3,
    -- filter=165 channel=2
    -5, -6, 0, 0, -4, -4, 2, -5, -6,
    -- filter=165 channel=3
    9, 2, -2, 5, 0, -2, 0, 13, -3,
    -- filter=165 channel=4
    -11, -9, -5, 3, -7, -7, 7, 5, -5,
    -- filter=165 channel=5
    -2, 6, 5, 2, 7, 1, 6, 10, 8,
    -- filter=165 channel=6
    -1, 0, -1, -3, -8, -4, -5, -6, -3,
    -- filter=165 channel=7
    3, -5, 1, 3, 2, -5, 0, 2, 6,
    -- filter=165 channel=8
    3, -2, 3, -10, 2, -7, -4, 0, -1,
    -- filter=165 channel=9
    -5, -4, 7, -7, 9, 9, -3, 4, 0,
    -- filter=165 channel=10
    -2, 0, 3, -4, -4, 6, -15, -11, 7,
    -- filter=165 channel=11
    -1, 1, -4, 6, 3, -9, -3, -6, -8,
    -- filter=165 channel=12
    -1, -6, 3, 5, 2, -7, -7, -5, 0,
    -- filter=165 channel=13
    2, 5, 1, -13, -7, -2, -15, -6, 2,
    -- filter=165 channel=14
    0, -4, -4, -6, 2, 2, -6, 7, -1,
    -- filter=165 channel=15
    -5, -3, -3, -7, 2, 1, -3, -9, -12,
    -- filter=165 channel=16
    -7, 4, 3, -7, 7, 3, 0, 5, 5,
    -- filter=165 channel=17
    -5, -6, 1, -6, 5, -3, -2, 4, 6,
    -- filter=165 channel=18
    5, -3, 0, -4, -10, -10, -4, -8, -13,
    -- filter=165 channel=19
    4, 3, -6, 0, 4, -6, 5, 3, 3,
    -- filter=165 channel=20
    -4, 7, -7, 4, 1, 0, 3, -3, 0,
    -- filter=165 channel=21
    -6, -4, 7, -7, 2, 5, -6, 1, 2,
    -- filter=165 channel=22
    0, -4, 0, 6, 4, -5, 7, 3, -5,
    -- filter=165 channel=23
    8, 13, 5, -5, -3, 7, -10, 0, -5,
    -- filter=165 channel=24
    0, 6, -4, 2, -6, 2, 5, 1, 3,
    -- filter=165 channel=25
    2, -1, 8, -6, -1, 6, -5, -15, 5,
    -- filter=165 channel=26
    6, -1, -2, 0, -2, -2, 5, -4, 3,
    -- filter=165 channel=27
    -3, 0, 14, -7, 1, 3, -18, -16, -3,
    -- filter=165 channel=28
    2, -1, 0, -2, 2, -4, 7, -7, -3,
    -- filter=165 channel=29
    7, -6, -8, -4, -8, -4, -4, -7, -7,
    -- filter=165 channel=30
    -5, 7, 7, 3, 7, 3, -5, 3, 3,
    -- filter=165 channel=31
    1, 10, 8, -1, 14, 24, -22, -6, 19,
    -- filter=165 channel=32
    2, 5, 5, -14, -8, 0, -6, -17, -13,
    -- filter=165 channel=33
    0, 8, 9, 2, -2, 6, -14, 2, -1,
    -- filter=165 channel=34
    -5, 10, 6, -10, 12, -4, -1, 4, 2,
    -- filter=165 channel=35
    -5, 1, -6, 7, -7, 6, -1, -2, 2,
    -- filter=165 channel=36
    -4, 0, 0, -5, 0, 8, -10, -3, 0,
    -- filter=165 channel=37
    4, 4, -3, 1, -1, 6, 3, -4, 0,
    -- filter=165 channel=38
    3, -2, -2, 3, -4, 9, -11, 3, 7,
    -- filter=165 channel=39
    4, 1, -4, -6, -8, -5, -2, -8, -1,
    -- filter=165 channel=40
    0, -3, 3, -5, 0, -3, 5, 0, 0,
    -- filter=165 channel=41
    -10, -3, -3, -12, -5, -11, -13, -14, -3,
    -- filter=165 channel=42
    -2, 5, 2, 6, 0, -1, -1, -2, 0,
    -- filter=165 channel=43
    4, 1, -3, 0, -7, 5, 2, -5, -3,
    -- filter=165 channel=44
    -5, 4, 3, 1, 7, 6, -9, -6, 7,
    -- filter=165 channel=45
    -3, 7, 0, 8, 4, 5, 9, -2, 3,
    -- filter=165 channel=46
    -4, 3, 5, -6, -7, 2, 1, -1, 4,
    -- filter=165 channel=47
    -2, 7, 11, -8, 1, 18, -14, 1, 13,
    -- filter=165 channel=48
    -5, 1, 2, -11, -7, 4, -11, -1, 4,
    -- filter=165 channel=49
    -7, -4, -3, 3, -6, -6, -8, 2, -12,
    -- filter=165 channel=50
    0, 3, 7, 1, 4, 11, -12, -4, 6,
    -- filter=165 channel=51
    5, -5, 7, -2, 6, 7, 7, -3, -2,
    -- filter=165 channel=52
    0, 6, 0, 0, 2, -6, -6, 1, -3,
    -- filter=165 channel=53
    -2, 3, 5, 4, -7, 3, 0, -7, 2,
    -- filter=165 channel=54
    4, 5, -4, 0, -5, 2, 0, 1, 6,
    -- filter=165 channel=55
    -2, 5, -6, -5, -3, 3, -13, -11, -11,
    -- filter=165 channel=56
    -7, 0, -1, 2, -7, 4, -6, 0, 0,
    -- filter=165 channel=57
    5, 1, 5, -3, -9, -3, -6, 4, 0,
    -- filter=165 channel=58
    8, 0, -5, 0, 4, -2, 3, 8, 0,
    -- filter=165 channel=59
    -1, -3, 7, -11, -2, 5, -19, -3, 1,
    -- filter=165 channel=60
    4, 3, -2, 1, 1, -7, -3, -2, 1,
    -- filter=165 channel=61
    -1, -5, 6, -9, -6, 0, -4, -4, -1,
    -- filter=165 channel=62
    1, 4, 0, 1, -2, -5, 0, 0, 3,
    -- filter=165 channel=63
    -2, -3, -10, -3, -5, -3, -6, 0, -4,
    -- filter=165 channel=64
    -5, 0, 3, 0, -2, -1, 1, 1, 2,
    -- filter=165 channel=65
    6, 2, -1, 4, -4, -2, -6, -2, 6,
    -- filter=165 channel=66
    -2, 2, -5, -6, 0, -1, 3, -11, -5,
    -- filter=165 channel=67
    2, 0, -6, 2, 0, -7, -5, -3, -4,
    -- filter=165 channel=68
    1, -6, -5, 0, 4, -2, -3, 3, 3,
    -- filter=165 channel=69
    1, -1, 0, -1, -1, 5, 1, 0, 5,
    -- filter=165 channel=70
    -4, 7, 9, -6, 2, 0, -13, -5, 3,
    -- filter=165 channel=71
    -2, 5, 2, 10, -2, 6, -4, 3, 2,
    -- filter=165 channel=72
    4, 0, 12, -4, 1, 15, -15, -3, 8,
    -- filter=165 channel=73
    3, 5, 3, -6, -1, -8, 0, -10, -1,
    -- filter=165 channel=74
    0, 12, 12, 0, 4, -3, -4, 6, 8,
    -- filter=165 channel=75
    -2, 1, 1, -2, 4, -2, 0, -4, -3,
    -- filter=165 channel=76
    2, -8, 0, -4, 1, 0, -4, -4, 0,
    -- filter=165 channel=77
    -2, -4, 1, -5, 0, 1, -6, 4, -5,
    -- filter=165 channel=78
    -1, 0, 3, 0, 1, 6, 3, 1, 0,
    -- filter=165 channel=79
    0, 1, -1, -10, -14, -8, -17, -17, -9,
    -- filter=165 channel=80
    3, 6, 6, -6, 8, 7, -17, -1, 6,
    -- filter=165 channel=81
    -4, -2, 5, 6, 7, -2, -1, 3, -6,
    -- filter=165 channel=82
    -1, 0, -1, -3, 5, -3, -7, -1, 7,
    -- filter=165 channel=83
    -2, -6, 0, -9, -7, -4, -8, -10, -3,
    -- filter=165 channel=84
    -8, -1, 5, -3, -10, -8, -3, -11, 0,
    -- filter=165 channel=85
    -2, 3, 0, 0, -3, 3, 6, -4, 2,
    -- filter=165 channel=86
    -8, 4, -4, 1, 1, 2, 0, 5, -3,
    -- filter=165 channel=87
    2, 1, -3, 0, 0, 0, 1, -5, -13,
    -- filter=165 channel=88
    1, 3, 3, 0, 2, 9, -6, 0, 4,
    -- filter=165 channel=89
    -6, 8, 2, -2, 0, 9, -16, -8, -2,
    -- filter=165 channel=90
    0, 4, 0, -3, 7, 1, -6, 4, 3,
    -- filter=165 channel=91
    -3, -5, 0, -11, -3, -3, -15, -5, -10,
    -- filter=165 channel=92
    7, 7, 2, -5, -4, 4, -3, 3, -4,
    -- filter=165 channel=93
    -7, -1, 2, -1, 0, 8, -10, -7, 11,
    -- filter=165 channel=94
    7, 0, -4, -3, 2, 0, 3, 1, 0,
    -- filter=165 channel=95
    3, 0, -1, -5, -3, 0, 4, 3, -1,
    -- filter=165 channel=96
    2, 6, 2, -5, 5, 0, -1, -7, -2,
    -- filter=165 channel=97
    0, 0, 5, 5, 7, 5, 2, 10, 8,
    -- filter=165 channel=98
    5, 13, 11, -13, 0, 12, -9, 0, 7,
    -- filter=165 channel=99
    2, 9, 8, -2, 0, 7, -13, -12, 6,
    -- filter=165 channel=100
    -3, 5, 0, 0, -7, -4, 1, 3, -9,
    -- filter=165 channel=101
    1, 0, 5, 5, -8, -5, 4, -1, -2,
    -- filter=165 channel=102
    2, 2, 1, -6, 0, 3, -2, -3, 2,
    -- filter=165 channel=103
    7, 11, 6, 5, 3, 7, -8, 0, 15,
    -- filter=165 channel=104
    -8, -2, 9, -6, -1, 15, -20, -3, 9,
    -- filter=165 channel=105
    0, 4, -10, 1, 3, 3, 6, -1, -2,
    -- filter=165 channel=106
    6, -2, -4, -1, -7, 3, -6, -4, 1,
    -- filter=165 channel=107
    -4, -5, 1, 3, -2, -4, -3, -3, -11,
    -- filter=165 channel=108
    2, 5, -9, -3, -4, -9, 4, 3, -1,
    -- filter=165 channel=109
    1, 0, 11, -11, -9, 5, -11, -5, -1,
    -- filter=165 channel=110
    7, -1, 6, -5, 5, 0, -9, 1, 8,
    -- filter=165 channel=111
    -3, 4, -4, 0, 0, -6, -3, 0, 0,
    -- filter=165 channel=112
    0, 7, 0, 3, 7, 3, -5, -4, 8,
    -- filter=165 channel=113
    0, 10, 3, 5, 6, 15, -3, -6, 8,
    -- filter=165 channel=114
    -4, 1, 4, -7, -8, -5, -6, -18, -11,
    -- filter=165 channel=115
    -6, 1, 5, -1, -3, 1, 6, 0, -1,
    -- filter=165 channel=116
    1, 0, -2, -7, -10, 4, -3, -7, -8,
    -- filter=165 channel=117
    -4, 0, -4, 0, -3, 2, 2, -1, 0,
    -- filter=165 channel=118
    2, -3, -1, -5, 6, -7, -1, -2, 4,
    -- filter=165 channel=119
    -4, 8, -1, 0, 7, 0, -4, 7, 2,
    -- filter=165 channel=120
    -3, 4, 4, -13, -2, 0, -10, 0, 0,
    -- filter=165 channel=121
    -7, -3, 0, -10, -4, 5, -4, -5, 0,
    -- filter=165 channel=122
    -4, 5, 11, -5, 3, 15, -14, -5, 20,
    -- filter=165 channel=123
    1, 2, 5, 0, -3, 0, -7, 4, -1,
    -- filter=165 channel=124
    -7, 0, -5, 1, -1, -3, -3, -4, -6,
    -- filter=165 channel=125
    -4, 1, 8, -16, 0, 11, -7, -4, 4,
    -- filter=165 channel=126
    -1, 6, 0, -9, 1, 8, -3, -4, 1,
    -- filter=165 channel=127
    -7, 4, -5, -7, 2, 0, -3, 1, -6,
    -- filter=166 channel=0
    1, -21, -17, 5, -2, 0, 22, 12, 3,
    -- filter=166 channel=1
    -11, -20, -12, 11, -7, 2, 19, 9, 4,
    -- filter=166 channel=2
    1, 1, 3, -2, -5, -6, -3, 0, 8,
    -- filter=166 channel=3
    5, 7, 7, 0, -5, 8, 0, 0, -4,
    -- filter=166 channel=4
    -1, 0, 10, 0, 3, -4, 5, -5, 0,
    -- filter=166 channel=5
    -9, -16, -11, 10, -9, -12, 24, 4, 6,
    -- filter=166 channel=6
    7, 1, 3, 4, 4, 7, -2, 0, -1,
    -- filter=166 channel=7
    -3, -6, 2, -2, 0, 6, -6, -1, -3,
    -- filter=166 channel=8
    -3, 0, 0, -5, 1, 0, -5, 3, 1,
    -- filter=166 channel=9
    0, -4, 2, -3, -5, 1, 10, 8, 1,
    -- filter=166 channel=10
    6, 9, -4, 0, 8, 2, 1, 2, 2,
    -- filter=166 channel=11
    10, 3, -3, 5, 1, 6, -6, 2, 3,
    -- filter=166 channel=12
    5, 0, 10, -3, 6, 0, -6, -6, 0,
    -- filter=166 channel=13
    7, 12, -1, -3, 3, 2, -4, -2, -5,
    -- filter=166 channel=14
    0, -4, 6, 3, 0, 3, -6, -1, -4,
    -- filter=166 channel=15
    3, 6, 6, 2, 10, 9, -12, -9, 8,
    -- filter=166 channel=16
    3, 0, 3, 5, 0, 0, 12, 0, 0,
    -- filter=166 channel=17
    -1, 3, 1, 3, -3, 1, 0, -1, -1,
    -- filter=166 channel=18
    5, 4, 5, -3, 6, 0, -2, 4, 3,
    -- filter=166 channel=19
    -4, 0, 5, 4, 0, -5, -7, -6, 0,
    -- filter=166 channel=20
    8, 13, -8, -4, 6, 4, -15, 0, 3,
    -- filter=166 channel=21
    -4, 2, -7, -2, 2, 2, -2, 0, 1,
    -- filter=166 channel=22
    6, -7, -6, -6, -1, -1, 5, 0, 6,
    -- filter=166 channel=23
    3, 1, -4, -7, 0, 7, -10, -4, -1,
    -- filter=166 channel=24
    -1, -3, -4, -1, 6, 2, 3, 6, 4,
    -- filter=166 channel=25
    0, -4, 5, 0, 0, -3, 7, 1, 6,
    -- filter=166 channel=26
    4, -9, 0, 2, -7, -5, 11, -4, -7,
    -- filter=166 channel=27
    -5, -8, -3, -11, 1, 0, -4, 4, -1,
    -- filter=166 channel=28
    3, 0, 1, 3, 3, -2, 5, 0, 7,
    -- filter=166 channel=29
    0, 1, -3, -3, -1, 2, -2, -7, 2,
    -- filter=166 channel=30
    3, -4, -5, 3, -1, -1, 12, 9, -2,
    -- filter=166 channel=31
    7, 1, -2, 5, 3, 0, -4, -1, 0,
    -- filter=166 channel=32
    3, 0, -2, 0, 4, -1, 0, 0, -3,
    -- filter=166 channel=33
    0, 0, -4, -3, 4, 0, 8, 0, 5,
    -- filter=166 channel=34
    7, -4, 5, -3, 8, 0, -4, 3, -5,
    -- filter=166 channel=35
    0, 0, -5, 0, 6, 5, 0, 2, -6,
    -- filter=166 channel=36
    0, 7, 8, 1, 1, -6, -3, -1, -2,
    -- filter=166 channel=37
    -11, -13, -7, 5, -3, -2, 16, 8, 1,
    -- filter=166 channel=38
    0, 8, 6, -6, 5, -4, 1, -7, -7,
    -- filter=166 channel=39
    8, -1, -7, -1, 9, 6, -1, -7, -1,
    -- filter=166 channel=40
    4, 2, -2, -5, -1, 8, -12, 2, -2,
    -- filter=166 channel=41
    1, 7, 1, -4, 0, 2, -1, 5, 9,
    -- filter=166 channel=42
    -7, 0, -7, 10, 3, 2, 7, 5, 8,
    -- filter=166 channel=43
    10, 3, 5, 0, 0, 4, -3, 0, 5,
    -- filter=166 channel=44
    0, -11, 0, 12, 0, 0, 6, 5, 0,
    -- filter=166 channel=45
    -6, 0, -9, 6, 1, 5, -5, -2, 3,
    -- filter=166 channel=46
    2, -6, 3, -3, -2, -2, 1, 0, -4,
    -- filter=166 channel=47
    -7, -8, -9, 7, 3, -10, 15, 5, -1,
    -- filter=166 channel=48
    -1, -3, 2, 7, -3, 1, 10, -1, -1,
    -- filter=166 channel=49
    -5, -4, 4, 4, 2, 3, -3, 1, 5,
    -- filter=166 channel=50
    6, -1, 2, -9, -6, -4, 5, -7, 3,
    -- filter=166 channel=51
    -5, 0, -7, -4, 5, -3, -4, -3, 2,
    -- filter=166 channel=52
    7, 1, -4, -1, 3, 3, -11, 2, 0,
    -- filter=166 channel=53
    8, -3, -1, -3, 6, 6, -9, 6, -2,
    -- filter=166 channel=54
    -1, -2, -3, -4, -4, 0, 5, 0, -1,
    -- filter=166 channel=55
    9, 15, -5, -6, 2, 4, -16, -11, 0,
    -- filter=166 channel=56
    -6, -1, 6, 5, 5, -2, 0, -5, -3,
    -- filter=166 channel=57
    1, -4, 0, -2, -2, 3, 0, 0, -2,
    -- filter=166 channel=58
    -5, -13, -7, 12, -3, -2, 10, 5, 6,
    -- filter=166 channel=59
    3, 1, 4, -9, -8, -4, 2, -7, 8,
    -- filter=166 channel=60
    -1, -1, -6, -4, -5, 1, -2, -4, 0,
    -- filter=166 channel=61
    -3, 6, 3, 5, 5, 6, -1, -4, 6,
    -- filter=166 channel=62
    -1, -6, -4, 2, 0, 4, 4, 5, 7,
    -- filter=166 channel=63
    -2, -4, -1, 8, -1, -9, 10, -2, -4,
    -- filter=166 channel=64
    6, 6, 4, -4, 8, -6, -1, 0, 0,
    -- filter=166 channel=65
    -2, -4, -4, 2, -5, -3, -6, -4, 3,
    -- filter=166 channel=66
    0, 8, 0, 2, -4, -3, -1, 0, 2,
    -- filter=166 channel=67
    1, 3, 4, -6, -3, -6, -1, -5, 5,
    -- filter=166 channel=68
    5, 1, 7, -6, 2, 0, -3, -7, 0,
    -- filter=166 channel=69
    4, 0, -4, 0, -2, -3, -4, 0, 7,
    -- filter=166 channel=70
    -5, 8, 4, -9, 0, -1, -4, 0, 0,
    -- filter=166 channel=71
    0, -3, -2, 0, -6, -5, -4, -4, 0,
    -- filter=166 channel=72
    -2, 13, -5, -5, 5, 3, -7, -4, -6,
    -- filter=166 channel=73
    5, 0, -1, -11, -3, -3, -8, 3, 0,
    -- filter=166 channel=74
    -4, 0, 1, -4, 0, -4, -2, 6, 5,
    -- filter=166 channel=75
    -7, -15, -2, 8, -9, -9, 23, 15, -3,
    -- filter=166 channel=76
    0, 13, 1, 0, 5, 0, -16, 0, 2,
    -- filter=166 channel=77
    -4, -3, -3, -3, -2, -3, -3, -4, 0,
    -- filter=166 channel=78
    8, 0, -5, 2, 4, 0, 9, 8, 5,
    -- filter=166 channel=79
    1, -3, -4, -12, 2, 11, -2, -4, -2,
    -- filter=166 channel=80
    4, 7, -2, 0, -2, -12, 0, -3, 3,
    -- filter=166 channel=81
    -7, -6, 2, -5, 6, -2, 4, -6, 2,
    -- filter=166 channel=82
    3, -3, 0, 7, 0, 3, -5, 2, 0,
    -- filter=166 channel=83
    -7, 0, -2, -6, -4, 0, 8, -6, -3,
    -- filter=166 channel=84
    0, -5, -3, -9, -1, 8, -1, -7, -2,
    -- filter=166 channel=85
    -6, 1, 6, 0, 6, -5, 3, -4, 5,
    -- filter=166 channel=86
    3, -4, -3, -2, 6, 5, 8, -1, 3,
    -- filter=166 channel=87
    6, -1, 4, 4, 3, -2, -10, 0, 0,
    -- filter=166 channel=88
    5, 2, -5, -4, 0, -2, 3, -4, 1,
    -- filter=166 channel=89
    10, 14, 0, -9, 1, 3, -12, -12, 2,
    -- filter=166 channel=90
    6, 0, 0, 4, 11, 5, -1, -6, -6,
    -- filter=166 channel=91
    3, 3, 4, -12, 7, 7, -9, 1, 3,
    -- filter=166 channel=92
    0, 0, -3, 4, 0, 7, -4, 4, 3,
    -- filter=166 channel=93
    -2, -8, 0, 13, -3, -11, 8, 7, 2,
    -- filter=166 channel=94
    2, 3, -3, 2, 0, 5, -4, 0, -4,
    -- filter=166 channel=95
    -1, 8, -6, 0, 5, 0, -5, 4, 2,
    -- filter=166 channel=96
    -4, -5, -6, -4, -2, -2, 6, 1, -3,
    -- filter=166 channel=97
    5, -4, 0, -1, -1, -3, 7, 4, 1,
    -- filter=166 channel=98
    -3, -1, -10, -3, -7, -4, 4, -3, 1,
    -- filter=166 channel=99
    12, 5, 6, -7, 8, -5, -8, 3, -2,
    -- filter=166 channel=100
    6, 7, 2, 3, -4, -3, -3, 7, 0,
    -- filter=166 channel=101
    3, 3, 0, 2, -3, -2, 1, -4, 0,
    -- filter=166 channel=102
    -5, -3, 0, 6, -2, 2, 0, 5, -6,
    -- filter=166 channel=103
    -2, 0, -8, 11, -5, 1, 17, 0, -6,
    -- filter=166 channel=104
    1, 5, 5, -1, -5, -7, 6, -5, 3,
    -- filter=166 channel=105
    5, 8, 2, 1, 1, 0, 1, -3, -2,
    -- filter=166 channel=106
    3, 2, -5, 5, -1, -5, -2, -6, 0,
    -- filter=166 channel=107
    9, 4, -3, 1, 3, 2, 0, 7, 2,
    -- filter=166 channel=108
    6, -8, -4, 0, 5, 3, 7, 2, 8,
    -- filter=166 channel=109
    -10, -4, -5, -11, -6, -1, -5, -6, 4,
    -- filter=166 channel=110
    1, 3, -6, 4, 1, -2, -6, -6, -1,
    -- filter=166 channel=111
    -4, -5, -1, -4, 1, -1, 5, -3, 7,
    -- filter=166 channel=112
    -5, 1, -4, -4, 4, -2, 8, 8, -3,
    -- filter=166 channel=113
    5, 8, 1, -6, 1, -6, -7, -6, 1,
    -- filter=166 channel=114
    -7, -14, -11, -7, -6, -4, 16, 0, 8,
    -- filter=166 channel=115
    2, -6, 3, 0, 0, 4, -6, 6, -5,
    -- filter=166 channel=116
    -4, 9, -4, -4, -2, -1, 0, -6, 4,
    -- filter=166 channel=117
    -6, 0, 6, 1, 0, 0, -1, 5, -6,
    -- filter=166 channel=118
    -6, -6, 4, -6, 3, 0, -7, 0, 0,
    -- filter=166 channel=119
    2, -2, 4, 1, 2, 0, -6, -4, 5,
    -- filter=166 channel=120
    6, 2, -2, -12, -6, 2, -14, -7, 5,
    -- filter=166 channel=121
    7, 0, 6, -3, 5, 0, 5, -1, 0,
    -- filter=166 channel=122
    -4, -3, 0, 16, 3, -2, 9, 0, 0,
    -- filter=166 channel=123
    3, 1, 0, 0, 6, -2, -2, 7, 0,
    -- filter=166 channel=124
    -1, -3, -5, 1, 4, 2, -5, -2, 3,
    -- filter=166 channel=125
    -2, 9, -3, -6, -2, 2, -1, 0, 0,
    -- filter=166 channel=126
    -5, 9, 7, -1, -6, 6, 3, -8, -4,
    -- filter=166 channel=127
    -2, -3, -1, 3, 3, 6, -1, 3, 4,
    -- filter=167 channel=0
    9, 4, -8, 6, -4, -3, 10, -9, -4,
    -- filter=167 channel=1
    6, 3, 0, 4, 4, -10, 2, -12, -15,
    -- filter=167 channel=2
    -7, 7, 3, -2, 2, -5, 6, 2, -2,
    -- filter=167 channel=3
    2, -14, -12, -8, -14, -11, 3, -4, 3,
    -- filter=167 channel=4
    -13, 0, -6, -11, -12, -7, 4, -15, -3,
    -- filter=167 channel=5
    26, 13, 9, 17, 6, -8, 15, -5, -6,
    -- filter=167 channel=6
    8, 3, 5, 10, -2, 7, 7, 1, 10,
    -- filter=167 channel=7
    -6, -1, -1, 0, 7, 3, 6, -4, -2,
    -- filter=167 channel=8
    -5, 1, -9, 7, 0, -8, 8, -10, 0,
    -- filter=167 channel=9
    6, 2, 1, -3, 9, 1, 7, 1, 0,
    -- filter=167 channel=10
    -14, -12, -3, -13, 9, 7, -2, 2, 4,
    -- filter=167 channel=11
    -8, -11, 8, -6, 11, 12, -3, -4, 14,
    -- filter=167 channel=12
    0, 0, 0, -8, -9, -1, -1, -5, 0,
    -- filter=167 channel=13
    -19, -16, -11, -20, 9, 12, -17, 3, 5,
    -- filter=167 channel=14
    -5, -3, 2, -5, -3, -1, -3, 1, -1,
    -- filter=167 channel=15
    -16, -14, -2, -11, 14, 11, 2, 13, 13,
    -- filter=167 channel=16
    3, 1, 0, 0, 3, -10, -2, -5, -3,
    -- filter=167 channel=17
    0, 6, -6, 6, -5, 0, -1, 2, 6,
    -- filter=167 channel=18
    -12, -24, -7, -19, 22, 26, -2, 9, 1,
    -- filter=167 channel=19
    -1, -4, -5, -4, 0, 2, 3, 2, 2,
    -- filter=167 channel=20
    -5, -5, 0, 1, 15, 18, 5, -1, 16,
    -- filter=167 channel=21
    7, 12, 1, 2, -3, -10, 2, 3, -3,
    -- filter=167 channel=22
    4, -5, -13, 3, -3, 1, -2, -5, 0,
    -- filter=167 channel=23
    -15, -34, -18, 5, 14, 2, 0, 7, 7,
    -- filter=167 channel=24
    2, -1, -6, 7, 3, -2, -3, 2, -3,
    -- filter=167 channel=25
    -12, -1, -10, -18, 22, 12, -3, 10, 8,
    -- filter=167 channel=26
    14, 13, -4, 9, 7, -5, 5, -7, -4,
    -- filter=167 channel=27
    -21, 0, 0, -2, 35, 10, 1, 7, 7,
    -- filter=167 channel=28
    5, 6, 4, -6, 1, 0, 3, -2, 2,
    -- filter=167 channel=29
    -8, 1, 2, -3, 14, 22, 2, 5, 15,
    -- filter=167 channel=30
    6, 15, 3, 1, 13, 3, 7, 2, 0,
    -- filter=167 channel=31
    -4, 3, -1, 0, 11, 5, 2, 1, 6,
    -- filter=167 channel=32
    -18, -9, -7, -6, 17, 18, -6, 9, -1,
    -- filter=167 channel=33
    -3, -24, -11, -18, 17, 13, -5, 12, 12,
    -- filter=167 channel=34
    -4, -15, -17, 9, -3, -11, 1, -1, -10,
    -- filter=167 channel=35
    -4, 0, -6, 0, 3, 0, 0, -1, 3,
    -- filter=167 channel=36
    0, -4, 4, 6, -2, -5, -7, -10, -5,
    -- filter=167 channel=37
    11, 7, -2, 8, 5, -9, 6, -4, -8,
    -- filter=167 channel=38
    4, -8, -7, -10, 5, 0, -2, 2, 2,
    -- filter=167 channel=39
    -8, 3, -2, -3, 4, 10, 5, 3, 8,
    -- filter=167 channel=40
    -10, -12, -8, 0, -1, 4, -5, -3, 6,
    -- filter=167 channel=41
    -9, -19, -13, -28, -14, 2, -26, -9, -9,
    -- filter=167 channel=42
    2, 1, 8, 0, 10, 1, 6, -6, 5,
    -- filter=167 channel=43
    -3, -17, -10, 2, -3, 0, 6, -2, 9,
    -- filter=167 channel=44
    11, 5, 0, 1, 0, -9, 0, -1, -8,
    -- filter=167 channel=45
    3, 8, 1, 10, 7, -4, 8, -4, -1,
    -- filter=167 channel=46
    -2, -2, 0, -1, -4, -5, -2, -3, -10,
    -- filter=167 channel=47
    9, 11, -4, 4, -5, -8, -3, 0, -9,
    -- filter=167 channel=48
    -8, 6, 0, -6, 21, 5, 5, 0, -8,
    -- filter=167 channel=49
    -10, 1, -2, 5, 13, 14, -1, -9, 7,
    -- filter=167 channel=50
    -9, -5, 0, 4, 18, 4, 0, 0, -2,
    -- filter=167 channel=51
    4, -5, 5, -1, -2, 5, 5, 6, 7,
    -- filter=167 channel=52
    0, -5, -11, 5, -8, -8, 6, -11, -4,
    -- filter=167 channel=53
    -2, -11, -1, 2, 10, 9, -5, -1, 0,
    -- filter=167 channel=54
    1, 7, -3, 0, -2, 5, -7, 2, 5,
    -- filter=167 channel=55
    -14, -14, -6, -4, 23, 11, -4, 13, 7,
    -- filter=167 channel=56
    5, 1, 0, 12, 1, -10, 2, -6, -2,
    -- filter=167 channel=57
    -10, -2, -3, -2, -1, 0, -5, 3, 5,
    -- filter=167 channel=58
    15, 12, -1, 15, -3, -3, 4, -4, 0,
    -- filter=167 channel=59
    -10, 1, -6, -21, 13, 7, -12, 11, -1,
    -- filter=167 channel=60
    -6, -3, -5, -6, -4, -3, 1, 2, 1,
    -- filter=167 channel=61
    -9, -4, 5, 2, -8, -3, 1, -1, -1,
    -- filter=167 channel=62
    -6, 3, -1, 0, 1, -4, 0, 3, -4,
    -- filter=167 channel=63
    15, 11, -2, 16, 0, 3, 14, 1, -4,
    -- filter=167 channel=64
    -5, 0, -5, 0, 4, -5, 5, -7, 0,
    -- filter=167 channel=65
    -5, 2, 0, 0, 0, -2, -1, -1, 6,
    -- filter=167 channel=66
    -1, -7, -2, -12, -6, 2, -9, -6, -4,
    -- filter=167 channel=67
    5, 2, -6, 9, -2, -6, 0, -3, -8,
    -- filter=167 channel=68
    -7, -6, 0, -10, -6, 5, -8, 1, -7,
    -- filter=167 channel=69
    1, -6, 0, 1, 2, 1, -7, 6, 3,
    -- filter=167 channel=70
    -20, -12, -11, -6, 6, 7, 0, -5, -5,
    -- filter=167 channel=71
    3, -16, -14, -11, -3, -8, 3, -3, -6,
    -- filter=167 channel=72
    -16, 2, 3, -5, 21, 14, -1, 8, 8,
    -- filter=167 channel=73
    -18, -4, 0, -8, 6, 12, 0, -8, -3,
    -- filter=167 channel=74
    0, 3, -6, 19, 8, -9, 0, 0, -2,
    -- filter=167 channel=75
    7, -4, -9, -1, -4, -8, 0, 5, 0,
    -- filter=167 channel=76
    -6, -17, 6, -1, 2, 8, -1, -2, 14,
    -- filter=167 channel=77
    0, -4, 2, -6, -7, -5, 3, 3, -3,
    -- filter=167 channel=78
    3, 4, 4, 13, 3, -3, 13, 0, 1,
    -- filter=167 channel=79
    -20, -24, -15, -16, 30, 20, -9, 11, 5,
    -- filter=167 channel=80
    -9, 10, 2, -18, 19, 9, -14, 10, 13,
    -- filter=167 channel=81
    3, -2, -6, 2, 1, 4, -2, 0, 7,
    -- filter=167 channel=82
    -6, -9, -10, -5, 1, -5, -5, -3, 0,
    -- filter=167 channel=83
    0, 13, -1, 5, 5, -1, -5, 2, 5,
    -- filter=167 channel=84
    -8, 3, -2, 3, 13, 4, -7, 1, 0,
    -- filter=167 channel=85
    0, -3, 4, 0, 3, -2, 4, 0, -4,
    -- filter=167 channel=86
    -1, -2, 0, 0, -6, -3, 6, -10, -7,
    -- filter=167 channel=87
    -3, -3, -1, 7, 4, 4, 2, 1, 1,
    -- filter=167 channel=88
    -5, 1, 1, 4, -4, -12, -4, -2, -6,
    -- filter=167 channel=89
    -28, -15, -13, -26, 10, 9, -13, 11, 8,
    -- filter=167 channel=90
    -5, -5, -13, 11, -12, -10, 0, 3, -6,
    -- filter=167 channel=91
    -19, -7, 0, -2, 21, 13, 0, -1, 1,
    -- filter=167 channel=92
    -9, -10, -11, -6, -11, 3, 5, -2, 1,
    -- filter=167 channel=93
    4, 9, 6, 8, 6, -15, 5, -2, -5,
    -- filter=167 channel=94
    2, 2, -1, -6, -1, 2, 0, -7, 0,
    -- filter=167 channel=95
    5, 0, -7, 0, 5, -3, -4, -1, -1,
    -- filter=167 channel=96
    0, 6, 6, -4, 1, 4, -9, 0, 6,
    -- filter=167 channel=97
    -10, -15, -4, -2, -10, -1, -7, 7, -4,
    -- filter=167 channel=98
    -11, -11, 2, 0, 27, 16, -7, 7, 9,
    -- filter=167 channel=99
    -17, -9, -1, 4, 13, -2, 8, 0, 0,
    -- filter=167 channel=100
    -7, -3, 2, -3, -10, -2, 9, -3, -11,
    -- filter=167 channel=101
    0, 0, -6, -4, -7, 2, -6, -12, -1,
    -- filter=167 channel=102
    -6, 6, 1, -5, -2, -2, 4, -1, 0,
    -- filter=167 channel=103
    4, -8, -8, -1, 0, -14, -5, 9, 0,
    -- filter=167 channel=104
    -8, 3, 4, -4, 13, 6, 1, 8, -1,
    -- filter=167 channel=105
    -7, 0, -1, 3, 5, 11, 10, -2, 10,
    -- filter=167 channel=106
    -7, -3, -6, -5, -3, 7, -4, 2, -6,
    -- filter=167 channel=107
    0, -7, 0, 3, 8, 1, 9, -1, 11,
    -- filter=167 channel=108
    0, 1, -5, -10, -5, -3, -8, 1, 2,
    -- filter=167 channel=109
    -17, -6, 1, -2, 30, 11, -5, 4, 8,
    -- filter=167 channel=110
    -8, -13, -14, -9, 9, 4, -3, 8, 3,
    -- filter=167 channel=111
    1, -2, -1, 1, 2, 3, -3, -1, -7,
    -- filter=167 channel=112
    3, 6, -6, 9, 10, 1, 3, 9, -2,
    -- filter=167 channel=113
    -15, -23, -13, -8, 7, -4, -8, 6, 6,
    -- filter=167 channel=114
    -10, -7, -6, 3, 25, 10, 0, -2, -2,
    -- filter=167 channel=115
    0, -5, 7, -6, 6, 2, 3, -3, -2,
    -- filter=167 channel=116
    -14, 6, -1, -17, 23, 9, -12, 5, 1,
    -- filter=167 channel=117
    -3, 3, 1, -9, -1, 8, -8, 6, -1,
    -- filter=167 channel=118
    1, -6, 0, -2, 1, 0, -4, 5, -3,
    -- filter=167 channel=119
    1, -13, -5, 20, -11, -6, 13, 0, 0,
    -- filter=167 channel=120
    -10, 4, -6, 19, 23, 9, 15, 6, -1,
    -- filter=167 channel=121
    -3, -11, -8, -3, -7, 2, -4, 3, -3,
    -- filter=167 channel=122
    6, 9, -5, 3, -6, -23, -5, -2, -5,
    -- filter=167 channel=123
    1, -14, -5, 2, 0, -12, 0, 0, -1,
    -- filter=167 channel=124
    0, -4, 2, 9, 7, 5, 7, -4, 5,
    -- filter=167 channel=125
    -16, 9, 3, -12, 29, 15, -6, 0, 3,
    -- filter=167 channel=126
    -16, -21, -6, -9, -3, -1, -1, 2, 8,
    -- filter=167 channel=127
    2, -4, -8, -1, -6, 2, -8, 2, 5,
    -- filter=168 channel=0
    -1, -7, -10, -2, -9, -10, 6, 13, 0,
    -- filter=168 channel=1
    -8, -10, -7, 0, 2, 1, -8, 17, 16,
    -- filter=168 channel=2
    5, 0, -3, 8, 1, 8, -2, -4, 6,
    -- filter=168 channel=3
    -4, 0, 11, 1, 2, 0, 13, 8, 2,
    -- filter=168 channel=4
    4, 0, 6, 5, 17, 16, 0, 5, 19,
    -- filter=168 channel=5
    0, -4, -2, -3, -3, -5, 8, 5, -2,
    -- filter=168 channel=6
    7, 0, 8, 7, -5, 5, 3, -8, -9,
    -- filter=168 channel=7
    0, 5, 7, -2, -3, 1, -5, -7, 1,
    -- filter=168 channel=8
    1, -7, 4, -1, 0, 3, -4, 3, 3,
    -- filter=168 channel=9
    3, -6, 3, 8, -1, 1, 6, 8, 0,
    -- filter=168 channel=10
    5, 1, -4, -3, -1, -14, 8, 9, 2,
    -- filter=168 channel=11
    7, 12, 17, -5, -1, -4, -2, -3, -13,
    -- filter=168 channel=12
    7, 0, 4, -7, -3, 0, -2, 0, 4,
    -- filter=168 channel=13
    -3, -1, -1, 0, 2, -3, -7, 10, -2,
    -- filter=168 channel=14
    -4, 7, 2, -3, -6, -1, 2, 6, 2,
    -- filter=168 channel=15
    9, 3, 17, 2, -13, -8, 2, -2, 1,
    -- filter=168 channel=16
    -7, -11, -3, -7, 0, 0, 1, 7, 4,
    -- filter=168 channel=17
    -1, 1, 1, -1, 0, 1, 3, 5, -1,
    -- filter=168 channel=18
    3, 0, 8, 8, -10, -8, 0, -4, 4,
    -- filter=168 channel=19
    6, 0, -4, -7, 6, -6, 0, 6, 0,
    -- filter=168 channel=20
    4, 10, 24, -12, -17, -8, -12, -8, -17,
    -- filter=168 channel=21
    -11, -19, -12, 5, 1, -6, -1, 8, 0,
    -- filter=168 channel=22
    -5, 6, 1, 3, -3, 0, 6, 0, 2,
    -- filter=168 channel=23
    -2, -2, 19, -10, -24, -17, 17, 6, -16,
    -- filter=168 channel=24
    -4, -1, -5, -2, 0, 6, -3, -1, -2,
    -- filter=168 channel=25
    -10, -5, -1, 10, 9, -18, 4, 27, 16,
    -- filter=168 channel=26
    -7, -7, -14, -4, -3, 0, 0, 0, -1,
    -- filter=168 channel=27
    -1, -5, -5, 7, -3, -25, 15, 30, 1,
    -- filter=168 channel=28
    1, -3, 6, 3, -2, -6, 4, -6, 7,
    -- filter=168 channel=29
    3, 9, 11, 0, 0, -4, -6, -15, 0,
    -- filter=168 channel=30
    -3, -15, 0, 4, -2, 0, -1, 6, 1,
    -- filter=168 channel=31
    -5, -13, -5, 0, -15, -15, 14, 24, 0,
    -- filter=168 channel=32
    -6, 3, 5, 3, -2, -18, -6, 18, -2,
    -- filter=168 channel=33
    -14, -9, 0, 2, -6, -13, 7, 16, -5,
    -- filter=168 channel=34
    -3, -5, 0, 0, -1, -1, 12, -1, -9,
    -- filter=168 channel=35
    0, 5, -4, 0, -4, 6, 2, -3, 5,
    -- filter=168 channel=36
    5, -2, -2, -6, -5, -1, -1, -6, -1,
    -- filter=168 channel=37
    -15, -13, -16, 2, 0, 4, -5, 1, 10,
    -- filter=168 channel=38
    -6, -6, 6, -2, -12, -3, 13, 3, -5,
    -- filter=168 channel=39
    3, -1, 13, 0, -9, 5, -9, -11, -10,
    -- filter=168 channel=40
    6, 0, 11, -2, -5, -4, -3, 1, -15,
    -- filter=168 channel=41
    12, 4, -4, 0, 13, -2, -10, -3, 6,
    -- filter=168 channel=42
    0, -7, 2, 4, 9, 7, 8, 11, 0,
    -- filter=168 channel=43
    -7, 7, 10, 0, -5, 5, 3, -4, -7,
    -- filter=168 channel=44
    -5, -6, -1, 2, 0, -3, 14, 15, 1,
    -- filter=168 channel=45
    2, 2, 4, 1, 4, 2, -9, 1, -6,
    -- filter=168 channel=46
    -4, 5, -6, 4, -5, 5, 0, 3, -1,
    -- filter=168 channel=47
    -10, -18, -15, 5, -1, -8, 14, 10, 3,
    -- filter=168 channel=48
    -7, -21, -14, 16, 3, -10, 10, 19, 14,
    -- filter=168 channel=49
    -5, 4, -3, 4, 4, 0, -9, 1, 3,
    -- filter=168 channel=50
    2, -11, 2, -3, -1, -15, -2, 18, 3,
    -- filter=168 channel=51
    -6, -2, 0, 7, -3, -7, 1, -2, 7,
    -- filter=168 channel=52
    -3, 8, 3, 3, -10, 0, -1, -1, -9,
    -- filter=168 channel=53
    9, -1, 10, 0, -10, 4, 2, -5, -10,
    -- filter=168 channel=54
    -5, 0, 0, 0, 2, 4, 0, 0, 4,
    -- filter=168 channel=55
    4, 14, 11, 3, -10, -15, -2, -5, -3,
    -- filter=168 channel=56
    -3, 3, -3, 7, -9, -3, -4, 0, -3,
    -- filter=168 channel=57
    0, 4, 3, 2, 8, 10, -6, 5, 8,
    -- filter=168 channel=58
    1, 0, -8, -4, -4, -3, 6, 2, -4,
    -- filter=168 channel=59
    1, -14, -16, 6, 0, -12, 7, 14, 11,
    -- filter=168 channel=60
    5, 2, 3, -5, 5, 1, -4, -7, -6,
    -- filter=168 channel=61
    1, -7, -5, 6, -5, -8, 1, -6, -3,
    -- filter=168 channel=62
    -2, 3, 5, 6, -5, -2, 7, -7, -4,
    -- filter=168 channel=63
    -8, -8, -11, -5, 0, 6, -5, 5, 3,
    -- filter=168 channel=64
    6, -4, 6, -4, -3, 0, 2, -7, -7,
    -- filter=168 channel=65
    3, -7, -3, -3, 2, 5, 0, 5, -3,
    -- filter=168 channel=66
    -2, -4, 5, 6, 9, 3, 3, 7, 1,
    -- filter=168 channel=67
    -4, 5, -1, -6, -2, -5, -6, -6, 3,
    -- filter=168 channel=68
    3, -5, -5, 3, 5, 0, -8, 3, 0,
    -- filter=168 channel=69
    0, 0, -2, -2, 2, -5, 6, 3, 6,
    -- filter=168 channel=70
    -11, 2, 1, 8, -8, -7, 3, 10, 0,
    -- filter=168 channel=71
    -1, -5, 4, 2, -6, -2, 3, -2, 4,
    -- filter=168 channel=72
    3, -6, 2, 4, 1, -17, 0, 10, 0,
    -- filter=168 channel=73
    3, 7, 3, 9, 5, 2, 3, 2, 7,
    -- filter=168 channel=74
    -7, -6, 0, 1, -5, -12, 3, 5, -1,
    -- filter=168 channel=75
    -9, -2, -4, -3, -2, -3, 5, 20, 11,
    -- filter=168 channel=76
    10, 11, 19, -14, -8, -6, -9, -12, -9,
    -- filter=168 channel=77
    5, 6, 1, -6, 1, 6, 0, 0, 5,
    -- filter=168 channel=78
    3, -3, -6, -3, 0, 0, -2, 5, 4,
    -- filter=168 channel=79
    -4, -7, -1, 5, -15, -22, 5, 12, 3,
    -- filter=168 channel=80
    -11, -20, -15, 9, -1, -13, 18, 29, 7,
    -- filter=168 channel=81
    0, -6, -7, -3, -1, -4, 6, 5, 0,
    -- filter=168 channel=82
    -5, -6, 4, 3, -6, 3, -3, -1, -5,
    -- filter=168 channel=83
    -1, -8, -10, 3, 5, -3, 0, 10, 0,
    -- filter=168 channel=84
    4, 0, 7, 0, -3, -2, 0, 0, -1,
    -- filter=168 channel=85
    0, 6, -2, 3, -7, 2, -6, 2, 5,
    -- filter=168 channel=86
    -1, 3, 7, -5, 1, -3, -7, 4, -5,
    -- filter=168 channel=87
    3, 9, 13, -4, -8, -4, -1, -8, -11,
    -- filter=168 channel=88
    0, -1, -2, -6, -10, 1, 2, -1, 2,
    -- filter=168 channel=89
    5, -5, -1, -1, -12, -15, 10, 4, 8,
    -- filter=168 channel=90
    -5, -5, 6, -5, -17, -2, 1, -3, -7,
    -- filter=168 channel=91
    -3, -2, 0, 3, 3, 0, -5, 6, 11,
    -- filter=168 channel=92
    2, 9, 1, -1, -6, 0, 12, -3, 4,
    -- filter=168 channel=93
    -17, -22, -12, 12, 8, -5, 9, 19, 21,
    -- filter=168 channel=94
    -7, -4, 2, 7, 2, 2, 4, -6, -5,
    -- filter=168 channel=95
    5, 3, -6, 3, -1, 3, 0, -6, -6,
    -- filter=168 channel=96
    1, 0, 0, 6, -1, -3, 0, 7, 2,
    -- filter=168 channel=97
    -4, 4, -1, -10, -7, -2, 3, 0, -9,
    -- filter=168 channel=98
    -7, -4, -8, 4, 0, -14, 7, 29, 0,
    -- filter=168 channel=99
    -5, -6, 6, 0, -12, -4, 12, 12, -4,
    -- filter=168 channel=100
    7, 4, -2, 0, -3, 6, 2, -3, 1,
    -- filter=168 channel=101
    -1, 4, -2, 2, 8, 3, 0, 1, 11,
    -- filter=168 channel=102
    6, -2, 1, -3, 0, -2, 1, 6, 0,
    -- filter=168 channel=103
    0, -17, 3, -2, -9, -9, 12, 24, 3,
    -- filter=168 channel=104
    -9, -19, -1, 4, 0, -10, 11, 15, 7,
    -- filter=168 channel=105
    1, 4, 19, -9, -4, 4, -10, -7, -7,
    -- filter=168 channel=106
    8, 0, 6, -6, 1, -2, -3, -8, -4,
    -- filter=168 channel=107
    3, 8, 20, -8, -4, 5, 3, -10, -17,
    -- filter=168 channel=108
    8, 1, 3, 0, 9, 0, 4, -8, 8,
    -- filter=168 channel=109
    -2, -14, 0, 15, -2, -12, 9, 20, 8,
    -- filter=168 channel=110
    1, 2, 8, 1, -1, 1, 4, 2, 0,
    -- filter=168 channel=111
    6, 1, 2, -5, 0, 2, -1, -1, 3,
    -- filter=168 channel=112
    0, -12, -4, 2, -7, -14, 3, 12, -9,
    -- filter=168 channel=113
    -7, -3, -1, -5, -14, -2, 17, 17, -5,
    -- filter=168 channel=114
    5, 5, 0, 7, 1, -15, -4, 4, -4,
    -- filter=168 channel=115
    -1, 1, 1, -8, 0, 0, -3, -4, 2,
    -- filter=168 channel=116
    3, -11, -9, 13, 7, -1, 1, 16, 14,
    -- filter=168 channel=117
    0, -1, 0, 5, 1, 1, -6, 4, -2,
    -- filter=168 channel=118
    0, 7, 0, 3, -2, 5, 1, 3, 1,
    -- filter=168 channel=119
    7, -6, 7, -3, -11, 3, 8, 2, -2,
    -- filter=168 channel=120
    0, -8, 10, 1, -6, -4, 1, 3, -2,
    -- filter=168 channel=121
    -5, 4, 3, -1, -1, -4, -2, -1, 2,
    -- filter=168 channel=122
    -11, -32, -16, 0, -3, -4, 8, 12, 12,
    -- filter=168 channel=123
    7, 0, 8, 1, -1, -4, 5, -1, 3,
    -- filter=168 channel=124
    1, 0, 13, -3, 1, 1, -4, -1, 0,
    -- filter=168 channel=125
    -9, -1, -8, 13, 0, -6, -4, 17, 7,
    -- filter=168 channel=126
    -5, -6, -4, 0, -2, -5, 0, -2, 3,
    -- filter=168 channel=127
    4, 3, -1, 1, 6, -5, -2, -4, -2,
    -- filter=169 channel=0
    -3, -1, 5, -18, -7, 8, -5, 0, 10,
    -- filter=169 channel=1
    -10, -6, 5, -7, 0, 10, -4, 5, 12,
    -- filter=169 channel=2
    -4, 1, -3, -6, -1, -10, 7, -7, 6,
    -- filter=169 channel=3
    -9, -12, -1, -4, -2, -4, 6, -6, -4,
    -- filter=169 channel=4
    -6, -3, -1, 3, -9, -8, 3, -3, 1,
    -- filter=169 channel=5
    -9, -8, -5, -6, -1, 2, 1, 1, -2,
    -- filter=169 channel=6
    -2, -5, 0, 3, 7, -4, -1, 2, 3,
    -- filter=169 channel=7
    0, -4, 1, 2, -1, 0, 3, 2, 0,
    -- filter=169 channel=8
    -2, 12, 1, -3, 1, -2, -5, 7, 6,
    -- filter=169 channel=9
    -6, 4, 4, -4, 6, 3, 1, 4, -8,
    -- filter=169 channel=10
    0, 3, 1, -6, 7, 7, 3, 5, -11,
    -- filter=169 channel=11
    8, -2, -10, 0, -5, -1, 1, -5, -8,
    -- filter=169 channel=12
    6, 4, 6, 4, 11, 10, 0, 6, 7,
    -- filter=169 channel=13
    6, -2, 0, 6, 2, -3, 3, 9, -2,
    -- filter=169 channel=14
    5, -2, 7, -2, 5, -7, 0, 0, 5,
    -- filter=169 channel=15
    -3, -6, -8, 2, -3, 0, 0, 10, -1,
    -- filter=169 channel=16
    4, -4, 2, -2, -3, 0, 5, 5, 6,
    -- filter=169 channel=17
    -2, 1, 3, -5, 2, 7, 3, 6, -4,
    -- filter=169 channel=18
    -8, -6, -2, 0, 4, -4, 3, 6, 5,
    -- filter=169 channel=19
    -4, -4, -4, 6, 1, 5, 5, -7, 1,
    -- filter=169 channel=20
    1, 0, -8, 4, -1, -14, 0, -5, 1,
    -- filter=169 channel=21
    -4, 1, 0, 0, -3, 6, 0, 6, 0,
    -- filter=169 channel=22
    -5, 0, -2, -9, 7, 0, -5, 1, 0,
    -- filter=169 channel=23
    -8, 13, 3, -20, 9, -9, 2, 1, -7,
    -- filter=169 channel=24
    3, -5, -7, 3, 0, -4, 1, -6, 1,
    -- filter=169 channel=25
    -3, 3, 9, -15, 5, 0, 0, 12, -5,
    -- filter=169 channel=26
    -5, 7, 5, 4, 6, 0, 0, 0, -3,
    -- filter=169 channel=27
    -15, 10, 9, -18, 20, 5, -5, 3, -3,
    -- filter=169 channel=28
    0, 2, 0, -4, 2, 0, 4, -5, 6,
    -- filter=169 channel=29
    9, -1, 0, 1, -4, -1, 0, 7, 2,
    -- filter=169 channel=30
    -5, -3, 6, -15, 10, 5, -2, 3, 6,
    -- filter=169 channel=31
    -17, -2, 6, -24, 7, -4, -8, 4, -10,
    -- filter=169 channel=32
    -12, -2, 9, -12, 6, -5, -8, 14, 2,
    -- filter=169 channel=33
    -12, 3, 9, -14, 12, 11, 2, 2, 2,
    -- filter=169 channel=34
    -1, 19, -1, -4, 14, -3, 2, 0, 4,
    -- filter=169 channel=35
    -6, -3, 2, -3, -6, 0, 4, 6, 3,
    -- filter=169 channel=36
    9, 4, -4, 3, -2, 0, -4, 3, -4,
    -- filter=169 channel=37
    0, -5, 0, -8, -2, 13, 2, 0, 9,
    -- filter=169 channel=38
    -7, -3, 0, -5, 9, -4, 0, 3, -1,
    -- filter=169 channel=39
    3, 1, -7, 6, 1, -8, -2, 0, -5,
    -- filter=169 channel=40
    -5, 4, 0, 3, -1, -4, 4, 4, -5,
    -- filter=169 channel=41
    14, 5, 1, 1, 10, 12, 8, 12, 3,
    -- filter=169 channel=42
    -3, -12, 8, -10, 0, 6, 5, -10, -5,
    -- filter=169 channel=43
    -4, 0, -8, -11, 4, 7, -1, -4, -8,
    -- filter=169 channel=44
    -14, -4, 2, -8, 4, 9, -4, 0, 2,
    -- filter=169 channel=45
    -4, -7, -7, 4, -1, 0, -1, -4, -5,
    -- filter=169 channel=46
    -3, 2, -2, 0, 3, -2, 5, -5, 1,
    -- filter=169 channel=47
    3, 1, 14, -11, -2, 6, 2, 4, 1,
    -- filter=169 channel=48
    -3, 2, 12, -12, -1, -1, 0, 0, 7,
    -- filter=169 channel=49
    -2, -4, 1, -5, 3, 0, -7, 5, 3,
    -- filter=169 channel=50
    -6, -5, 5, -8, 2, -9, -5, 1, 0,
    -- filter=169 channel=51
    6, 4, -5, -6, -3, 4, 0, 5, 6,
    -- filter=169 channel=52
    4, 4, 4, 1, 5, 4, -5, 4, -7,
    -- filter=169 channel=53
    6, 0, 0, -4, -2, -11, -3, -1, -6,
    -- filter=169 channel=54
    4, 0, -6, 0, 3, 2, -3, 7, 0,
    -- filter=169 channel=55
    -4, 8, -2, 0, 12, -13, 4, 5, -5,
    -- filter=169 channel=56
    -5, 16, -4, 9, 8, -4, -3, 0, 1,
    -- filter=169 channel=57
    -1, -7, 2, 1, -7, -1, -4, -5, -3,
    -- filter=169 channel=58
    2, -5, 4, -1, 0, -3, -1, -3, 1,
    -- filter=169 channel=59
    -5, -6, 14, -14, 8, 7, 5, 3, -5,
    -- filter=169 channel=60
    -4, 5, 6, -5, 4, 0, 5, -1, 0,
    -- filter=169 channel=61
    6, 6, 4, 8, 10, -2, -6, 9, -6,
    -- filter=169 channel=62
    -2, -3, 3, 0, 6, 2, 0, 4, -5,
    -- filter=169 channel=63
    -5, 2, -3, -6, 3, -2, 0, 4, 0,
    -- filter=169 channel=64
    0, -3, 0, -2, -4, -3, 2, -5, 3,
    -- filter=169 channel=65
    -6, 5, 5, -2, 0, 5, 1, 6, 5,
    -- filter=169 channel=66
    19, 0, 3, 9, 8, 11, 1, 15, 0,
    -- filter=169 channel=67
    2, -4, -2, 2, 5, -2, -1, 0, 7,
    -- filter=169 channel=68
    -4, -8, -4, -2, -4, -1, 4, -6, -4,
    -- filter=169 channel=69
    7, -5, -4, 0, -2, 7, 0, 7, 6,
    -- filter=169 channel=70
    -6, 10, -5, -2, 0, 3, 0, -4, 4,
    -- filter=169 channel=71
    -2, -5, -2, -1, -4, -3, -8, 0, 3,
    -- filter=169 channel=72
    1, -9, 0, -11, -2, 1, 0, 2, -12,
    -- filter=169 channel=73
    -5, 1, 6, -2, 14, 0, -2, -2, -6,
    -- filter=169 channel=74
    -13, 22, -5, 2, 15, -6, 4, 5, 0,
    -- filter=169 channel=75
    -3, -14, 2, -16, -2, 17, -6, 3, 1,
    -- filter=169 channel=76
    11, 0, -11, 5, 0, -12, 2, 7, -9,
    -- filter=169 channel=77
    3, 3, 5, -5, 5, 5, 7, -2, -5,
    -- filter=169 channel=78
    -6, -4, 2, -2, -1, -1, 1, 5, -3,
    -- filter=169 channel=79
    -6, -1, 12, -5, 17, 0, 0, 9, -6,
    -- filter=169 channel=80
    -13, -5, 8, -14, 11, 4, -2, 1, -4,
    -- filter=169 channel=81
    4, 5, -6, -5, -1, -3, 4, 5, 1,
    -- filter=169 channel=82
    2, -6, 1, -6, -2, 0, -6, -4, 3,
    -- filter=169 channel=83
    -5, 2, -3, -9, 0, 2, 4, -1, -1,
    -- filter=169 channel=84
    0, 11, -6, -7, 6, -7, 6, 13, 0,
    -- filter=169 channel=85
    -6, -7, -3, -6, -1, 0, 2, 5, 2,
    -- filter=169 channel=86
    7, 0, 2, 4, 8, 0, 8, 8, -1,
    -- filter=169 channel=87
    4, 12, -10, 3, 2, -1, 7, 1, -7,
    -- filter=169 channel=88
    -4, 12, -6, -2, -1, -11, -2, 0, 0,
    -- filter=169 channel=89
    6, -12, -2, -10, 5, -3, -9, 12, 0,
    -- filter=169 channel=90
    1, 7, -9, 2, 8, 0, -7, -2, -2,
    -- filter=169 channel=91
    -13, 8, -6, -8, 12, -7, -3, 2, 4,
    -- filter=169 channel=92
    -9, -4, -5, 5, 7, -2, -2, 2, -1,
    -- filter=169 channel=93
    -1, -8, 11, -9, 4, 1, 1, 2, 2,
    -- filter=169 channel=94
    1, -4, 1, 6, -4, -4, 1, 1, -1,
    -- filter=169 channel=95
    3, -6, 3, 5, 0, -2, 0, -2, -5,
    -- filter=169 channel=96
    -8, -4, -5, 4, -7, 0, -6, -3, 5,
    -- filter=169 channel=97
    2, -11, 1, 0, -11, -3, -2, -5, -5,
    -- filter=169 channel=98
    -9, -6, 14, -15, 7, -2, 0, 14, -8,
    -- filter=169 channel=99
    -11, 6, -5, -15, 15, -9, 3, 2, -7,
    -- filter=169 channel=100
    -5, -1, 4, 9, -4, -2, 2, 3, 7,
    -- filter=169 channel=101
    -2, -10, -2, -5, -5, -5, 0, -1, 0,
    -- filter=169 channel=102
    6, 4, 1, 5, 7, -6, 1, -5, 1,
    -- filter=169 channel=103
    -8, -12, 0, -4, -4, 16, -5, 1, -5,
    -- filter=169 channel=104
    -4, -7, 0, -14, -1, 1, -6, -1, -9,
    -- filter=169 channel=105
    5, -4, 0, 9, -5, -7, 5, 4, 3,
    -- filter=169 channel=106
    -1, -4, 3, -2, -6, -1, -8, 0, -3,
    -- filter=169 channel=107
    -3, 0, -9, -8, -4, 0, -6, 0, -10,
    -- filter=169 channel=108
    -1, 1, -4, -6, 4, 6, 6, 1, 2,
    -- filter=169 channel=109
    -16, 12, 11, -5, 25, -4, -8, 7, 0,
    -- filter=169 channel=110
    1, 2, 3, -6, -2, -9, 6, -5, -1,
    -- filter=169 channel=111
    -2, -4, 5, 2, -1, 5, -7, 2, -1,
    -- filter=169 channel=112
    -5, 7, -1, -5, 11, -4, -1, 6, -4,
    -- filter=169 channel=113
    0, -8, 4, -8, 0, 3, -1, 1, -8,
    -- filter=169 channel=114
    -5, 2, 5, -13, 19, 5, 0, 12, 4,
    -- filter=169 channel=115
    -1, -1, 6, -4, -6, 2, -7, -6, -1,
    -- filter=169 channel=116
    -1, 2, -2, -8, 11, -9, -6, 9, -1,
    -- filter=169 channel=117
    -3, 4, 3, 6, 6, 2, 0, 6, 2,
    -- filter=169 channel=118
    3, 3, 0, 6, 2, 5, -3, 2, 3,
    -- filter=169 channel=119
    -3, 13, 6, 7, 12, 6, 3, -1, 3,
    -- filter=169 channel=120
    -21, 16, -2, -2, 16, -5, 0, -1, -1,
    -- filter=169 channel=121
    9, 5, -1, 3, 4, 6, 0, 2, 3,
    -- filter=169 channel=122
    -2, 7, 7, -3, 9, 5, 6, -4, -9,
    -- filter=169 channel=123
    0, 2, -5, 4, 0, 6, -5, -5, -3,
    -- filter=169 channel=124
    3, -2, -4, -3, -1, -3, -6, -5, 3,
    -- filter=169 channel=125
    0, 4, 11, -15, 15, 2, -8, 1, -9,
    -- filter=169 channel=126
    5, -12, -4, -9, 3, 3, -9, -2, 5,
    -- filter=169 channel=127
    -1, -4, -4, 0, 5, 0, -3, 4, 4,
    -- filter=170 channel=0
    -1, -13, -1, -10, -28, -16, -4, -13, -15,
    -- filter=170 channel=1
    -4, -6, 8, -3, -19, -19, 0, 0, -5,
    -- filter=170 channel=2
    -4, 6, 7, 2, 2, -4, -4, 6, -3,
    -- filter=170 channel=3
    10, 13, 5, 3, -1, 8, -6, -2, -3,
    -- filter=170 channel=4
    3, 4, 6, 0, -6, -10, 4, -5, 5,
    -- filter=170 channel=5
    4, -1, -4, -6, -10, -2, -12, -8, -7,
    -- filter=170 channel=6
    5, 0, 0, -4, 0, -7, -5, 3, -9,
    -- filter=170 channel=7
    -6, 4, -1, 0, -3, -2, 5, 4, 1,
    -- filter=170 channel=8
    -5, -3, 4, 3, -1, -6, 2, 3, 5,
    -- filter=170 channel=9
    -5, 1, -4, -8, 0, 1, -3, -1, 3,
    -- filter=170 channel=10
    11, 11, 1, 1, 3, -2, -9, 0, -8,
    -- filter=170 channel=11
    -8, 3, -1, -2, -6, -4, 4, 1, -1,
    -- filter=170 channel=12
    0, 0, 6, 6, 0, -6, 7, -2, 0,
    -- filter=170 channel=13
    0, 6, 4, -5, -12, 6, 5, 0, -8,
    -- filter=170 channel=14
    -7, 0, 2, 2, 5, 5, -1, 4, 7,
    -- filter=170 channel=15
    -2, -5, -1, -2, -17, 4, -6, -7, -11,
    -- filter=170 channel=16
    5, 9, 8, -5, 7, 3, -10, -3, -1,
    -- filter=170 channel=17
    -3, 0, 4, 0, 4, 2, 1, -6, 4,
    -- filter=170 channel=18
    -2, -17, 5, -4, -28, -12, 6, -6, -15,
    -- filter=170 channel=19
    2, -5, -3, 2, 3, 3, -4, -4, -5,
    -- filter=170 channel=20
    -6, 7, 3, 7, 0, -3, 11, 2, -3,
    -- filter=170 channel=21
    0, 15, -3, 5, 14, 10, -3, 11, -1,
    -- filter=170 channel=22
    1, 3, 6, -10, -8, -9, -3, 0, -4,
    -- filter=170 channel=23
    6, 14, 9, -7, -4, 4, -4, -10, 6,
    -- filter=170 channel=24
    -1, -4, 5, 0, -2, -7, 5, -6, 0,
    -- filter=170 channel=25
    0, -4, 7, -4, -19, 1, 0, -7, -7,
    -- filter=170 channel=26
    -2, 8, 5, 4, -2, 0, -3, 1, 9,
    -- filter=170 channel=27
    1, 6, 3, -14, -18, -2, 2, -12, -11,
    -- filter=170 channel=28
    3, 2, -1, -5, 7, -5, 6, -5, 6,
    -- filter=170 channel=29
    5, 5, 0, -3, 1, 0, 10, 8, -9,
    -- filter=170 channel=30
    -2, 1, 7, -3, -20, -9, -5, -9, -2,
    -- filter=170 channel=31
    8, 26, 6, 4, 20, 5, -3, 0, 3,
    -- filter=170 channel=32
    -5, -1, 10, -18, -22, -7, 1, -7, -3,
    -- filter=170 channel=33
    -4, 1, 1, -13, -6, 0, -9, -11, -5,
    -- filter=170 channel=34
    0, 1, 5, 0, 2, 1, -2, -5, 8,
    -- filter=170 channel=35
    -7, -7, 1, 5, 2, 6, -2, -2, 2,
    -- filter=170 channel=36
    7, 1, -1, 9, 6, 1, 8, 4, 4,
    -- filter=170 channel=37
    5, 1, -1, -10, -14, -2, -8, -12, 6,
    -- filter=170 channel=38
    5, 5, 8, 1, 4, 4, -7, -7, 2,
    -- filter=170 channel=39
    3, 4, 4, 4, -4, 2, -2, 4, 5,
    -- filter=170 channel=40
    0, 2, 8, -1, -5, 5, 7, 0, -4,
    -- filter=170 channel=41
    10, -9, 1, 14, -5, -16, 1, -2, -4,
    -- filter=170 channel=42
    5, 2, -4, -3, -8, -6, -6, 0, -9,
    -- filter=170 channel=43
    8, 0, 1, -1, 0, 5, -5, -5, -4,
    -- filter=170 channel=44
    2, 6, 7, 1, 1, -1, -9, -11, 7,
    -- filter=170 channel=45
    -7, -7, 0, -2, -7, 3, -7, 5, -5,
    -- filter=170 channel=46
    6, -5, -1, -4, -6, 0, -2, -7, 3,
    -- filter=170 channel=47
    10, 8, -4, 0, 3, -2, -10, 1, -5,
    -- filter=170 channel=48
    -2, 0, 2, 0, -11, -10, -3, 0, 1,
    -- filter=170 channel=49
    -1, -2, -2, -11, -7, 0, 8, -8, -10,
    -- filter=170 channel=50
    2, 0, 0, -11, 1, -5, -5, 3, 0,
    -- filter=170 channel=51
    -2, -3, 0, -4, 4, -3, 0, -6, -6,
    -- filter=170 channel=52
    -1, -1, 8, 2, 0, 3, 6, -8, -1,
    -- filter=170 channel=53
    -7, -6, 6, 3, 6, 2, -2, 6, 4,
    -- filter=170 channel=54
    -7, -1, 3, -7, 4, 7, -3, 6, 0,
    -- filter=170 channel=55
    6, -3, 2, -3, 0, 7, -1, 2, -11,
    -- filter=170 channel=56
    3, 5, 2, 0, -8, 1, 0, 0, 8,
    -- filter=170 channel=57
    2, -4, -2, -6, 3, 4, 0, 1, 3,
    -- filter=170 channel=58
    -3, -3, 1, -3, -11, -4, -3, -10, -5,
    -- filter=170 channel=59
    -7, 2, -1, -9, 2, -1, -7, -8, 0,
    -- filter=170 channel=60
    -1, 4, 0, -4, -3, 2, -4, 3, -1,
    -- filter=170 channel=61
    4, 4, 8, 10, -3, 5, -1, 5, -2,
    -- filter=170 channel=62
    0, 1, 0, 3, -5, -3, -3, 4, 5,
    -- filter=170 channel=63
    0, -2, -8, 3, -1, -3, 0, -3, -3,
    -- filter=170 channel=64
    3, 6, 2, 9, 11, 0, -2, 0, 2,
    -- filter=170 channel=65
    0, 5, 4, -3, 7, 3, 0, -2, -4,
    -- filter=170 channel=66
    -2, -6, 5, 9, -5, -7, 8, -4, -7,
    -- filter=170 channel=67
    3, 5, -3, 0, 7, -1, -3, -4, 3,
    -- filter=170 channel=68
    0, 4, 6, 2, 6, 1, 6, 0, 5,
    -- filter=170 channel=69
    6, -2, 1, -6, -2, -4, 0, -4, 0,
    -- filter=170 channel=70
    -4, -2, 13, -5, -19, -2, -7, -14, 0,
    -- filter=170 channel=71
    3, 11, 3, 2, 0, 14, 4, -4, 1,
    -- filter=170 channel=72
    2, 9, 4, -4, 11, -2, 6, 0, -10,
    -- filter=170 channel=73
    -6, 1, -2, -8, -10, 3, 6, -6, -8,
    -- filter=170 channel=74
    -1, 0, 10, -4, -11, 0, -3, 0, 0,
    -- filter=170 channel=75
    4, -1, 4, -5, -25, -7, -11, -15, -6,
    -- filter=170 channel=76
    -6, -6, -3, 1, 2, 0, 10, 5, -3,
    -- filter=170 channel=77
    -4, 2, 1, 8, -4, -2, 8, -6, 2,
    -- filter=170 channel=78
    -2, 5, 1, 4, -5, 5, 0, -6, 5,
    -- filter=170 channel=79
    -3, 0, 2, -16, -23, -9, 0, -17, -10,
    -- filter=170 channel=80
    8, 15, 3, -9, 2, 0, -7, 2, -13,
    -- filter=170 channel=81
    -3, 0, -2, -3, -7, -6, 2, -4, 4,
    -- filter=170 channel=82
    8, 6, 6, -7, 4, 5, 0, -5, 1,
    -- filter=170 channel=83
    0, 4, 0, -5, -1, 1, -1, 4, 1,
    -- filter=170 channel=84
    -1, 1, 0, 2, -12, -3, -3, -10, -2,
    -- filter=170 channel=85
    -3, 3, 4, 1, -3, 6, 5, -1, 6,
    -- filter=170 channel=86
    0, 2, 6, 3, -16, 0, -6, -8, 0,
    -- filter=170 channel=87
    4, -4, 9, 9, -5, 0, 9, 0, 8,
    -- filter=170 channel=88
    1, 7, 0, 15, 20, 8, 6, 2, 7,
    -- filter=170 channel=89
    2, -3, -1, -4, 1, 0, 0, -2, -1,
    -- filter=170 channel=90
    11, 4, 3, 13, 19, 19, -2, 2, 7,
    -- filter=170 channel=91
    -11, 0, 5, -4, -5, 2, 0, -4, -8,
    -- filter=170 channel=92
    3, 3, 4, -2, 0, 3, 2, -4, 5,
    -- filter=170 channel=93
    5, 1, 6, -5, -11, -16, -4, 0, -2,
    -- filter=170 channel=94
    1, -3, 3, 2, 7, -1, -6, 7, -3,
    -- filter=170 channel=95
    7, 0, -2, -2, 3, 5, 4, -5, -4,
    -- filter=170 channel=96
    -4, -4, 3, -1, -2, 3, -1, 6, 3,
    -- filter=170 channel=97
    10, 3, 2, -2, 0, 6, -9, -7, -3,
    -- filter=170 channel=98
    5, 5, 7, -13, -6, -9, 2, -11, -15,
    -- filter=170 channel=99
    11, 7, 7, 0, 14, 18, -4, 5, 0,
    -- filter=170 channel=100
    7, 3, -4, 0, 5, -4, -1, 4, 7,
    -- filter=170 channel=101
    -6, 4, -2, 7, -3, -1, 11, 0, 4,
    -- filter=170 channel=102
    -3, -1, 1, 1, 0, -4, -7, 0, 3,
    -- filter=170 channel=103
    3, 14, 4, 4, 10, 0, -14, -1, -6,
    -- filter=170 channel=104
    4, 2, 0, -6, 13, 5, 0, -5, 0,
    -- filter=170 channel=105
    -5, 2, -4, 8, 6, -5, 4, -4, 5,
    -- filter=170 channel=106
    3, 3, -5, 6, 8, -5, 10, -3, 4,
    -- filter=170 channel=107
    -5, -8, 6, -12, -17, -6, -1, -6, -7,
    -- filter=170 channel=108
    1, -9, -6, 0, 0, -9, 2, 4, -9,
    -- filter=170 channel=109
    -3, 2, 3, -16, -19, 0, 0, -6, 0,
    -- filter=170 channel=110
    7, 11, 1, 10, 8, 9, -2, 3, 3,
    -- filter=170 channel=111
    0, 1, 0, 7, 3, 3, 7, 7, -3,
    -- filter=170 channel=112
    4, 2, -1, 0, -6, 9, -8, -14, 0,
    -- filter=170 channel=113
    -1, 8, 1, -6, 0, 15, -9, -3, 2,
    -- filter=170 channel=114
    -14, -13, -2, -20, -25, -26, -5, -14, -19,
    -- filter=170 channel=115
    6, 1, 0, -1, -2, 0, 0, -5, 0,
    -- filter=170 channel=116
    1, -3, -1, -9, -8, 0, 9, 0, -3,
    -- filter=170 channel=117
    -8, 0, 2, -8, -5, -4, 0, 7, 5,
    -- filter=170 channel=118
    4, 3, 1, 1, 3, 5, 5, -2, -1,
    -- filter=170 channel=119
    3, 6, 6, 10, 5, -6, 5, -1, 2,
    -- filter=170 channel=120
    -4, 6, 0, -5, -18, 3, -2, -6, 3,
    -- filter=170 channel=121
    -2, -2, -1, -3, 5, 4, -2, -3, 0,
    -- filter=170 channel=122
    15, 8, 0, 9, 20, 12, -10, -2, 5,
    -- filter=170 channel=123
    -3, 9, 11, -2, -3, 10, 0, -5, 0,
    -- filter=170 channel=124
    -6, -3, 5, 3, 0, -1, 7, 7, -7,
    -- filter=170 channel=125
    -9, 12, -3, -4, 8, 6, -1, 2, -9,
    -- filter=170 channel=126
    2, 3, 6, 4, 0, -4, -10, -9, -14,
    -- filter=170 channel=127
    2, 0, 3, 7, 3, -3, 3, 0, -1,
    -- filter=171 channel=0
    5, 8, 0, 12, 0, 4, 5, -9, 1,
    -- filter=171 channel=1
    5, 7, -2, 9, -4, -8, 5, 4, -5,
    -- filter=171 channel=2
    -5, 0, -5, -6, 1, -8, 5, -5, -6,
    -- filter=171 channel=3
    -1, 9, -3, -4, 5, -5, -4, 1, 0,
    -- filter=171 channel=4
    4, 3, -4, -1, -13, 0, -9, -1, -7,
    -- filter=171 channel=5
    5, 13, 1, 7, 14, 10, -5, 2, 8,
    -- filter=171 channel=6
    -4, 0, 0, 2, 4, -2, -5, 2, 0,
    -- filter=171 channel=7
    5, 2, 0, -6, 7, 4, -6, 3, -2,
    -- filter=171 channel=8
    5, 1, -7, 3, 3, 1, 0, 3, 6,
    -- filter=171 channel=9
    6, 9, 8, -2, 3, 4, 3, 5, -2,
    -- filter=171 channel=10
    -3, 8, 4, 4, -4, -1, 0, -4, -3,
    -- filter=171 channel=11
    2, 0, -8, 2, 0, -4, -4, 0, -1,
    -- filter=171 channel=12
    2, -5, 2, -4, 0, -11, -1, -11, 0,
    -- filter=171 channel=13
    -4, 0, 2, -10, -11, -13, -2, -9, -15,
    -- filter=171 channel=14
    1, 0, 4, -6, -1, -3, 4, 3, -4,
    -- filter=171 channel=15
    0, -1, -8, -14, -12, -4, -12, -6, -2,
    -- filter=171 channel=16
    0, 0, -2, 6, 9, -3, 5, 7, 0,
    -- filter=171 channel=17
    2, 4, -6, 1, -4, 7, 7, -3, -5,
    -- filter=171 channel=18
    -5, -6, -1, -12, -9, -16, -4, -6, -16,
    -- filter=171 channel=19
    -2, 2, 3, -2, -5, -5, 0, 1, 5,
    -- filter=171 channel=20
    2, -9, -9, -3, 0, -11, -2, -4, -2,
    -- filter=171 channel=21
    -1, 3, 4, 9, 12, 7, 1, 8, 6,
    -- filter=171 channel=22
    3, -4, 4, -2, -7, -8, 5, 1, -4,
    -- filter=171 channel=23
    0, 2, -8, -2, -17, -18, -10, -8, -3,
    -- filter=171 channel=24
    0, 5, 5, 6, 7, -6, -2, -3, 6,
    -- filter=171 channel=25
    6, 3, -3, -5, -5, -13, 3, 0, 0,
    -- filter=171 channel=26
    7, 5, -3, 10, 2, 0, -4, 6, 3,
    -- filter=171 channel=27
    3, 2, 4, -3, -18, -5, -5, -11, -9,
    -- filter=171 channel=28
    -6, -1, 0, -2, 1, -3, -3, -6, 5,
    -- filter=171 channel=29
    -4, 5, 0, -8, -7, -3, -1, -7, 2,
    -- filter=171 channel=30
    -3, 3, 8, -1, 4, -3, 5, 4, -2,
    -- filter=171 channel=31
    0, -1, 7, 3, -12, 2, 4, -5, 3,
    -- filter=171 channel=32
    -5, 1, -4, 0, -18, -8, 2, -11, -9,
    -- filter=171 channel=33
    3, 0, 0, -7, -8, -5, -3, -5, -7,
    -- filter=171 channel=34
    1, -4, 0, -4, -9, -3, 0, -2, 1,
    -- filter=171 channel=35
    4, 4, -5, 3, -6, -6, 0, 1, -3,
    -- filter=171 channel=36
    -1, -10, -1, -8, -4, 0, -6, -8, -5,
    -- filter=171 channel=37
    7, 6, 3, 0, 2, 9, 0, 1, 6,
    -- filter=171 channel=38
    6, 2, 5, 5, -7, -5, 2, 2, 4,
    -- filter=171 channel=39
    5, -5, 0, 6, -3, 2, 0, -7, -5,
    -- filter=171 channel=40
    -4, 0, -2, -8, -3, -10, 0, -1, 2,
    -- filter=171 channel=41
    -4, -2, -6, -6, -9, -18, -4, -16, -5,
    -- filter=171 channel=42
    1, 7, 2, -6, -2, 7, -5, 4, 3,
    -- filter=171 channel=43
    3, -7, -6, -1, -2, -7, -5, -9, -10,
    -- filter=171 channel=44
    5, 0, 2, 2, -6, 10, -4, 1, 7,
    -- filter=171 channel=45
    1, -6, 1, 5, -1, -3, 0, -2, 6,
    -- filter=171 channel=46
    -5, 2, -4, -3, -7, 2, -5, 4, -3,
    -- filter=171 channel=47
    3, 5, 10, 8, 6, 12, 0, 12, 15,
    -- filter=171 channel=48
    0, 0, -4, 3, 4, 2, -5, -2, 9,
    -- filter=171 channel=49
    0, 3, -3, -3, -3, -5, -1, 1, -7,
    -- filter=171 channel=50
    0, -7, 10, -2, -15, 4, -7, 0, 2,
    -- filter=171 channel=51
    3, 1, 6, 2, -2, -3, -3, 4, 3,
    -- filter=171 channel=52
    4, 3, -5, 0, -6, -9, -1, -12, 2,
    -- filter=171 channel=53
    -5, -8, -5, 4, -1, 4, -1, -9, 1,
    -- filter=171 channel=54
    0, 4, 5, 6, -7, 2, -6, -4, -1,
    -- filter=171 channel=55
    -6, 1, 0, -16, -14, -10, -3, -15, -12,
    -- filter=171 channel=56
    0, 3, -5, 2, -8, 5, -8, 3, 3,
    -- filter=171 channel=57
    -1, 0, -1, 4, -2, -6, 5, -2, 4,
    -- filter=171 channel=58
    -2, 3, 4, 0, 3, 10, -3, 2, 7,
    -- filter=171 channel=59
    -5, -4, -2, -8, -2, -9, 0, -7, -3,
    -- filter=171 channel=60
    6, 4, 4, -3, -2, 6, 2, -2, 0,
    -- filter=171 channel=61
    -6, -4, 3, 0, 3, -9, -1, -4, -2,
    -- filter=171 channel=62
    1, -5, 3, 0, -2, 4, 6, 1, 6,
    -- filter=171 channel=63
    6, 1, 0, 10, 2, 3, 7, 0, 5,
    -- filter=171 channel=64
    -6, -3, -7, -7, -9, -9, 4, 0, 0,
    -- filter=171 channel=65
    -5, -2, 0, -5, -7, 7, 0, 3, 1,
    -- filter=171 channel=66
    3, -2, -5, -3, -12, -7, 5, -13, 2,
    -- filter=171 channel=67
    3, -6, 0, 0, -4, 4, -4, 1, 3,
    -- filter=171 channel=68
    0, -1, 2, -8, 2, -7, 5, 2, -5,
    -- filter=171 channel=69
    -1, 7, 4, 1, 4, -2, 0, -6, 5,
    -- filter=171 channel=70
    5, -5, 5, -12, -18, -14, -6, -5, -10,
    -- filter=171 channel=71
    -6, 5, 0, -1, 0, 1, -2, 2, 4,
    -- filter=171 channel=72
    0, -8, 1, 3, -11, 0, -2, -2, 0,
    -- filter=171 channel=73
    1, 0, -2, -8, -11, -6, 2, -5, -5,
    -- filter=171 channel=74
    -3, 0, 5, -6, -3, -5, 3, -3, 1,
    -- filter=171 channel=75
    -3, 16, 8, -1, 12, 1, 1, -3, 2,
    -- filter=171 channel=76
    -2, -1, -11, -1, -5, -3, -4, -4, -6,
    -- filter=171 channel=77
    -1, 1, 0, 6, 3, -6, 2, 2, -3,
    -- filter=171 channel=78
    6, 9, 1, 9, 0, 5, 4, 2, 3,
    -- filter=171 channel=79
    -2, -13, -11, -14, -18, -19, -14, -13, -19,
    -- filter=171 channel=80
    3, -2, -2, 3, 4, 0, -1, 0, 14,
    -- filter=171 channel=81
    -7, -3, 4, -5, -7, -7, 5, 0, 0,
    -- filter=171 channel=82
    -5, -6, 0, -1, 3, 0, 1, -8, 1,
    -- filter=171 channel=83
    -5, 0, -2, -1, 2, 2, -8, -5, -1,
    -- filter=171 channel=84
    -6, -1, 3, 0, -5, -5, -3, -2, -7,
    -- filter=171 channel=85
    2, 1, 2, 3, 5, -5, 2, -4, -7,
    -- filter=171 channel=86
    -5, -6, -3, 0, 1, -2, 6, -8, 6,
    -- filter=171 channel=87
    3, 3, -10, -4, -1, -2, 5, -6, -1,
    -- filter=171 channel=88
    -2, 0, -5, -5, 2, -2, 0, 1, 4,
    -- filter=171 channel=89
    -8, -3, 2, -16, -5, -12, -4, -6, -8,
    -- filter=171 channel=90
    -3, -10, 5, -3, -7, -3, -6, -4, -1,
    -- filter=171 channel=91
    1, -2, -3, -1, -6, 0, 0, 0, -7,
    -- filter=171 channel=92
    -3, 0, -7, -7, 0, -6, -2, 2, 1,
    -- filter=171 channel=93
    0, 5, 11, 12, 3, 0, -2, 10, 7,
    -- filter=171 channel=94
    0, -6, 1, 0, -1, 4, 7, 6, -1,
    -- filter=171 channel=95
    -7, 3, -3, -8, -1, 0, 5, 5, -4,
    -- filter=171 channel=96
    2, 4, -3, 1, 3, 1, -3, -3, -7,
    -- filter=171 channel=97
    7, 7, 0, 4, 1, -3, 0, 0, -2,
    -- filter=171 channel=98
    6, 2, 12, -2, 0, 3, -2, -5, 0,
    -- filter=171 channel=99
    -4, 0, -1, -6, -14, 3, -1, -9, 5,
    -- filter=171 channel=100
    2, 0, 5, 2, -4, 4, -4, 3, -2,
    -- filter=171 channel=101
    -6, -9, 2, -7, -9, -3, 0, -2, -7,
    -- filter=171 channel=102
    7, 1, -1, 1, 5, -6, 6, -3, 0,
    -- filter=171 channel=103
    3, 10, 12, 0, 11, 13, 7, -2, 7,
    -- filter=171 channel=104
    -3, -1, 8, -4, 3, 0, -6, -2, 7,
    -- filter=171 channel=105
    1, 3, -2, 3, -5, 4, -3, -4, -8,
    -- filter=171 channel=106
    -4, -7, -2, -7, 3, -1, -1, -7, -8,
    -- filter=171 channel=107
    -7, -5, 3, -6, -5, -11, -5, -11, -2,
    -- filter=171 channel=108
    -3, -1, -1, 0, -3, -4, 7, 5, -8,
    -- filter=171 channel=109
    -2, -8, 7, -9, -17, -11, -10, -11, 1,
    -- filter=171 channel=110
    -5, 0, 3, 6, 4, -4, -3, -3, 4,
    -- filter=171 channel=111
    -5, -1, 3, 1, -7, 3, 2, 7, -6,
    -- filter=171 channel=112
    8, -5, 3, 0, -3, -2, -7, 1, -3,
    -- filter=171 channel=113
    -2, 1, 3, -7, -5, 2, -7, 1, 4,
    -- filter=171 channel=114
    2, -9, -6, 3, -13, -6, 0, -9, -13,
    -- filter=171 channel=115
    7, -5, 3, -5, 6, -3, -5, -4, 1,
    -- filter=171 channel=116
    4, -2, 1, -8, -11, -4, 6, 0, 4,
    -- filter=171 channel=117
    -5, 2, -3, -5, 4, 2, 6, -6, -8,
    -- filter=171 channel=118
    4, 5, 1, -3, -1, 4, -5, -2, 2,
    -- filter=171 channel=119
    -1, 0, -5, -4, -7, -3, 2, -12, -5,
    -- filter=171 channel=120
    5, -8, 5, -7, -15, -1, -5, -9, 0,
    -- filter=171 channel=121
    -3, 5, -7, -8, -4, 2, -1, 2, -8,
    -- filter=171 channel=122
    1, -2, 1, 13, 13, 7, 1, 13, 16,
    -- filter=171 channel=123
    0, -1, -1, -6, -8, -7, 3, -6, -3,
    -- filter=171 channel=124
    -2, 1, 2, -3, -4, -1, -5, -6, -9,
    -- filter=171 channel=125
    -2, 4, -2, 0, -2, -1, -6, -2, -4,
    -- filter=171 channel=126
    0, 7, -7, -3, 1, -5, -3, -7, 2,
    -- filter=171 channel=127
    -7, 2, -6, 0, -8, 3, -3, -3, 1,
    -- filter=172 channel=0
    21, 18, 8, 19, -2, -1, 6, -12, -14,
    -- filter=172 channel=1
    11, 16, 2, 6, -13, -12, 5, -21, -13,
    -- filter=172 channel=2
    3, -2, 6, -7, -6, 4, -3, -8, 3,
    -- filter=172 channel=3
    -8, 3, 0, -11, 1, -2, -6, -2, -2,
    -- filter=172 channel=4
    -7, -10, 0, -12, -16, -5, -7, -2, 12,
    -- filter=172 channel=5
    7, 18, 11, 9, 0, -9, -1, -21, -18,
    -- filter=172 channel=6
    -12, -13, -4, -8, -1, -1, 5, 12, 7,
    -- filter=172 channel=7
    -7, -6, 1, -7, 3, -6, -4, -6, -6,
    -- filter=172 channel=8
    0, 4, 0, -9, 0, -8, -10, 2, -3,
    -- filter=172 channel=9
    8, 14, 5, 9, 2, 8, -6, -3, 1,
    -- filter=172 channel=10
    2, -4, 6, 6, 6, 3, -5, -6, -2,
    -- filter=172 channel=11
    -10, -11, -15, -1, 2, 9, 5, 20, 11,
    -- filter=172 channel=12
    -8, -10, 0, 0, -9, -2, -5, -8, -3,
    -- filter=172 channel=13
    -5, -8, -4, -6, -2, 7, 5, -4, 8,
    -- filter=172 channel=14
    0, 7, -1, 7, -4, 6, 2, 0, 4,
    -- filter=172 channel=15
    -15, -12, -11, 0, 9, 3, 6, 19, 19,
    -- filter=172 channel=16
    10, 14, 5, 9, -8, 1, -15, -25, -17,
    -- filter=172 channel=17
    -5, -7, 6, 6, -6, -4, -2, 7, 6,
    -- filter=172 channel=18
    -14, -11, -7, 1, -5, 4, 24, 25, 4,
    -- filter=172 channel=19
    3, 6, 0, 0, -3, -2, 5, -1, -1,
    -- filter=172 channel=20
    -26, -26, -19, -12, -7, 9, 15, 25, 18,
    -- filter=172 channel=21
    17, 20, 14, 17, -4, -2, -10, -26, -9,
    -- filter=172 channel=22
    -4, -3, -4, -11, -7, -5, 0, -3, 10,
    -- filter=172 channel=23
    -15, -15, 0, -7, 8, 12, -5, 12, 6,
    -- filter=172 channel=24
    -1, -5, 6, -6, -6, 6, 3, 4, 0,
    -- filter=172 channel=25
    8, 7, 3, 0, 0, -4, 3, -15, -5,
    -- filter=172 channel=26
    14, 4, 7, 12, -8, -7, 1, -9, -11,
    -- filter=172 channel=27
    11, 4, -13, 0, 4, -2, 0, 5, 8,
    -- filter=172 channel=28
    -2, -1, 6, 6, 2, 5, -3, 6, -2,
    -- filter=172 channel=29
    -12, -28, -12, -3, -3, 6, 15, 29, 5,
    -- filter=172 channel=30
    15, 4, 6, 8, -6, -2, 0, -2, -9,
    -- filter=172 channel=31
    22, 24, 10, 12, 11, 10, -16, -14, -12,
    -- filter=172 channel=32
    -8, -9, -5, -13, -11, 0, -1, 3, 10,
    -- filter=172 channel=33
    9, 8, 6, 0, -5, 3, 1, -1, -5,
    -- filter=172 channel=34
    -18, -9, -1, -24, -9, -6, -19, -5, -1,
    -- filter=172 channel=35
    0, -6, -6, -2, 1, 6, 3, -3, 5,
    -- filter=172 channel=36
    -10, 1, 8, 2, 1, -4, 0, 0, 9,
    -- filter=172 channel=37
    16, 22, 4, 11, -6, -8, -3, -25, -22,
    -- filter=172 channel=38
    6, 3, -1, 2, 4, 3, 1, 3, -4,
    -- filter=172 channel=39
    -10, -4, -9, -1, 1, 4, 9, 9, 9,
    -- filter=172 channel=40
    0, -9, -3, -9, 3, 6, 0, 9, 3,
    -- filter=172 channel=41
    -22, -29, -6, -25, -21, -15, 0, -19, 1,
    -- filter=172 channel=42
    9, 4, -2, 3, 0, -2, 11, 4, -11,
    -- filter=172 channel=43
    -8, 0, 4, -3, -2, 5, 3, 9, 1,
    -- filter=172 channel=44
    10, 25, 14, 6, 3, -5, -1, -28, -11,
    -- filter=172 channel=45
    9, 8, -5, 9, -5, -2, -1, 8, 1,
    -- filter=172 channel=46
    -7, 2, 3, 3, 0, -2, -2, 1, -5,
    -- filter=172 channel=47
    21, 22, 10, 11, 6, 0, -10, -33, -16,
    -- filter=172 channel=48
    24, 24, 0, 7, 0, -4, -7, -24, -9,
    -- filter=172 channel=49
    0, -3, -11, 2, 0, 1, 0, 13, 7,
    -- filter=172 channel=50
    13, 12, 0, 1, 11, 6, 2, 0, -6,
    -- filter=172 channel=51
    -6, 0, 0, 4, -4, 1, -5, -6, -3,
    -- filter=172 channel=52
    -9, -18, -5, -17, -11, 0, -9, -4, 11,
    -- filter=172 channel=53
    -15, -10, -1, 1, 1, -1, 0, 4, 10,
    -- filter=172 channel=54
    1, -1, 0, 4, 5, -4, 1, 1, 0,
    -- filter=172 channel=55
    -23, -15, -11, 0, -2, 8, 14, 17, 16,
    -- filter=172 channel=56
    -4, -7, 1, -13, -1, -4, -7, -9, 1,
    -- filter=172 channel=57
    0, -7, 2, -8, -8, 3, 0, -6, -3,
    -- filter=172 channel=58
    7, 4, 7, 8, -2, -7, -9, -11, -7,
    -- filter=172 channel=59
    5, 2, 7, 12, 0, 7, 3, -18, -9,
    -- filter=172 channel=60
    -5, 6, 0, 2, 0, 3, -4, -1, -5,
    -- filter=172 channel=61
    -6, -1, -6, -2, -7, 5, 0, -4, -2,
    -- filter=172 channel=62
    -4, 0, 2, 2, -1, -1, 0, 0, -5,
    -- filter=172 channel=63
    -3, 9, -2, 3, 4, -6, -4, -11, -7,
    -- filter=172 channel=64
    -2, -11, 0, 4, -3, -5, 4, 1, 2,
    -- filter=172 channel=65
    0, 2, -4, -1, 0, 0, -2, 4, 5,
    -- filter=172 channel=66
    -6, -15, 1, -15, -18, -1, -11, -4, 7,
    -- filter=172 channel=67
    3, -1, 6, -2, -5, 6, 6, 8, -2,
    -- filter=172 channel=68
    0, -2, -1, 4, 0, -1, 8, 2, -1,
    -- filter=172 channel=69
    -7, 0, 3, 6, 6, 1, -3, -9, -3,
    -- filter=172 channel=70
    -6, -10, -11, -5, -8, -4, -3, 3, 10,
    -- filter=172 channel=71
    -6, 5, 6, 4, 6, -7, -7, -4, 5,
    -- filter=172 channel=72
    11, 7, 9, 11, 8, 6, 7, -8, -4,
    -- filter=172 channel=73
    2, -3, 1, -3, -9, 8, 6, 8, 8,
    -- filter=172 channel=74
    10, 8, 2, -3, -1, 1, -6, 3, 12,
    -- filter=172 channel=75
    10, 15, 5, -1, -14, -13, -1, -35, -18,
    -- filter=172 channel=76
    -18, -16, -11, -13, -5, 0, 15, 24, 16,
    -- filter=172 channel=77
    4, -7, -4, 2, 3, 5, -2, 0, -4,
    -- filter=172 channel=78
    -2, 7, 0, -2, -5, 2, 0, -11, -10,
    -- filter=172 channel=79
    -9, -12, -8, -3, 1, 7, 23, 14, 4,
    -- filter=172 channel=80
    20, 26, 8, 23, -4, 1, -3, -21, -9,
    -- filter=172 channel=81
    -1, 4, 7, -4, -6, -4, -7, 1, -2,
    -- filter=172 channel=82
    1, -3, -2, -2, -2, 0, -7, -1, -6,
    -- filter=172 channel=83
    9, 11, 7, 5, 5, 3, 7, -2, -4,
    -- filter=172 channel=84
    -11, -8, 0, -6, -10, -8, 1, 5, 7,
    -- filter=172 channel=85
    2, 0, 5, -6, -5, -4, 5, 0, 5,
    -- filter=172 channel=86
    -3, -8, 0, -9, -11, -6, 1, -3, 5,
    -- filter=172 channel=87
    -21, -19, -6, -20, -11, -1, -7, 0, 0,
    -- filter=172 channel=88
    3, 0, 9, 0, 0, -1, -9, -8, 7,
    -- filter=172 channel=89
    -9, -5, 3, 5, 1, 9, 13, 10, 4,
    -- filter=172 channel=90
    -5, 2, 7, -5, -9, 5, -12, -10, 6,
    -- filter=172 channel=91
    -5, -7, -10, 0, -2, -3, 2, 1, -1,
    -- filter=172 channel=92
    -11, -7, -3, -14, -10, -5, -1, 1, 6,
    -- filter=172 channel=93
    14, 28, 12, 15, -3, -5, -3, -16, -21,
    -- filter=172 channel=94
    -5, 4, 2, 4, 1, -4, 5, 4, 3,
    -- filter=172 channel=95
    -1, 1, -1, -1, 3, 0, 4, -2, -6,
    -- filter=172 channel=96
    0, -3, 2, 3, 0, -1, 1, 6, 5,
    -- filter=172 channel=97
    -1, 2, 8, -1, 0, -6, -2, 0, -9,
    -- filter=172 channel=98
    8, 15, 1, 14, 0, 6, 7, -12, -4,
    -- filter=172 channel=99
    -1, -7, 7, -13, 0, 14, 1, 2, 7,
    -- filter=172 channel=100
    -1, -3, 4, -8, -8, -5, 0, 0, 3,
    -- filter=172 channel=101
    -3, -2, 3, -6, 0, -3, 0, -7, 2,
    -- filter=172 channel=102
    -3, 0, -1, 7, -5, -2, -3, -6, 1,
    -- filter=172 channel=103
    8, 19, 11, 10, 8, 4, -9, -36, -13,
    -- filter=172 channel=104
    19, 18, 15, 8, 1, 6, 1, -11, -5,
    -- filter=172 channel=105
    -15, -11, -4, -5, -8, 9, 15, 22, 10,
    -- filter=172 channel=106
    -12, -5, -8, -6, 5, -6, 13, 13, 9,
    -- filter=172 channel=107
    -21, -22, -9, -9, -6, 7, 13, 18, 16,
    -- filter=172 channel=108
    3, -2, -3, -3, -7, 5, -3, 0, -5,
    -- filter=172 channel=109
    -3, -2, -6, -4, -11, -2, -1, -7, 0,
    -- filter=172 channel=110
    2, -1, 12, -1, -6, 1, -1, -1, 4,
    -- filter=172 channel=111
    -8, -2, -5, -1, 3, 7, -7, 0, 2,
    -- filter=172 channel=112
    10, 7, -4, 0, -5, 5, -4, 1, -4,
    -- filter=172 channel=113
    4, 1, 9, -10, -7, 3, -7, -5, 3,
    -- filter=172 channel=114
    -4, -8, -7, 4, -8, 0, 21, 12, 15,
    -- filter=172 channel=115
    -2, -5, 0, -7, -7, 6, 0, -3, -7,
    -- filter=172 channel=116
    8, 4, -5, 0, 3, -2, 1, 7, 4,
    -- filter=172 channel=117
    -3, 0, 1, -3, 0, 4, 5, -2, -4,
    -- filter=172 channel=118
    -1, 5, 6, 1, 5, 0, -5, -1, 0,
    -- filter=172 channel=119
    -14, -17, 1, -16, -19, 2, -18, -11, 7,
    -- filter=172 channel=120
    4, -9, -3, -6, 11, 11, 8, 12, 15,
    -- filter=172 channel=121
    1, -3, 2, -3, -3, -5, -7, -10, 6,
    -- filter=172 channel=122
    23, 36, 30, 14, 3, -3, -21, -47, -24,
    -- filter=172 channel=123
    -11, -5, -4, -9, -6, 1, -12, 0, 0,
    -- filter=172 channel=124
    -5, -4, -12, -1, 4, 3, 1, 7, 6,
    -- filter=172 channel=125
    13, 7, -3, -1, -2, 9, 0, 1, -5,
    -- filter=172 channel=126
    -3, 2, -4, -1, -7, -4, 0, 5, -4,
    -- filter=172 channel=127
    -4, 1, 5, 0, 0, 1, -3, 4, 0,
    -- filter=173 channel=0
    -4, 6, -2, 0, 11, 7, -11, -19, -10,
    -- filter=173 channel=1
    0, 8, -5, 12, -1, -5, -4, -27, -20,
    -- filter=173 channel=2
    1, 3, -1, 3, -8, -5, 4, -8, -3,
    -- filter=173 channel=3
    -4, -6, -1, -9, 11, 12, -10, 9, 2,
    -- filter=173 channel=4
    -4, 11, 7, 2, -5, 2, 0, 1, 4,
    -- filter=173 channel=5
    5, 11, -3, 10, 18, 8, 0, -2, -1,
    -- filter=173 channel=6
    4, -4, -4, 0, 4, -2, 6, -1, 4,
    -- filter=173 channel=7
    6, 4, 0, -1, 3, -3, 6, 0, 5,
    -- filter=173 channel=8
    -4, 6, 1, -4, -3, -6, 3, -10, 3,
    -- filter=173 channel=9
    4, -1, 9, 1, 0, 2, 0, 0, -9,
    -- filter=173 channel=10
    -1, 5, 1, 2, 1, 9, 6, 0, 2,
    -- filter=173 channel=11
    -10, -14, -1, -1, -11, 0, 7, 4, 4,
    -- filter=173 channel=12
    0, 0, -8, -5, 5, -3, 5, 0, -4,
    -- filter=173 channel=13
    -9, -7, -4, 0, 2, 1, 0, 0, 0,
    -- filter=173 channel=14
    -3, -1, 0, 4, -6, 1, -6, 6, 0,
    -- filter=173 channel=15
    -7, -7, -7, 2, 2, 11, 12, 3, -1,
    -- filter=173 channel=16
    1, -2, -9, 3, 5, 1, -8, 3, -2,
    -- filter=173 channel=17
    -3, -3, 6, -6, -1, -6, 5, 0, -1,
    -- filter=173 channel=18
    6, -3, 5, 0, 0, 4, 5, 0, -3,
    -- filter=173 channel=19
    4, -2, 6, 4, 5, -3, -5, -2, 4,
    -- filter=173 channel=20
    -3, -17, -13, -2, -9, 1, 8, 13, 18,
    -- filter=173 channel=21
    1, 0, 2, -4, 8, -5, -1, 0, -2,
    -- filter=173 channel=22
    -2, 1, -9, 5, 0, -3, 2, -6, 0,
    -- filter=173 channel=23
    -10, -9, 5, -8, 5, 8, 0, -2, -5,
    -- filter=173 channel=24
    -5, 3, -5, -4, 0, -4, 7, -1, -3,
    -- filter=173 channel=25
    -4, 4, 6, 11, 12, 6, -6, -21, -12,
    -- filter=173 channel=26
    -6, 2, 0, 0, 1, -2, 3, -2, -3,
    -- filter=173 channel=27
    0, 13, 10, 7, 12, 2, -1, -27, -22,
    -- filter=173 channel=28
    3, 0, 6, 1, 1, 3, 7, 6, -5,
    -- filter=173 channel=29
    -2, -17, -11, 0, -8, 1, 20, 12, 19,
    -- filter=173 channel=30
    -6, 8, 2, 8, 7, -3, -4, -15, -5,
    -- filter=173 channel=31
    -7, 2, 3, 3, 12, -2, 0, -20, -18,
    -- filter=173 channel=32
    0, 0, 7, 2, 0, 11, 3, -9, 0,
    -- filter=173 channel=33
    -8, 10, 11, -1, 3, 7, 3, -8, -11,
    -- filter=173 channel=34
    3, -1, -3, -2, 11, -6, 0, 1, 7,
    -- filter=173 channel=35
    1, -3, -6, -5, 1, 4, -3, -1, -6,
    -- filter=173 channel=36
    -1, -7, -10, -2, 0, -6, 0, 5, 1,
    -- filter=173 channel=37
    3, 11, 2, 13, 7, -4, -11, -24, -14,
    -- filter=173 channel=38
    4, 8, 2, 0, 10, 8, -1, -8, -2,
    -- filter=173 channel=39
    2, -13, -11, 3, 0, 0, 3, 5, 12,
    -- filter=173 channel=40
    -8, 0, -1, -4, -6, -2, 8, -4, -5,
    -- filter=173 channel=41
    -6, 10, 0, 8, -2, -1, 16, 13, -13,
    -- filter=173 channel=42
    0, 3, 8, 0, 5, 8, 1, -14, -6,
    -- filter=173 channel=43
    -4, -2, 6, 3, 3, 4, -1, 7, 1,
    -- filter=173 channel=44
    8, 5, 4, 8, 15, 2, -9, -14, -15,
    -- filter=173 channel=45
    -7, -8, 2, -3, 3, -4, -10, -8, 2,
    -- filter=173 channel=46
    -4, 7, 6, 1, 5, -5, 3, -4, -1,
    -- filter=173 channel=47
    -6, 14, 9, 5, 7, 14, -3, -11, -17,
    -- filter=173 channel=48
    1, 18, 13, 8, 2, 9, -11, -26, -24,
    -- filter=173 channel=49
    1, -2, 6, -9, -12, -7, -6, -8, 3,
    -- filter=173 channel=50
    0, 2, 9, 3, 1, -3, 3, -18, -5,
    -- filter=173 channel=51
    -4, 2, 0, 3, 2, -1, 7, 7, -1,
    -- filter=173 channel=52
    4, 4, -8, 2, 2, -8, -5, -1, 3,
    -- filter=173 channel=53
    4, -5, -6, -2, -5, -2, 14, 2, 5,
    -- filter=173 channel=54
    -4, -7, -2, -1, 0, -3, 7, -3, 0,
    -- filter=173 channel=55
    7, -12, -2, -1, 3, 0, 19, 11, 6,
    -- filter=173 channel=56
    5, -2, 0, -3, 2, 2, 2, -9, -2,
    -- filter=173 channel=57
    4, 7, 6, -3, -7, 0, 3, -2, 0,
    -- filter=173 channel=58
    5, 9, -2, 1, 2, 5, -4, 0, 0,
    -- filter=173 channel=59
    0, 5, 10, -1, 5, 9, -3, -7, -11,
    -- filter=173 channel=60
    1, 7, 1, 4, -1, -5, 4, 5, -1,
    -- filter=173 channel=61
    3, -4, -3, 0, 3, -4, 0, -5, 8,
    -- filter=173 channel=62
    -5, 0, 0, -6, 0, 2, -3, 6, -2,
    -- filter=173 channel=63
    3, -1, 1, 2, 4, 0, -6, 0, -8,
    -- filter=173 channel=64
    0, -1, -11, -2, -9, -7, -1, 1, 6,
    -- filter=173 channel=65
    2, 3, 0, 4, -3, -6, 7, 6, 1,
    -- filter=173 channel=66
    1, 0, -2, -3, -3, 0, 5, 9, -6,
    -- filter=173 channel=67
    6, -2, -5, 0, 0, 0, 5, 6, 3,
    -- filter=173 channel=68
    -5, -5, 1, -6, -5, 0, 3, 2, -9,
    -- filter=173 channel=69
    -1, 5, -5, 5, 4, -6, -3, -7, -5,
    -- filter=173 channel=70
    -3, 0, 8, -1, 0, -1, -15, -11, -1,
    -- filter=173 channel=71
    0, 3, 0, -6, -3, 2, -3, 8, 6,
    -- filter=173 channel=72
    -8, 3, 8, 6, 5, 5, 1, 0, -18,
    -- filter=173 channel=73
    -4, 0, 4, 3, 0, 2, -2, -10, 0,
    -- filter=173 channel=74
    0, 6, -2, 4, 13, 0, 0, -17, -6,
    -- filter=173 channel=75
    1, 7, 2, 16, 11, 12, -14, -22, -10,
    -- filter=173 channel=76
    -10, -17, -6, -4, -16, 7, 4, 9, 2,
    -- filter=173 channel=77
    0, 1, 2, -6, 1, 5, 7, -3, -3,
    -- filter=173 channel=78
    -5, 0, -2, 4, 12, 0, -1, 3, -7,
    -- filter=173 channel=79
    -5, -5, 10, -2, 8, 16, 9, -15, -11,
    -- filter=173 channel=80
    3, 7, 0, 3, 16, 12, 1, -19, -21,
    -- filter=173 channel=81
    4, -4, -4, 6, -7, 3, -5, 5, -5,
    -- filter=173 channel=82
    4, 3, -1, 0, -6, 2, -5, 0, -5,
    -- filter=173 channel=83
    1, 6, 6, 2, -1, -8, -6, -13, -2,
    -- filter=173 channel=84
    4, 9, 5, 2, -2, 1, 3, -14, -9,
    -- filter=173 channel=85
    7, 5, 1, 1, 0, -5, 0, 4, -1,
    -- filter=173 channel=86
    -4, 0, 3, -2, 0, -4, -9, 1, 3,
    -- filter=173 channel=87
    0, -2, -7, 1, 3, 0, -1, 0, 13,
    -- filter=173 channel=88
    1, 0, 2, 0, -6, -14, 3, -2, -8,
    -- filter=173 channel=89
    -6, 0, -2, -2, 4, 15, 12, 0, -12,
    -- filter=173 channel=90
    -4, -5, -9, -9, 2, 0, 3, 4, -2,
    -- filter=173 channel=91
    -4, 3, 6, -3, 3, 1, -3, -24, -6,
    -- filter=173 channel=92
    2, -4, -2, 3, -6, -6, -1, -6, 3,
    -- filter=173 channel=93
    -1, 20, 2, 3, 7, 3, -5, -12, -17,
    -- filter=173 channel=94
    7, 2, -3, -2, -5, -2, -5, -1, -6,
    -- filter=173 channel=95
    -6, -1, 8, -1, 1, 7, 4, 11, 1,
    -- filter=173 channel=96
    3, -2, 6, 2, 2, 4, 0, 5, -6,
    -- filter=173 channel=97
    5, -4, -1, -1, -2, 3, -3, 3, -2,
    -- filter=173 channel=98
    -3, 4, 17, 6, 15, 14, 2, -7, -13,
    -- filter=173 channel=99
    -4, -1, 1, 4, 15, 1, 5, -11, -3,
    -- filter=173 channel=100
    -5, 0, -2, 5, 7, 2, 7, 5, 3,
    -- filter=173 channel=101
    3, 5, 0, 4, -6, 1, 0, -4, -4,
    -- filter=173 channel=102
    -1, -7, -1, -1, -1, -3, -2, 0, 4,
    -- filter=173 channel=103
    0, 0, 9, 11, 21, 6, -10, -9, -10,
    -- filter=173 channel=104
    -5, 14, 3, 2, 11, 8, -2, -14, -18,
    -- filter=173 channel=105
    -7, -14, -3, -4, 1, -3, 2, 2, 11,
    -- filter=173 channel=106
    -6, 1, -11, -4, -8, -7, 0, 1, 6,
    -- filter=173 channel=107
    0, -9, -2, -5, -8, -4, 4, -3, 13,
    -- filter=173 channel=108
    3, 0, -10, -3, -3, -2, 3, 7, -7,
    -- filter=173 channel=109
    10, 17, 7, 6, 8, 4, -2, -19, -18,
    -- filter=173 channel=110
    -1, 8, 4, 0, 7, -1, -2, 8, -4,
    -- filter=173 channel=111
    4, 0, -9, 2, -3, 4, 6, 9, -1,
    -- filter=173 channel=112
    -4, 6, 0, 5, 6, 3, -11, -17, -4,
    -- filter=173 channel=113
    1, 0, 4, -4, 7, 10, 0, -2, 1,
    -- filter=173 channel=114
    2, 1, 5, 7, -4, -5, 0, -27, -10,
    -- filter=173 channel=115
    -1, 1, -4, -4, 4, 0, 5, -1, -1,
    -- filter=173 channel=116
    5, 11, 4, 1, 8, 2, -1, -8, -19,
    -- filter=173 channel=117
    -2, -5, -5, -6, -2, 0, 2, -10, -3,
    -- filter=173 channel=118
    -5, 6, 6, -1, 1, 3, 7, -4, -7,
    -- filter=173 channel=119
    11, 6, -3, 7, 3, -15, -1, -2, 0,
    -- filter=173 channel=120
    1, 1, 7, -3, 9, -5, 7, -17, -10,
    -- filter=173 channel=121
    6, 5, -2, 0, 10, 8, 0, -1, 3,
    -- filter=173 channel=122
    -9, 16, 11, 0, 12, 1, -16, -6, -20,
    -- filter=173 channel=123
    6, 5, 0, 0, 2, 2, -1, 1, 5,
    -- filter=173 channel=124
    4, -9, 2, 3, 0, 0, 0, 10, 1,
    -- filter=173 channel=125
    0, 12, 5, 6, 7, 1, 4, -13, -16,
    -- filter=173 channel=126
    -6, 6, -4, 0, 11, 17, 6, 5, 4,
    -- filter=173 channel=127
    -1, 1, 3, 4, 8, -3, 7, 5, -8,
    -- filter=174 channel=0
    3, 6, 8, -5, 13, 2, -13, -1, 4,
    -- filter=174 channel=1
    1, 8, 4, -2, 14, -3, -9, 2, 9,
    -- filter=174 channel=2
    1, -7, -2, 1, -2, 6, 3, 0, -2,
    -- filter=174 channel=3
    -1, 5, -2, -6, 6, 3, 7, 0, 9,
    -- filter=174 channel=4
    6, 2, -7, 3, 7, 7, 0, 5, 21,
    -- filter=174 channel=5
    11, 14, 2, 11, 5, -11, 0, 1, -7,
    -- filter=174 channel=6
    0, -7, 0, 0, 1, 10, 1, -3, -2,
    -- filter=174 channel=7
    2, 1, -2, -4, -5, -2, -6, -6, -4,
    -- filter=174 channel=8
    1, -7, 5, 0, 4, 3, 6, 7, 3,
    -- filter=174 channel=9
    5, -4, -4, 4, 0, -10, 3, 3, 5,
    -- filter=174 channel=10
    -7, -13, -11, 5, -6, -11, 10, 4, -1,
    -- filter=174 channel=11
    -4, 6, 0, 1, 0, -6, 2, 0, -4,
    -- filter=174 channel=12
    4, 4, -4, -9, 5, 0, 0, 3, -3,
    -- filter=174 channel=13
    3, -3, -14, 3, -5, -11, 3, 6, -3,
    -- filter=174 channel=14
    3, 7, 1, 2, 5, 2, 2, 0, 5,
    -- filter=174 channel=15
    1, -6, -5, 11, -3, -6, 12, 0, -1,
    -- filter=174 channel=16
    -3, 4, -4, 7, 5, -6, 7, 0, -10,
    -- filter=174 channel=17
    -1, 1, -6, -4, 7, -4, 0, 2, -2,
    -- filter=174 channel=18
    10, -13, -11, 9, 1, -12, -1, 12, 7,
    -- filter=174 channel=19
    2, 5, -6, 3, 7, -5, -6, 4, -6,
    -- filter=174 channel=20
    5, -5, -4, 5, 3, -4, 2, -6, -11,
    -- filter=174 channel=21
    7, 5, -14, 10, -9, -19, 18, 1, -8,
    -- filter=174 channel=22
    -4, 3, 4, 3, 5, 2, -6, 4, -1,
    -- filter=174 channel=23
    -4, -16, -9, 0, -5, -18, 17, 2, -10,
    -- filter=174 channel=24
    -4, -6, -4, 0, 0, 0, 5, 3, 0,
    -- filter=174 channel=25
    -2, -14, -11, 11, 5, -11, 2, 12, -3,
    -- filter=174 channel=26
    1, 3, -2, -4, 8, 2, -1, 0, 1,
    -- filter=174 channel=27
    -7, -15, -22, 16, -10, -24, 11, 18, -6,
    -- filter=174 channel=28
    1, 2, 4, 2, 5, -5, 7, 0, 1,
    -- filter=174 channel=29
    4, -6, 0, 6, 7, -5, 7, 4, -4,
    -- filter=174 channel=30
    6, -3, -7, 10, 3, -8, 1, 15, 4,
    -- filter=174 channel=31
    -3, -12, -25, 9, -15, -34, 13, 18, -11,
    -- filter=174 channel=32
    -4, -14, -17, 11, 4, -16, 8, 12, 2,
    -- filter=174 channel=33
    2, -6, -11, 3, 0, -17, -2, 3, -5,
    -- filter=174 channel=34
    -10, -12, 2, 0, -7, -4, 3, -6, -1,
    -- filter=174 channel=35
    2, 4, -4, -2, -6, 1, 0, -4, 5,
    -- filter=174 channel=36
    10, -3, -3, -2, 6, -6, 10, 6, 5,
    -- filter=174 channel=37
    -4, 2, -3, -7, 15, 0, -8, 8, 2,
    -- filter=174 channel=38
    8, -1, -14, 4, -8, -6, 3, 5, 1,
    -- filter=174 channel=39
    5, 6, 6, 4, 7, 0, 10, 4, 2,
    -- filter=174 channel=40
    8, 3, 0, 0, -6, 2, 10, 5, 0,
    -- filter=174 channel=41
    5, -8, 5, 1, 5, 12, -6, 2, 11,
    -- filter=174 channel=42
    4, 7, 6, 6, 4, 6, -7, -1, 10,
    -- filter=174 channel=43
    4, 0, 6, -4, -6, 6, 0, 6, 2,
    -- filter=174 channel=44
    2, -4, -15, 6, -1, -12, -1, 5, -2,
    -- filter=174 channel=45
    2, -2, 8, 6, -2, -4, -5, 6, 3,
    -- filter=174 channel=46
    -3, 7, 9, 2, 5, 0, 2, -6, 1,
    -- filter=174 channel=47
    6, 13, -6, 5, -3, -16, 11, 2, -11,
    -- filter=174 channel=48
    0, 2, -9, 4, -5, -10, 9, 9, 0,
    -- filter=174 channel=49
    6, -4, -10, -1, 1, 6, 8, 7, 11,
    -- filter=174 channel=50
    3, -4, -17, 2, -4, -10, 13, 10, 2,
    -- filter=174 channel=51
    5, -6, -6, 2, 4, -4, -5, 0, -7,
    -- filter=174 channel=52
    4, -10, 4, -3, -1, -5, 6, -1, 1,
    -- filter=174 channel=53
    4, -5, 0, 8, -7, -4, 6, 6, -3,
    -- filter=174 channel=54
    -5, -5, -4, -2, 5, 0, 0, 6, -4,
    -- filter=174 channel=55
    2, -11, -11, 9, 1, -20, 17, 11, 0,
    -- filter=174 channel=56
    -3, -3, -7, 0, -8, -1, -2, -7, 0,
    -- filter=174 channel=57
    6, 2, -3, 1, 8, -1, 0, 9, 8,
    -- filter=174 channel=58
    -3, 11, -2, -2, 11, 0, 0, 8, 3,
    -- filter=174 channel=59
    6, -7, -23, 7, 6, -19, 6, 16, 5,
    -- filter=174 channel=60
    0, -6, 5, 0, 7, 7, -1, -1, 6,
    -- filter=174 channel=61
    5, -8, 5, 7, -3, 2, 7, -2, 2,
    -- filter=174 channel=62
    -4, 4, -2, 5, -6, -1, -3, -2, -2,
    -- filter=174 channel=63
    2, 0, 1, 8, 9, -2, -4, 4, 1,
    -- filter=174 channel=64
    -3, 5, -4, -2, 1, 1, -1, -1, -3,
    -- filter=174 channel=65
    -6, 0, -1, -6, 0, -2, 0, -3, -3,
    -- filter=174 channel=66
    2, -10, -1, -5, 10, 0, 1, 0, 0,
    -- filter=174 channel=67
    0, -3, -1, -5, -4, 4, 5, 3, -1,
    -- filter=174 channel=68
    3, -3, -6, -6, -4, 7, 3, 0, 4,
    -- filter=174 channel=69
    7, 7, 4, 3, -2, 2, 0, 2, -4,
    -- filter=174 channel=70
    -7, -16, -6, -7, -1, -5, 0, 10, -2,
    -- filter=174 channel=71
    -6, 3, -5, 0, 5, -5, 4, 7, 0,
    -- filter=174 channel=72
    9, -6, -17, 9, -5, -22, 17, 11, -8,
    -- filter=174 channel=73
    -1, -11, -11, -2, 5, -9, 6, 7, 2,
    -- filter=174 channel=74
    -8, -14, -14, 4, -7, -1, 4, 1, -10,
    -- filter=174 channel=75
    5, 6, 0, 1, 2, -9, -5, 6, 7,
    -- filter=174 channel=76
    6, 4, 5, 11, 9, 7, 5, 0, 7,
    -- filter=174 channel=77
    4, 6, -6, 4, 1, -6, 3, -6, -1,
    -- filter=174 channel=78
    3, 6, 0, 0, -3, -2, 5, -2, 4,
    -- filter=174 channel=79
    -6, -11, -18, 9, 2, -22, -4, 3, 0,
    -- filter=174 channel=80
    10, 0, -14, 16, 2, -36, 18, 16, 0,
    -- filter=174 channel=81
    3, 1, -4, 0, -5, -1, -2, 5, 4,
    -- filter=174 channel=82
    -2, 0, 7, 0, -1, 1, -2, -2, 5,
    -- filter=174 channel=83
    -1, -4, -3, 2, 7, -11, 2, 9, 6,
    -- filter=174 channel=84
    7, -8, -13, -3, 4, 0, -2, 8, 0,
    -- filter=174 channel=85
    -5, -4, 4, -6, -1, 6, 3, 0, 1,
    -- filter=174 channel=86
    -7, 3, -7, 4, -5, -7, 1, -6, 2,
    -- filter=174 channel=87
    7, -1, 7, 5, 0, 6, 8, 3, -6,
    -- filter=174 channel=88
    -1, -11, 0, -3, -1, 0, 7, 5, -4,
    -- filter=174 channel=89
    0, -15, -19, 11, -11, -15, 13, 0, -10,
    -- filter=174 channel=90
    -2, 2, -4, 4, -5, -11, 1, -2, -8,
    -- filter=174 channel=91
    8, -12, -19, 4, -2, -11, 1, 3, -4,
    -- filter=174 channel=92
    -8, -5, -6, 3, 0, 6, 0, 1, 3,
    -- filter=174 channel=93
    8, 9, -5, -4, -2, -13, -3, 8, 2,
    -- filter=174 channel=94
    2, 4, 3, 2, 0, 0, 4, 7, -6,
    -- filter=174 channel=95
    -4, 5, -2, 4, -7, -5, 4, 3, 2,
    -- filter=174 channel=96
    4, 0, 4, -2, 2, -6, 1, 2, 8,
    -- filter=174 channel=97
    7, 2, 0, -6, 3, 5, 1, -5, 4,
    -- filter=174 channel=98
    3, -8, -18, 6, -3, -15, 7, 5, 4,
    -- filter=174 channel=99
    5, -21, -19, 7, -11, -25, 21, 5, -16,
    -- filter=174 channel=100
    0, 5, -4, -2, -8, 5, 4, -2, 5,
    -- filter=174 channel=101
    8, -7, -8, -4, -2, 9, 9, 9, 5,
    -- filter=174 channel=102
    6, -2, -5, 0, 1, -6, 1, 4, 7,
    -- filter=174 channel=103
    10, 12, -10, 3, 0, -14, 8, 10, -10,
    -- filter=174 channel=104
    2, 0, -26, 15, -8, -25, 13, 5, -10,
    -- filter=174 channel=105
    1, 8, 5, 8, -2, 5, -4, 4, -6,
    -- filter=174 channel=106
    -2, 2, 6, 8, 3, 9, 5, 5, 7,
    -- filter=174 channel=107
    -3, -2, -4, 7, 7, 8, 0, -7, -2,
    -- filter=174 channel=108
    9, 1, 4, -3, 5, 0, 5, 0, 0,
    -- filter=174 channel=109
    5, -15, -17, 2, 3, -23, 14, 2, -9,
    -- filter=174 channel=110
    -2, 1, -9, 6, -4, -7, 7, 4, -2,
    -- filter=174 channel=111
    8, -3, -4, 8, -1, 6, 3, 0, -3,
    -- filter=174 channel=112
    -6, -5, -9, 2, 2, -6, 0, 8, 1,
    -- filter=174 channel=113
    0, -1, 0, 8, -2, -17, 9, 8, 1,
    -- filter=174 channel=114
    -4, -9, -17, -2, 14, -6, -1, 8, 9,
    -- filter=174 channel=115
    7, -4, 7, 6, 4, -2, 0, 0, -5,
    -- filter=174 channel=116
    2, -15, -21, 8, 7, -21, 16, 7, 9,
    -- filter=174 channel=117
    -4, -4, 1, 0, -4, -8, 7, -3, 5,
    -- filter=174 channel=118
    0, -4, 3, -1, 7, -2, -5, -1, 8,
    -- filter=174 channel=119
    -6, -11, -4, -7, -5, 4, 2, -2, -10,
    -- filter=174 channel=120
    0, -10, -18, 2, -6, -19, 2, 9, -12,
    -- filter=174 channel=121
    2, -6, -1, -2, -1, -5, 0, -4, -6,
    -- filter=174 channel=122
    8, 10, -21, 6, -10, -31, 15, 1, -9,
    -- filter=174 channel=123
    3, -5, 7, -4, -3, -1, 2, -6, -1,
    -- filter=174 channel=124
    6, -5, -3, -3, 0, -2, -5, 0, -3,
    -- filter=174 channel=125
    5, -5, -21, 14, -2, -19, 17, 3, -13,
    -- filter=174 channel=126
    3, 0, -1, -5, 1, -13, -2, 4, 3,
    -- filter=174 channel=127
    1, -6, -5, -1, 6, -1, 5, 0, 4,
    -- filter=175 channel=0
    -3, 8, -9, 2, 13, 3, 0, 8, 0,
    -- filter=175 channel=1
    3, -3, 0, 2, 2, 0, 5, 4, 2,
    -- filter=175 channel=2
    1, -5, 8, -5, -5, 2, -6, -5, -6,
    -- filter=175 channel=3
    -4, -10, 3, -9, -3, 8, 6, 4, 6,
    -- filter=175 channel=4
    2, -7, 6, 3, 0, 5, -7, 3, 7,
    -- filter=175 channel=5
    -6, -8, -6, 9, 9, 3, -2, 1, -1,
    -- filter=175 channel=6
    3, -6, -7, 10, 7, 0, 5, 9, -1,
    -- filter=175 channel=7
    -5, 3, -5, 2, -3, 7, 2, 6, 5,
    -- filter=175 channel=8
    2, -7, 0, 3, -5, 9, 2, 2, -2,
    -- filter=175 channel=9
    3, -1, 0, -5, -5, 4, 0, -5, -4,
    -- filter=175 channel=10
    10, 3, 3, 2, 2, 0, -12, -10, 2,
    -- filter=175 channel=11
    2, 0, -4, 2, 0, -4, 4, 3, -5,
    -- filter=175 channel=12
    0, -3, -3, -2, 0, 8, -3, -2, -1,
    -- filter=175 channel=13
    -3, -4, -2, 2, -7, 6, 3, 1, 3,
    -- filter=175 channel=14
    0, -2, -1, 0, 5, -7, 0, -3, -6,
    -- filter=175 channel=15
    0, 0, -12, 10, 6, 0, 9, 11, -6,
    -- filter=175 channel=16
    -10, 0, 7, -1, -10, -4, -6, -7, 2,
    -- filter=175 channel=17
    -3, 5, 7, 7, -3, 1, -2, 2, -4,
    -- filter=175 channel=18
    0, 3, -8, 3, 16, -5, 14, 20, 2,
    -- filter=175 channel=19
    0, -2, 0, 0, 5, -5, 6, -2, 5,
    -- filter=175 channel=20
    0, -12, -15, 11, -6, -8, 3, 9, -5,
    -- filter=175 channel=21
    -4, -13, 7, -15, -20, 6, -11, -24, -1,
    -- filter=175 channel=22
    0, 5, 5, 7, 4, 4, 8, 2, 7,
    -- filter=175 channel=23
    5, 0, -9, 6, -7, -3, 6, 0, 6,
    -- filter=175 channel=24
    -2, 4, 1, -4, -6, -5, 5, 4, 2,
    -- filter=175 channel=25
    -3, -5, 2, -3, -3, 7, 4, 1, -5,
    -- filter=175 channel=26
    -9, -6, 0, 1, -10, -4, -3, -3, -6,
    -- filter=175 channel=27
    8, 3, 9, -2, 2, 13, -5, 0, 12,
    -- filter=175 channel=28
    2, 5, 0, -3, 3, 1, -4, 3, -3,
    -- filter=175 channel=29
    -9, -15, -19, 0, 7, -19, 10, 1, -14,
    -- filter=175 channel=30
    0, -7, -2, -3, 2, -4, -2, -7, 2,
    -- filter=175 channel=31
    -9, -9, 6, -30, -20, 5, -22, -25, -4,
    -- filter=175 channel=32
    -4, -3, -1, -1, 6, -3, 0, 9, -5,
    -- filter=175 channel=33
    4, -1, -8, 4, 1, 0, 0, 9, 7,
    -- filter=175 channel=34
    13, 8, 0, 9, 6, 11, 5, 3, 9,
    -- filter=175 channel=35
    4, 1, 7, 7, 1, -6, 7, 3, -1,
    -- filter=175 channel=36
    5, -2, 3, -5, -3, 7, -4, -10, 6,
    -- filter=175 channel=37
    -4, 0, -4, 1, 8, 3, 3, -5, 0,
    -- filter=175 channel=38
    2, -4, 1, -2, -4, -1, -8, 0, 7,
    -- filter=175 channel=39
    -7, -8, -5, 2, 2, -14, 1, 5, -8,
    -- filter=175 channel=40
    3, 1, -4, 6, -4, -5, 4, 9, 4,
    -- filter=175 channel=41
    9, 8, -7, 10, -6, 0, 7, -5, 5,
    -- filter=175 channel=42
    -6, 5, -8, -10, 1, -5, -1, -3, 2,
    -- filter=175 channel=43
    -1, -7, -4, 11, 2, -3, 0, 4, 8,
    -- filter=175 channel=44
    -2, -5, 3, -2, -13, -1, -8, -10, 3,
    -- filter=175 channel=45
    -8, -4, -5, 2, 3, -5, 4, 2, -2,
    -- filter=175 channel=46
    7, 6, 7, 4, 7, 2, -1, 6, 4,
    -- filter=175 channel=47
    -3, -14, -1, -12, -17, 2, -21, -16, -13,
    -- filter=175 channel=48
    -12, 0, 11, -10, -16, -2, -9, -9, 1,
    -- filter=175 channel=49
    -6, 1, -6, -2, 5, 0, 7, 1, -10,
    -- filter=175 channel=50
    6, -2, 10, -2, 0, -2, -7, 0, 2,
    -- filter=175 channel=51
    4, 5, 3, -3, 0, 4, -1, -2, 3,
    -- filter=175 channel=52
    -5, 4, -3, 8, 3, 8, 6, -5, 6,
    -- filter=175 channel=53
    -3, 1, 0, -2, -3, -8, 5, 2, 2,
    -- filter=175 channel=54
    -5, -1, -5, -3, 4, 6, -7, 4, 6,
    -- filter=175 channel=55
    1, 0, -8, 7, 8, -10, 4, 5, -4,
    -- filter=175 channel=56
    5, 6, 0, -1, -3, 7, 4, 0, -1,
    -- filter=175 channel=57
    0, -3, -7, -1, -1, -1, 6, 5, -4,
    -- filter=175 channel=58
    0, -2, 0, 0, 3, -7, 6, 1, 6,
    -- filter=175 channel=59
    -6, 2, 9, -2, -6, 8, -5, -5, 5,
    -- filter=175 channel=60
    1, -6, -1, -6, -7, 0, -6, -6, -6,
    -- filter=175 channel=61
    -2, 5, -5, 2, 1, 4, 6, -2, 5,
    -- filter=175 channel=62
    0, 2, 6, -5, -1, 0, 1, -6, 0,
    -- filter=175 channel=63
    -4, -5, -1, -1, -1, 2, -6, -3, 0,
    -- filter=175 channel=64
    5, -1, 2, -3, -1, 0, -6, 5, 8,
    -- filter=175 channel=65
    -1, 0, 5, 0, 4, -4, 7, -3, 4,
    -- filter=175 channel=66
    -3, -2, 6, -2, -5, 0, 0, 7, 0,
    -- filter=175 channel=67
    -2, -5, -2, 2, 5, -2, -1, 1, -1,
    -- filter=175 channel=68
    3, -6, -5, 2, 1, 0, -5, 4, -5,
    -- filter=175 channel=69
    -5, 2, 1, -7, 6, 0, 1, -1, -1,
    -- filter=175 channel=70
    11, 9, 13, 3, 12, 5, -2, 4, 3,
    -- filter=175 channel=71
    2, -6, -4, 0, -1, 0, 0, -1, 3,
    -- filter=175 channel=72
    0, 5, 5, -15, -5, 3, -10, -9, -2,
    -- filter=175 channel=73
    -1, -4, -6, 4, 1, 4, -3, 5, 2,
    -- filter=175 channel=74
    -1, -2, 6, 0, 0, 4, 3, -11, 13,
    -- filter=175 channel=75
    -8, -6, -4, 5, 9, 5, -4, -1, -6,
    -- filter=175 channel=76
    -3, -3, -17, 0, 10, -8, -1, 4, -10,
    -- filter=175 channel=77
    6, 0, -2, -1, -2, 1, 0, -1, -1,
    -- filter=175 channel=78
    6, 0, -6, 7, -9, -3, -6, -8, -2,
    -- filter=175 channel=79
    2, 7, -12, 12, 21, -3, 11, 17, 7,
    -- filter=175 channel=80
    -11, -1, 14, -21, -16, -2, -21, -20, 0,
    -- filter=175 channel=81
    4, -1, 3, -5, 6, -1, -6, 6, -4,
    -- filter=175 channel=82
    -3, 0, 6, 3, 0, -6, -3, 0, 6,
    -- filter=175 channel=83
    -6, 3, 4, -7, -2, 3, -6, -1, 1,
    -- filter=175 channel=84
    2, -3, 0, 4, 9, 2, 7, 2, -1,
    -- filter=175 channel=85
    0, 7, -5, 1, -6, -2, -3, 6, 3,
    -- filter=175 channel=86
    0, 0, -2, 4, -3, 4, 12, 3, 0,
    -- filter=175 channel=87
    -1, -11, -5, -1, 7, 0, 10, -3, -1,
    -- filter=175 channel=88
    5, 3, 14, -3, -9, 3, 0, -9, 6,
    -- filter=175 channel=89
    0, -1, -2, -9, -5, 2, -2, -1, 5,
    -- filter=175 channel=90
    -7, 6, 13, -6, -6, 10, 0, -4, 1,
    -- filter=175 channel=91
    2, 2, -4, 0, 7, -4, 6, -3, 0,
    -- filter=175 channel=92
    4, -7, 8, 0, -1, -1, 6, 2, 6,
    -- filter=175 channel=93
    -8, 0, 7, 0, -8, -7, -2, -1, 5,
    -- filter=175 channel=94
    -5, -1, 1, 0, 1, 0, 2, -6, 0,
    -- filter=175 channel=95
    -6, 6, 2, -4, 1, 0, -1, 6, 6,
    -- filter=175 channel=96
    4, 1, 0, 0, -2, -8, -6, 7, 2,
    -- filter=175 channel=97
    5, -6, 5, -3, -7, 2, 0, 2, 6,
    -- filter=175 channel=98
    3, 0, -5, -10, -10, 4, -12, -1, 2,
    -- filter=175 channel=99
    -7, -2, 7, -2, -15, 0, -5, -10, -1,
    -- filter=175 channel=100
    5, 5, 1, 8, 8, 9, 0, 2, 0,
    -- filter=175 channel=101
    -1, -3, 1, -9, -3, 8, -3, -8, 4,
    -- filter=175 channel=102
    0, 3, -2, 1, 2, -4, -3, -2, -1,
    -- filter=175 channel=103
    0, -3, 5, -14, -7, 1, -23, -10, -12,
    -- filter=175 channel=104
    -2, 0, 6, -17, -21, -2, -8, -15, -6,
    -- filter=175 channel=105
    1, -10, -12, 3, 8, -13, 10, 7, -7,
    -- filter=175 channel=106
    -7, 0, -5, 3, 0, 1, 3, -4, 5,
    -- filter=175 channel=107
    0, -3, -15, 5, 2, -9, 16, 6, 5,
    -- filter=175 channel=108
    7, 0, -3, 0, 0, 5, 9, 6, -1,
    -- filter=175 channel=109
    1, 3, -1, -4, -4, 1, 2, -2, 10,
    -- filter=175 channel=110
    0, 4, -7, 0, -8, 4, -7, -7, 0,
    -- filter=175 channel=111
    -3, -1, -6, 8, 4, -2, 2, 0, 3,
    -- filter=175 channel=112
    -2, -4, 2, -6, 3, -1, -2, -8, 0,
    -- filter=175 channel=113
    9, 3, 0, 4, 5, 9, 2, -9, 10,
    -- filter=175 channel=114
    -4, 6, -6, 19, 24, -9, 14, 26, 1,
    -- filter=175 channel=115
    -1, 0, -5, 1, -6, -4, 8, 0, 0,
    -- filter=175 channel=116
    -1, -8, 3, -9, 2, 1, 0, -8, -2,
    -- filter=175 channel=117
    -4, 1, 1, 2, -2, 3, -6, -3, 6,
    -- filter=175 channel=118
    -4, -1, 1, 6, -3, 0, -3, -3, -4,
    -- filter=175 channel=119
    10, 0, 12, 1, 3, 18, 12, 8, 16,
    -- filter=175 channel=120
    -12, -9, 1, -8, -8, 6, 4, 0, 8,
    -- filter=175 channel=121
    4, 1, -2, -1, -4, 8, 3, 4, 0,
    -- filter=175 channel=122
    -21, -19, 12, -26, -27, 0, -25, -21, -13,
    -- filter=175 channel=123
    5, 4, 10, -4, 6, 12, -5, 0, 10,
    -- filter=175 channel=124
    -3, -2, -5, 2, 0, -4, 5, 1, -3,
    -- filter=175 channel=125
    -2, -8, 5, -2, -15, 8, -12, -14, 1,
    -- filter=175 channel=126
    0, 5, 2, 0, -7, 4, -1, -4, 5,
    -- filter=175 channel=127
    -2, 4, 1, -4, -5, -1, -2, 1, 5,
    -- filter=176 channel=0
    -17, 21, 12, -35, 20, 19, -38, -15, -2,
    -- filter=176 channel=1
    -10, 20, 4, -29, 15, 18, -20, -14, -11,
    -- filter=176 channel=2
    -4, -3, 4, -1, -6, -4, 4, 5, -2,
    -- filter=176 channel=3
    -19, -11, 9, -7, -3, 0, -12, 0, 10,
    -- filter=176 channel=4
    -6, -5, 14, -19, -10, 1, -7, 9, 19,
    -- filter=176 channel=5
    -9, 29, 3, -17, 32, 17, -32, 4, -5,
    -- filter=176 channel=6
    1, 1, 3, -4, -3, 3, 3, -1, 13,
    -- filter=176 channel=7
    4, 6, 0, 6, 0, -4, -2, 6, 0,
    -- filter=176 channel=8
    -6, 0, -5, 1, -4, 5, 1, -9, 6,
    -- filter=176 channel=9
    -1, -1, 4, 4, 13, 1, -8, 0, -6,
    -- filter=176 channel=10
    4, 0, -4, 6, -6, 0, 6, -2, 9,
    -- filter=176 channel=11
    -7, -18, -1, -5, -10, 6, 4, 16, 16,
    -- filter=176 channel=12
    8, -4, 0, 4, 0, -9, -7, 1, -4,
    -- filter=176 channel=13
    0, -14, 0, 3, -10, -10, -1, 2, 7,
    -- filter=176 channel=14
    5, 0, -1, -3, 3, 3, -1, -1, -2,
    -- filter=176 channel=15
    -1, -2, 0, 5, -9, -12, 14, 2, 7,
    -- filter=176 channel=16
    -4, 1, 5, -12, 13, 11, -18, -10, -9,
    -- filter=176 channel=17
    3, -3, 1, 0, 5, 0, -4, 4, 5,
    -- filter=176 channel=18
    10, 9, -10, -2, -9, -13, 10, -1, 2,
    -- filter=176 channel=19
    -1, 1, 6, -1, -6, -6, 6, -6, 4,
    -- filter=176 channel=20
    3, -14, 4, 6, -20, -3, 20, 6, 34,
    -- filter=176 channel=21
    -4, 3, 7, -5, 19, 2, -6, 0, -15,
    -- filter=176 channel=22
    -2, 4, -3, 1, 6, -9, 0, 5, -1,
    -- filter=176 channel=23
    0, -13, -5, 4, -27, -11, 9, -4, 14,
    -- filter=176 channel=24
    -3, -1, -5, -7, 2, 0, 1, -6, 5,
    -- filter=176 channel=25
    8, 13, 3, -6, 15, 0, -1, 0, -12,
    -- filter=176 channel=26
    1, 7, 10, -10, 12, 4, -17, 3, -6,
    -- filter=176 channel=27
    -6, 10, -3, -6, 12, -8, -2, -2, -5,
    -- filter=176 channel=28
    -3, 6, 5, 5, 3, 6, -4, 2, -2,
    -- filter=176 channel=29
    -10, -8, 1, 3, -18, -4, 13, 20, 36,
    -- filter=176 channel=30
    0, 3, 10, -13, 17, 12, -11, -2, -2,
    -- filter=176 channel=31
    0, -5, 2, 4, 0, 11, -6, -2, 7,
    -- filter=176 channel=32
    0, -3, -5, -10, 3, -11, 4, 5, 7,
    -- filter=176 channel=33
    -3, 10, 3, -1, 3, 0, -9, -11, -6,
    -- filter=176 channel=34
    0, 3, -5, 4, 0, -3, 7, -5, -16,
    -- filter=176 channel=35
    -7, 0, 6, -4, -5, 4, -7, -2, 5,
    -- filter=176 channel=36
    -1, -21, -12, -4, -5, 0, 4, -8, -1,
    -- filter=176 channel=37
    -12, 21, 4, -35, 13, 15, -33, -10, -15,
    -- filter=176 channel=38
    -2, 6, -6, -3, 2, -2, -7, 0, -2,
    -- filter=176 channel=39
    4, -1, -2, -5, -13, -1, 4, 11, 20,
    -- filter=176 channel=40
    -10, -10, 1, 2, -4, -11, 0, 2, 7,
    -- filter=176 channel=41
    1, 4, 2, 7, 10, -14, -1, 2, -16,
    -- filter=176 channel=42
    0, 2, 13, -15, 2, 8, -15, -3, 6,
    -- filter=176 channel=43
    -8, 0, -5, -7, 3, -6, 0, -2, 3,
    -- filter=176 channel=44
    -12, 14, 9, -21, 15, 11, -19, -13, -9,
    -- filter=176 channel=45
    -8, 0, 7, 1, 5, 9, -3, 5, 3,
    -- filter=176 channel=46
    -4, -2, -2, 7, 0, -8, -5, -4, -4,
    -- filter=176 channel=47
    -12, 5, 0, -9, 26, 10, -22, 1, -14,
    -- filter=176 channel=48
    0, 6, 11, -11, 19, 9, -11, -1, -2,
    -- filter=176 channel=49
    3, -9, 0, 3, -14, -4, 7, 8, 10,
    -- filter=176 channel=50
    -5, 6, 1, 0, 5, -2, -3, 5, -9,
    -- filter=176 channel=51
    7, 1, 5, 6, -3, -7, 0, -4, 4,
    -- filter=176 channel=52
    1, -6, -6, -4, -10, -10, 3, 2, 5,
    -- filter=176 channel=53
    1, 0, -5, 5, -12, -2, 10, -1, 19,
    -- filter=176 channel=54
    0, 3, -2, 0, -6, 0, -4, 3, 7,
    -- filter=176 channel=55
    1, -7, -17, 15, -21, -24, 21, 13, 12,
    -- filter=176 channel=56
    -2, 0, 0, -2, 3, -5, -5, -2, -11,
    -- filter=176 channel=57
    4, -4, 0, 4, -3, 2, 3, 5, 5,
    -- filter=176 channel=58
    -9, 15, 15, -16, 12, 17, -12, -6, 7,
    -- filter=176 channel=59
    10, 11, 4, 0, 18, -1, -6, 3, -7,
    -- filter=176 channel=60
    2, 5, 7, -4, 7, 7, -7, 5, -5,
    -- filter=176 channel=61
    -1, -2, -4, 0, -2, 4, 0, 4, 1,
    -- filter=176 channel=62
    -8, 0, 6, 0, -7, -3, -7, 0, 6,
    -- filter=176 channel=63
    -3, 13, 16, -4, 9, 17, -17, -7, -5,
    -- filter=176 channel=64
    1, -6, -10, -5, -5, -7, 10, 11, 2,
    -- filter=176 channel=65
    0, 0, 0, -5, 6, 6, -1, -3, 6,
    -- filter=176 channel=66
    8, 3, 0, 0, 6, -1, 0, -5, 5,
    -- filter=176 channel=67
    -1, -2, 2, -1, -5, -5, -1, -1, -5,
    -- filter=176 channel=68
    -3, -8, -6, 3, -11, 0, 6, -5, 1,
    -- filter=176 channel=69
    1, 3, 3, -3, 6, 0, 5, 0, 4,
    -- filter=176 channel=70
    -6, 4, -6, 6, -16, -12, 0, -9, -12,
    -- filter=176 channel=71
    4, 2, -5, -3, 3, 1, -3, -8, -3,
    -- filter=176 channel=72
    -2, -14, -4, 15, -5, 5, 7, -2, -1,
    -- filter=176 channel=73
    -4, 0, -1, 4, -15, -15, 11, 5, 2,
    -- filter=176 channel=74
    -6, 8, -4, 5, -5, 0, -7, -5, -10,
    -- filter=176 channel=75
    -8, 24, 20, -22, 24, 18, -27, -11, -11,
    -- filter=176 channel=76
    9, -11, -3, 9, -9, -14, 14, 16, 24,
    -- filter=176 channel=77
    2, -2, 5, 1, -1, 7, -5, 0, 7,
    -- filter=176 channel=78
    -13, 8, 10, -13, 2, 8, -8, 3, 6,
    -- filter=176 channel=79
    7, 6, -6, 6, -9, -9, -5, 7, 1,
    -- filter=176 channel=80
    1, 2, 10, -3, 22, 14, 0, 2, 9,
    -- filter=176 channel=81
    6, -2, 6, 4, 4, 0, -7, 0, 3,
    -- filter=176 channel=82
    0, 0, 0, 4, -3, 2, -5, -7, -1,
    -- filter=176 channel=83
    1, 2, 3, 7, 9, -4, 3, 11, 7,
    -- filter=176 channel=84
    7, -5, -2, -3, -11, -9, 3, 2, 6,
    -- filter=176 channel=85
    3, 2, -4, 5, 2, 5, -6, 0, 4,
    -- filter=176 channel=86
    1, 2, -7, -6, 2, -2, -1, -10, -7,
    -- filter=176 channel=87
    -3, -11, 4, 2, -16, -7, 0, 4, 8,
    -- filter=176 channel=88
    -7, -9, -12, 5, 1, -1, 0, 2, 4,
    -- filter=176 channel=89
    -2, -12, -1, 5, -13, -10, 0, 0, -4,
    -- filter=176 channel=90
    -2, -6, -10, -4, -19, -4, 0, -4, -6,
    -- filter=176 channel=91
    4, -7, -10, 0, -19, -12, 6, 0, -2,
    -- filter=176 channel=92
    -4, 3, 0, -3, -7, -7, 0, -8, 1,
    -- filter=176 channel=93
    -16, 14, 16, -14, 15, 25, -29, -6, -2,
    -- filter=176 channel=94
    4, -4, 4, -1, -5, 5, -2, -4, -4,
    -- filter=176 channel=95
    0, -4, -4, 2, 0, -5, 3, -6, 5,
    -- filter=176 channel=96
    -7, -5, 8, -4, -2, 0, -5, -4, -1,
    -- filter=176 channel=97
    -8, 5, 1, -1, -9, 1, -4, -1, 2,
    -- filter=176 channel=98
    -1, 9, 9, -1, 17, 9, -13, 0, 4,
    -- filter=176 channel=99
    -1, -9, -5, 15, -3, -1, 6, -2, 6,
    -- filter=176 channel=100
    0, -1, -6, -2, -3, -1, -4, -4, -2,
    -- filter=176 channel=101
    0, -10, 1, -14, -15, 3, 0, 0, 8,
    -- filter=176 channel=102
    -2, 1, 4, 6, 5, 2, 1, 1, 5,
    -- filter=176 channel=103
    -15, 5, 2, -18, 22, 20, -24, -8, -14,
    -- filter=176 channel=104
    1, 3, -1, 7, 12, 2, 3, 9, 0,
    -- filter=176 channel=105
    -4, 0, 6, 5, -13, 6, 7, 7, 20,
    -- filter=176 channel=106
    1, -4, 0, -1, -6, -1, 11, -3, 9,
    -- filter=176 channel=107
    -13, -4, -4, -5, -14, -13, -1, 1, 5,
    -- filter=176 channel=108
    -1, 0, 6, 0, 10, 0, -5, 2, 2,
    -- filter=176 channel=109
    8, 17, -3, 6, 11, -13, 0, 6, -5,
    -- filter=176 channel=110
    0, -1, -1, -6, -11, 10, 3, -2, 10,
    -- filter=176 channel=111
    1, 9, 4, 3, -1, 0, 6, 9, 4,
    -- filter=176 channel=112
    -5, 11, 3, -6, 9, 6, -9, -5, -14,
    -- filter=176 channel=113
    -4, -1, -3, -3, 5, 2, 2, -7, -7,
    -- filter=176 channel=114
    0, 26, 5, -22, 12, -4, -8, 0, -3,
    -- filter=176 channel=115
    -1, 6, 2, 0, 5, 0, 0, 6, 1,
    -- filter=176 channel=116
    -2, -5, -6, -3, 5, -7, 13, 7, 10,
    -- filter=176 channel=117
    -2, 3, 3, 1, -5, -1, 2, -3, -6,
    -- filter=176 channel=118
    -2, -5, 4, -2, 2, 3, 1, -4, 0,
    -- filter=176 channel=119
    6, 6, -10, 5, 0, -21, 0, -6, -20,
    -- filter=176 channel=120
    -7, 0, -3, 8, -9, -7, 14, 15, 6,
    -- filter=176 channel=121
    4, -2, -4, 2, 0, -12, 3, -4, -11,
    -- filter=176 channel=122
    -16, 14, 2, -14, 28, 9, -26, -13, -31,
    -- filter=176 channel=123
    -3, 0, -6, 6, 1, -1, 4, 4, 0,
    -- filter=176 channel=124
    -3, -3, 7, 0, -12, -4, 0, 9, 21,
    -- filter=176 channel=125
    -2, -3, 4, 1, 6, 8, 9, 7, 11,
    -- filter=176 channel=126
    2, 1, 5, 2, 7, -2, -8, 0, 0,
    -- filter=176 channel=127
    -5, 1, 2, 0, 5, 1, 6, 0, -6,
    -- filter=177 channel=0
    3, 0, 6, 0, -16, 11, 2, -7, 9,
    -- filter=177 channel=1
    3, 5, 1, -6, -12, 6, -2, 3, 2,
    -- filter=177 channel=2
    1, -7, -2, 0, -5, -3, -7, -9, -7,
    -- filter=177 channel=3
    -13, -13, 6, -13, -5, -2, 3, -6, 3,
    -- filter=177 channel=4
    -3, 0, -2, -17, -20, -10, -6, -12, -2,
    -- filter=177 channel=5
    -2, -9, -4, -12, -3, 3, -13, -4, 0,
    -- filter=177 channel=6
    -2, 0, 8, 0, -9, 4, -11, -12, -1,
    -- filter=177 channel=7
    1, 2, 1, 3, 5, -4, -4, 7, -1,
    -- filter=177 channel=8
    5, 1, -3, -13, -12, -5, -1, 0, -7,
    -- filter=177 channel=9
    6, 0, -7, 11, 4, -8, -4, 5, 2,
    -- filter=177 channel=10
    -5, -2, -3, 14, 2, -3, 8, 0, 0,
    -- filter=177 channel=11
    0, -7, 11, 6, -2, 7, 4, -6, 5,
    -- filter=177 channel=12
    -3, -7, 4, -2, -8, 1, -8, 0, 3,
    -- filter=177 channel=13
    3, 0, 11, 6, -11, 11, 3, -13, -4,
    -- filter=177 channel=14
    -7, -1, 0, -3, 5, -2, -1, 1, 5,
    -- filter=177 channel=15
    6, -4, 8, 7, -8, 12, 0, -11, 6,
    -- filter=177 channel=16
    1, -4, 1, 0, -3, -4, 0, -3, 2,
    -- filter=177 channel=17
    6, -5, 2, -3, 2, -4, 1, -6, -7,
    -- filter=177 channel=18
    0, -11, 7, 9, -13, 14, 5, -11, 16,
    -- filter=177 channel=19
    3, -4, 6, 0, 7, -3, 1, 7, -2,
    -- filter=177 channel=20
    -10, -7, 2, -8, -16, 5, -7, -10, 4,
    -- filter=177 channel=21
    3, 13, -12, 19, 18, -3, 10, 11, -11,
    -- filter=177 channel=22
    -8, -8, 8, -11, -1, 5, -3, -1, 9,
    -- filter=177 channel=23
    -1, 4, 11, 13, -14, 13, -7, -1, 7,
    -- filter=177 channel=24
    1, -4, 0, 3, -6, 1, 0, 0, -4,
    -- filter=177 channel=25
    7, -11, 0, 18, -12, -3, -5, -2, -3,
    -- filter=177 channel=26
    4, -4, 1, 3, -2, -11, 1, 0, 2,
    -- filter=177 channel=27
    7, 2, 14, 16, -8, 9, -7, -5, 10,
    -- filter=177 channel=28
    -1, -6, 4, 0, -4, -4, 6, 0, 4,
    -- filter=177 channel=29
    0, -12, 10, -4, -22, -12, -5, -11, -3,
    -- filter=177 channel=30
    -5, -1, 2, 8, -11, -4, 2, -3, -2,
    -- filter=177 channel=31
    11, 13, -7, 20, 9, 0, 0, 3, -19,
    -- filter=177 channel=32
    0, -4, 8, 3, -15, 14, -2, -14, 2,
    -- filter=177 channel=33
    5, 1, 1, 3, -3, 7, 6, 0, 12,
    -- filter=177 channel=34
    -9, -4, 11, -11, -18, -6, -10, -10, 6,
    -- filter=177 channel=35
    -2, -6, 3, 1, 2, -7, -1, -1, 6,
    -- filter=177 channel=36
    5, 3, 1, 5, -1, -13, -6, -8, -12,
    -- filter=177 channel=37
    -1, 1, 7, -5, -12, 0, -2, 6, 16,
    -- filter=177 channel=38
    5, 3, -3, 13, 0, 3, 5, -1, 0,
    -- filter=177 channel=39
    -8, -5, -4, -5, 1, -1, 1, -6, 0,
    -- filter=177 channel=40
    0, -2, 7, 2, 7, 4, -1, 0, 8,
    -- filter=177 channel=41
    -4, -2, 2, -9, -7, -17, 0, -24, 3,
    -- filter=177 channel=42
    5, 7, -5, 5, 0, 4, 0, 7, 3,
    -- filter=177 channel=43
    -13, -7, 3, -8, -5, 7, 0, -7, 9,
    -- filter=177 channel=44
    4, 0, -5, 9, 3, 1, 0, -6, 7,
    -- filter=177 channel=45
    -1, 5, 2, 4, -5, 5, 4, 4, 7,
    -- filter=177 channel=46
    -2, 4, 4, -1, -4, -5, 5, -1, 3,
    -- filter=177 channel=47
    0, 9, -2, 11, 7, -13, -5, 3, -10,
    -- filter=177 channel=48
    9, 1, 0, 10, 10, -6, -6, 3, 1,
    -- filter=177 channel=49
    -5, 1, 2, -3, -3, 2, -1, -1, 3,
    -- filter=177 channel=50
    11, -6, 0, 11, 0, 11, 6, 1, 2,
    -- filter=177 channel=51
    5, -4, 1, 2, -5, 2, -4, -6, -7,
    -- filter=177 channel=52
    -3, 0, 11, -9, -5, 2, 0, 1, 7,
    -- filter=177 channel=53
    -3, 3, -1, -1, 0, -3, -2, -6, -7,
    -- filter=177 channel=54
    3, 3, 3, 2, -1, 7, -3, 6, -6,
    -- filter=177 channel=55
    3, -12, 4, 8, -8, -1, 9, -4, 7,
    -- filter=177 channel=56
    1, -2, 1, -2, 2, 4, -10, 4, -6,
    -- filter=177 channel=57
    -5, 6, 1, 0, -2, -7, 3, -7, -1,
    -- filter=177 channel=58
    -12, 0, -3, -10, 0, -3, -11, -4, 4,
    -- filter=177 channel=59
    11, 1, -6, 15, 1, -5, 5, -9, -1,
    -- filter=177 channel=60
    -5, -2, 7, 5, -3, 1, 5, -6, 0,
    -- filter=177 channel=61
    6, -5, 2, 2, -1, -1, -3, 1, -6,
    -- filter=177 channel=62
    0, -3, -1, -8, 0, 3, 0, -4, -5,
    -- filter=177 channel=63
    -2, 4, -7, -1, 0, -8, -6, -10, 1,
    -- filter=177 channel=64
    -6, -6, 2, 0, 7, -2, 0, 7, 4,
    -- filter=177 channel=65
    2, -2, -2, -1, 1, -5, -1, -6, -3,
    -- filter=177 channel=66
    -10, -5, 2, 1, -16, -7, -7, -9, 3,
    -- filter=177 channel=67
    -7, -6, 4, -2, -2, 0, 3, -2, 5,
    -- filter=177 channel=68
    -1, -6, -6, 3, 5, 0, -2, 6, 4,
    -- filter=177 channel=69
    -1, -2, 3, 2, -3, -6, 0, -8, 5,
    -- filter=177 channel=70
    10, -1, 12, 5, -4, 18, 1, -3, 18,
    -- filter=177 channel=71
    2, 0, -2, -3, 0, 5, 9, 7, 2,
    -- filter=177 channel=72
    11, 0, -7, 26, 6, 0, 14, -7, -4,
    -- filter=177 channel=73
    -3, 0, 4, 4, -7, 5, -6, 0, 0,
    -- filter=177 channel=74
    4, 5, -3, 1, -16, 9, -9, -5, 4,
    -- filter=177 channel=75
    -9, 1, 7, 0, -3, 1, -5, -6, 1,
    -- filter=177 channel=76
    1, -5, 0, 2, -6, 4, -6, -8, 0,
    -- filter=177 channel=77
    3, -2, 5, 2, 2, 3, 5, 3, 0,
    -- filter=177 channel=78
    -3, 0, 1, -7, 0, -6, -10, -1, -3,
    -- filter=177 channel=79
    2, -17, 17, 10, -18, 21, -2, -12, 16,
    -- filter=177 channel=80
    5, -1, -14, 23, 7, -4, 11, -4, -8,
    -- filter=177 channel=81
    3, 1, 0, -1, 0, 0, 7, -4, -7,
    -- filter=177 channel=82
    4, 0, 8, 0, 3, 3, -4, 3, 6,
    -- filter=177 channel=83
    7, -3, 3, 0, 4, 1, 1, 5, -2,
    -- filter=177 channel=84
    4, -1, 8, -2, -9, 11, -10, -12, -2,
    -- filter=177 channel=85
    6, 0, 4, 2, -7, -4, 5, 2, 3,
    -- filter=177 channel=86
    -12, -1, 2, -12, -5, 4, -9, -1, -2,
    -- filter=177 channel=87
    -13, -8, 5, -12, -15, -4, -13, -8, 2,
    -- filter=177 channel=88
    2, 3, 4, 0, 10, -7, 1, -1, -1,
    -- filter=177 channel=89
    11, -5, -3, 21, -1, 0, 12, -8, 0,
    -- filter=177 channel=90
    -7, 7, -2, 2, 9, -2, -6, 5, -6,
    -- filter=177 channel=91
    10, -6, 10, 11, -7, 16, 0, 3, -1,
    -- filter=177 channel=92
    -7, 7, -2, -10, -4, -1, -2, 5, -5,
    -- filter=177 channel=93
    6, 0, -6, 6, 5, -3, -12, -9, 0,
    -- filter=177 channel=94
    -2, -4, 7, 2, -6, 7, -4, 3, 5,
    -- filter=177 channel=95
    -8, 3, 0, -2, -2, 6, -3, -3, 4,
    -- filter=177 channel=96
    0, 3, 5, 6, 7, -4, 4, -5, -6,
    -- filter=177 channel=97
    -2, 8, 2, 0, 0, 7, 3, -1, -2,
    -- filter=177 channel=98
    0, -16, -2, 17, -15, -1, 3, -5, -4,
    -- filter=177 channel=99
    -3, -5, -1, 11, 1, -3, -4, -4, -9,
    -- filter=177 channel=100
    3, -2, 7, -5, 8, -3, -9, 0, -8,
    -- filter=177 channel=101
    -3, 0, 0, -2, -4, -3, -7, -1, -5,
    -- filter=177 channel=102
    -2, 2, 0, 1, 0, 0, 0, -2, 0,
    -- filter=177 channel=103
    0, 9, -1, 9, 9, -12, -2, -2, -9,
    -- filter=177 channel=104
    11, 7, -13, 16, 16, -13, 6, 2, -20,
    -- filter=177 channel=105
    -2, -5, -3, -6, -16, -1, -11, -16, 5,
    -- filter=177 channel=106
    4, 0, 5, 0, 0, -5, 8, -3, -8,
    -- filter=177 channel=107
    -9, -2, 18, -3, -22, 12, -2, -11, 17,
    -- filter=177 channel=108
    0, 1, 0, 2, -7, -11, 1, -6, -6,
    -- filter=177 channel=109
    -1, -3, 9, 0, -6, 0, 1, -6, 1,
    -- filter=177 channel=110
    -1, 2, 0, 0, 8, 0, -6, -9, -12,
    -- filter=177 channel=111
    5, 5, -8, -7, -4, 2, -6, -5, -4,
    -- filter=177 channel=112
    0, -4, -3, -3, -8, 10, -6, -2, 10,
    -- filter=177 channel=113
    1, 5, -2, 12, 6, 6, 3, -1, -1,
    -- filter=177 channel=114
    -8, -20, 17, -5, -22, 10, -4, -22, 8,
    -- filter=177 channel=115
    -4, -6, 0, -2, 6, -5, 5, -5, -5,
    -- filter=177 channel=116
    3, -3, -3, 7, -8, -8, 0, -13, -2,
    -- filter=177 channel=117
    4, 6, 0, 6, 10, -3, -2, 0, 6,
    -- filter=177 channel=118
    4, -5, 6, 0, 1, -3, -1, 5, -6,
    -- filter=177 channel=119
    -5, -8, 10, -8, -8, 0, -16, 2, -6,
    -- filter=177 channel=120
    1, -3, 4, 3, -20, 12, -2, -9, -2,
    -- filter=177 channel=121
    10, 4, 1, -2, -8, -4, 6, -2, 2,
    -- filter=177 channel=122
    6, 18, -11, 15, 17, -20, 4, 7, -15,
    -- filter=177 channel=123
    -9, 1, 2, 3, -3, -1, -10, -5, -8,
    -- filter=177 channel=124
    -12, 2, 3, -7, -9, -1, -7, -7, 2,
    -- filter=177 channel=125
    7, 0, 2, 15, -3, -6, 2, -8, -13,
    -- filter=177 channel=126
    3, -13, -8, 13, 1, 1, 10, -10, 1,
    -- filter=177 channel=127
    -4, 1, 2, 4, -7, 0, -4, 3, 6,
    -- filter=178 channel=0
    -14, 2, 6, -11, 13, 3, -12, -3, 2,
    -- filter=178 channel=1
    -17, 10, -8, -16, 5, 7, -10, 5, 9,
    -- filter=178 channel=2
    0, -2, 6, 2, 3, 0, -5, -6, -2,
    -- filter=178 channel=3
    -7, -8, 5, -2, 0, 1, -2, -8, -4,
    -- filter=178 channel=4
    -8, -4, 6, -11, -12, 2, -9, -8, 8,
    -- filter=178 channel=5
    -5, 6, -2, -10, 6, 7, -14, 11, 7,
    -- filter=178 channel=6
    3, -5, 1, 3, -7, 6, -2, -2, -2,
    -- filter=178 channel=7
    0, 5, -7, 2, -2, 2, 6, -5, 0,
    -- filter=178 channel=8
    2, -5, -2, 4, -3, 0, 1, -1, 0,
    -- filter=178 channel=9
    -4, 7, 3, 6, 0, -2, 5, 5, 4,
    -- filter=178 channel=10
    -1, 6, 0, 4, -2, -4, -6, 5, -6,
    -- filter=178 channel=11
    1, -7, 2, 10, -12, 5, -1, -4, 4,
    -- filter=178 channel=12
    -3, 7, -2, -9, 3, 8, -8, 0, -7,
    -- filter=178 channel=13
    2, 9, -8, 0, -1, -8, -8, -1, -11,
    -- filter=178 channel=14
    4, 4, -3, -1, -4, -5, 2, 0, 2,
    -- filter=178 channel=15
    4, -5, -10, 2, -5, -14, 11, 2, -13,
    -- filter=178 channel=16
    0, 7, 4, -15, 2, 1, -1, 5, -6,
    -- filter=178 channel=17
    -5, 6, -2, 0, -6, 0, -7, -1, 0,
    -- filter=178 channel=18
    -2, -4, -12, -2, 2, -8, -1, 7, -4,
    -- filter=178 channel=19
    5, 3, -5, 7, -1, -2, -1, 5, -6,
    -- filter=178 channel=20
    10, -4, 2, 3, -8, 0, 12, 2, -7,
    -- filter=178 channel=21
    -2, 8, 2, -2, 7, -8, 0, 2, 0,
    -- filter=178 channel=22
    7, 2, 4, 1, 7, -4, -2, 1, -7,
    -- filter=178 channel=23
    12, 0, -5, 12, -8, -4, 1, -2, 0,
    -- filter=178 channel=24
    7, 7, 3, 5, -6, 0, -2, 5, -2,
    -- filter=178 channel=25
    -9, 6, -1, -4, 18, -17, -4, 17, -14,
    -- filter=178 channel=26
    -10, 6, -3, 2, -2, -3, -4, -3, 0,
    -- filter=178 channel=27
    4, 12, -7, -5, 7, -16, -1, 20, -17,
    -- filter=178 channel=28
    0, -6, 6, 6, 4, 4, -2, 1, -3,
    -- filter=178 channel=29
    12, 1, 2, 4, -5, 3, 12, 3, -2,
    -- filter=178 channel=30
    -5, 0, 2, -6, 1, -8, 0, 0, 2,
    -- filter=178 channel=31
    -1, 5, -4, 4, 15, -16, -6, 15, -7,
    -- filter=178 channel=32
    6, 3, -5, -5, 15, -4, -9, 9, -8,
    -- filter=178 channel=33
    0, 1, -8, -5, 12, -3, -3, 17, -11,
    -- filter=178 channel=34
    2, 1, 11, 5, 4, 13, 3, 2, 7,
    -- filter=178 channel=35
    6, 6, 7, 6, 1, -3, 5, -2, -4,
    -- filter=178 channel=36
    -1, -3, 0, -6, -7, -7, 0, 2, -1,
    -- filter=178 channel=37
    -12, 4, 2, -23, 3, 9, -16, -1, 1,
    -- filter=178 channel=38
    -4, 0, -9, -7, 8, -2, -7, 10, -3,
    -- filter=178 channel=39
    1, 1, 2, -4, -1, 3, 7, 2, 0,
    -- filter=178 channel=40
    -1, -5, -5, 6, -3, -3, 1, -3, 0,
    -- filter=178 channel=41
    3, 7, -2, 1, 13, 0, 11, -5, 1,
    -- filter=178 channel=42
    0, -4, 1, -4, -1, 5, 0, 0, 9,
    -- filter=178 channel=43
    1, 1, -7, 0, 1, 0, 0, -9, 0,
    -- filter=178 channel=44
    -11, 8, -6, -8, 10, -7, -1, 0, -5,
    -- filter=178 channel=45
    -3, 6, 0, -4, 5, -6, -7, 0, 3,
    -- filter=178 channel=46
    1, -1, -3, -1, -1, 3, -2, -4, -3,
    -- filter=178 channel=47
    0, 7, 4, -6, 8, -11, -15, 15, 0,
    -- filter=178 channel=48
    0, 10, 0, -11, 7, -12, -3, 13, -7,
    -- filter=178 channel=49
    -4, -5, -3, 0, -3, -10, -8, 6, -2,
    -- filter=178 channel=50
    -4, 7, -9, -4, 10, -5, -2, 12, -2,
    -- filter=178 channel=51
    1, -4, -3, 2, 1, 5, 3, 0, -3,
    -- filter=178 channel=52
    0, 0, -3, -1, 0, 3, 6, 1, -9,
    -- filter=178 channel=53
    9, -9, 4, -1, -8, -2, 5, -7, 1,
    -- filter=178 channel=54
    1, -5, 3, -1, 6, 6, 0, -7, 5,
    -- filter=178 channel=55
    7, 1, -5, 11, -3, -15, 8, -3, -14,
    -- filter=178 channel=56
    1, -6, 0, 8, 6, 7, -2, 6, 1,
    -- filter=178 channel=57
    -1, 6, 1, 7, -4, 0, 0, 2, -2,
    -- filter=178 channel=58
    0, -5, 7, -13, -3, 5, -6, -6, 8,
    -- filter=178 channel=59
    -8, 17, -7, -8, 20, -3, -11, 18, -9,
    -- filter=178 channel=60
    0, 2, 5, 0, -4, 3, 3, 4, -2,
    -- filter=178 channel=61
    -4, -2, 5, 4, 6, 2, 2, -5, -6,
    -- filter=178 channel=62
    3, 0, -4, 0, 1, -4, -1, -3, -3,
    -- filter=178 channel=63
    -1, 7, -2, -10, 0, -3, -5, 3, 7,
    -- filter=178 channel=64
    1, 4, 6, 5, -9, -5, -3, -5, -4,
    -- filter=178 channel=65
    -2, -6, 0, 4, -3, 1, -6, -1, 1,
    -- filter=178 channel=66
    0, 7, -6, -2, 16, -1, 1, 7, -5,
    -- filter=178 channel=67
    2, 0, -6, -3, 4, 4, 5, 3, 0,
    -- filter=178 channel=68
    0, 1, -2, -8, -9, 2, 6, -1, -6,
    -- filter=178 channel=69
    0, 9, -5, -2, 6, 2, 4, 4, 3,
    -- filter=178 channel=70
    0, 3, -7, 0, -2, -7, 2, 7, 0,
    -- filter=178 channel=71
    -2, 4, -3, -8, -4, 4, -6, -4, 4,
    -- filter=178 channel=72
    -4, 6, 2, 2, 4, -5, -8, 0, -12,
    -- filter=178 channel=73
    5, -1, -3, 7, -4, -1, 6, -3, -6,
    -- filter=178 channel=74
    0, -7, 5, 9, 1, 1, -5, 6, -6,
    -- filter=178 channel=75
    -8, 10, 5, -22, 13, 6, -9, 3, 0,
    -- filter=178 channel=76
    -1, -1, 1, 4, -7, -2, 0, -12, -7,
    -- filter=178 channel=77
    -7, -3, -7, 4, 0, -3, -1, 2, -5,
    -- filter=178 channel=78
    6, -1, 6, -6, -2, -3, -6, 2, 8,
    -- filter=178 channel=79
    -1, 1, -7, -2, 11, -15, -5, 15, -9,
    -- filter=178 channel=80
    -7, 16, -3, -11, 23, -15, -15, 10, -3,
    -- filter=178 channel=81
    -6, 1, -5, -2, 0, -6, 1, -6, 4,
    -- filter=178 channel=82
    4, -3, 1, 6, -3, -6, 0, -3, 2,
    -- filter=178 channel=83
    -7, 5, 4, -5, 8, 2, -3, 0, 3,
    -- filter=178 channel=84
    -3, 6, 1, 0, 0, -10, 0, 9, -4,
    -- filter=178 channel=85
    7, -2, -3, -2, 0, 0, 0, 6, -6,
    -- filter=178 channel=86
    2, 4, 8, -5, 1, -1, 0, 1, 5,
    -- filter=178 channel=87
    2, -2, 4, 2, -3, 4, -1, -4, -7,
    -- filter=178 channel=88
    -4, -7, 2, 3, -7, -8, 0, 1, -7,
    -- filter=178 channel=89
    -2, 4, -11, 5, 1, -4, -2, -1, 0,
    -- filter=178 channel=90
    -2, 3, -5, -4, -4, 1, 7, 4, -5,
    -- filter=178 channel=91
    -2, -7, -1, -4, 6, -14, 0, 3, -5,
    -- filter=178 channel=92
    4, 3, -4, 5, -1, 2, 9, 4, 8,
    -- filter=178 channel=93
    0, 13, 6, -10, 13, -4, -8, 5, 5,
    -- filter=178 channel=94
    7, -3, -4, 1, 2, 3, 3, 4, 2,
    -- filter=178 channel=95
    0, -2, 5, -4, -3, 1, 1, -6, 2,
    -- filter=178 channel=96
    4, 0, 1, 2, -1, 5, -6, 0, -5,
    -- filter=178 channel=97
    -4, 1, -6, 0, -5, -4, 4, -3, 3,
    -- filter=178 channel=98
    -1, 19, -2, -7, 9, -2, -8, 18, 1,
    -- filter=178 channel=99
    10, 5, -5, 6, 3, -18, 1, 6, -14,
    -- filter=178 channel=100
    -2, 7, -3, 10, 5, 2, 6, -4, 0,
    -- filter=178 channel=101
    3, -3, -7, 0, -9, -3, 1, -4, -6,
    -- filter=178 channel=102
    -6, -5, -6, 5, -3, 6, 3, 4, 4,
    -- filter=178 channel=103
    -4, 19, 4, -3, 15, -12, -12, 5, 3,
    -- filter=178 channel=104
    -6, 15, -1, -3, 12, -18, -13, 16, -3,
    -- filter=178 channel=105
    7, -2, 6, 2, -10, -5, 4, 2, -4,
    -- filter=178 channel=106
    3, -10, 4, -2, -6, 6, 3, -9, 5,
    -- filter=178 channel=107
    8, -8, -4, -3, -11, -1, 7, -10, -6,
    -- filter=178 channel=108
    4, -1, 1, 5, 0, 0, 6, -6, 6,
    -- filter=178 channel=109
    9, 4, -7, 6, 8, -12, 2, 19, -11,
    -- filter=178 channel=110
    0, -3, -3, 2, -3, -4, 6, -6, 3,
    -- filter=178 channel=111
    -2, -1, -8, 3, 4, 4, 4, 0, -5,
    -- filter=178 channel=112
    -1, 9, -1, 1, 4, -6, 1, 8, -2,
    -- filter=178 channel=113
    1, 1, -7, 6, 4, 0, -6, 12, -9,
    -- filter=178 channel=114
    -3, 2, -5, -3, 3, -3, 0, 3, -6,
    -- filter=178 channel=115
    5, -3, 4, 0, 0, -2, 2, 6, -5,
    -- filter=178 channel=116
    5, 10, -10, 0, 9, -12, -3, 10, -7,
    -- filter=178 channel=117
    -4, -6, -6, -6, -1, -9, -4, 1, 0,
    -- filter=178 channel=118
    0, -1, 6, -3, -2, 2, 5, -2, -2,
    -- filter=178 channel=119
    12, -2, -2, 9, 2, 7, 11, 2, 1,
    -- filter=178 channel=120
    15, 1, -3, 2, -2, -9, 0, 12, -3,
    -- filter=178 channel=121
    -5, 6, 2, 0, 7, -5, -7, 4, 4,
    -- filter=178 channel=122
    -18, 15, -7, -10, 18, -16, -8, 16, -4,
    -- filter=178 channel=123
    1, -4, -3, 0, -3, -4, -3, -3, 0,
    -- filter=178 channel=124
    8, -2, -6, 6, -8, -5, 6, -6, 0,
    -- filter=178 channel=125
    2, 7, -3, -1, 8, -17, -13, 9, -12,
    -- filter=178 channel=126
    5, 8, -5, -10, 8, -8, 1, 3, -9,
    -- filter=178 channel=127
    3, 3, -5, 1, 3, 0, 0, 4, -1,
    -- filter=179 channel=0
    0, 7, -6, 7, -6, 4, -6, -1, 3,
    -- filter=179 channel=1
    6, 5, -5, -3, -2, 0, -1, -3, -2,
    -- filter=179 channel=2
    3, -3, 5, -6, 6, -1, 1, -2, 1,
    -- filter=179 channel=3
    7, 5, 6, 3, -7, 4, 7, -5, 6,
    -- filter=179 channel=4
    7, -4, -6, 0, 5, 5, 5, 1, 6,
    -- filter=179 channel=5
    3, -5, 7, 1, 0, 8, 0, 0, 7,
    -- filter=179 channel=6
    2, -4, 0, 2, 2, -4, 0, 0, -2,
    -- filter=179 channel=7
    1, -4, 0, -5, 3, -5, 3, 1, 2,
    -- filter=179 channel=8
    -2, 4, 3, 6, 6, -3, 2, -6, 2,
    -- filter=179 channel=9
    -1, 3, -1, -6, -1, 0, -1, 7, -7,
    -- filter=179 channel=10
    4, 6, -7, 3, -4, -2, -4, -5, -5,
    -- filter=179 channel=11
    0, -1, -4, 0, 3, -5, 2, 1, -5,
    -- filter=179 channel=12
    -4, 1, -3, 1, 5, 5, -3, 5, -6,
    -- filter=179 channel=13
    -2, 3, 2, 1, 0, -3, -6, -7, -4,
    -- filter=179 channel=14
    3, -2, 1, -5, -7, 0, -3, 2, 0,
    -- filter=179 channel=15
    -1, 2, -6, -2, -1, 1, 0, 5, 6,
    -- filter=179 channel=16
    -3, -5, -2, -3, 6, 5, -4, -2, -4,
    -- filter=179 channel=17
    2, 3, -7, 0, 0, 0, -1, 3, 1,
    -- filter=179 channel=18
    0, -7, -7, 3, 6, -6, 2, -4, -6,
    -- filter=179 channel=19
    0, -4, 6, -4, -5, 0, 4, 0, -3,
    -- filter=179 channel=20
    -4, -3, -5, -1, 8, 7, 5, 5, 4,
    -- filter=179 channel=21
    5, -4, -3, -3, 7, -3, 2, 7, 1,
    -- filter=179 channel=22
    -3, 6, -3, -1, 0, 5, 4, 2, 3,
    -- filter=179 channel=23
    0, 0, 0, 3, -1, -6, 2, -4, -2,
    -- filter=179 channel=24
    3, 7, 1, 0, -1, 4, -7, 3, 2,
    -- filter=179 channel=25
    -6, 5, -4, 5, -3, 0, -1, -4, -7,
    -- filter=179 channel=26
    -4, 7, 1, 3, -2, -1, 1, 7, -1,
    -- filter=179 channel=27
    -6, 1, -3, -7, 4, 4, -5, -8, -6,
    -- filter=179 channel=28
    7, 0, 2, 3, -3, 2, 2, -6, -3,
    -- filter=179 channel=29
    4, -5, -2, 7, 5, 7, 0, 8, -6,
    -- filter=179 channel=30
    5, -7, 0, -3, 2, 0, -3, 3, -3,
    -- filter=179 channel=31
    3, -7, 1, 2, -4, -4, 6, -1, 5,
    -- filter=179 channel=32
    -7, 1, -7, 2, 0, -1, -7, -6, -3,
    -- filter=179 channel=33
    -5, 3, -5, 3, -1, -2, 6, 2, 2,
    -- filter=179 channel=34
    3, 3, -4, -1, -1, 2, -1, -2, 4,
    -- filter=179 channel=35
    -5, -5, 1, 5, -2, 7, 1, 1, 1,
    -- filter=179 channel=36
    -3, 0, -3, 0, -6, 0, 0, 0, 0,
    -- filter=179 channel=37
    -1, -1, 3, 1, -4, -5, -4, -1, -2,
    -- filter=179 channel=38
    0, 4, 6, 0, 3, 5, -5, -6, -4,
    -- filter=179 channel=39
    1, 6, -6, 2, 3, 0, 7, 6, 5,
    -- filter=179 channel=40
    0, -6, 5, 5, -3, -6, -3, 3, 7,
    -- filter=179 channel=41
    7, 2, -4, 2, 1, 0, 2, 5, -1,
    -- filter=179 channel=42
    -1, -3, 0, 0, 4, -6, -3, -6, -6,
    -- filter=179 channel=43
    3, 1, 0, -6, 6, 2, 1, 5, 4,
    -- filter=179 channel=44
    1, 7, 6, -3, -7, -5, 4, -1, 0,
    -- filter=179 channel=45
    1, -2, 0, -2, 0, -1, 5, -3, 7,
    -- filter=179 channel=46
    0, 0, -6, -2, -7, 5, 3, -2, 6,
    -- filter=179 channel=47
    -2, 0, 4, -2, 2, 0, -2, -3, 4,
    -- filter=179 channel=48
    -6, -6, -3, -5, -5, -3, -1, -1, -3,
    -- filter=179 channel=49
    0, -7, 1, 7, 7, -6, 4, -2, -6,
    -- filter=179 channel=50
    4, 0, -6, 3, -7, 3, -3, 4, 4,
    -- filter=179 channel=51
    -7, -2, 5, 6, 0, 0, 7, -2, -6,
    -- filter=179 channel=52
    -4, -3, 1, 7, -5, 5, -1, -3, -6,
    -- filter=179 channel=53
    -2, 6, 0, -1, 3, 4, 0, -1, 5,
    -- filter=179 channel=54
    0, 3, -6, 5, 6, -3, -4, 0, 3,
    -- filter=179 channel=55
    4, 3, -5, 6, -8, 4, 0, -1, -2,
    -- filter=179 channel=56
    -3, -2, 3, -4, 3, 0, 1, 2, 4,
    -- filter=179 channel=57
    4, 0, 0, -2, 0, 0, -6, 1, 5,
    -- filter=179 channel=58
    6, -6, 2, 6, 0, 6, 5, 2, 7,
    -- filter=179 channel=59
    0, -2, 1, 6, -8, 4, 5, -4, -4,
    -- filter=179 channel=60
    7, -4, 4, 0, -4, 5, -1, -2, -5,
    -- filter=179 channel=61
    0, -2, -6, 0, -6, 3, -5, 0, 1,
    -- filter=179 channel=62
    2, -2, 6, 6, 1, -3, -2, -6, -1,
    -- filter=179 channel=63
    0, 5, 7, -6, 7, -6, 2, 0, -2,
    -- filter=179 channel=64
    -4, 3, 4, 0, -1, -5, 2, 7, -3,
    -- filter=179 channel=65
    -2, 3, -6, 7, -3, 4, 1, 0, 5,
    -- filter=179 channel=66
    7, 1, -2, -5, -1, 3, -7, 6, -3,
    -- filter=179 channel=67
    6, 7, -6, -2, 1, 0, 1, -5, 5,
    -- filter=179 channel=68
    4, 4, 1, -2, -3, 0, -4, -6, 7,
    -- filter=179 channel=69
    -1, -4, 1, 0, 3, -7, -1, -4, 3,
    -- filter=179 channel=70
    6, 0, -2, -6, 0, -4, 0, -7, -2,
    -- filter=179 channel=71
    -3, 4, -6, 6, -4, -4, -5, -4, 5,
    -- filter=179 channel=72
    -3, 3, -4, -2, -3, 4, 5, 0, 6,
    -- filter=179 channel=73
    -3, 3, -2, -2, -4, -1, -5, -2, 2,
    -- filter=179 channel=74
    3, 1, -3, 0, -2, 1, -2, -3, -6,
    -- filter=179 channel=75
    0, -4, 0, 5, 6, 7, 4, 2, 0,
    -- filter=179 channel=76
    2, 0, 2, 7, -3, 2, 6, -3, -2,
    -- filter=179 channel=77
    -1, -5, -4, 5, 0, 1, -2, -2, -2,
    -- filter=179 channel=78
    -5, -2, 1, 3, -1, 0, -5, 2, 5,
    -- filter=179 channel=79
    7, 0, -1, 4, -1, -5, 4, -2, -8,
    -- filter=179 channel=80
    0, -4, 0, 3, 0, 6, 2, -4, -4,
    -- filter=179 channel=81
    -3, -6, 0, 4, -4, -2, -6, -5, -7,
    -- filter=179 channel=82
    2, 5, -3, -6, -3, -2, -4, -4, 1,
    -- filter=179 channel=83
    -6, 6, -4, -3, 4, -6, -5, 0, 0,
    -- filter=179 channel=84
    1, 0, -6, 4, 3, 0, -4, -1, -7,
    -- filter=179 channel=85
    7, 5, 1, -4, -7, 0, -1, -2, -7,
    -- filter=179 channel=86
    7, 0, 1, 6, 5, 1, -5, 3, 6,
    -- filter=179 channel=87
    5, 0, 7, 5, -5, -5, -1, 1, 0,
    -- filter=179 channel=88
    -4, 1, -3, 5, 2, -6, -5, -4, -1,
    -- filter=179 channel=89
    -5, 4, -8, 2, 4, -7, 3, -5, -2,
    -- filter=179 channel=90
    -1, -6, -3, 4, -2, 5, -6, 6, -1,
    -- filter=179 channel=91
    -7, -7, -7, 1, 0, -1, -3, 5, -2,
    -- filter=179 channel=92
    -6, 6, 4, 0, -7, 5, -2, 2, -2,
    -- filter=179 channel=93
    -5, -2, 0, 4, 6, 0, -6, 0, 0,
    -- filter=179 channel=94
    1, -3, -1, 5, -5, 2, -4, 0, 2,
    -- filter=179 channel=95
    4, 2, 5, 2, 2, 5, -2, -6, 6,
    -- filter=179 channel=96
    -4, -4, 7, 2, 1, 0, 4, 2, -4,
    -- filter=179 channel=97
    -2, 4, 3, 1, 6, 0, 1, -4, 0,
    -- filter=179 channel=98
    -2, 5, 0, 7, 0, 1, 1, 0, -3,
    -- filter=179 channel=99
    5, 0, 6, 1, -6, 0, -5, 0, -4,
    -- filter=179 channel=100
    -1, -4, 3, 0, 2, -7, 0, -6, 2,
    -- filter=179 channel=101
    -7, -3, 2, 4, 7, 3, -1, -4, 3,
    -- filter=179 channel=102
    -7, -4, 6, 6, 0, 0, -2, -4, -1,
    -- filter=179 channel=103
    -5, 0, -6, 1, 2, 0, -6, -3, -6,
    -- filter=179 channel=104
    0, -3, -2, -4, -6, -3, -2, 6, -7,
    -- filter=179 channel=105
    -6, 0, 5, 8, 0, 3, 1, -4, -2,
    -- filter=179 channel=106
    -3, 1, 0, 1, 6, 0, 1, -3, 7,
    -- filter=179 channel=107
    -2, -7, 1, 1, 6, 5, -4, 1, 6,
    -- filter=179 channel=108
    0, 7, 3, 4, 0, 6, 3, 6, 2,
    -- filter=179 channel=109
    -5, -3, -7, -5, -6, 0, -5, 5, -3,
    -- filter=179 channel=110
    -5, 0, 1, 1, -7, 0, 0, -4, 5,
    -- filter=179 channel=111
    5, -1, 0, -3, 3, -4, -4, 0, 1,
    -- filter=179 channel=112
    5, 2, 4, 6, -6, 0, 4, -7, 1,
    -- filter=179 channel=113
    -4, 3, 0, 1, -7, -3, 6, 0, 0,
    -- filter=179 channel=114
    5, -6, -3, 0, -8, 1, 0, -5, -3,
    -- filter=179 channel=115
    3, 0, -2, 6, 0, -3, -1, -2, -3,
    -- filter=179 channel=116
    4, 5, -4, 6, -7, 4, -5, 3, -3,
    -- filter=179 channel=117
    -5, 2, -6, -4, -7, 6, 3, -7, 0,
    -- filter=179 channel=118
    -2, 4, 3, 5, 1, -7, 2, 0, 6,
    -- filter=179 channel=119
    1, -1, 4, 3, 1, -1, 0, 5, 2,
    -- filter=179 channel=120
    4, 5, 7, -3, 0, 6, -6, -6, 1,
    -- filter=179 channel=121
    -2, 3, -3, -7, -2, 5, 5, -4, 4,
    -- filter=179 channel=122
    0, 0, 2, 8, 3, 3, 7, -4, 1,
    -- filter=179 channel=123
    1, 4, -6, -7, 4, 0, 2, 5, 2,
    -- filter=179 channel=124
    3, 5, 5, 2, 3, 4, -2, 7, 1,
    -- filter=179 channel=125
    -6, -6, -4, -2, -5, -2, 4, 1, 4,
    -- filter=179 channel=126
    -1, 0, 0, -1, 5, -5, 4, 2, 2,
    -- filter=179 channel=127
    2, -3, -6, 2, 2, -2, 4, 3, -6,
    -- filter=180 channel=0
    -2, -5, 4, 11, 0, -1, 11, -2, 0,
    -- filter=180 channel=1
    3, 0, -1, 8, 3, 0, 1, -3, -1,
    -- filter=180 channel=2
    -1, -5, 6, 3, 0, 3, -2, -3, -6,
    -- filter=180 channel=3
    5, 6, 5, 15, 5, 10, 7, 4, 7,
    -- filter=180 channel=4
    3, 0, -4, 8, 3, -1, 0, 8, 9,
    -- filter=180 channel=5
    0, -9, 3, 8, -4, -6, -2, -5, -9,
    -- filter=180 channel=6
    4, -7, -7, -4, -8, 2, 2, -7, 0,
    -- filter=180 channel=7
    -1, -7, -4, 4, 4, 4, 6, 4, 3,
    -- filter=180 channel=8
    4, -1, 3, -2, -5, -6, 0, -3, 4,
    -- filter=180 channel=9
    3, -3, 1, 4, -6, -7, 0, 0, -1,
    -- filter=180 channel=10
    2, 3, 2, -6, 5, 5, -1, -8, -2,
    -- filter=180 channel=11
    -1, -3, -8, 2, 3, -1, -7, -8, -1,
    -- filter=180 channel=12
    5, 0, -5, -8, -8, 6, 1, -9, 4,
    -- filter=180 channel=13
    7, 6, 5, 0, -2, -2, 3, -4, -10,
    -- filter=180 channel=14
    7, -7, 4, -3, -2, 4, -3, -6, 5,
    -- filter=180 channel=15
    12, 10, -5, 2, 4, 0, -10, -9, -12,
    -- filter=180 channel=16
    6, -1, 1, 3, 5, 8, 5, -5, 0,
    -- filter=180 channel=17
    -3, -4, 0, 6, -6, -2, 1, 4, 3,
    -- filter=180 channel=18
    6, 14, -8, -12, 4, -9, -4, -7, -2,
    -- filter=180 channel=19
    4, -2, 0, 0, 0, -3, 7, -2, 2,
    -- filter=180 channel=20
    -4, -5, 0, -10, -6, 2, -6, 3, -2,
    -- filter=180 channel=21
    4, 9, 3, 9, 9, 3, -8, -4, 1,
    -- filter=180 channel=22
    8, -2, 3, 0, 7, 4, 4, 3, -9,
    -- filter=180 channel=23
    15, 1, -8, 3, -4, -3, -10, -10, -15,
    -- filter=180 channel=24
    4, -3, -5, 2, 0, 5, 3, -1, 2,
    -- filter=180 channel=25
    3, 3, -2, -3, 3, -9, -4, -13, -2,
    -- filter=180 channel=26
    0, -5, 3, 0, -6, -5, 7, -5, 2,
    -- filter=180 channel=27
    18, 3, -6, -14, 3, -12, -9, -2, -14,
    -- filter=180 channel=28
    -5, -4, 6, -3, 4, 5, 0, -1, -7,
    -- filter=180 channel=29
    5, 0, -2, -11, -11, -4, 3, 4, 5,
    -- filter=180 channel=30
    10, -3, 1, -5, 1, -9, -4, 0, -10,
    -- filter=180 channel=31
    20, 14, 8, -2, -5, 2, -11, -16, -12,
    -- filter=180 channel=32
    6, 8, -11, -14, 4, -14, -11, -9, -4,
    -- filter=180 channel=33
    10, 10, 0, -2, -1, -9, -8, -9, -2,
    -- filter=180 channel=34
    6, 0, -2, 2, -4, -9, -12, 3, -11,
    -- filter=180 channel=35
    3, 2, -4, -2, -6, 7, -3, 0, 6,
    -- filter=180 channel=36
    8, 9, 10, 4, -1, -3, -3, -3, 5,
    -- filter=180 channel=37
    7, 4, 1, 12, 7, -9, 9, 4, 2,
    -- filter=180 channel=38
    6, 4, 0, 3, 7, -5, -10, -8, 1,
    -- filter=180 channel=39
    1, 0, -5, -3, 2, -6, 4, -3, -2,
    -- filter=180 channel=40
    9, 3, 3, 7, -1, 3, 4, 0, 0,
    -- filter=180 channel=41
    0, 6, 0, -3, -10, 9, 7, -2, -4,
    -- filter=180 channel=42
    0, 0, 6, -4, 2, -8, 5, -1, 2,
    -- filter=180 channel=43
    7, -1, 1, 1, -1, 7, 6, -2, 0,
    -- filter=180 channel=44
    11, 4, 7, 0, -2, -10, -1, -2, -4,
    -- filter=180 channel=45
    7, 1, -4, 3, 3, -4, -2, -4, 1,
    -- filter=180 channel=46
    7, -1, 3, 3, 4, 1, 8, 0, 1,
    -- filter=180 channel=47
    6, 0, 0, 9, 6, 7, -10, 0, -2,
    -- filter=180 channel=48
    11, 13, 8, -3, -1, 0, -12, -9, 0,
    -- filter=180 channel=49
    8, 1, -9, 1, 1, -3, -4, -5, 0,
    -- filter=180 channel=50
    6, -2, -4, 3, -1, 2, -6, 0, -6,
    -- filter=180 channel=51
    4, 1, -6, 2, 2, 7, -1, 5, -4,
    -- filter=180 channel=52
    3, 0, 0, -8, 5, -2, -7, -5, 2,
    -- filter=180 channel=53
    -3, 2, -5, 3, -4, -8, -7, 2, -6,
    -- filter=180 channel=54
    -6, -7, -6, 3, 7, -5, 0, 0, 7,
    -- filter=180 channel=55
    3, 13, -3, -2, 3, -4, -12, -9, 1,
    -- filter=180 channel=56
    2, 0, -3, -7, -8, 2, 1, 2, -5,
    -- filter=180 channel=57
    -2, 2, 3, 1, 4, -2, 0, -4, 6,
    -- filter=180 channel=58
    4, 4, 4, -1, 6, -3, -3, 6, 4,
    -- filter=180 channel=59
    12, 4, 1, 0, -2, -9, -3, -17, -13,
    -- filter=180 channel=60
    2, 1, -2, -5, 0, 0, 2, -1, 3,
    -- filter=180 channel=61
    -5, 0, -3, -8, -7, -1, -8, 5, 0,
    -- filter=180 channel=62
    4, -3, -3, 2, 3, 4, -5, 2, 0,
    -- filter=180 channel=63
    4, -8, 2, 2, 4, 4, 4, -8, -2,
    -- filter=180 channel=64
    -2, -3, -5, 2, -2, 6, 1, 5, 5,
    -- filter=180 channel=65
    6, -6, -2, 1, 2, 6, -5, 3, 5,
    -- filter=180 channel=66
    5, 10, 8, 0, -4, -4, -6, -9, 7,
    -- filter=180 channel=67
    3, 3, 4, -5, 6, 2, 7, 0, 7,
    -- filter=180 channel=68
    -3, -3, 3, 7, 2, 4, -4, 8, 0,
    -- filter=180 channel=69
    -6, 7, 7, 7, 0, 5, -3, -4, 7,
    -- filter=180 channel=70
    8, 1, -8, -6, 0, -2, 0, -6, 0,
    -- filter=180 channel=71
    3, 0, 2, 1, 8, 7, 1, 6, 4,
    -- filter=180 channel=72
    16, 6, 9, 0, 2, 2, -11, -7, -11,
    -- filter=180 channel=73
    -3, 1, 0, -6, -8, -9, -11, 0, -6,
    -- filter=180 channel=74
    7, -7, 2, -1, 3, -5, -12, 3, 1,
    -- filter=180 channel=75
    11, 3, 1, 8, 3, -4, 7, -2, -3,
    -- filter=180 channel=76
    8, 1, -3, -10, -6, 3, 0, 0, -1,
    -- filter=180 channel=77
    0, 1, -3, 4, 6, 0, -2, -3, 3,
    -- filter=180 channel=78
    0, -6, 2, -4, -7, 5, -8, 1, -9,
    -- filter=180 channel=79
    15, 6, 0, -6, 7, -2, -6, -9, -6,
    -- filter=180 channel=80
    9, 12, 9, 2, 0, -2, -13, -19, -3,
    -- filter=180 channel=81
    3, 3, 2, 6, -1, -5, 3, -3, 5,
    -- filter=180 channel=82
    -3, 2, 7, -2, -2, -4, 1, 7, -6,
    -- filter=180 channel=83
    0, 4, -3, -8, -1, -8, -6, -5, 5,
    -- filter=180 channel=84
    5, 9, 0, -4, -1, -10, 1, -10, -5,
    -- filter=180 channel=85
    4, -7, 4, -6, 7, 5, 4, 0, 1,
    -- filter=180 channel=86
    -1, -6, -7, 0, 3, -5, 4, 3, -4,
    -- filter=180 channel=87
    8, 5, 3, -6, -5, -3, -5, 3, -7,
    -- filter=180 channel=88
    9, 5, 5, -3, -7, -2, -1, -4, 0,
    -- filter=180 channel=89
    15, 5, 1, -5, 4, -6, -8, -10, -5,
    -- filter=180 channel=90
    7, -4, 5, -1, 9, 7, -8, 0, 2,
    -- filter=180 channel=91
    -2, 7, 3, -9, -8, -8, -1, 0, 0,
    -- filter=180 channel=92
    1, 0, 4, 0, -6, -4, 5, 6, 1,
    -- filter=180 channel=93
    5, -3, -2, -3, -3, -12, 0, -3, -10,
    -- filter=180 channel=94
    0, 0, -2, 7, 3, -2, 0, 3, 7,
    -- filter=180 channel=95
    3, 7, 6, -3, 0, 1, -6, -4, 2,
    -- filter=180 channel=96
    0, -3, 5, 3, -2, 5, 7, 0, 6,
    -- filter=180 channel=97
    8, -5, 1, 10, 10, 2, 2, 0, 0,
    -- filter=180 channel=98
    10, 10, -5, -6, 7, -2, -15, -8, -9,
    -- filter=180 channel=99
    18, 7, 0, -1, -3, -11, -19, -12, -15,
    -- filter=180 channel=100
    -7, -1, -4, 0, 4, 3, -4, -5, -4,
    -- filter=180 channel=101
    -1, 0, 0, 0, -3, 5, 7, 5, 0,
    -- filter=180 channel=102
    3, 4, -6, -5, -3, 3, -5, 4, -3,
    -- filter=180 channel=103
    14, 4, 3, 5, 2, 9, 4, -4, -5,
    -- filter=180 channel=104
    8, 9, 5, 2, -8, -2, -3, -9, -10,
    -- filter=180 channel=105
    -2, 0, -4, -2, -1, -7, 0, -1, 6,
    -- filter=180 channel=106
    0, 0, 5, -6, -6, -2, -1, -5, 7,
    -- filter=180 channel=107
    -5, 0, -8, 2, 0, -3, -3, 0, 0,
    -- filter=180 channel=108
    0, 3, 6, -3, -3, -3, -1, 3, 0,
    -- filter=180 channel=109
    0, 4, 0, -13, -10, -11, -16, -4, -15,
    -- filter=180 channel=110
    0, 2, 0, 6, -3, -6, -12, -4, 4,
    -- filter=180 channel=111
    -8, 0, -5, 0, 0, 5, 1, 1, 2,
    -- filter=180 channel=112
    0, -3, -2, 0, -1, 1, -6, 5, -6,
    -- filter=180 channel=113
    5, 7, 4, 0, 6, -5, -8, 2, -11,
    -- filter=180 channel=114
    6, 5, -8, -1, -11, -7, 0, 0, -12,
    -- filter=180 channel=115
    3, -1, -3, -3, -3, 2, 6, -7, -7,
    -- filter=180 channel=116
    10, 8, 6, -11, -7, -2, -16, -15, -8,
    -- filter=180 channel=117
    -1, 3, 5, -5, -3, 7, 1, -4, -3,
    -- filter=180 channel=118
    1, 3, 0, 5, 1, 5, -7, 0, 1,
    -- filter=180 channel=119
    6, -7, 6, -2, -6, -5, -5, 0, 4,
    -- filter=180 channel=120
    4, -5, -13, -3, -6, -17, -7, -10, -11,
    -- filter=180 channel=121
    7, 3, 2, 4, 0, 3, -8, -11, -6,
    -- filter=180 channel=122
    20, 12, 9, 13, 4, 0, -3, -6, -5,
    -- filter=180 channel=123
    9, 2, 0, 0, 1, 2, 1, 0, 2,
    -- filter=180 channel=124
    -5, 3, 1, -3, -4, -1, -4, -4, -3,
    -- filter=180 channel=125
    8, 7, 7, -11, -8, 0, -16, -9, -10,
    -- filter=180 channel=126
    0, 12, -3, -1, 9, 6, -6, -1, 0,
    -- filter=180 channel=127
    3, -6, 4, 0, 1, -7, 0, -1, -7,
    -- filter=181 channel=0
    3, 7, 6, 6, 3, -1, 6, 2, 3,
    -- filter=181 channel=1
    -1, -2, 0, 4, 3, -3, -4, 1, 1,
    -- filter=181 channel=2
    1, 4, 0, 0, 1, -5, 0, 0, 0,
    -- filter=181 channel=3
    -6, -8, 0, -6, -10, -10, -1, 1, -4,
    -- filter=181 channel=4
    -9, -2, -12, 0, -6, -3, 0, 2, 2,
    -- filter=181 channel=5
    2, -7, 3, 0, -1, -1, 0, -2, -7,
    -- filter=181 channel=6
    0, 3, 3, 2, 0, 0, 0, 1, -7,
    -- filter=181 channel=7
    0, -5, 6, 0, -5, -6, 3, 0, 0,
    -- filter=181 channel=8
    -7, -5, -5, -5, -8, -5, 1, 0, 4,
    -- filter=181 channel=9
    -2, 6, 4, 6, 2, 4, 6, 0, 4,
    -- filter=181 channel=10
    -15, 2, 0, -4, 4, -7, 3, 4, 7,
    -- filter=181 channel=11
    -4, 4, -7, 4, 10, 4, -3, 6, -5,
    -- filter=181 channel=12
    0, -8, 0, -12, 0, -2, -1, 3, 0,
    -- filter=181 channel=13
    -2, -5, 1, -9, 4, 7, -7, 2, 7,
    -- filter=181 channel=14
    -7, -5, -4, 6, 0, 6, -1, 5, 2,
    -- filter=181 channel=15
    -1, 3, -7, -6, 8, -6, 1, 8, -6,
    -- filter=181 channel=16
    2, -7, 4, -5, -13, -8, 0, -10, 0,
    -- filter=181 channel=17
    0, -5, 0, 6, -6, 5, -5, -6, 1,
    -- filter=181 channel=18
    -2, 0, 0, -2, 12, -4, 3, 7, -2,
    -- filter=181 channel=19
    -5, 4, 2, -2, 2, -1, -1, 3, -4,
    -- filter=181 channel=20
    -14, 0, -5, -8, 3, -2, -11, 1, -11,
    -- filter=181 channel=21
    -2, -1, 9, 4, -6, 5, 0, 3, 0,
    -- filter=181 channel=22
    1, -3, 6, 0, -3, -4, 6, -6, -6,
    -- filter=181 channel=23
    -1, 0, -10, -3, -5, -3, 8, 0, 0,
    -- filter=181 channel=24
    3, 0, 5, 3, 3, 0, -3, 2, 2,
    -- filter=181 channel=25
    -2, 2, 2, -1, -2, 7, -6, 3, 6,
    -- filter=181 channel=26
    -4, 3, 3, 0, 3, 0, 5, 0, -9,
    -- filter=181 channel=27
    0, 4, 4, -3, 7, -2, 7, 18, -2,
    -- filter=181 channel=28
    5, 0, 3, 3, -2, -4, 2, -4, 3,
    -- filter=181 channel=29
    -1, -3, -2, -6, -5, -2, -6, -4, -5,
    -- filter=181 channel=30
    5, 2, -2, 7, -4, -4, 9, 0, 6,
    -- filter=181 channel=31
    3, -2, 9, 0, -4, 5, 10, 9, 0,
    -- filter=181 channel=32
    0, 6, -9, -4, 0, -8, -1, 6, -1,
    -- filter=181 channel=33
    1, -5, 0, -5, 4, 0, 2, 6, 7,
    -- filter=181 channel=34
    -7, -14, -6, -8, -14, -7, -4, -19, 2,
    -- filter=181 channel=35
    0, 4, -7, 6, 6, 2, -2, 5, 4,
    -- filter=181 channel=36
    -8, -3, -3, -8, 2, 1, -7, -3, 5,
    -- filter=181 channel=37
    10, 2, 3, 7, -1, -1, 1, 0, -3,
    -- filter=181 channel=38
    -7, -3, 4, -1, 0, -8, 3, 7, 4,
    -- filter=181 channel=39
    0, -1, -1, -1, -4, 0, -4, 2, -5,
    -- filter=181 channel=40
    -3, 4, -1, 0, 6, -5, -2, 6, 5,
    -- filter=181 channel=41
    -22, -17, -2, -19, -25, -5, -15, -10, 8,
    -- filter=181 channel=42
    0, 0, 4, 7, 5, 5, 7, 8, 3,
    -- filter=181 channel=43
    1, -8, -9, -13, 0, -8, 1, -1, 0,
    -- filter=181 channel=44
    8, -5, 4, 0, -6, 0, -2, 6, -2,
    -- filter=181 channel=45
    0, -3, 5, 3, 6, -3, 8, -3, 4,
    -- filter=181 channel=46
    -3, -1, -3, 5, -9, -5, 3, -2, 5,
    -- filter=181 channel=47
    0, -7, -1, 2, -8, 9, 7, 7, 13,
    -- filter=181 channel=48
    6, -4, 2, 6, 0, 0, 9, 13, 2,
    -- filter=181 channel=49
    3, 8, -11, 2, 0, -9, 9, 6, -8,
    -- filter=181 channel=50
    0, 9, 7, 0, 2, -3, 11, 6, 8,
    -- filter=181 channel=51
    3, -3, 5, -7, -1, 1, 0, 0, -2,
    -- filter=181 channel=52
    -10, -4, -6, -4, -3, -4, -9, 2, -6,
    -- filter=181 channel=53
    0, 0, -3, 3, 1, -6, 0, -4, 0,
    -- filter=181 channel=54
    6, -5, 0, -2, 5, 0, 0, -6, -5,
    -- filter=181 channel=55
    -11, 0, 2, 0, -3, -1, 5, 9, -7,
    -- filter=181 channel=56
    -9, -8, -3, -11, -12, -4, -1, -3, 0,
    -- filter=181 channel=57
    2, -5, 0, -2, -1, 6, -9, -4, -4,
    -- filter=181 channel=58
    3, 1, -5, -1, 3, -5, 3, 0, -7,
    -- filter=181 channel=59
    -5, 0, 5, -1, 11, 4, 4, 4, 10,
    -- filter=181 channel=60
    0, 4, 0, -4, -1, 4, -1, 4, -5,
    -- filter=181 channel=61
    -2, -10, 4, -7, -8, 5, 0, -7, -4,
    -- filter=181 channel=62
    3, 3, 5, -6, -3, 2, -7, -6, -7,
    -- filter=181 channel=63
    -5, 4, 0, 4, -6, -7, 0, -7, -5,
    -- filter=181 channel=64
    -6, -7, -1, 5, 3, -6, 3, -2, 6,
    -- filter=181 channel=65
    6, -3, -6, 4, 1, -6, -5, 1, -2,
    -- filter=181 channel=66
    -10, -4, -8, -14, -17, 4, -6, -13, -6,
    -- filter=181 channel=67
    0, -4, 1, -5, -6, -3, 0, -6, 2,
    -- filter=181 channel=68
    2, -4, -6, 2, -1, -5, 2, 7, -5,
    -- filter=181 channel=69
    1, 3, 0, 3, 1, 3, 4, -1, 1,
    -- filter=181 channel=70
    0, 9, -3, -5, 6, 2, 0, 3, 4,
    -- filter=181 channel=71
    3, -5, -1, -6, -8, 2, -3, 3, 3,
    -- filter=181 channel=72
    0, -3, 5, 0, 3, 5, 2, 7, 3,
    -- filter=181 channel=73
    -8, -5, 1, -3, -2, -1, 5, 0, 0,
    -- filter=181 channel=74
    -2, 0, 1, -4, -4, -6, 8, -3, 0,
    -- filter=181 channel=75
    -4, -2, -7, -2, -9, -3, 5, -2, 9,
    -- filter=181 channel=76
    -4, 0, 0, -9, 3, -8, -5, -5, -12,
    -- filter=181 channel=77
    5, 2, 6, -5, 0, 4, 4, -4, -7,
    -- filter=181 channel=78
    -3, -2, 1, 3, 2, -6, -2, 1, -2,
    -- filter=181 channel=79
    -4, -4, 0, -9, 4, 2, 1, 7, -6,
    -- filter=181 channel=80
    -8, 0, 4, -3, 4, -1, 6, 18, 4,
    -- filter=181 channel=81
    -6, 2, 3, 5, 3, 1, -6, 0, -6,
    -- filter=181 channel=82
    -7, 0, 1, -2, 1, 4, 6, 1, -8,
    -- filter=181 channel=83
    0, 8, -1, 0, -1, 1, 4, 1, 11,
    -- filter=181 channel=84
    -2, -6, -8, -1, -1, 0, 3, -4, 3,
    -- filter=181 channel=85
    0, 0, -2, 2, 2, 1, -1, 3, -1,
    -- filter=181 channel=86
    6, 0, -6, 3, -13, -5, -9, -13, -8,
    -- filter=181 channel=87
    -12, -1, -9, -8, -8, -1, -13, -8, -10,
    -- filter=181 channel=88
    -9, -7, 6, -3, -11, -2, 4, 2, 3,
    -- filter=181 channel=89
    -7, -1, 4, 0, 2, 8, -2, 12, 3,
    -- filter=181 channel=90
    -7, -4, -2, -11, -13, -5, 0, -9, 0,
    -- filter=181 channel=91
    3, 4, 0, 9, 5, -2, 8, 12, 4,
    -- filter=181 channel=92
    -6, 0, -2, -7, 0, 4, -9, -6, -2,
    -- filter=181 channel=93
    -2, -7, 3, 6, -5, 5, 8, 0, -1,
    -- filter=181 channel=94
    0, 7, -5, 4, -1, 4, 0, 5, 2,
    -- filter=181 channel=95
    -3, -2, 2, -5, -7, -4, -4, -6, 3,
    -- filter=181 channel=96
    -6, -5, -5, 7, -4, 4, -2, 8, 3,
    -- filter=181 channel=97
    -8, 3, -9, 3, -4, 0, 0, 0, -3,
    -- filter=181 channel=98
    0, 5, 5, 5, 6, -6, 0, 15, -2,
    -- filter=181 channel=99
    -14, -10, 4, -5, 3, 0, 4, -1, 0,
    -- filter=181 channel=100
    0, -8, -7, -9, -7, -2, 2, -9, -6,
    -- filter=181 channel=101
    0, -9, -9, 3, -11, -6, -6, 0, -1,
    -- filter=181 channel=102
    -1, -4, -1, 7, 3, -2, -4, 5, -3,
    -- filter=181 channel=103
    2, -11, 10, -2, 0, 5, -2, 6, 0,
    -- filter=181 channel=104
    -1, -1, -1, -4, 4, 6, 3, 1, 5,
    -- filter=181 channel=105
    -11, -2, -8, 1, 1, -12, 1, -2, -11,
    -- filter=181 channel=106
    -6, -6, -1, 5, 3, -5, -4, -6, -8,
    -- filter=181 channel=107
    6, -6, -7, -3, 0, -4, -2, 3, -7,
    -- filter=181 channel=108
    0, 0, 3, -12, -7, 3, -10, -2, 2,
    -- filter=181 channel=109
    0, 3, -8, -1, 8, 9, 1, 17, 4,
    -- filter=181 channel=110
    -11, -7, 6, 2, -7, 0, 6, 0, -4,
    -- filter=181 channel=111
    -1, 2, 2, -5, -7, 0, -3, -4, 4,
    -- filter=181 channel=112
    1, -3, -3, 9, 5, 4, 3, 7, 6,
    -- filter=181 channel=113
    0, -11, 3, -1, 3, 4, 6, 7, 6,
    -- filter=181 channel=114
    7, -2, 0, -1, 0, -6, 0, 13, -8,
    -- filter=181 channel=115
    -4, 1, -1, -6, 0, 5, 0, 7, 5,
    -- filter=181 channel=116
    -7, 5, 4, -4, 1, 2, -2, 5, 0,
    -- filter=181 channel=117
    4, -6, -4, 1, 4, -1, 4, 5, -6,
    -- filter=181 channel=118
    -3, -6, 2, 6, 5, 0, 4, 2, -3,
    -- filter=181 channel=119
    -15, -6, 4, -9, -13, -5, 0, -4, 3,
    -- filter=181 channel=120
    4, -2, 2, 4, 4, -6, 14, 13, -2,
    -- filter=181 channel=121
    -6, -10, 2, -2, -6, 7, -4, -3, 9,
    -- filter=181 channel=122
    -8, -12, 5, 0, -4, 4, -3, 0, 10,
    -- filter=181 channel=123
    0, -2, -2, -1, -8, 1, 3, 1, -3,
    -- filter=181 channel=124
    -4, 0, -1, -6, 6, 0, -2, -3, -8,
    -- filter=181 channel=125
    0, 4, -5, -1, 7, 0, 6, 4, 6,
    -- filter=181 channel=126
    -5, 0, -4, -12, -3, -2, -1, 0, 0,
    -- filter=181 channel=127
    -2, -12, -2, -2, 1, 2, -9, -5, -4,
    -- filter=182 channel=0
    -16, -6, 13, -5, 0, 0, 9, -3, 1,
    -- filter=182 channel=1
    -1, -1, 6, 5, 0, 6, 9, -4, 4,
    -- filter=182 channel=2
    10, 6, -5, 0, -8, 0, -11, 1, -3,
    -- filter=182 channel=3
    -6, 0, 13, -4, 16, -2, 7, 5, 0,
    -- filter=182 channel=4
    2, 1, -6, 4, 1, 8, -12, 0, 5,
    -- filter=182 channel=5
    -10, -9, 4, 7, -2, -8, 0, -6, -4,
    -- filter=182 channel=6
    -9, -7, 0, 4, 0, 8, -5, -3, -2,
    -- filter=182 channel=7
    -6, 0, 3, -3, 1, 2, -7, 1, -1,
    -- filter=182 channel=8
    10, 12, 2, 11, 1, -2, -1, 13, 6,
    -- filter=182 channel=9
    -2, 0, -1, 3, -8, -2, -2, -11, -1,
    -- filter=182 channel=10
    7, 9, 0, 15, 9, -10, 7, -11, -4,
    -- filter=182 channel=11
    -7, -6, -7, 1, 1, 1, 0, -1, 8,
    -- filter=182 channel=12
    -4, -4, 7, 0, 12, -5, 7, -1, 4,
    -- filter=182 channel=13
    6, 6, 4, 4, 13, -2, 8, -5, 3,
    -- filter=182 channel=14
    0, 0, 0, -2, -2, -3, 0, -1, 7,
    -- filter=182 channel=15
    -5, -10, 6, -7, 2, -1, 2, 2, 6,
    -- filter=182 channel=16
    7, -3, 4, 15, 9, -2, 8, -2, -17,
    -- filter=182 channel=17
    -2, 0, 4, 3, -4, -6, 6, -4, 3,
    -- filter=182 channel=18
    -5, -6, 2, 4, 5, 3, 3, -12, -2,
    -- filter=182 channel=19
    -5, 0, -5, 0, 3, -4, -3, -3, -3,
    -- filter=182 channel=20
    5, -13, -4, 2, -3, 0, 5, 6, 10,
    -- filter=182 channel=21
    13, 5, 1, 10, 6, -12, 12, -6, -18,
    -- filter=182 channel=22
    -8, 0, -5, -2, 0, 7, -3, -3, 4,
    -- filter=182 channel=23
    0, 8, -12, 0, -2, 4, 1, -11, -1,
    -- filter=182 channel=24
    -3, 5, 4, 5, 1, 1, 0, -1, 2,
    -- filter=182 channel=25
    -2, -4, -2, 15, 0, -14, -5, -20, -1,
    -- filter=182 channel=26
    6, 4, -8, 8, -5, -5, 3, -2, -7,
    -- filter=182 channel=27
    -8, 9, -2, 6, -16, -15, -10, -23, 7,
    -- filter=182 channel=28
    -5, -2, -2, 2, 3, 3, 0, -3, 3,
    -- filter=182 channel=29
    -5, -3, 2, -3, -3, 0, 0, -3, 6,
    -- filter=182 channel=30
    -5, 6, 8, 2, 2, -5, -11, -11, 0,
    -- filter=182 channel=31
    14, 6, -12, 26, -7, -21, -7, -31, -17,
    -- filter=182 channel=32
    -4, 2, 2, 9, 0, -8, 0, -11, 4,
    -- filter=182 channel=33
    -1, 4, -2, 10, 8, -5, 5, -6, -10,
    -- filter=182 channel=34
    -3, 4, -10, 4, -1, -3, 0, 11, 6,
    -- filter=182 channel=35
    6, -6, -1, 0, 0, -2, 1, 1, -1,
    -- filter=182 channel=36
    16, 7, -10, 1, 3, -4, 3, 2, -2,
    -- filter=182 channel=37
    -4, 4, 1, 1, 0, -3, -4, 6, 5,
    -- filter=182 channel=38
    -1, 3, 2, 9, 0, -2, 4, -14, -8,
    -- filter=182 channel=39
    -7, -9, -10, -5, 0, 4, 0, 8, 7,
    -- filter=182 channel=40
    0, -1, 5, 4, 0, 10, 0, -3, 7,
    -- filter=182 channel=41
    8, -9, 1, 7, 5, 5, 22, 8, -4,
    -- filter=182 channel=42
    -7, -5, 0, 2, -6, -2, -2, -8, -3,
    -- filter=182 channel=43
    0, -7, 8, 0, 13, 9, 0, 12, 5,
    -- filter=182 channel=44
    1, 6, -1, 14, -1, 0, -7, -2, 5,
    -- filter=182 channel=45
    3, -5, -1, -4, -7, 5, 0, -7, 6,
    -- filter=182 channel=46
    -5, -5, 0, 2, -2, 3, 4, 5, 1,
    -- filter=182 channel=47
    12, -2, -3, 22, 6, -19, 2, -21, -9,
    -- filter=182 channel=48
    5, 14, -4, 11, 1, -8, -14, -24, 5,
    -- filter=182 channel=49
    -3, -5, -3, -4, -12, -7, -10, 0, 12,
    -- filter=182 channel=50
    4, 2, 0, 11, -14, 1, -4, -6, 0,
    -- filter=182 channel=51
    0, 4, -5, -4, 0, -4, 7, 7, -5,
    -- filter=182 channel=52
    3, 4, -8, 8, -8, 9, 4, 0, 3,
    -- filter=182 channel=53
    0, -8, -4, 0, -5, -3, -5, 0, -1,
    -- filter=182 channel=54
    -2, 0, -1, -4, 3, 1, -6, -3, 5,
    -- filter=182 channel=55
    -2, -1, -6, -1, 0, 0, 2, -7, -3,
    -- filter=182 channel=56
    12, 2, -8, 0, -3, 10, -5, 14, -2,
    -- filter=182 channel=57
    0, -2, 4, 1, 5, -2, 1, -9, 0,
    -- filter=182 channel=58
    -7, -1, -5, 0, -3, 0, 6, 0, -2,
    -- filter=182 channel=59
    8, 2, 1, 11, -2, -14, 0, -13, -8,
    -- filter=182 channel=60
    0, 0, 1, 3, -6, -6, 6, -2, 7,
    -- filter=182 channel=61
    8, 2, -4, 5, -3, 1, -2, -3, 0,
    -- filter=182 channel=62
    6, 0, 4, 5, 3, 5, -3, 4, -3,
    -- filter=182 channel=63
    -5, -1, 4, -1, 1, 0, 8, -8, -2,
    -- filter=182 channel=64
    3, 0, -7, 8, -5, 3, -1, 9, -7,
    -- filter=182 channel=65
    -1, -2, 0, 4, 0, 6, 0, 5, 4,
    -- filter=182 channel=66
    5, -3, -3, 1, 12, -5, 10, 3, -3,
    -- filter=182 channel=67
    -7, 0, 4, -2, 1, -5, 4, 1, 4,
    -- filter=182 channel=68
    3, 2, 0, -2, 4, 5, -3, -2, -3,
    -- filter=182 channel=69
    3, -4, 0, 1, 7, 0, 1, 4, -6,
    -- filter=182 channel=70
    0, 9, -3, -4, -6, 2, -5, 1, 10,
    -- filter=182 channel=71
    -1, -5, 1, -4, -3, -1, 10, 4, -2,
    -- filter=182 channel=72
    5, 7, 4, 14, -2, -12, -5, -22, -16,
    -- filter=182 channel=73
    6, -1, 1, 9, -5, -3, -10, -13, 0,
    -- filter=182 channel=74
    3, 0, -8, 11, -7, 3, 1, 5, 0,
    -- filter=182 channel=75
    -3, -3, 18, 6, 18, 3, 15, 4, -3,
    -- filter=182 channel=76
    0, -8, 0, -6, -2, 10, 10, 5, -1,
    -- filter=182 channel=77
    6, 6, -6, 0, -3, -7, 0, 4, -5,
    -- filter=182 channel=78
    -5, 0, -1, -2, 5, -2, 0, -4, 3,
    -- filter=182 channel=79
    -17, -10, 0, 7, 1, -4, 2, -8, 7,
    -- filter=182 channel=80
    3, 5, 8, 20, -4, -26, 9, -28, -13,
    -- filter=182 channel=81
    6, 5, 0, -3, 6, -7, 0, -6, -1,
    -- filter=182 channel=82
    3, 0, -6, -4, 0, 0, -3, -4, -6,
    -- filter=182 channel=83
    9, 0, -3, 7, -6, 4, -4, -4, 5,
    -- filter=182 channel=84
    2, -4, 2, 0, -6, 5, -8, -8, 3,
    -- filter=182 channel=85
    -5, -6, -1, 7, 4, 1, -5, -4, 3,
    -- filter=182 channel=86
    3, -1, 0, 0, 5, 0, 10, 8, 7,
    -- filter=182 channel=87
    6, -6, -2, 7, 0, 1, 6, 9, 0,
    -- filter=182 channel=88
    10, 1, -2, 3, 0, -10, 2, 0, 2,
    -- filter=182 channel=89
    3, 7, 11, 7, 13, -15, 13, -14, -14,
    -- filter=182 channel=90
    14, 9, -6, 9, -2, 0, 0, 8, -8,
    -- filter=182 channel=91
    6, 8, -11, 7, -15, 1, -14, -10, 7,
    -- filter=182 channel=92
    -7, 0, -3, -3, 6, -1, 0, -3, 8,
    -- filter=182 channel=93
    4, 7, -2, 12, 2, -15, -4, -9, 0,
    -- filter=182 channel=94
    7, -7, -3, 4, 2, 7, 0, 0, -5,
    -- filter=182 channel=95
    7, 2, -2, -2, -2, 5, 1, -2, -6,
    -- filter=182 channel=96
    0, -9, 8, 5, 1, 2, 3, 2, -4,
    -- filter=182 channel=97
    0, 0, 5, -4, 9, 7, 12, -2, -6,
    -- filter=182 channel=98
    -4, -6, 0, 6, 1, -11, -3, -15, 0,
    -- filter=182 channel=99
    15, 4, -7, 13, -5, -11, -10, -21, 3,
    -- filter=182 channel=100
    -1, -2, -6, -2, 3, 6, -2, 0, -7,
    -- filter=182 channel=101
    8, 8, 0, 5, -6, -6, -5, 0, 5,
    -- filter=182 channel=102
    5, 0, -1, 7, 4, 2, 4, 0, 7,
    -- filter=182 channel=103
    0, -3, -5, 17, 0, -5, 16, -10, -10,
    -- filter=182 channel=104
    11, 6, -3, 10, 0, -7, 3, -13, -16,
    -- filter=182 channel=105
    0, -2, 1, -2, 0, 5, 9, 9, 6,
    -- filter=182 channel=106
    -6, -4, -5, 0, -2, 5, 5, 7, 5,
    -- filter=182 channel=107
    -8, 0, -8, -3, 0, 7, -8, 6, 3,
    -- filter=182 channel=108
    -3, 1, 0, -1, 6, 0, 6, 3, 0,
    -- filter=182 channel=109
    -3, -1, -11, 12, -4, -9, -6, -20, -3,
    -- filter=182 channel=110
    1, 0, -9, 4, 3, -2, 5, 1, -8,
    -- filter=182 channel=111
    -4, -8, -6, -1, -1, -2, 4, 0, -5,
    -- filter=182 channel=112
    3, 0, -2, 5, -6, 0, -5, -7, 3,
    -- filter=182 channel=113
    2, -6, 7, 0, -2, -9, 5, -1, -7,
    -- filter=182 channel=114
    -19, -2, 0, -2, -6, -10, -9, -5, 10,
    -- filter=182 channel=115
    1, -3, -7, 7, -5, -4, -5, 2, 3,
    -- filter=182 channel=116
    2, -1, -4, 3, -10, -5, -4, -22, 2,
    -- filter=182 channel=117
    -3, 8, -5, 8, -2, -5, -5, -3, -4,
    -- filter=182 channel=118
    -2, 0, -7, 3, 1, -5, 3, -1, 4,
    -- filter=182 channel=119
    7, -1, -3, 10, 1, 7, -5, 6, 1,
    -- filter=182 channel=120
    0, 9, -9, 6, -12, -3, -17, 0, 11,
    -- filter=182 channel=121
    9, -3, 7, 13, 4, 3, 6, -5, -7,
    -- filter=182 channel=122
    26, 3, -6, 33, 3, -16, 17, -15, -21,
    -- filter=182 channel=123
    -5, 2, -2, 0, 0, 5, 5, 5, -3,
    -- filter=182 channel=124
    -9, -9, 4, -2, -1, 2, 5, 1, 3,
    -- filter=182 channel=125
    10, 7, 1, 20, -10, -9, -3, -24, -1,
    -- filter=182 channel=126
    -10, -1, 9, 8, 11, -9, 16, 1, -3,
    -- filter=182 channel=127
    -3, 0, 0, 7, -3, 2, 11, 5, 4,
    -- filter=183 channel=0
    -8, -18, -10, -4, -19, -21, 7, -15, -5,
    -- filter=183 channel=1
    -7, -18, -15, 4, -17, -24, 4, -11, -17,
    -- filter=183 channel=2
    -6, 0, -5, -6, 6, 0, -5, 7, 3,
    -- filter=183 channel=3
    -1, -12, -5, -5, -3, -13, 5, -4, 3,
    -- filter=183 channel=4
    0, -13, -12, -10, -12, -14, -7, -6, 0,
    -- filter=183 channel=5
    -2, -3, 0, -1, -3, -8, -1, -10, 0,
    -- filter=183 channel=6
    2, 6, -1, -5, 1, 6, 3, 1, -3,
    -- filter=183 channel=7
    -4, 0, 4, 1, 6, -7, 2, -2, -5,
    -- filter=183 channel=8
    0, 1, -1, 4, -10, 5, -2, 2, 4,
    -- filter=183 channel=9
    0, 0, -4, 4, 1, 0, 5, -5, 7,
    -- filter=183 channel=10
    0, 6, 5, -3, -6, 5, -3, 4, 2,
    -- filter=183 channel=11
    2, 3, 15, 0, 16, 13, -5, 7, 15,
    -- filter=183 channel=12
    -6, 4, 3, -2, -2, -2, -6, -9, 5,
    -- filter=183 channel=13
    4, 0, -1, 7, -3, 2, -6, -7, 2,
    -- filter=183 channel=14
    7, 1, 6, 0, 0, -7, 5, -1, 2,
    -- filter=183 channel=15
    4, -8, 8, -8, -5, 3, -9, -2, 3,
    -- filter=183 channel=16
    -7, -5, 0, 3, 0, -1, -2, 0, -8,
    -- filter=183 channel=17
    -5, -3, 5, -2, 7, 0, 0, 3, 0,
    -- filter=183 channel=18
    5, -6, 1, -10, 2, -4, 6, -9, 6,
    -- filter=183 channel=19
    -1, -4, 0, 5, 1, 6, -3, 0, 6,
    -- filter=183 channel=20
    -4, 9, 19, -17, 16, 17, -15, 2, 14,
    -- filter=183 channel=21
    -3, 2, -4, 0, -8, -8, 4, -9, -10,
    -- filter=183 channel=22
    0, -9, 2, -8, -12, -3, -6, 0, 0,
    -- filter=183 channel=23
    1, -4, 16, 4, 0, 23, -1, -5, 21,
    -- filter=183 channel=24
    0, 2, 4, 1, 7, 7, -2, -1, 5,
    -- filter=183 channel=25
    9, -12, -6, 12, -6, -7, 1, -2, 0,
    -- filter=183 channel=26
    1, -4, -3, 5, -2, 5, -4, -8, 5,
    -- filter=183 channel=27
    8, -10, 4, 3, -10, 8, 4, -14, 5,
    -- filter=183 channel=28
    5, -6, -6, 1, 1, -1, 6, 2, -3,
    -- filter=183 channel=29
    -8, 9, 17, -11, 14, 27, -17, -3, 16,
    -- filter=183 channel=30
    0, -11, 0, 7, -15, -4, 3, -5, -4,
    -- filter=183 channel=31
    7, 1, 0, 12, -8, 1, 6, -2, 1,
    -- filter=183 channel=32
    3, -11, 0, 5, -15, 8, -1, -9, 2,
    -- filter=183 channel=33
    10, -3, 4, 4, -15, -1, 7, 0, -2,
    -- filter=183 channel=34
    4, -4, 0, -10, -1, -2, -4, -2, -6,
    -- filter=183 channel=35
    -3, -6, -6, 7, 6, -3, -1, 6, -4,
    -- filter=183 channel=36
    -1, 0, 10, 1, -1, 12, -3, -7, -2,
    -- filter=183 channel=37
    0, -17, -18, 8, -14, -21, -1, -6, -22,
    -- filter=183 channel=38
    9, -2, -2, 4, -1, 1, 9, -1, 11,
    -- filter=183 channel=39
    -3, 2, 0, 3, 2, 5, -3, -3, 2,
    -- filter=183 channel=40
    -5, 4, -3, -7, 4, 7, -1, 1, 5,
    -- filter=183 channel=41
    14, 2, 3, -3, 15, -14, 0, 3, -8,
    -- filter=183 channel=42
    1, 1, -5, 4, -4, -10, 3, 6, -3,
    -- filter=183 channel=43
    -6, -4, 0, 0, -11, -7, -2, 0, -2,
    -- filter=183 channel=44
    6, -16, -9, 0, -12, -15, 4, -8, -10,
    -- filter=183 channel=45
    -1, -4, -1, 3, -7, 1, -2, -6, 5,
    -- filter=183 channel=46
    -5, -6, -1, 0, 2, -3, 7, 2, -7,
    -- filter=183 channel=47
    -2, -7, -3, 8, -12, -14, 2, -12, -2,
    -- filter=183 channel=48
    6, -9, -7, 6, -10, -9, 12, -4, 1,
    -- filter=183 channel=49
    -1, 2, 2, -1, -5, -3, -6, 7, 6,
    -- filter=183 channel=50
    -1, -5, 2, 3, -12, 6, 10, -1, 13,
    -- filter=183 channel=51
    -5, -1, -5, -3, -1, -1, 5, -4, 0,
    -- filter=183 channel=52
    -9, 0, 9, -12, -10, 8, -11, 0, -4,
    -- filter=183 channel=53
    -7, 4, 0, 1, 5, 14, 0, 0, 2,
    -- filter=183 channel=54
    7, -5, -5, -1, 2, 4, 5, 4, 5,
    -- filter=183 channel=55
    -4, -6, 7, -8, 0, 17, -7, -3, 13,
    -- filter=183 channel=56
    5, 4, -1, -4, 5, -5, -6, 8, -5,
    -- filter=183 channel=57
    -5, 4, 1, -4, -2, 3, 6, 4, 0,
    -- filter=183 channel=58
    -1, -3, -5, 6, -4, -6, -3, 0, -2,
    -- filter=183 channel=59
    9, 0, 2, 6, -3, -6, 11, -1, -3,
    -- filter=183 channel=60
    -4, 0, 2, -7, 0, 5, 5, -6, 2,
    -- filter=183 channel=61
    -6, -1, -1, -1, 4, 6, -10, -2, 3,
    -- filter=183 channel=62
    2, 0, -7, -4, 0, -5, -7, -6, 5,
    -- filter=183 channel=63
    -2, 6, -3, 2, 6, 0, -1, -4, -6,
    -- filter=183 channel=64
    0, 3, 9, -4, 9, -2, -6, -4, 1,
    -- filter=183 channel=65
    -5, -4, 0, 3, -2, 5, 6, 0, 2,
    -- filter=183 channel=66
    -6, 3, 5, -2, 9, -1, -7, -2, 0,
    -- filter=183 channel=67
    6, -6, 0, 1, 4, 5, -3, 1, 7,
    -- filter=183 channel=68
    -4, 4, -2, 1, 0, -6, 5, 1, -5,
    -- filter=183 channel=69
    -3, -1, 2, -4, -4, -3, 4, 0, 5,
    -- filter=183 channel=70
    3, -8, 6, 6, -7, 1, -5, 2, 5,
    -- filter=183 channel=71
    -2, -2, -1, -1, -3, -4, 3, -6, 0,
    -- filter=183 channel=72
    15, 3, 2, 5, 4, 9, 6, -2, 10,
    -- filter=183 channel=73
    2, -4, 6, 2, -5, 4, -7, -7, 8,
    -- filter=183 channel=74
    7, -13, 10, 2, -3, 0, 1, 0, 2,
    -- filter=183 channel=75
    -2, -16, -22, -4, -18, -19, 0, -12, -3,
    -- filter=183 channel=76
    -5, -2, 13, -9, 3, 19, -7, 0, 5,
    -- filter=183 channel=77
    -6, -4, -7, 0, -5, 0, -1, -4, 2,
    -- filter=183 channel=78
    -2, 5, -6, 2, -1, 4, 0, 2, -4,
    -- filter=183 channel=79
    0, -11, -5, 2, -12, 0, 4, -8, 12,
    -- filter=183 channel=80
    13, 0, 4, 8, -10, -7, 14, -9, -3,
    -- filter=183 channel=81
    1, 0, -6, 3, -4, 0, 4, 7, 0,
    -- filter=183 channel=82
    0, 7, -6, 2, 7, 3, -2, -3, 4,
    -- filter=183 channel=83
    9, -1, 4, 7, -7, -3, -4, 0, 1,
    -- filter=183 channel=84
    -5, -11, 9, 2, -1, 7, 0, -6, 7,
    -- filter=183 channel=85
    4, 6, -4, 3, 0, 5, -3, -1, 3,
    -- filter=183 channel=86
    -6, -10, 5, 6, -6, 1, 5, -2, -3,
    -- filter=183 channel=87
    -5, 2, 6, -14, -3, 7, -5, 4, 7,
    -- filter=183 channel=88
    -5, 9, 11, 0, 9, 0, -5, -6, 10,
    -- filter=183 channel=89
    13, -5, 9, 9, 0, 10, 13, 4, 2,
    -- filter=183 channel=90
    -7, -4, 3, 0, -1, 10, -5, 3, 0,
    -- filter=183 channel=91
    6, -10, 9, 5, -3, 13, -8, 0, 8,
    -- filter=183 channel=92
    -7, -1, 4, 4, -6, -3, 0, 3, 1,
    -- filter=183 channel=93
    2, -7, -14, 0, -14, -19, -4, -13, -5,
    -- filter=183 channel=94
    -6, -7, -2, -6, 2, 2, 2, 4, -7,
    -- filter=183 channel=95
    4, 2, 6, -1, -1, -6, 4, 2, -5,
    -- filter=183 channel=96
    8, 0, 1, -3, 4, -2, -2, 5, -6,
    -- filter=183 channel=97
    0, -10, -8, -3, -5, -13, -1, -3, 3,
    -- filter=183 channel=98
    3, -12, 3, 14, -18, 2, 9, -12, -3,
    -- filter=183 channel=99
    -1, 1, 16, 2, -3, 20, -12, 2, 17,
    -- filter=183 channel=100
    0, 11, 3, 2, 2, 2, -5, 10, 3,
    -- filter=183 channel=101
    0, -1, -8, -6, -6, -8, -4, 2, -2,
    -- filter=183 channel=102
    -3, 4, 0, -1, 0, -3, -3, -1, 5,
    -- filter=183 channel=103
    0, 0, -12, 0, -19, -17, 6, -9, -5,
    -- filter=183 channel=104
    7, -1, 3, 7, -7, 0, 1, -4, -2,
    -- filter=183 channel=105
    -5, 0, 9, 0, 4, 9, -14, -4, 8,
    -- filter=183 channel=106
    2, 8, 3, -3, 5, -4, 0, 8, 6,
    -- filter=183 channel=107
    -1, -9, 1, -9, -2, 1, -4, 3, 6,
    -- filter=183 channel=108
    6, 4, 1, 0, 8, -5, -1, 6, 0,
    -- filter=183 channel=109
    5, -11, 6, -1, -5, 0, 3, -13, 10,
    -- filter=183 channel=110
    -1, 7, 6, 6, -5, 5, -4, 1, 0,
    -- filter=183 channel=111
    2, 3, -3, -2, -5, 2, 1, 5, -4,
    -- filter=183 channel=112
    1, -11, 0, 1, -15, 8, 9, -5, 2,
    -- filter=183 channel=113
    1, -7, -3, 8, -6, -6, 7, -4, 5,
    -- filter=183 channel=114
    2, -10, -9, -8, -10, -2, 1, -11, 2,
    -- filter=183 channel=115
    -5, -1, 0, -2, 4, 6, -2, 4, 3,
    -- filter=183 channel=116
    11, 0, 1, 4, 3, 1, 4, -3, 4,
    -- filter=183 channel=117
    9, -1, -2, -2, 3, -3, 7, -3, 0,
    -- filter=183 channel=118
    -5, 6, 0, 6, 0, -5, -1, 1, -1,
    -- filter=183 channel=119
    3, 8, 8, -10, 7, 10, -2, 4, 7,
    -- filter=183 channel=120
    7, -9, 19, 0, -10, 22, -5, -10, 22,
    -- filter=183 channel=121
    0, 1, 1, 0, -4, 4, -5, 1, -1,
    -- filter=183 channel=122
    -3, -10, -5, 4, -8, -16, -9, -10, -11,
    -- filter=183 channel=123
    -3, 5, 3, 4, 2, -5, -1, 3, -2,
    -- filter=183 channel=124
    0, 2, 7, 2, 4, 4, -1, -6, 2,
    -- filter=183 channel=125
    0, -6, 12, 16, -5, 12, 4, -12, 10,
    -- filter=183 channel=126
    0, -5, 2, 0, 7, -6, 6, 2, 5,
    -- filter=183 channel=127
    2, 9, -5, 1, 9, 5, -1, -4, 1,
    -- filter=184 channel=0
    -3, -1, 6, 4, 8, 9, -1, 7, 7,
    -- filter=184 channel=1
    11, 0, 5, -1, 7, 6, 0, 10, 7,
    -- filter=184 channel=2
    1, -4, -1, -4, 3, 0, -4, -5, 3,
    -- filter=184 channel=3
    -10, -10, 0, -7, -2, -1, -3, -3, -7,
    -- filter=184 channel=4
    11, -9, 1, -9, -6, -11, 3, -5, -2,
    -- filter=184 channel=5
    0, 12, 6, -3, 8, 8, 0, 11, 8,
    -- filter=184 channel=6
    7, 5, -2, 4, -7, -6, 4, 4, 1,
    -- filter=184 channel=7
    2, 0, -4, 5, 6, 2, -4, 0, 5,
    -- filter=184 channel=8
    6, -8, -9, -5, -9, 4, 1, -7, -7,
    -- filter=184 channel=9
    -2, -8, -5, 9, 6, -3, 5, 5, 0,
    -- filter=184 channel=10
    -6, -5, -2, -5, 3, 0, 0, 2, -2,
    -- filter=184 channel=11
    4, -7, 3, 0, 7, -2, 7, 0, -3,
    -- filter=184 channel=12
    1, -3, 1, -6, -7, -2, 0, -4, -2,
    -- filter=184 channel=13
    5, -6, -15, 1, -8, -12, 9, -1, -6,
    -- filter=184 channel=14
    -6, -1, 2, 1, -2, 0, 3, 0, -4,
    -- filter=184 channel=15
    0, -8, -11, 0, -8, -16, 6, -9, -19,
    -- filter=184 channel=16
    0, 12, 0, 6, 6, 4, 6, 9, 12,
    -- filter=184 channel=17
    -1, -4, 0, -3, 5, 1, 4, -2, 0,
    -- filter=184 channel=18
    -3, -6, -24, 0, -9, -27, 1, -10, -19,
    -- filter=184 channel=19
    0, 2, 3, -3, 5, -5, -2, 0, -4,
    -- filter=184 channel=20
    10, -10, -10, 12, -1, 1, 7, 1, -8,
    -- filter=184 channel=21
    -2, 8, 9, 6, 23, 8, 1, 8, 7,
    -- filter=184 channel=22
    5, -4, -10, -1, -2, -2, -4, 4, -9,
    -- filter=184 channel=23
    -6, -17, -21, -1, -18, -26, -3, -23, -15,
    -- filter=184 channel=24
    1, 6, -1, 6, -4, 7, 0, 4, -4,
    -- filter=184 channel=25
    -6, 0, -17, 11, -3, -19, 6, -5, -3,
    -- filter=184 channel=26
    3, 9, 5, 8, 7, 11, 4, 6, 11,
    -- filter=184 channel=27
    3, -14, -29, 10, -14, -27, 7, -10, -25,
    -- filter=184 channel=28
    -4, 6, -3, 0, -5, 1, 0, -1, 2,
    -- filter=184 channel=29
    1, -3, -7, 0, 6, 1, 9, 0, -3,
    -- filter=184 channel=30
    -6, 2, -3, 3, -7, -8, 9, 1, 0,
    -- filter=184 channel=31
    -18, -9, -14, -2, -4, -3, 0, -5, 0,
    -- filter=184 channel=32
    5, -15, -22, 0, -5, -22, 6, -6, -13,
    -- filter=184 channel=33
    -5, -15, -20, 9, -7, -17, 10, -14, -13,
    -- filter=184 channel=34
    -4, 2, 2, -8, -7, -14, -6, -12, -10,
    -- filter=184 channel=35
    -6, -6, 4, 0, 3, 7, -3, -6, -2,
    -- filter=184 channel=36
    -4, 0, 3, -4, 2, 8, 1, 8, 0,
    -- filter=184 channel=37
    -2, 0, 10, -1, 5, 1, 0, 4, 12,
    -- filter=184 channel=38
    -7, -8, 0, 8, -4, -1, 7, -6, -5,
    -- filter=184 channel=39
    -2, 6, -2, 6, -4, 0, 1, 3, 6,
    -- filter=184 channel=40
    7, 1, -5, -4, -6, 1, -3, -5, -5,
    -- filter=184 channel=41
    7, 2, -8, 0, 6, 3, 5, 4, -5,
    -- filter=184 channel=42
    -2, 6, -6, -3, 3, -4, 1, 4, -5,
    -- filter=184 channel=43
    2, -4, 0, -7, -6, -9, 1, 4, -2,
    -- filter=184 channel=44
    0, -7, -5, 4, 4, 0, -4, -1, 0,
    -- filter=184 channel=45
    1, 2, -1, 7, 2, -4, -3, 9, 0,
    -- filter=184 channel=46
    -6, -2, -5, -4, 8, 0, 1, -5, -1,
    -- filter=184 channel=47
    -8, 10, 4, -5, 22, 17, 4, 7, 15,
    -- filter=184 channel=48
    7, 3, -14, 6, 7, -4, 7, 9, 0,
    -- filter=184 channel=49
    3, -12, -15, -2, -15, -10, -3, 1, -9,
    -- filter=184 channel=50
    0, -13, -9, 2, -3, -10, 1, -4, -11,
    -- filter=184 channel=51
    -2, 6, 0, 2, -2, -1, -7, 6, -3,
    -- filter=184 channel=52
    -1, 0, 0, 5, -7, -6, -1, -2, -10,
    -- filter=184 channel=53
    -6, -9, -1, -4, -6, 3, 0, -7, -9,
    -- filter=184 channel=54
    6, -5, -7, 3, 0, 0, 1, 3, 0,
    -- filter=184 channel=55
    -5, -13, -17, 6, -10, -23, 9, -19, -24,
    -- filter=184 channel=56
    0, -6, -8, 2, 2, 4, -5, 0, 2,
    -- filter=184 channel=57
    -1, 3, 6, -7, 6, -6, -4, 4, -3,
    -- filter=184 channel=58
    0, 2, 12, 1, 0, 2, 4, 12, 10,
    -- filter=184 channel=59
    -3, 0, -13, 1, 7, -3, 3, -4, -9,
    -- filter=184 channel=60
    7, -2, 8, -3, -6, 7, -2, -3, -2,
    -- filter=184 channel=61
    3, 0, -8, -2, 0, -5, 0, 0, 5,
    -- filter=184 channel=62
    -3, -7, 2, 5, -4, -1, -3, -6, 0,
    -- filter=184 channel=63
    -6, 14, 11, 0, 9, 12, 7, 11, 12,
    -- filter=184 channel=64
    -3, -6, 0, -2, -1, -6, 0, -5, 5,
    -- filter=184 channel=65
    0, 1, 4, -4, -4, 3, -1, 4, 7,
    -- filter=184 channel=66
    1, -2, -9, 6, -3, 4, -4, 2, -2,
    -- filter=184 channel=67
    0, -6, -2, 6, 1, -2, 7, 7, -1,
    -- filter=184 channel=68
    -4, -3, 4, 4, -6, -4, -1, 6, -3,
    -- filter=184 channel=69
    0, 8, 1, 5, 0, 9, 4, 9, 1,
    -- filter=184 channel=70
    3, -13, -20, 5, -16, -22, -3, -8, -11,
    -- filter=184 channel=71
    3, 4, 0, 4, 7, 5, -4, 4, 1,
    -- filter=184 channel=72
    -10, 1, -12, 9, -7, -9, 4, -3, -7,
    -- filter=184 channel=73
    7, -10, -10, -3, -11, -11, -4, 0, -3,
    -- filter=184 channel=74
    -1, -13, -9, 6, -13, -11, 6, -14, -14,
    -- filter=184 channel=75
    5, 11, 0, 5, 11, -1, 3, 9, 6,
    -- filter=184 channel=76
    -2, 5, 4, 2, -4, -4, 9, 6, -1,
    -- filter=184 channel=77
    3, 6, 8, 0, -3, 8, 1, -6, -1,
    -- filter=184 channel=78
    -4, 9, 10, -8, 0, 12, -8, -1, -1,
    -- filter=184 channel=79
    3, -13, -17, 8, -22, -27, 6, -17, -19,
    -- filter=184 channel=80
    -1, 3, -10, 12, 16, -5, 11, 9, -9,
    -- filter=184 channel=81
    -7, 0, -6, -6, 3, 1, -3, -5, -1,
    -- filter=184 channel=82
    -4, 2, 1, -2, 3, -2, 6, -4, 0,
    -- filter=184 channel=83
    4, 5, -3, 3, 8, -5, -6, -2, 6,
    -- filter=184 channel=84
    -3, -3, -4, 2, -3, -11, 0, -12, -9,
    -- filter=184 channel=85
    -1, 0, 2, 5, 5, -4, 1, 4, -6,
    -- filter=184 channel=86
    -1, -1, 3, -6, -8, -6, 4, 0, 0,
    -- filter=184 channel=87
    5, -9, 3, 8, -5, 2, -3, -5, -8,
    -- filter=184 channel=88
    -2, 5, 6, 1, 9, 6, 1, 8, -5,
    -- filter=184 channel=89
    -8, -12, -13, -2, -9, -17, 1, -3, -13,
    -- filter=184 channel=90
    -11, -3, 0, 1, 6, 0, 4, 3, 2,
    -- filter=184 channel=91
    9, -10, -17, 4, -9, -20, -4, -5, -4,
    -- filter=184 channel=92
    5, -1, 7, -3, -6, 0, 2, -1, -5,
    -- filter=184 channel=93
    -3, 4, -7, 9, 12, 10, 1, 14, 9,
    -- filter=184 channel=94
    0, 3, 5, -3, 3, 0, 0, 0, -5,
    -- filter=184 channel=95
    2, -2, 4, -7, -3, -8, 3, -1, 3,
    -- filter=184 channel=96
    3, 5, -4, 3, -5, -7, 8, 6, 6,
    -- filter=184 channel=97
    1, -6, -2, 1, 0, -5, 4, 6, 1,
    -- filter=184 channel=98
    -8, -13, -15, 8, -5, -11, 0, -7, -15,
    -- filter=184 channel=99
    -5, -20, -11, 4, -10, -6, -5, -5, -6,
    -- filter=184 channel=100
    -8, -8, -6, -2, -8, -4, -4, -7, -3,
    -- filter=184 channel=101
    8, -10, -9, -5, -1, 0, -7, -5, -6,
    -- filter=184 channel=102
    -4, -3, -5, 0, -3, 1, 4, -6, 0,
    -- filter=184 channel=103
    -5, 0, 6, 5, 18, 8, 6, 13, 12,
    -- filter=184 channel=104
    -10, -8, -12, 1, 3, -2, 0, 2, 0,
    -- filter=184 channel=105
    4, -8, -1, 5, 3, 0, -1, 4, -1,
    -- filter=184 channel=106
    -4, 2, -6, 0, 5, 5, 6, -1, 0,
    -- filter=184 channel=107
    8, -9, -8, 0, -9, -6, -5, -7, 0,
    -- filter=184 channel=108
    -2, 10, 0, -4, 1, 5, 4, 3, 12,
    -- filter=184 channel=109
    4, -21, -18, 5, -12, -16, 0, -12, -17,
    -- filter=184 channel=110
    1, -5, -4, -5, 2, -2, 2, -5, -8,
    -- filter=184 channel=111
    3, -1, 1, -5, 9, 3, 0, 5, 8,
    -- filter=184 channel=112
    -6, -13, -5, -2, -14, -14, -1, -14, -10,
    -- filter=184 channel=113
    0, -8, -10, -4, -10, -15, 4, -7, -12,
    -- filter=184 channel=114
    4, -6, -20, 11, -5, -17, 0, -13, -17,
    -- filter=184 channel=115
    3, 0, 5, -1, -4, 0, 0, -3, 1,
    -- filter=184 channel=116
    8, -6, -22, 7, -3, -8, 7, -4, -10,
    -- filter=184 channel=117
    6, 2, -8, 3, 5, -2, 1, 7, 2,
    -- filter=184 channel=118
    -3, -1, 3, 4, 0, -2, -3, -2, 7,
    -- filter=184 channel=119
    -1, -12, -7, -2, -4, -8, 5, -5, 2,
    -- filter=184 channel=120
    0, -17, -22, 2, -16, -25, 5, -19, -22,
    -- filter=184 channel=121
    0, 0, -5, -5, -5, -6, 9, -3, 1,
    -- filter=184 channel=122
    -14, 6, 7, 11, 29, 19, 3, 27, 18,
    -- filter=184 channel=123
    0, -4, -3, 4, 2, -9, -6, -3, -6,
    -- filter=184 channel=124
    0, -6, -4, 1, -7, -1, -3, -2, -6,
    -- filter=184 channel=125
    -10, -2, -18, 0, 2, -2, 6, -8, -13,
    -- filter=184 channel=126
    0, 0, -11, 3, 8, -10, 0, 0, -7,
    -- filter=184 channel=127
    -2, -1, 1, 2, -2, -1, 1, 4, -6,
    -- filter=185 channel=0
    -19, -12, 0, -15, -12, 7, -8, -6, 0,
    -- filter=185 channel=1
    -14, -9, -4, -10, -13, 8, 2, -1, 4,
    -- filter=185 channel=2
    -6, 8, -3, -3, -3, -6, -5, 0, 0,
    -- filter=185 channel=3
    0, 0, 1, -11, -2, -4, 0, 2, -7,
    -- filter=185 channel=4
    3, 0, 0, -3, -2, -2, 6, 1, 3,
    -- filter=185 channel=5
    -5, 4, -4, -1, -1, 7, -7, 0, 5,
    -- filter=185 channel=6
    0, 1, -8, 0, -9, -2, 3, 6, 8,
    -- filter=185 channel=7
    3, 4, 3, 0, 3, -2, -6, -5, 2,
    -- filter=185 channel=8
    -3, 7, 0, -1, 4, 0, -4, 3, -3,
    -- filter=185 channel=9
    -2, 1, -2, 7, 2, -2, -2, -2, 5,
    -- filter=185 channel=10
    -1, -1, -1, 3, -4, -1, 4, -2, 4,
    -- filter=185 channel=11
    0, -3, 0, 4, 2, 3, -1, 9, 2,
    -- filter=185 channel=12
    -6, 1, 7, -11, -6, 2, 0, 6, -5,
    -- filter=185 channel=13
    -7, -14, -6, -9, -1, 2, -1, -4, 5,
    -- filter=185 channel=14
    5, -7, -1, -2, -3, 3, 0, -1, 2,
    -- filter=185 channel=15
    -2, -16, 0, -4, -11, 4, 3, 1, 10,
    -- filter=185 channel=16
    -3, -6, 4, 4, 1, 8, 0, 1, -3,
    -- filter=185 channel=17
    6, 2, -3, -5, -7, 7, 2, -4, -4,
    -- filter=185 channel=18
    -10, -24, 8, -5, -8, 8, 5, 0, 9,
    -- filter=185 channel=19
    5, -6, 3, 5, 4, 1, -2, -3, 5,
    -- filter=185 channel=20
    3, -16, -11, -2, -7, 0, 6, 1, 7,
    -- filter=185 channel=21
    -4, 7, 2, -2, 8, 3, -3, -8, -12,
    -- filter=185 channel=22
    -5, -10, 2, -10, -6, 6, -1, -1, 10,
    -- filter=185 channel=23
    -9, -12, 1, -9, -4, 5, -4, 7, 14,
    -- filter=185 channel=24
    7, -5, -1, 4, 0, 1, 5, -1, -5,
    -- filter=185 channel=25
    -10, -9, 3, 6, -1, 14, 10, -1, -3,
    -- filter=185 channel=26
    -6, 10, 0, 5, 0, 0, 5, 3, -2,
    -- filter=185 channel=27
    -24, -2, 15, 1, -1, 20, 4, 2, 14,
    -- filter=185 channel=28
    -2, 5, 4, -3, -3, -2, 3, 0, 0,
    -- filter=185 channel=29
    -8, -11, 0, -2, -10, -12, 0, -4, 1,
    -- filter=185 channel=30
    -8, 2, 10, -2, -3, 0, -1, -9, 2,
    -- filter=185 channel=31
    -1, 13, 8, 7, 20, 7, 1, -9, -10,
    -- filter=185 channel=32
    -17, -9, 1, -3, -6, 7, 10, 4, 1,
    -- filter=185 channel=33
    -13, -18, 10, -9, -8, 14, 4, 5, 0,
    -- filter=185 channel=34
    -13, -1, 0, -8, -10, 4, -6, -6, 16,
    -- filter=185 channel=35
    -3, 1, -3, 3, 0, 2, -6, 6, -5,
    -- filter=185 channel=36
    -3, 3, 1, 8, 10, -6, -1, 3, -2,
    -- filter=185 channel=37
    -3, 8, 3, -11, -1, 4, 2, -4, 3,
    -- filter=185 channel=38
    -4, -7, -4, 0, -4, -2, 0, -2, 7,
    -- filter=185 channel=39
    -1, -7, 1, 5, -4, -8, 0, 0, 1,
    -- filter=185 channel=40
    -4, -1, -5, -6, -1, -5, -4, 0, 2,
    -- filter=185 channel=41
    -4, -14, -1, -8, -22, 0, 0, 0, -1,
    -- filter=185 channel=42
    -9, -5, -2, 1, 6, -3, -4, 5, -7,
    -- filter=185 channel=43
    -12, -6, -7, -8, -13, -2, 1, 3, 3,
    -- filter=185 channel=44
    -13, 2, 10, -6, -1, 0, 0, 3, -2,
    -- filter=185 channel=45
    2, -1, 1, 0, 4, -2, 3, -3, -7,
    -- filter=185 channel=46
    -8, 2, -5, 0, -7, 7, 7, 2, 5,
    -- filter=185 channel=47
    -7, 3, 1, -1, 0, 7, 0, -8, -13,
    -- filter=185 channel=48
    -2, 7, 2, 6, 5, 11, -1, 3, 7,
    -- filter=185 channel=49
    -4, -2, -2, 1, -6, 0, 1, 0, 7,
    -- filter=185 channel=50
    -8, 1, -2, 0, -1, 0, 3, 5, 2,
    -- filter=185 channel=51
    1, 0, 5, 5, 5, 0, 5, 4, -4,
    -- filter=185 channel=52
    -10, -1, -5, 2, 0, 3, -5, 6, 1,
    -- filter=185 channel=53
    -1, -4, 2, 1, 0, 3, -1, -1, -5,
    -- filter=185 channel=54
    2, 6, 3, 1, -4, 6, 3, -3, -1,
    -- filter=185 channel=55
    -13, -20, 3, -3, -7, -5, 5, -1, 11,
    -- filter=185 channel=56
    -7, 6, 9, -1, 4, 4, -7, -7, 1,
    -- filter=185 channel=57
    -8, -10, 3, 2, -6, 0, -6, -5, 0,
    -- filter=185 channel=58
    -9, -4, -2, -5, 4, 3, -8, 0, 0,
    -- filter=185 channel=59
    -1, -14, 8, -1, 5, 6, 3, -1, 6,
    -- filter=185 channel=60
    1, 1, 6, 2, 6, 2, -1, 0, -1,
    -- filter=185 channel=61
    0, 0, 1, -5, 0, 2, -6, 0, 6,
    -- filter=185 channel=62
    1, -6, -5, 5, -7, 4, 5, 6, -3,
    -- filter=185 channel=63
    0, -3, -6, 4, 7, 0, -4, -3, -6,
    -- filter=185 channel=64
    1, 1, 5, -1, 4, 2, -5, 1, -7,
    -- filter=185 channel=65
    6, -5, -4, -1, -7, 2, -5, -2, -3,
    -- filter=185 channel=66
    2, -17, -2, -2, -13, 6, 2, -5, 3,
    -- filter=185 channel=67
    1, 0, -7, -7, 0, 1, 1, -3, 4,
    -- filter=185 channel=68
    6, 6, -2, 0, -3, 1, -5, -2, -8,
    -- filter=185 channel=69
    -6, -10, -2, -8, -8, 6, -5, 5, 2,
    -- filter=185 channel=70
    -13, -2, 12, -3, 2, 12, 4, 5, 17,
    -- filter=185 channel=71
    2, 1, -4, -8, -3, 1, -8, 3, -5,
    -- filter=185 channel=72
    -1, -3, 3, 5, 1, 8, -3, 4, -7,
    -- filter=185 channel=73
    -13, -5, 3, -5, 2, 4, 7, 9, 12,
    -- filter=185 channel=74
    -8, 2, 14, -6, 10, 1, 4, 3, 8,
    -- filter=185 channel=75
    -9, -14, 1, -13, -16, 4, -12, -7, -5,
    -- filter=185 channel=76
    5, -7, 1, -9, -7, -6, 11, -4, 4,
    -- filter=185 channel=77
    2, 3, -2, 3, -5, -1, -5, 0, 2,
    -- filter=185 channel=78
    -6, 6, 4, 2, 1, 3, 0, 2, 0,
    -- filter=185 channel=79
    -19, -30, 11, -14, -8, 1, 15, -3, 10,
    -- filter=185 channel=80
    -11, -2, 8, -1, 8, 8, 0, -5, -3,
    -- filter=185 channel=81
    4, 1, 3, 6, 6, 4, 4, 6, -1,
    -- filter=185 channel=82
    -4, 2, 3, 3, -1, 0, -7, -4, 2,
    -- filter=185 channel=83
    5, -1, -1, 4, 0, 7, -3, 4, 1,
    -- filter=185 channel=84
    -6, -9, -5, 0, 0, 1, 2, 1, 14,
    -- filter=185 channel=85
    3, 1, -1, -5, 1, 2, 0, -4, 4,
    -- filter=185 channel=86
    -5, 0, -4, 0, -8, 9, -4, 1, 2,
    -- filter=185 channel=87
    -2, -8, -4, -11, -11, -3, -5, -8, 9,
    -- filter=185 channel=88
    -2, 7, 7, 10, 12, -7, -7, -6, -6,
    -- filter=185 channel=89
    -12, -18, 9, -6, 4, 9, 9, 3, -5,
    -- filter=185 channel=90
    3, 6, 0, -8, 2, 1, 0, -3, 2,
    -- filter=185 channel=91
    -6, -9, 11, 0, -3, 10, 8, 3, 5,
    -- filter=185 channel=92
    0, -6, 6, -5, -8, 0, 6, -2, 10,
    -- filter=185 channel=93
    -3, 8, 7, 1, 8, 4, 3, -11, -7,
    -- filter=185 channel=94
    0, -7, -6, 0, 7, 7, 0, -5, -2,
    -- filter=185 channel=95
    3, 4, 1, -6, -3, -1, 3, 0, -1,
    -- filter=185 channel=96
    0, 0, -6, -3, 4, 1, -5, 5, 4,
    -- filter=185 channel=97
    2, 1, -1, 1, -9, 2, -6, -4, -7,
    -- filter=185 channel=98
    -10, -15, 11, 1, 2, 8, 5, -4, 3,
    -- filter=185 channel=99
    -3, 1, 11, -1, 5, -3, 1, 10, 4,
    -- filter=185 channel=100
    2, -1, 5, -4, 4, 0, -2, 6, 1,
    -- filter=185 channel=101
    -5, 5, -1, -2, 0, 0, 7, 1, -3,
    -- filter=185 channel=102
    -7, -6, -2, 6, -3, 0, -7, 0, 1,
    -- filter=185 channel=103
    0, -5, -1, -6, 0, -4, -4, -12, -6,
    -- filter=185 channel=104
    -6, 9, -3, 3, 10, 7, 1, 5, -3,
    -- filter=185 channel=105
    3, -7, -7, -7, 1, 2, 8, 6, -2,
    -- filter=185 channel=106
    4, -7, -4, -3, 4, 0, 7, -3, 0,
    -- filter=185 channel=107
    -3, -8, 0, -6, -1, -5, 0, -8, 5,
    -- filter=185 channel=108
    -7, -5, 2, -1, -1, 0, 0, -3, 0,
    -- filter=185 channel=109
    -16, -8, 15, 2, -4, 11, 9, 1, 17,
    -- filter=185 channel=110
    0, -6, 0, -3, -1, -6, 5, 2, -2,
    -- filter=185 channel=111
    2, 3, -9, -2, 0, -2, -2, 3, -1,
    -- filter=185 channel=112
    -5, 6, 11, 0, 0, 5, -4, -1, 8,
    -- filter=185 channel=113
    -9, -6, -5, -3, 0, 6, 3, -4, -4,
    -- filter=185 channel=114
    -22, -14, 2, -9, -12, 7, 9, 7, 17,
    -- filter=185 channel=115
    4, 0, -7, -2, -6, 3, 4, 3, -3,
    -- filter=185 channel=116
    -6, -4, 0, 10, -2, -3, 13, 6, -1,
    -- filter=185 channel=117
    -3, 2, 4, 0, 5, 0, -3, -2, -10,
    -- filter=185 channel=118
    0, 1, -3, 1, -6, -6, -6, 3, -4,
    -- filter=185 channel=119
    -9, 5, 9, -2, -4, 9, 1, -1, 10,
    -- filter=185 channel=120
    -23, 6, 11, -4, 4, 15, 1, 7, 14,
    -- filter=185 channel=121
    5, -2, -3, -7, 0, 1, 0, 7, 6,
    -- filter=185 channel=122
    -5, 15, 5, -1, 6, 11, -12, -11, -14,
    -- filter=185 channel=123
    -6, -2, -6, -1, 5, 6, 0, -4, 5,
    -- filter=185 channel=124
    4, -9, -5, -7, 1, 0, 3, 5, 1,
    -- filter=185 channel=125
    0, 6, 5, 0, 12, 0, 2, 2, 5,
    -- filter=185 channel=126
    -4, -8, -8, -4, -13, -4, 5, 3, -1,
    -- filter=185 channel=127
    -1, 0, 1, 4, -3, -5, 6, -7, 5,
    -- filter=186 channel=0
    -4, -4, -2, 3, 3, 9, 8, 4, -1,
    -- filter=186 channel=1
    -4, 0, 0, 7, 5, -6, -4, 1, 0,
    -- filter=186 channel=2
    -4, 1, -3, 6, 1, 5, -6, -6, 5,
    -- filter=186 channel=3
    5, 0, -5, 2, 7, 3, 5, 2, -6,
    -- filter=186 channel=4
    8, -4, 1, -3, 0, -5, 3, 2, 6,
    -- filter=186 channel=5
    -7, 4, 0, -4, -1, -3, 4, -2, -5,
    -- filter=186 channel=6
    -7, -3, 0, -4, -3, 4, 8, 0, -2,
    -- filter=186 channel=7
    2, 3, 3, -7, 3, 0, 4, 3, -7,
    -- filter=186 channel=8
    0, 2, 6, -1, -4, -7, 3, 3, 3,
    -- filter=186 channel=9
    -5, 0, -4, -8, -2, 3, -8, 4, -7,
    -- filter=186 channel=10
    1, 1, 0, 7, -1, -6, 0, -3, -3,
    -- filter=186 channel=11
    5, -7, 2, -5, 7, 1, -4, -4, -5,
    -- filter=186 channel=12
    0, 0, 0, -3, 0, 0, 3, -4, -6,
    -- filter=186 channel=13
    8, -3, 3, -3, -7, -2, 4, -8, 0,
    -- filter=186 channel=14
    1, 0, -6, 6, -3, -6, 2, 1, 0,
    -- filter=186 channel=15
    -2, 2, 3, -4, -2, -7, 2, 1, 2,
    -- filter=186 channel=16
    -5, 7, 4, -4, -1, 0, 4, -3, -4,
    -- filter=186 channel=17
    1, 6, -1, 1, -3, -6, 3, 2, 4,
    -- filter=186 channel=18
    -4, -2, 2, 4, 0, -4, -2, 2, 4,
    -- filter=186 channel=19
    -7, -4, -3, -5, 5, -6, -3, 0, 5,
    -- filter=186 channel=20
    -2, 1, -4, 0, -4, 0, 1, 2, 2,
    -- filter=186 channel=21
    2, 9, -5, -3, -4, 0, -2, 1, -3,
    -- filter=186 channel=22
    -4, 2, -7, 2, 1, 0, -3, 2, 3,
    -- filter=186 channel=23
    -5, -7, 5, -8, 6, -2, -4, 2, 5,
    -- filter=186 channel=24
    -2, 3, -5, -1, -1, 6, 1, -2, -4,
    -- filter=186 channel=25
    9, -5, -7, 4, 3, -7, 4, -5, -8,
    -- filter=186 channel=26
    -2, -3, 4, 2, -1, 3, 1, -3, -1,
    -- filter=186 channel=27
    4, -7, -3, -4, -11, -3, 2, -2, 4,
    -- filter=186 channel=28
    2, -1, 6, -2, 6, -6, -2, 6, -7,
    -- filter=186 channel=29
    0, -6, 4, -5, 6, 3, 2, 7, -5,
    -- filter=186 channel=30
    3, -2, -3, 5, 3, -3, 0, -1, -3,
    -- filter=186 channel=31
    8, -4, 9, 2, 2, 3, 1, -3, -4,
    -- filter=186 channel=32
    5, 3, -4, -4, -7, -7, 0, -5, -6,
    -- filter=186 channel=33
    3, 7, 6, 2, 0, 1, 4, -9, -3,
    -- filter=186 channel=34
    -2, 0, -1, -3, 4, -3, -2, -6, -4,
    -- filter=186 channel=35
    2, 4, 0, 0, 6, 3, -3, -4, -1,
    -- filter=186 channel=36
    1, 4, -6, -4, 6, -5, 2, -3, -5,
    -- filter=186 channel=37
    -1, 4, 8, 6, 3, 3, 0, 7, 1,
    -- filter=186 channel=38
    2, -2, -7, 7, -4, 3, 5, -6, -4,
    -- filter=186 channel=39
    5, 1, -2, 5, 2, -6, 3, 0, 4,
    -- filter=186 channel=40
    -1, 0, -3, 5, 1, 1, 2, 5, -2,
    -- filter=186 channel=41
    -5, 0, -5, 0, 1, -7, -1, 3, -6,
    -- filter=186 channel=42
    -1, 6, 6, 5, -3, 6, 0, 1, 3,
    -- filter=186 channel=43
    0, 1, -7, -5, 1, -1, 7, -3, 0,
    -- filter=186 channel=44
    4, 0, -5, 1, 3, -2, -4, -1, 5,
    -- filter=186 channel=45
    -4, 0, 3, 4, 0, -2, 4, 8, 2,
    -- filter=186 channel=46
    -1, -4, 2, -2, 6, -1, -5, -6, -6,
    -- filter=186 channel=47
    4, 0, 4, -2, 1, 0, -4, 2, 1,
    -- filter=186 channel=48
    6, 7, 0, -2, 0, 0, -2, 0, -2,
    -- filter=186 channel=49
    0, -4, 4, 1, 6, -5, 5, 5, 1,
    -- filter=186 channel=50
    5, 0, -3, 5, 0, -5, -8, -1, -6,
    -- filter=186 channel=51
    6, -7, 4, 5, -2, 2, -3, 0, -6,
    -- filter=186 channel=52
    6, 5, 1, 0, -5, 1, 2, 0, 6,
    -- filter=186 channel=53
    1, 0, -6, -2, 5, 2, 5, 6, -5,
    -- filter=186 channel=54
    1, 7, 5, -1, 1, 4, 3, 0, 0,
    -- filter=186 channel=55
    -4, -6, 4, -3, 1, 5, 5, 1, -6,
    -- filter=186 channel=56
    -7, 2, -2, -7, 4, 0, 2, 0, -5,
    -- filter=186 channel=57
    5, 4, 5, 5, -1, 3, 3, -5, 6,
    -- filter=186 channel=58
    -6, 0, 5, 6, 3, 7, -6, 1, 5,
    -- filter=186 channel=59
    6, -6, -3, 4, -8, -5, -7, -6, 3,
    -- filter=186 channel=60
    5, 0, -1, -3, 0, 6, 7, 0, 0,
    -- filter=186 channel=61
    3, -1, 4, -7, -2, 3, 4, 0, -5,
    -- filter=186 channel=62
    6, 0, -1, 3, 4, 2, 0, 0, 4,
    -- filter=186 channel=63
    0, -3, -3, 2, -2, -4, 5, 5, -3,
    -- filter=186 channel=64
    2, -2, 3, 4, -7, -4, 3, 3, 1,
    -- filter=186 channel=65
    5, 5, -1, 7, -4, 6, 5, 5, -2,
    -- filter=186 channel=66
    5, -7, -4, 10, -7, -2, 5, -1, 0,
    -- filter=186 channel=67
    -3, -6, 4, 3, 4, -6, 3, 4, 5,
    -- filter=186 channel=68
    7, -3, 7, -5, -1, 0, 3, -4, -7,
    -- filter=186 channel=69
    -2, 4, 3, 5, -2, 2, 6, 6, 0,
    -- filter=186 channel=70
    7, -8, 1, -4, -6, 0, -2, -3, 0,
    -- filter=186 channel=71
    7, 2, 3, 7, 3, 0, -4, -6, -4,
    -- filter=186 channel=72
    -1, -4, 0, -6, -8, -5, 0, -1, 5,
    -- filter=186 channel=73
    0, -3, 1, -3, -4, 2, 6, -1, 0,
    -- filter=186 channel=74
    7, 2, 4, 1, -4, -7, -3, 0, -1,
    -- filter=186 channel=75
    -7, -4, 1, 6, 5, 1, 1, 6, 4,
    -- filter=186 channel=76
    -6, 0, 0, -4, 6, -4, 0, 7, -5,
    -- filter=186 channel=77
    4, -5, -4, -4, 6, 3, 5, 2, -6,
    -- filter=186 channel=78
    3, 2, -6, 4, 4, 6, 1, -3, -7,
    -- filter=186 channel=79
    -3, 4, -7, -5, -5, -1, 2, -4, 5,
    -- filter=186 channel=80
    3, -3, 1, 5, -2, -8, -4, -11, -2,
    -- filter=186 channel=81
    0, 7, 5, -4, -3, 1, -5, -4, 1,
    -- filter=186 channel=82
    3, 5, -6, -2, -2, 2, -3, 0, -5,
    -- filter=186 channel=83
    -1, 0, -5, -4, -5, -3, -8, -8, -4,
    -- filter=186 channel=84
    -3, -2, 0, 2, -3, 3, 6, -5, 3,
    -- filter=186 channel=85
    -6, -4, 6, -3, 4, 6, 2, -1, 6,
    -- filter=186 channel=86
    -3, 0, -1, 3, 0, 2, 0, 5, -2,
    -- filter=186 channel=87
    6, 1, -6, -6, 5, 5, -6, -6, -6,
    -- filter=186 channel=88
    0, -5, -4, 3, 2, -6, -6, 4, -6,
    -- filter=186 channel=89
    3, 3, 3, 0, -8, 3, 0, -10, -5,
    -- filter=186 channel=90
    -4, -3, 3, -5, 0, 0, -3, -6, -5,
    -- filter=186 channel=91
    0, -1, 0, 2, 0, -1, -1, -1, -6,
    -- filter=186 channel=92
    -4, 3, 2, 2, 4, -6, 0, -4, 6,
    -- filter=186 channel=93
    5, 5, -6, -5, 3, -6, -4, 4, -7,
    -- filter=186 channel=94
    6, -6, 5, -3, 6, 2, 5, 3, 3,
    -- filter=186 channel=95
    1, 4, 0, 1, -1, 7, 1, 1, 3,
    -- filter=186 channel=96
    -3, -1, 2, 3, 2, -7, 0, 5, -4,
    -- filter=186 channel=97
    1, -2, 0, 5, 8, 1, 2, -6, 3,
    -- filter=186 channel=98
    6, -4, -3, -4, -7, -5, -2, -3, -3,
    -- filter=186 channel=99
    0, -7, -5, -1, -1, -3, -2, -3, 3,
    -- filter=186 channel=100
    3, 5, 6, -7, 2, -3, -4, 0, 0,
    -- filter=186 channel=101
    4, 4, 1, 0, 3, -2, -2, 7, 1,
    -- filter=186 channel=102
    0, 0, 0, 4, -4, -4, 2, -5, -5,
    -- filter=186 channel=103
    -1, 3, 5, 0, 3, 8, -6, -7, -1,
    -- filter=186 channel=104
    -2, -5, 0, -1, -6, -5, 0, 4, -1,
    -- filter=186 channel=105
    1, -4, -3, -3, -4, -2, 5, 1, 6,
    -- filter=186 channel=106
    0, 6, -3, -5, 1, -1, 8, 5, -1,
    -- filter=186 channel=107
    0, 4, -5, -6, 1, -4, 1, -3, 6,
    -- filter=186 channel=108
    -1, 0, 1, -2, 1, 4, 2, -2, 5,
    -- filter=186 channel=109
    5, 0, 0, -6, -8, -6, -4, -11, -8,
    -- filter=186 channel=110
    6, 6, 3, 0, 5, 0, 5, 4, 0,
    -- filter=186 channel=111
    2, 4, -1, 2, 1, -3, 0, 0, -1,
    -- filter=186 channel=112
    -1, -2, 0, 5, 0, 0, -2, 4, -4,
    -- filter=186 channel=113
    8, 3, -2, -4, 5, 0, -5, -6, -6,
    -- filter=186 channel=114
    4, -8, 3, 7, -8, 0, -2, 6, 7,
    -- filter=186 channel=115
    -4, 4, -4, -4, 2, -4, 6, 2, -2,
    -- filter=186 channel=116
    8, -6, -5, 1, 2, -2, -5, 4, 5,
    -- filter=186 channel=117
    2, 6, 0, -2, 2, 6, 6, -5, 0,
    -- filter=186 channel=118
    -5, -6, -6, -6, -6, 1, -6, 1, 2,
    -- filter=186 channel=119
    -4, -8, -6, 1, -1, -6, -3, -3, 4,
    -- filter=186 channel=120
    -2, 2, -1, -9, 0, -5, -7, -9, -6,
    -- filter=186 channel=121
    0, 5, 1, 1, -2, -3, 3, -6, 1,
    -- filter=186 channel=122
    8, 3, 3, -5, -5, -5, 0, -3, 1,
    -- filter=186 channel=123
    5, -5, -5, 6, 2, -2, -5, 5, 0,
    -- filter=186 channel=124
    -4, -1, 1, 7, -5, 7, -6, 7, -5,
    -- filter=186 channel=125
    -1, -7, 5, -5, 2, -8, 0, -3, 5,
    -- filter=186 channel=126
    3, 8, -5, 4, -7, 0, 0, -8, 0,
    -- filter=186 channel=127
    -6, 0, 2, 7, 2, -5, -3, 2, -5,
    -- filter=187 channel=0
    5, 17, 3, 7, 22, 12, 10, 14, 9,
    -- filter=187 channel=1
    13, 18, -3, 3, 20, 6, 9, 12, -4,
    -- filter=187 channel=2
    -1, -2, 2, 8, 2, 7, -4, -4, 6,
    -- filter=187 channel=3
    1, -4, 6, -2, -2, -2, 8, 8, 8,
    -- filter=187 channel=4
    -3, -3, 6, 9, 10, -3, 0, 0, -1,
    -- filter=187 channel=5
    3, 1, -3, 8, 9, -5, 6, 6, -7,
    -- filter=187 channel=6
    -1, 7, 5, -4, 7, 2, -4, 1, 10,
    -- filter=187 channel=7
    0, -1, 0, 4, -6, 2, 0, -1, -3,
    -- filter=187 channel=8
    0, 6, -7, 8, -1, -7, 3, 0, -6,
    -- filter=187 channel=9
    4, 3, 0, 6, -8, -11, -4, 0, -4,
    -- filter=187 channel=10
    4, -7, 3, 0, 0, 0, 3, 3, -5,
    -- filter=187 channel=11
    -10, -3, 0, -7, 4, -3, -6, 7, 13,
    -- filter=187 channel=12
    -1, -3, -2, 4, 6, -1, 4, 7, -1,
    -- filter=187 channel=13
    0, -8, -3, 1, -4, 4, 0, 6, 6,
    -- filter=187 channel=14
    0, 6, 6, -3, -6, -6, 4, 3, -3,
    -- filter=187 channel=15
    -11, -1, -8, 1, -2, -7, 1, 6, 3,
    -- filter=187 channel=16
    7, -8, 0, 5, 0, -9, 0, -8, -7,
    -- filter=187 channel=17
    0, 6, 6, 5, -6, -1, -4, 3, -4,
    -- filter=187 channel=18
    -6, -1, 0, 5, 0, -5, 1, -1, -2,
    -- filter=187 channel=19
    -1, 7, 4, 4, 7, -5, -1, 0, -5,
    -- filter=187 channel=20
    3, 2, -2, -1, 10, 8, 6, 6, 22,
    -- filter=187 channel=21
    -4, -5, -2, 1, -3, -1, -9, -10, -9,
    -- filter=187 channel=22
    2, 0, -4, 8, 9, 0, 8, 5, 6,
    -- filter=187 channel=23
    -2, -3, -12, -9, -13, -16, -1, -3, 0,
    -- filter=187 channel=24
    -1, 6, 1, 6, 0, -4, 4, 0, 7,
    -- filter=187 channel=25
    -6, -1, 1, -2, -5, -11, -1, -6, -14,
    -- filter=187 channel=26
    7, -1, 4, 2, 5, 2, 4, 6, 0,
    -- filter=187 channel=27
    -1, -6, -14, 1, -10, -13, 3, -6, -7,
    -- filter=187 channel=28
    1, -6, 4, 0, -6, 4, -3, -2, 3,
    -- filter=187 channel=29
    0, 3, 2, -2, 5, 6, -2, 0, 12,
    -- filter=187 channel=30
    3, 3, -7, -2, 4, -5, 8, 2, -8,
    -- filter=187 channel=31
    3, -4, -6, -1, -16, -9, -3, -7, -13,
    -- filter=187 channel=32
    -6, 1, -6, 7, -1, 0, 3, 7, 2,
    -- filter=187 channel=33
    -5, 0, -4, 2, -8, -5, 2, 0, 0,
    -- filter=187 channel=34
    8, 3, -3, 10, -6, -2, 11, 4, 3,
    -- filter=187 channel=35
    -3, -5, -6, 4, -3, -4, 6, 7, 6,
    -- filter=187 channel=36
    0, 6, 0, -2, 4, 10, -5, -3, 2,
    -- filter=187 channel=37
    7, 15, 1, 3, 11, 1, 2, 7, -4,
    -- filter=187 channel=38
    -1, -9, 0, -4, 0, -10, -5, -8, -2,
    -- filter=187 channel=39
    2, -3, 0, -1, -3, -2, 5, 6, 7,
    -- filter=187 channel=40
    6, -2, 0, -4, 5, 5, -5, 0, 5,
    -- filter=187 channel=41
    0, 5, -4, 1, 10, 1, -2, 0, 5,
    -- filter=187 channel=42
    -8, 2, 1, -6, 1, -1, -1, -4, 2,
    -- filter=187 channel=43
    3, 0, 2, -3, 0, 3, -1, 10, 3,
    -- filter=187 channel=44
    -4, 2, 2, -2, 2, -6, 4, 0, -14,
    -- filter=187 channel=45
    4, 7, -3, -5, 2, -4, 3, -3, -5,
    -- filter=187 channel=46
    1, -1, -5, -5, 5, -4, -2, 8, 2,
    -- filter=187 channel=47
    0, 3, 2, -1, -3, -14, -6, -2, -10,
    -- filter=187 channel=48
    1, -4, -12, -4, -3, -9, 2, -2, -11,
    -- filter=187 channel=49
    -3, -7, -4, -4, 4, -9, 0, -2, -4,
    -- filter=187 channel=50
    -10, 0, -6, -11, -2, -14, 3, -10, -15,
    -- filter=187 channel=51
    6, 4, -2, 0, -5, 0, 3, 6, -6,
    -- filter=187 channel=52
    5, 4, 2, 0, -4, 2, 9, -3, 5,
    -- filter=187 channel=53
    -8, -2, -6, -5, 4, 0, 6, 0, 8,
    -- filter=187 channel=54
    -4, -6, -4, 0, 4, -4, -3, -3, -4,
    -- filter=187 channel=55
    -4, -7, 0, 4, -3, -7, 1, 3, -1,
    -- filter=187 channel=56
    4, -4, -3, 3, -3, -1, 7, 1, -5,
    -- filter=187 channel=57
    5, -8, -1, 1, 2, 0, 3, -3, -2,
    -- filter=187 channel=58
    -1, 12, 7, 10, 14, -1, 7, 6, 7,
    -- filter=187 channel=59
    -3, -5, 0, -2, -1, -5, -9, -13, -9,
    -- filter=187 channel=60
    8, 4, 0, -3, -2, 7, -5, 6, -4,
    -- filter=187 channel=61
    6, -4, 1, -2, 0, 6, -3, -4, -2,
    -- filter=187 channel=62
    3, 2, -1, -4, -5, 6, 6, 6, 2,
    -- filter=187 channel=63
    7, 1, -1, 7, 7, 2, 9, 0, 1,
    -- filter=187 channel=64
    -5, 7, -3, 6, -3, 5, 0, 5, 8,
    -- filter=187 channel=65
    -3, 1, 6, -4, 4, -5, 0, 2, 4,
    -- filter=187 channel=66
    -1, -7, -4, 6, -3, 2, -7, 7, -2,
    -- filter=187 channel=67
    2, -4, -3, 1, 8, -3, -4, -5, 5,
    -- filter=187 channel=68
    -3, 5, 5, 7, -4, -4, 0, 2, 3,
    -- filter=187 channel=69
    5, 1, 6, 1, 5, -3, -7, -3, -4,
    -- filter=187 channel=70
    -8, -3, -4, 5, 0, -9, -3, 1, -14,
    -- filter=187 channel=71
    -1, 0, -3, -6, -4, -6, 6, 0, -4,
    -- filter=187 channel=72
    -10, -5, -6, -5, -14, 1, 0, -12, 1,
    -- filter=187 channel=73
    -6, 1, 2, -1, 0, -3, 1, -1, 1,
    -- filter=187 channel=74
    6, 0, -10, -1, -3, -12, -4, -13, -11,
    -- filter=187 channel=75
    5, 10, 5, -4, 6, 4, 1, 13, -3,
    -- filter=187 channel=76
    -3, 2, 1, 5, 9, 12, 6, 6, 19,
    -- filter=187 channel=77
    5, 3, 7, 1, -6, 0, 3, -4, 6,
    -- filter=187 channel=78
    -7, 2, 0, -5, 0, -7, 2, 0, 0,
    -- filter=187 channel=79
    -7, 0, -8, 5, 4, -1, -2, 10, 5,
    -- filter=187 channel=80
    -12, -2, -7, 1, -7, -13, -6, -15, -13,
    -- filter=187 channel=81
    -1, -5, -3, -3, -2, 0, 5, 3, -3,
    -- filter=187 channel=82
    -3, -3, 3, 5, 0, 1, 6, 5, -2,
    -- filter=187 channel=83
    6, 0, -2, 1, -7, -7, 0, -4, 2,
    -- filter=187 channel=84
    1, 3, 0, 7, -1, 1, -3, -3, -2,
    -- filter=187 channel=85
    5, 2, 2, 4, -7, -3, -1, 4, -6,
    -- filter=187 channel=86
    4, 9, -3, 13, -2, -4, 3, 4, -4,
    -- filter=187 channel=87
    4, -2, 7, 8, -3, 0, -1, 10, 8,
    -- filter=187 channel=88
    11, 0, 1, 5, -6, 0, 10, 5, -4,
    -- filter=187 channel=89
    -7, -8, 0, -7, -4, 0, -11, -8, 1,
    -- filter=187 channel=90
    8, 0, -1, 6, 0, 7, 2, 0, 3,
    -- filter=187 channel=91
    1, -6, -2, -1, -9, -10, 2, -12, -11,
    -- filter=187 channel=92
    -2, -1, -4, -2, 7, -1, -3, 6, 2,
    -- filter=187 channel=93
    0, 4, -4, -6, 0, -6, -7, -4, 0,
    -- filter=187 channel=94
    3, 4, 1, 5, 3, 1, 4, -3, -6,
    -- filter=187 channel=95
    0, 2, -1, -7, 1, -2, -1, -6, 0,
    -- filter=187 channel=96
    -4, 0, -1, 4, -4, 1, -7, -5, 4,
    -- filter=187 channel=97
    -3, -3, 7, 4, -2, 3, 4, 1, 6,
    -- filter=187 channel=98
    -9, -10, -2, -5, -5, -7, -3, -5, -13,
    -- filter=187 channel=99
    -5, 0, -6, 0, -1, -13, 0, -11, 3,
    -- filter=187 channel=100
    -3, 0, -2, 0, -1, 0, -6, 0, 5,
    -- filter=187 channel=101
    4, 0, 3, 2, -3, 9, 0, -4, 7,
    -- filter=187 channel=102
    -1, 0, 6, 0, 0, 0, -2, -7, -7,
    -- filter=187 channel=103
    -10, 0, -9, -1, 0, 0, -4, 0, -15,
    -- filter=187 channel=104
    -2, -9, 0, 0, 0, -5, 0, -9, -12,
    -- filter=187 channel=105
    -7, 0, -1, 7, 8, 6, 5, 6, 14,
    -- filter=187 channel=106
    -1, -5, 5, -2, 6, 8, -4, 6, -2,
    -- filter=187 channel=107
    -1, 0, -1, 9, 8, 9, 8, 0, 8,
    -- filter=187 channel=108
    7, -1, 0, 4, 13, 0, 5, 1, 9,
    -- filter=187 channel=109
    -7, -7, -15, 2, -7, -12, 0, -1, -13,
    -- filter=187 channel=110
    4, 1, 7, 2, -4, 7, 0, 3, -6,
    -- filter=187 channel=111
    5, 3, 0, 4, -5, -2, 6, -5, 8,
    -- filter=187 channel=112
    5, -3, -6, -4, -2, -7, 0, -5, -2,
    -- filter=187 channel=113
    3, -10, 2, -4, -10, -5, 0, -3, -10,
    -- filter=187 channel=114
    9, 11, -4, 2, 21, 1, 3, 12, 2,
    -- filter=187 channel=115
    1, -1, 5, 2, 5, -6, -2, -3, -4,
    -- filter=187 channel=116
    -7, -10, 1, 6, -4, -11, -8, -11, -6,
    -- filter=187 channel=117
    -3, 5, -5, -7, -5, -5, 4, 2, -6,
    -- filter=187 channel=118
    -5, 5, -1, 0, 5, 7, 6, 5, -6,
    -- filter=187 channel=119
    -5, 1, -1, 6, -4, -10, 5, -8, -6,
    -- filter=187 channel=120
    -2, -5, -7, -3, -17, -14, 0, -11, -6,
    -- filter=187 channel=121
    -2, -9, 2, 1, -9, -3, 0, -5, 2,
    -- filter=187 channel=122
    -2, -4, -12, 5, -13, -7, 1, -14, -19,
    -- filter=187 channel=123
    -7, 0, 0, 5, 0, -5, -3, -4, -1,
    -- filter=187 channel=124
    6, -5, 5, 4, 2, -2, 6, 2, 6,
    -- filter=187 channel=125
    -7, -10, -7, 3, -5, -2, -2, -8, -10,
    -- filter=187 channel=126
    2, 5, -4, 3, 7, 1, 0, -1, -1,
    -- filter=187 channel=127
    4, 0, 0, -5, 5, 4, -2, 1, -2,
    -- filter=188 channel=0
    -3, 13, -16, -12, 9, -9, 0, 6, -12,
    -- filter=188 channel=1
    6, 15, -1, -2, 12, -10, 2, 3, 0,
    -- filter=188 channel=2
    -1, 8, 0, -1, -11, -6, 0, 0, 8,
    -- filter=188 channel=3
    -16, -12, -11, -10, -16, -18, -14, -18, -11,
    -- filter=188 channel=4
    -17, -15, -12, -11, -13, 6, -16, -16, 0,
    -- filter=188 channel=5
    -1, 13, -7, -7, 11, -21, 3, 2, -8,
    -- filter=188 channel=6
    1, 1, 5, -1, 1, -1, -1, 4, 1,
    -- filter=188 channel=7
    -5, -7, -5, -6, -1, 7, -5, -3, 5,
    -- filter=188 channel=8
    -6, 15, 8, -6, 8, 13, 2, 4, 9,
    -- filter=188 channel=9
    -10, 3, -5, 3, 0, -3, 2, 2, 3,
    -- filter=188 channel=10
    0, 7, 5, 3, 9, -9, -2, 5, 0,
    -- filter=188 channel=11
    5, -5, -7, -6, -6, 0, -2, -4, 7,
    -- filter=188 channel=12
    9, 14, -3, 9, 18, -6, 13, 20, 7,
    -- filter=188 channel=13
    0, 9, -4, -1, 13, 1, 8, 8, 2,
    -- filter=188 channel=14
    -4, -6, -3, -6, 2, -7, 6, 4, 0,
    -- filter=188 channel=15
    -8, 1, -5, -4, -3, -2, -4, 0, 0,
    -- filter=188 channel=16
    -2, 14, -1, 6, 15, -15, -6, 7, -2,
    -- filter=188 channel=17
    7, 2, 4, 6, -3, 4, 5, -7, -6,
    -- filter=188 channel=18
    0, 1, -7, 2, 0, 0, 5, -4, 4,
    -- filter=188 channel=19
    4, -6, -2, -8, 0, 2, -7, -7, 1,
    -- filter=188 channel=20
    6, -6, -12, -3, 1, -9, -1, -11, 0,
    -- filter=188 channel=21
    0, 10, -8, 5, 14, -13, -5, 9, 0,
    -- filter=188 channel=22
    -3, 13, 3, -2, 6, 3, -4, -2, 3,
    -- filter=188 channel=23
    -12, 8, -12, -16, 22, -14, -2, -8, 8,
    -- filter=188 channel=24
    1, -2, -7, -1, 3, 3, 5, -4, 7,
    -- filter=188 channel=25
    3, 16, -9, 4, 27, -26, 0, 8, -7,
    -- filter=188 channel=26
    8, 0, 0, 1, 0, -2, -5, 5, 2,
    -- filter=188 channel=27
    -11, 18, -9, -5, 24, -18, -3, -3, 9,
    -- filter=188 channel=28
    6, 0, 7, 6, 6, 0, -6, 0, -6,
    -- filter=188 channel=29
    5, -8, -10, 6, -8, -5, 0, -16, 7,
    -- filter=188 channel=30
    -1, 9, -17, -3, 5, -6, 2, -3, -5,
    -- filter=188 channel=31
    -11, 15, -16, -17, 21, -31, -1, 12, 0,
    -- filter=188 channel=32
    0, 6, -3, -5, 22, -14, 11, 3, -4,
    -- filter=188 channel=33
    1, 6, -9, 2, 16, -15, 7, 5, -5,
    -- filter=188 channel=34
    1, 39, 11, 7, 35, 26, -6, 25, 22,
    -- filter=188 channel=35
    0, -5, -2, -5, 3, -4, -6, -6, -6,
    -- filter=188 channel=36
    0, 1, 0, 6, 0, -4, 4, 13, 1,
    -- filter=188 channel=37
    -3, 25, -7, 0, 23, -12, -4, 2, -1,
    -- filter=188 channel=38
    -4, 6, -14, -5, 8, -16, 4, 2, 0,
    -- filter=188 channel=39
    -1, -1, -9, 4, -14, 2, -5, 0, 3,
    -- filter=188 channel=40
    1, 0, 4, -6, 0, -3, -2, -6, 2,
    -- filter=188 channel=41
    20, -7, 30, 15, 1, 37, -6, 9, 14,
    -- filter=188 channel=42
    0, -9, 0, 0, -4, -3, -6, -10, 2,
    -- filter=188 channel=43
    -6, -6, 1, -2, -2, 2, -3, 1, 2,
    -- filter=188 channel=44
    -2, 20, -17, -7, 15, -13, 5, 1, -6,
    -- filter=188 channel=45
    -1, -7, -12, 0, -7, -6, -3, -2, -8,
    -- filter=188 channel=46
    -2, -2, 2, 0, -5, 6, 3, -3, 9,
    -- filter=188 channel=47
    2, 11, -19, -6, 18, -26, 3, 9, -12,
    -- filter=188 channel=48
    -5, 17, -7, -7, 11, -18, -9, 6, 0,
    -- filter=188 channel=49
    -6, 4, -5, -12, -7, 1, -4, -11, 5,
    -- filter=188 channel=50
    -3, 5, -11, -7, 0, -7, -2, -7, -4,
    -- filter=188 channel=51
    5, 4, -3, 0, -2, -7, 0, -3, -5,
    -- filter=188 channel=52
    3, 24, 3, 0, 17, 6, 5, 9, 14,
    -- filter=188 channel=53
    -6, 0, 3, 4, -8, 4, 4, -9, 2,
    -- filter=188 channel=54
    5, 0, 0, -5, 1, 4, -7, 6, -5,
    -- filter=188 channel=55
    2, 9, -6, 6, 7, -8, 6, -8, 1,
    -- filter=188 channel=56
    -7, 10, 3, -2, 13, 20, 0, 7, 11,
    -- filter=188 channel=57
    0, -7, 6, -3, 3, 9, -7, 6, -3,
    -- filter=188 channel=58
    3, 9, 0, 4, 5, 0, 0, -4, 4,
    -- filter=188 channel=59
    -6, 14, -7, 3, 10, -17, 5, 6, -11,
    -- filter=188 channel=60
    0, -3, 3, 6, 0, -4, -3, 0, -7,
    -- filter=188 channel=61
    1, 14, -7, 6, 17, -5, 1, 4, 0,
    -- filter=188 channel=62
    4, 3, 7, 3, 2, 0, -3, 4, -3,
    -- filter=188 channel=63
    0, 4, -4, 4, 8, -4, 9, 8, -1,
    -- filter=188 channel=64
    -3, -2, 3, 4, 3, 6, 5, -2, 0,
    -- filter=188 channel=65
    -1, 0, 2, -2, -1, 5, 1, 3, -6,
    -- filter=188 channel=66
    21, 13, 1, 19, 23, 0, 0, 5, -9,
    -- filter=188 channel=67
    0, 7, 6, 4, -8, 0, 5, -5, -6,
    -- filter=188 channel=68
    0, 0, -7, -3, -10, 2, 0, -10, 3,
    -- filter=188 channel=69
    9, 1, -5, -4, 8, -6, -3, -1, -2,
    -- filter=188 channel=70
    -11, 15, 0, -11, 17, 5, -2, 7, 8,
    -- filter=188 channel=71
    0, -5, -10, 0, -11, -10, -7, -8, -5,
    -- filter=188 channel=72
    -7, 1, -6, -8, 5, -19, 3, 0, -7,
    -- filter=188 channel=73
    -7, 5, -5, 0, 2, -9, 0, -2, 3,
    -- filter=188 channel=74
    -7, 32, -1, -3, 22, 1, 6, 12, 15,
    -- filter=188 channel=75
    -8, 5, 3, -6, 28, -7, 7, 8, -12,
    -- filter=188 channel=76
    -3, -6, 5, 5, -2, -2, -4, -7, 5,
    -- filter=188 channel=77
    3, 2, -2, -4, -4, -5, 0, 3, 6,
    -- filter=188 channel=78
    2, 6, -6, 6, 0, -8, -5, -1, 0,
    -- filter=188 channel=79
    -7, 11, -6, 0, 19, -4, 4, -5, -2,
    -- filter=188 channel=80
    -11, 0, -22, 0, 12, -22, -3, 6, -16,
    -- filter=188 channel=81
    6, 6, -4, 1, 5, 0, -6, 3, -4,
    -- filter=188 channel=82
    2, -4, -3, -1, 4, -5, -1, -3, 2,
    -- filter=188 channel=83
    -11, -3, 0, 4, -2, 1, -5, 6, -1,
    -- filter=188 channel=84
    -4, 12, -5, 7, 12, -4, 1, -1, 12,
    -- filter=188 channel=85
    -4, 3, -1, -5, 0, 6, -7, 1, 2,
    -- filter=188 channel=86
    10, 19, -8, 5, 30, 3, -2, 16, 1,
    -- filter=188 channel=87
    7, 19, 0, 0, 15, 15, 0, 2, 14,
    -- filter=188 channel=88
    -9, 12, -6, -1, 3, 3, 5, 10, 4,
    -- filter=188 channel=89
    -3, 0, -6, -9, 2, -20, -2, 0, -6,
    -- filter=188 channel=90
    3, 13, 4, 0, 6, 9, -2, 5, 13,
    -- filter=188 channel=91
    -1, 13, -11, -9, 6, 1, 1, -6, 10,
    -- filter=188 channel=92
    -10, 6, 3, -5, 5, 5, -10, 4, 4,
    -- filter=188 channel=93
    -7, 20, -9, -8, 11, -22, 1, 14, 2,
    -- filter=188 channel=94
    5, -1, -4, -7, -3, -6, 1, 2, 1,
    -- filter=188 channel=95
    0, 3, 0, 0, -4, -3, 2, 5, -5,
    -- filter=188 channel=96
    -6, -10, 2, -1, -7, 3, -1, -2, 1,
    -- filter=188 channel=97
    -9, -12, -5, -5, -5, 0, -5, -6, 2,
    -- filter=188 channel=98
    -12, 3, -14, -10, 19, -32, 0, 5, -5,
    -- filter=188 channel=99
    -2, 32, -17, -8, 25, -25, 2, 14, 10,
    -- filter=188 channel=100
    6, 13, 19, -2, 13, 13, -5, 11, 17,
    -- filter=188 channel=101
    -6, -2, -13, -7, -13, -1, -12, -6, -6,
    -- filter=188 channel=102
    -2, 3, 4, -6, 7, -3, 4, 2, -3,
    -- filter=188 channel=103
    -9, 5, -21, -4, 20, -36, 2, 9, -1,
    -- filter=188 channel=104
    -8, 13, -21, -1, 9, -13, -4, 8, 3,
    -- filter=188 channel=105
    -3, 0, 2, -8, -9, 3, -1, -13, 2,
    -- filter=188 channel=106
    -6, 0, 12, 3, -1, 13, 2, -9, 0,
    -- filter=188 channel=107
    3, 7, -2, -3, 9, -7, 2, 5, 7,
    -- filter=188 channel=108
    -2, -5, 11, 0, 4, 9, 3, -2, -6,
    -- filter=188 channel=109
    2, 23, -19, 5, 27, -18, 6, 0, 6,
    -- filter=188 channel=110
    -10, 0, -1, -1, 18, 3, 0, 3, 2,
    -- filter=188 channel=111
    6, -7, 5, 1, -1, 2, -8, 6, -3,
    -- filter=188 channel=112
    -10, 16, -11, 2, 7, -11, -7, 4, 4,
    -- filter=188 channel=113
    -8, 8, -3, -3, 15, -11, -2, 9, 5,
    -- filter=188 channel=114
    -5, 14, -14, -1, 22, -16, 0, -3, -6,
    -- filter=188 channel=115
    2, 0, -6, -4, 1, 7, 0, 7, 7,
    -- filter=188 channel=116
    -11, 3, -10, -5, 0, -7, -4, -8, -1,
    -- filter=188 channel=117
    1, 2, -5, -3, 0, 3, -8, 3, -1,
    -- filter=188 channel=118
    -5, -3, -6, -5, 6, 7, -7, -2, 0,
    -- filter=188 channel=119
    2, 34, 14, 7, 31, 35, -8, 23, 14,
    -- filter=188 channel=120
    -11, 30, -19, -5, 12, -24, -8, -6, 0,
    -- filter=188 channel=121
    5, 8, 7, 0, 15, 1, 7, 12, -4,
    -- filter=188 channel=122
    -6, 23, -26, 1, 34, -25, 0, 14, -13,
    -- filter=188 channel=123
    2, 5, 1, 0, 15, 9, 5, 11, 9,
    -- filter=188 channel=124
    6, 2, 3, 5, -2, -7, 1, -3, -5,
    -- filter=188 channel=125
    -10, 22, -20, 4, 22, -22, 0, 1, -6,
    -- filter=188 channel=126
    3, -5, -1, 0, 3, 4, -12, -7, -16,
    -- filter=188 channel=127
    0, 0, 14, 3, 3, 7, -3, 3, 9,
    -- filter=189 channel=0
    -7, -12, 1, -2, -1, 10, -11, -4, 0,
    -- filter=189 channel=1
    -6, 0, -4, -10, 6, 13, -2, -5, -1,
    -- filter=189 channel=2
    0, 1, 0, 4, 7, 8, -6, 3, -3,
    -- filter=189 channel=3
    -7, 3, -1, -1, 2, 0, 0, -4, -3,
    -- filter=189 channel=4
    -1, 12, 0, -4, -1, 8, 1, -7, 0,
    -- filter=189 channel=5
    -7, -1, -2, 2, 4, 5, 2, 9, 1,
    -- filter=189 channel=6
    5, 3, 13, -2, 1, 9, -11, -4, 5,
    -- filter=189 channel=7
    1, -3, 6, 1, -2, 3, 6, 6, -7,
    -- filter=189 channel=8
    -1, -9, -5, 2, 0, 5, -6, -4, -8,
    -- filter=189 channel=9
    2, -4, -4, -3, -1, 8, 2, 3, 2,
    -- filter=189 channel=10
    -1, -8, -10, 3, 11, -3, 1, 6, 5,
    -- filter=189 channel=11
    8, 2, 6, 3, 4, -4, -2, -5, -11,
    -- filter=189 channel=12
    3, 0, 4, 3, -3, 1, 1, 0, 0,
    -- filter=189 channel=13
    2, -4, 1, -6, 11, 7, -3, 1, -2,
    -- filter=189 channel=14
    -1, 5, 2, -2, 4, 5, -3, 2, -3,
    -- filter=189 channel=15
    2, 0, 6, -2, 11, 5, -12, -10, -10,
    -- filter=189 channel=16
    -6, -10, -8, 0, 0, -6, 7, 5, 3,
    -- filter=189 channel=17
    0, 2, 5, -4, 1, -1, 2, -7, -6,
    -- filter=189 channel=18
    4, 11, -1, 0, 16, 14, -13, -3, 0,
    -- filter=189 channel=19
    0, 0, 4, 0, 0, 0, -3, -1, 3,
    -- filter=189 channel=20
    7, 9, 16, 5, -1, 3, -15, -16, -12,
    -- filter=189 channel=21
    -5, -16, -15, 7, -4, -13, 5, 17, 10,
    -- filter=189 channel=22
    -8, -5, 5, -2, 8, 3, -1, 0, 2,
    -- filter=189 channel=23
    0, -11, 1, 3, -2, -5, -13, -6, -2,
    -- filter=189 channel=24
    3, -1, -4, 1, 4, -2, 4, -6, 6,
    -- filter=189 channel=25
    0, -5, -8, -7, 12, 11, 0, 4, 4,
    -- filter=189 channel=26
    1, -3, -1, -5, 0, 2, -3, 6, 2,
    -- filter=189 channel=27
    5, -17, -5, 5, 16, 8, -6, 2, 9,
    -- filter=189 channel=28
    -6, -3, -1, -5, -4, 5, -5, -5, 0,
    -- filter=189 channel=29
    5, 20, 20, -6, 6, 10, -15, -18, -9,
    -- filter=189 channel=30
    0, -10, 0, 0, 2, 0, 4, 5, -2,
    -- filter=189 channel=31
    -5, -12, -9, 0, 8, -12, 8, 20, 6,
    -- filter=189 channel=32
    4, 5, -5, -1, 10, 11, -8, -5, -5,
    -- filter=189 channel=33
    -4, -9, -10, -3, 13, 8, -9, 0, 12,
    -- filter=189 channel=34
    -6, -17, 2, 0, -8, -9, -5, -5, -11,
    -- filter=189 channel=35
    4, 3, -7, -3, -7, -2, -3, -3, 7,
    -- filter=189 channel=36
    4, 8, 2, 9, 3, -10, 9, 5, -8,
    -- filter=189 channel=37
    -10, -2, -15, -2, 2, 3, -5, -1, 11,
    -- filter=189 channel=38
    6, -7, 0, 1, 1, 4, 3, 3, -3,
    -- filter=189 channel=39
    9, 0, 6, 0, 7, -3, 2, -7, -6,
    -- filter=189 channel=40
    3, 8, 0, 4, 2, -8, -6, 2, -9,
    -- filter=189 channel=41
    -2, 10, -4, -11, 0, -16, 2, -3, -14,
    -- filter=189 channel=42
    0, 1, 1, 0, 5, 2, 6, 5, 3,
    -- filter=189 channel=43
    -14, -5, 7, -8, -1, 0, -12, -9, -6,
    -- filter=189 channel=44
    -10, -7, -13, 0, 6, -1, 0, 13, 12,
    -- filter=189 channel=45
    0, -3, -2, -5, 7, 2, -3, 6, 2,
    -- filter=189 channel=46
    1, 0, -6, -1, -4, -2, -5, 1, 6,
    -- filter=189 channel=47
    0, -4, -16, -3, 1, -3, 12, 10, 5,
    -- filter=189 channel=48
    3, -5, -15, -6, 2, 11, 12, 1, 12,
    -- filter=189 channel=49
    4, 13, 4, -7, 10, 15, -5, -10, -6,
    -- filter=189 channel=50
    0, -5, -9, 5, 10, 9, -1, 8, 2,
    -- filter=189 channel=51
    -5, 0, 4, -3, 1, 2, 3, 0, 3,
    -- filter=189 channel=52
    -3, -10, -1, 7, -5, 5, -2, 3, -3,
    -- filter=189 channel=53
    4, 6, -2, 7, 2, 4, -4, -12, 0,
    -- filter=189 channel=54
    7, -7, 2, -7, 3, 7, 7, 0, 3,
    -- filter=189 channel=55
    8, 8, 7, -6, 0, -3, -15, -10, -6,
    -- filter=189 channel=56
    6, -10, 2, 2, -3, -6, 4, 1, -3,
    -- filter=189 channel=57
    -7, -2, 3, -5, 0, -6, -4, -2, 4,
    -- filter=189 channel=58
    3, -4, -4, 0, -3, -1, -4, 7, 6,
    -- filter=189 channel=59
    -1, -7, -5, -5, 0, -1, 4, 0, 12,
    -- filter=189 channel=60
    5, -2, 0, -1, 4, 2, 5, 0, 4,
    -- filter=189 channel=61
    3, -4, 2, 2, -2, 0, -4, 2, -9,
    -- filter=189 channel=62
    6, -4, 0, 6, 0, -1, 1, -8, -1,
    -- filter=189 channel=63
    -3, 2, -5, -2, 4, 4, 0, 5, 5,
    -- filter=189 channel=64
    0, 2, 2, 2, 2, -10, -1, 3, -10,
    -- filter=189 channel=65
    6, -5, 6, -5, -4, 2, 4, -1, 5,
    -- filter=189 channel=66
    -3, 0, 5, 0, -1, -3, -6, 1, -8,
    -- filter=189 channel=67
    -4, 6, 3, 0, -7, 0, 2, 0, 0,
    -- filter=189 channel=68
    -7, -2, 3, 4, -2, -5, 3, -6, -1,
    -- filter=189 channel=69
    6, 1, -7, 0, -5, 6, -7, -7, 0,
    -- filter=189 channel=70
    5, -10, 5, 0, 3, 0, -11, -1, 8,
    -- filter=189 channel=71
    -5, -4, 4, 1, -3, -8, 0, -1, 2,
    -- filter=189 channel=72
    -2, -5, -13, 3, 1, -4, 4, 2, 2,
    -- filter=189 channel=73
    -1, -1, -1, -7, 0, 6, -6, -6, 6,
    -- filter=189 channel=74
    3, -8, -4, 5, 3, -1, 0, -2, 1,
    -- filter=189 channel=75
    -4, -8, -15, 7, 0, 4, -4, 10, 6,
    -- filter=189 channel=76
    8, 5, 13, 3, -6, -6, -11, -14, -16,
    -- filter=189 channel=77
    -4, -1, -4, -4, 4, 1, -4, -1, -5,
    -- filter=189 channel=78
    -3, 4, 5, 9, -6, -1, 6, 0, 7,
    -- filter=189 channel=79
    3, 3, -2, -1, 15, 19, -8, -2, 4,
    -- filter=189 channel=80
    5, -15, -21, 0, 8, -6, 6, 14, 2,
    -- filter=189 channel=81
    7, 4, -7, 0, -2, -5, -6, -6, -3,
    -- filter=189 channel=82
    -6, 4, 0, -2, -5, -4, 5, 1, -6,
    -- filter=189 channel=83
    -6, -2, -5, 3, 0, 5, -4, -7, 1,
    -- filter=189 channel=84
    9, -1, 10, -1, 10, 14, -2, -9, -3,
    -- filter=189 channel=85
    1, -2, 3, -4, 4, 4, 0, 5, -7,
    -- filter=189 channel=86
    2, -8, 0, 0, 5, -5, -1, -4, -3,
    -- filter=189 channel=87
    -6, 6, 5, -2, -2, 3, -2, -6, 0,
    -- filter=189 channel=88
    -1, -2, -8, 4, -1, 0, 7, -2, 0,
    -- filter=189 channel=89
    1, -2, -8, 6, 13, 0, -9, 0, -5,
    -- filter=189 channel=90
    -4, 2, 2, 0, -7, -1, 2, 6, -8,
    -- filter=189 channel=91
    4, -5, 3, -5, 9, 6, -1, -7, 6,
    -- filter=189 channel=92
    -2, -3, 1, 5, -7, -8, 3, 4, 2,
    -- filter=189 channel=93
    -2, -4, -20, 2, 0, 4, 0, -1, 0,
    -- filter=189 channel=94
    -2, 3, 2, -5, 4, 0, 0, 0, -1,
    -- filter=189 channel=95
    -2, -6, -6, -4, 5, -5, -2, -2, 0,
    -- filter=189 channel=96
    1, -5, -5, -1, 0, 5, -7, -1, -2,
    -- filter=189 channel=97
    -5, -8, -5, 1, 0, -6, -2, 0, 1,
    -- filter=189 channel=98
    3, -4, -11, 5, 14, 10, 0, -1, 0,
    -- filter=189 channel=99
    4, -13, -9, 13, 0, -1, -3, 3, -4,
    -- filter=189 channel=100
    6, -7, -6, 0, -5, -7, 4, -8, 3,
    -- filter=189 channel=101
    -2, -2, 7, 1, 2, 4, 6, -4, -5,
    -- filter=189 channel=102
    2, 3, 6, -5, 0, 0, -7, 6, 5,
    -- filter=189 channel=103
    -9, -8, -5, -2, 2, -9, 8, 18, 16,
    -- filter=189 channel=104
    -5, -11, -19, -2, 0, 2, 13, 14, 9,
    -- filter=189 channel=105
    -3, 11, 13, -5, -5, 5, -12, -11, -10,
    -- filter=189 channel=106
    0, 0, 0, 0, 7, 3, 5, -3, 1,
    -- filter=189 channel=107
    3, 11, 9, 0, 0, 6, -14, -11, 0,
    -- filter=189 channel=108
    -1, 1, -1, -7, 0, -2, -6, 2, -8,
    -- filter=189 channel=109
    -5, -7, -11, 6, 8, 10, -8, -3, 1,
    -- filter=189 channel=110
    2, -11, 0, 5, 2, -9, -2, 7, 0,
    -- filter=189 channel=111
    0, -1, 4, -4, -4, 0, -4, -4, 0,
    -- filter=189 channel=112
    -3, -6, -7, 1, 8, 7, 3, -3, 3,
    -- filter=189 channel=113
    0, -4, -8, 2, 2, 0, 1, 6, 4,
    -- filter=189 channel=114
    4, 6, 2, -14, 4, 27, -7, -2, 8,
    -- filter=189 channel=115
    4, -2, 5, 0, 5, -2, -5, 0, -1,
    -- filter=189 channel=116
    -2, 2, -11, -5, 13, -1, 5, -1, 3,
    -- filter=189 channel=117
    -6, 0, 3, 1, 9, 6, 1, 7, 0,
    -- filter=189 channel=118
    2, 3, 6, 1, 3, 0, -3, 1, 1,
    -- filter=189 channel=119
    -9, -3, 0, 4, -11, -6, -8, -3, -9,
    -- filter=189 channel=120
    -4, -7, 6, 7, 0, 12, -5, -1, 2,
    -- filter=189 channel=121
    5, 4, -7, 4, 7, -9, 8, -3, -1,
    -- filter=189 channel=122
    -9, -18, -32, 7, 5, -1, 10, 14, 7,
    -- filter=189 channel=123
    -2, -8, 5, 0, -9, -5, -5, -6, -6,
    -- filter=189 channel=124
    5, 0, 0, 1, -3, 1, -2, -8, -11,
    -- filter=189 channel=125
    8, 2, -7, 1, 4, 2, 3, 0, 0,
    -- filter=189 channel=126
    3, -1, -6, 0, 3, -5, 2, 1, 1,
    -- filter=189 channel=127
    0, -3, -8, 3, 0, -9, 2, -6, 4,
    -- filter=190 channel=0
    0, 0, 1, 7, 3, -4, -2, 4, -2,
    -- filter=190 channel=1
    4, 0, -2, -5, 5, -1, -5, -7, 2,
    -- filter=190 channel=2
    3, 3, -2, 1, 4, -1, -5, 5, -5,
    -- filter=190 channel=3
    -2, 0, 1, -3, 1, -1, 1, 1, 8,
    -- filter=190 channel=4
    1, 3, -2, -3, -6, 5, -2, -5, -5,
    -- filter=190 channel=5
    -1, 10, 0, 0, 5, 8, 3, 0, 0,
    -- filter=190 channel=6
    1, 2, -3, -3, -3, 4, 7, -2, -2,
    -- filter=190 channel=7
    1, 2, 7, 0, -1, -5, -2, -7, -2,
    -- filter=190 channel=8
    1, 6, 1, 6, -2, -2, -3, -3, -4,
    -- filter=190 channel=9
    2, 4, 0, 3, -5, -4, -7, 1, -1,
    -- filter=190 channel=10
    -2, -8, -6, 2, 0, 0, 1, -5, -6,
    -- filter=190 channel=11
    -2, -2, 2, 7, 0, -3, 0, 3, 5,
    -- filter=190 channel=12
    6, 4, -8, -2, -6, 2, 0, -4, 0,
    -- filter=190 channel=13
    -4, -3, -2, -6, -5, -7, 6, -2, -5,
    -- filter=190 channel=14
    5, -5, -5, 2, -7, 3, 7, 5, -2,
    -- filter=190 channel=15
    -1, 2, -1, 6, 3, 1, 4, 0, 7,
    -- filter=190 channel=16
    3, 3, 3, 0, -3, 0, 3, 1, 4,
    -- filter=190 channel=17
    -4, -6, -6, -1, 3, -6, -1, 1, -1,
    -- filter=190 channel=18
    3, -2, -5, -2, -3, -1, 1, -6, -7,
    -- filter=190 channel=19
    -1, 0, 4, 5, -5, 3, -2, 6, -3,
    -- filter=190 channel=20
    5, -5, -1, 2, 0, 7, 11, 14, 7,
    -- filter=190 channel=21
    0, 1, 9, 4, -1, 0, -3, 7, -2,
    -- filter=190 channel=22
    1, -2, 2, -3, 5, -5, 6, -5, -5,
    -- filter=190 channel=23
    -5, -4, 6, -7, 6, -3, 0, 1, -6,
    -- filter=190 channel=24
    -5, -3, 3, -1, -3, 0, 3, -6, 3,
    -- filter=190 channel=25
    -7, -4, -5, -4, 1, -9, 1, -9, -6,
    -- filter=190 channel=26
    -1, 1, 8, 8, 7, -2, 5, -1, -3,
    -- filter=190 channel=27
    1, -3, 3, -10, -4, -4, -1, -5, 4,
    -- filter=190 channel=28
    -3, -1, 1, -6, 5, -7, -4, 0, 4,
    -- filter=190 channel=29
    2, -9, 0, -1, 5, -6, 4, 0, 9,
    -- filter=190 channel=30
    4, 3, 4, -1, -4, 6, -1, -1, 0,
    -- filter=190 channel=31
    5, 1, 1, 3, -7, 1, -5, -5, -4,
    -- filter=190 channel=32
    -2, 2, 4, 1, -3, 0, -2, -1, -3,
    -- filter=190 channel=33
    0, -7, -8, -4, -1, 3, -3, 2, -2,
    -- filter=190 channel=34
    0, -7, -5, 4, -6, 0, 0, 3, -1,
    -- filter=190 channel=35
    3, 0, -2, 2, -1, 0, -4, -5, -6,
    -- filter=190 channel=36
    -3, -5, -3, 8, -2, -2, 3, 7, -5,
    -- filter=190 channel=37
    7, 9, 3, 0, 7, 6, -4, -4, -1,
    -- filter=190 channel=38
    0, 5, 4, 3, 6, -6, -8, 3, -2,
    -- filter=190 channel=39
    5, 1, 7, 0, 4, -2, 9, -1, 6,
    -- filter=190 channel=40
    9, 0, 8, 1, 0, 1, 9, 0, 4,
    -- filter=190 channel=41
    4, -4, -9, 12, -12, -11, 0, -11, -2,
    -- filter=190 channel=42
    -5, -1, -6, -6, 4, 0, 5, -6, -5,
    -- filter=190 channel=43
    0, 0, 7, 2, 8, -2, 8, 7, 5,
    -- filter=190 channel=44
    -1, 6, 8, -8, -6, 7, -1, 1, 2,
    -- filter=190 channel=45
    4, 3, 5, -1, 6, 4, 1, -2, 7,
    -- filter=190 channel=46
    0, -3, 4, 7, 5, 5, 0, 7, -5,
    -- filter=190 channel=47
    -7, 4, -2, 4, -6, 6, -3, -7, 0,
    -- filter=190 channel=48
    -2, 0, 0, -4, 4, -2, -5, -5, -6,
    -- filter=190 channel=49
    -4, -7, -7, 1, 1, 1, -2, -3, 5,
    -- filter=190 channel=50
    -1, 3, 3, 1, 6, 6, -3, -1, 3,
    -- filter=190 channel=51
    4, 3, -5, -1, 3, -5, 3, -2, 0,
    -- filter=190 channel=52
    -3, -1, -5, 0, 2, 7, 5, 6, 4,
    -- filter=190 channel=53
    1, -7, -3, 2, -7, -6, 4, 0, 1,
    -- filter=190 channel=54
    0, -6, 2, 0, -5, -5, -7, -3, 7,
    -- filter=190 channel=55
    2, -6, -8, -1, -7, -3, -2, 6, -4,
    -- filter=190 channel=56
    -4, 0, -1, 1, 4, 0, -5, -3, -2,
    -- filter=190 channel=57
    4, -5, -1, 7, 3, -2, 0, -1, 0,
    -- filter=190 channel=58
    0, -1, 7, 3, -5, 3, 3, 7, -4,
    -- filter=190 channel=59
    -1, -4, 2, -9, 3, 3, -3, -5, 2,
    -- filter=190 channel=60
    1, 5, 2, 7, 2, -6, 0, -1, -6,
    -- filter=190 channel=61
    -1, 6, 6, -4, 0, -7, -5, -1, -1,
    -- filter=190 channel=62
    3, 5, -7, 5, 4, 4, -2, -2, 3,
    -- filter=190 channel=63
    3, 2, 0, -1, 7, 2, -1, -3, 0,
    -- filter=190 channel=64
    -4, 4, -2, -4, 2, -3, -3, -2, -1,
    -- filter=190 channel=65
    -7, 2, 5, 1, -4, 0, 0, 2, 7,
    -- filter=190 channel=66
    6, -7, -4, 8, 1, -6, -4, 4, -4,
    -- filter=190 channel=67
    -1, 7, -6, 0, -1, -5, -5, 0, 6,
    -- filter=190 channel=68
    0, 6, 7, 5, 2, -2, 3, 6, -2,
    -- filter=190 channel=69
    -3, 7, 3, 3, -5, 4, 3, 3, -5,
    -- filter=190 channel=70
    4, 3, -4, -6, -7, 5, -3, 4, -1,
    -- filter=190 channel=71
    -3, 0, 5, -3, 8, -3, 4, -4, 7,
    -- filter=190 channel=72
    -6, -6, -5, -6, -3, 6, -6, -5, -4,
    -- filter=190 channel=73
    -4, -1, -6, -5, 1, 3, -5, 6, 0,
    -- filter=190 channel=74
    6, 6, 3, -2, 2, 4, -1, 3, -4,
    -- filter=190 channel=75
    4, 0, -3, 0, -3, 3, 2, -2, 3,
    -- filter=190 channel=76
    -2, -1, 2, 5, 9, 0, 12, 0, 10,
    -- filter=190 channel=77
    6, -7, -2, -4, 3, 3, 0, 7, -6,
    -- filter=190 channel=78
    -6, 4, -2, 4, 4, -3, -7, -6, -4,
    -- filter=190 channel=79
    2, -8, 0, -1, -3, -3, 0, -9, -9,
    -- filter=190 channel=80
    2, -3, 6, -4, 0, 0, 0, 0, 4,
    -- filter=190 channel=81
    -5, 3, -3, -6, 5, 0, -3, 1, 5,
    -- filter=190 channel=82
    -6, 2, 7, -3, 5, 5, 3, 5, 2,
    -- filter=190 channel=83
    -2, -7, -3, -8, -2, -2, 0, -2, -6,
    -- filter=190 channel=84
    0, -2, -1, -5, -3, -6, -7, 1, -2,
    -- filter=190 channel=85
    5, 3, -6, -3, 0, 3, 0, 7, 0,
    -- filter=190 channel=86
    -2, -1, 0, -3, -7, -4, 0, 0, -5,
    -- filter=190 channel=87
    0, 3, -7, 6, -5, 7, 8, -2, -1,
    -- filter=190 channel=88
    0, -4, 6, 1, 3, 6, 4, 2, 0,
    -- filter=190 channel=89
    -3, 0, 0, 0, -8, -5, -4, 1, -2,
    -- filter=190 channel=90
    3, 9, 10, -3, 1, 8, 6, 8, -1,
    -- filter=190 channel=91
    -9, 1, -6, 5, 5, -4, 1, -6, 3,
    -- filter=190 channel=92
    0, 0, -3, 1, -6, 0, -5, 5, 4,
    -- filter=190 channel=93
    -3, 3, 9, -4, 1, -3, -9, -4, -3,
    -- filter=190 channel=94
    2, -2, 1, -3, 6, 3, -2, -4, 6,
    -- filter=190 channel=95
    1, -7, 0, 3, -3, -3, -6, 5, 1,
    -- filter=190 channel=96
    6, 5, -3, 3, 0, 0, -6, -5, 5,
    -- filter=190 channel=97
    8, 5, -1, 3, -4, 8, 8, -6, 6,
    -- filter=190 channel=98
    -3, 0, 4, 1, -8, 0, 2, -9, -7,
    -- filter=190 channel=99
    4, -7, 3, -6, 1, 6, 0, -9, -1,
    -- filter=190 channel=100
    0, -6, -2, -6, 1, -5, 0, -1, -5,
    -- filter=190 channel=101
    1, 0, -2, 5, -3, -5, -6, 8, -5,
    -- filter=190 channel=102
    0, 2, -5, 0, -6, 0, -4, -4, 1,
    -- filter=190 channel=103
    -1, 2, 6, -3, -1, 5, -5, 0, 4,
    -- filter=190 channel=104
    -6, 7, -1, -8, -7, -7, 4, -3, 3,
    -- filter=190 channel=105
    5, 4, -5, -3, -4, -6, 6, 10, -1,
    -- filter=190 channel=106
    -3, 0, -4, 5, -2, -3, -2, -2, 6,
    -- filter=190 channel=107
    -3, 4, 7, 7, 5, 7, 4, 4, 0,
    -- filter=190 channel=108
    4, 4, -2, 0, -2, 0, 5, -2, 5,
    -- filter=190 channel=109
    -7, 0, 0, -4, 4, -3, -2, -9, 4,
    -- filter=190 channel=110
    2, -6, 0, -7, -1, 5, -4, -5, 3,
    -- filter=190 channel=111
    -2, 4, 4, 7, -2, -4, -4, 0, 0,
    -- filter=190 channel=112
    5, 7, -2, 0, 5, 5, 0, 2, 6,
    -- filter=190 channel=113
    2, -2, 1, -8, -6, 2, -1, 5, -7,
    -- filter=190 channel=114
    -9, -5, -1, 0, 2, -8, -8, -7, 1,
    -- filter=190 channel=115
    -3, -1, 4, 5, 2, -5, -5, 5, -6,
    -- filter=190 channel=116
    3, -9, -8, 0, 2, -4, 4, -6, -2,
    -- filter=190 channel=117
    -4, -6, 3, 0, -2, -6, -3, 2, -4,
    -- filter=190 channel=118
    0, 3, 0, 1, -4, -3, 7, 4, 4,
    -- filter=190 channel=119
    -4, 6, 6, 1, -7, 2, -5, 1, 6,
    -- filter=190 channel=120
    -8, -5, 5, -3, 2, 0, 4, 2, -3,
    -- filter=190 channel=121
    5, -4, 3, 7, 3, 1, -4, -5, -5,
    -- filter=190 channel=122
    -3, 8, 1, -1, 7, 3, -6, 4, 7,
    -- filter=190 channel=123
    -1, 5, 5, 6, 3, -3, 1, -5, 4,
    -- filter=190 channel=124
    -1, 0, -7, -5, 7, -4, 3, -5, 0,
    -- filter=190 channel=125
    -8, 1, 1, -10, 0, -8, 1, -3, -1,
    -- filter=190 channel=126
    -6, -6, -4, -1, -2, -6, -1, 4, -7,
    -- filter=190 channel=127
    -6, -8, 1, 1, -4, 0, -4, 2, -1,
    -- filter=191 channel=0
    -12, -18, -17, -14, -16, -12, 2, -15, -16,
    -- filter=191 channel=1
    -15, -17, -1, -18, -19, -8, -17, -13, -11,
    -- filter=191 channel=2
    1, 7, -6, 3, 3, -1, 5, -2, -4,
    -- filter=191 channel=3
    -3, -9, -10, -7, -5, -9, 1, -7, -2,
    -- filter=191 channel=4
    -4, 0, -6, 0, -6, 0, -5, -3, -8,
    -- filter=191 channel=5
    -12, -22, -3, -5, -9, -3, -4, -17, -7,
    -- filter=191 channel=6
    6, -1, -10, 9, 5, -11, 5, 6, -14,
    -- filter=191 channel=7
    5, -2, -2, -4, 0, 7, 1, -7, -7,
    -- filter=191 channel=8
    6, 4, -1, 0, -5, -3, -4, 3, 3,
    -- filter=191 channel=9
    -11, -8, 1, -4, 4, 3, -5, -3, 0,
    -- filter=191 channel=10
    -7, -3, 0, -4, 9, 15, 0, -5, 6,
    -- filter=191 channel=11
    8, 15, -11, 12, 6, -12, 9, -1, -6,
    -- filter=191 channel=12
    -1, 9, 8, -2, 5, 4, -6, -1, 11,
    -- filter=191 channel=13
    -4, -2, 2, 2, 11, 10, -2, 0, -3,
    -- filter=191 channel=14
    -1, -4, 3, 2, -5, -1, 5, 0, -5,
    -- filter=191 channel=15
    3, 4, -19, 10, 11, -10, -4, 4, -9,
    -- filter=191 channel=16
    -12, -6, 11, -15, 0, 14, -12, -3, 6,
    -- filter=191 channel=17
    7, -4, 6, 0, 0, 6, 0, 7, -6,
    -- filter=191 channel=18
    -12, -4, -16, -8, 4, -27, -7, 0, -17,
    -- filter=191 channel=19
    -6, -5, -1, 5, -1, 1, 6, 3, 3,
    -- filter=191 channel=20
    17, 10, -17, 16, 18, -5, 12, 12, -8,
    -- filter=191 channel=21
    -4, -2, 18, -1, -5, 13, -13, -4, 8,
    -- filter=191 channel=22
    0, -9, -9, 2, -10, -8, -3, 6, 0,
    -- filter=191 channel=23
    0, 0, 1, 13, 18, -10, 0, 10, -3,
    -- filter=191 channel=24
    6, 0, 6, 6, -6, 4, 4, 4, 2,
    -- filter=191 channel=25
    -12, 0, -1, -16, 5, 6, -18, -3, 2,
    -- filter=191 channel=26
    3, -1, 4, -8, -8, 7, 1, 0, -2,
    -- filter=191 channel=27
    -14, 2, -5, -2, 7, -7, -11, -2, -2,
    -- filter=191 channel=28
    -5, -2, -5, 7, 4, 5, 3, 1, 7,
    -- filter=191 channel=29
    11, 6, -17, 5, 15, -13, 0, 8, -17,
    -- filter=191 channel=30
    -10, 0, 3, -5, 1, -2, -7, -2, -2,
    -- filter=191 channel=31
    -4, 5, 20, -1, 15, 19, -10, -2, 11,
    -- filter=191 channel=32
    -9, 1, -8, 0, 10, -14, -7, -5, -11,
    -- filter=191 channel=33
    -12, -9, 3, -15, -6, -1, -7, 6, 2,
    -- filter=191 channel=34
    6, -3, 6, -1, -6, 5, -1, 8, 5,
    -- filter=191 channel=35
    4, -1, -1, 2, 3, -2, -7, -7, -5,
    -- filter=191 channel=36
    11, 9, 16, 0, 14, 17, -4, 2, 13,
    -- filter=191 channel=37
    -19, -16, -10, -20, -23, -11, -19, -15, -5,
    -- filter=191 channel=38
    -2, -1, 1, -8, 3, 7, -4, 0, 0,
    -- filter=191 channel=39
    1, 1, -2, 2, 9, -10, 2, -3, -12,
    -- filter=191 channel=40
    3, 4, 5, 0, 0, -9, 0, 8, -3,
    -- filter=191 channel=41
    0, -4, 0, -10, -5, 1, -12, -3, 2,
    -- filter=191 channel=42
    -6, -10, 0, -9, -8, -8, -9, -9, 0,
    -- filter=191 channel=43
    8, 2, -8, 3, -2, -14, 10, 9, -13,
    -- filter=191 channel=44
    -18, -4, 4, -21, -6, 0, -11, -12, 5,
    -- filter=191 channel=45
    -2, -3, -2, 0, 0, 0, -2, 7, -4,
    -- filter=191 channel=46
    -1, -8, 2, -2, 4, 4, 3, -10, 1,
    -- filter=191 channel=47
    -9, -8, 9, -18, -2, 9, -26, -6, 10,
    -- filter=191 channel=48
    -14, -4, 12, -17, -8, 7, -14, -6, 4,
    -- filter=191 channel=49
    7, -5, -12, -2, 1, -10, -1, 2, -17,
    -- filter=191 channel=50
    -5, 0, 5, -1, 0, -2, 1, 0, 0,
    -- filter=191 channel=51
    2, 1, 5, 0, -1, -3, -3, 2, 0,
    -- filter=191 channel=52
    3, 2, 6, 6, 0, 5, 4, 9, 6,
    -- filter=191 channel=53
    5, 7, -7, 10, 14, -1, 4, 0, -8,
    -- filter=191 channel=54
    -6, -7, -3, -1, -2, -3, 1, 4, -6,
    -- filter=191 channel=55
    -1, 9, 4, 1, 16, -3, 0, 14, -7,
    -- filter=191 channel=56
    -6, 0, 4, 6, -3, 5, -1, -1, 2,
    -- filter=191 channel=57
    -3, -6, 0, 1, 5, -2, 1, -5, 3,
    -- filter=191 channel=58
    -2, -13, -10, -6, -11, -6, 0, -10, -7,
    -- filter=191 channel=59
    -17, -7, 8, -16, -3, 17, -17, 0, 0,
    -- filter=191 channel=60
    -2, 1, 0, 5, 0, -1, 7, 7, -4,
    -- filter=191 channel=61
    0, -1, 7, 3, 3, 11, -5, 2, 6,
    -- filter=191 channel=62
    -6, 0, -1, -5, -1, -1, 5, 0, -5,
    -- filter=191 channel=63
    2, -2, -5, -1, -2, 2, -5, -10, -1,
    -- filter=191 channel=64
    1, 5, 7, 0, 9, 2, 1, 1, -2,
    -- filter=191 channel=65
    4, 4, 5, -1, 6, -2, 2, 2, 0,
    -- filter=191 channel=66
    -2, 3, 9, -6, 8, 8, 6, 8, 3,
    -- filter=191 channel=67
    -2, 1, 3, -4, -4, -7, 5, 4, 4,
    -- filter=191 channel=68
    3, -1, 4, -2, 3, 2, -4, 6, 6,
    -- filter=191 channel=69
    -5, 0, 3, 1, 5, 0, 4, 4, 2,
    -- filter=191 channel=70
    -10, -8, -11, -3, -4, -2, -7, -3, 0,
    -- filter=191 channel=71
    -5, -8, 8, -6, -4, -3, 5, -6, 6,
    -- filter=191 channel=72
    -8, 4, 18, -9, 4, 22, -2, -4, 5,
    -- filter=191 channel=73
    2, 2, 1, -2, 0, -4, -7, 8, -5,
    -- filter=191 channel=74
    0, 2, 13, -5, -3, 5, 0, 0, 1,
    -- filter=191 channel=75
    -20, -23, -11, -19, -17, -12, -4, -7, -13,
    -- filter=191 channel=76
    5, 17, -1, 6, 15, -4, 1, 15, -14,
    -- filter=191 channel=77
    6, 3, -3, 0, 7, 0, 1, -4, -5,
    -- filter=191 channel=78
    1, 3, -3, 4, -3, -2, 3, -6, 2,
    -- filter=191 channel=79
    -17, -6, -18, -8, -5, -21, -4, -3, -15,
    -- filter=191 channel=80
    -8, -8, 21, -17, 2, 18, -14, -4, 15,
    -- filter=191 channel=81
    -5, 0, 3, 3, 0, -6, 0, 6, -6,
    -- filter=191 channel=82
    0, 7, 3, 0, -5, -5, 0, 1, 1,
    -- filter=191 channel=83
    -3, -3, 8, -4, 7, -2, -8, -5, 7,
    -- filter=191 channel=84
    -1, -1, -13, 8, 6, -11, 0, 2, -1,
    -- filter=191 channel=85
    6, 6, 1, -1, 0, 3, 3, 0, 0,
    -- filter=191 channel=86
    0, -7, 1, 0, -2, 6, -2, 1, 7,
    -- filter=191 channel=87
    0, 9, -2, 14, 14, -5, 0, 3, 2,
    -- filter=191 channel=88
    7, 14, 21, 5, 3, 14, -6, 4, 16,
    -- filter=191 channel=89
    -13, -1, 6, -12, 19, 10, -2, 0, 1,
    -- filter=191 channel=90
    9, 4, 11, 12, 4, 11, 6, 3, 5,
    -- filter=191 channel=91
    3, 5, -3, 7, 1, -2, 1, 2, -4,
    -- filter=191 channel=92
    4, -6, 7, 3, -5, 8, 1, 3, 2,
    -- filter=191 channel=93
    -4, -7, 9, -13, -8, 0, -10, -22, -5,
    -- filter=191 channel=94
    -1, 1, 3, 6, 1, -6, -4, -4, 3,
    -- filter=191 channel=95
    -5, 0, 1, 5, -2, 0, -5, 0, 3,
    -- filter=191 channel=96
    -4, -5, -6, 0, -9, 4, -7, 0, -5,
    -- filter=191 channel=97
    -11, -10, -5, 2, -7, 0, -3, 0, 7,
    -- filter=191 channel=98
    -10, -9, 5, -11, 9, -2, -17, -4, 7,
    -- filter=191 channel=99
    3, 14, 10, 13, 18, 18, 0, 9, 8,
    -- filter=191 channel=100
    1, 1, 0, 1, 2, -4, -2, -3, -4,
    -- filter=191 channel=101
    -1, 4, 7, 3, -1, -4, -2, -8, 6,
    -- filter=191 channel=102
    0, -6, -7, -3, -5, 7, -4, 0, 5,
    -- filter=191 channel=103
    -16, -16, 12, -17, -9, 6, -16, -5, 13,
    -- filter=191 channel=104
    -1, -3, 16, -3, 11, 18, -18, -8, 19,
    -- filter=191 channel=105
    11, 12, -16, 7, 5, -7, 8, 6, -13,
    -- filter=191 channel=106
    -3, -2, 3, 8, 0, -4, 0, -3, -8,
    -- filter=191 channel=107
    11, -2, -20, 15, 7, -13, 11, 1, -21,
    -- filter=191 channel=108
    -5, -3, 2, 0, -8, -9, -2, -4, 6,
    -- filter=191 channel=109
    -12, 6, 1, -10, 9, -2, -6, 0, -1,
    -- filter=191 channel=110
    6, -3, 12, -3, 1, 12, -1, -3, 1,
    -- filter=191 channel=111
    -6, 0, 8, -5, 5, -3, 1, 6, -1,
    -- filter=191 channel=112
    -8, -6, -4, -12, -6, -2, -4, -6, -2,
    -- filter=191 channel=113
    -1, 0, 0, -11, -1, 11, -2, 2, -2,
    -- filter=191 channel=114
    -16, -11, -20, 2, -7, -31, 1, -5, -31,
    -- filter=191 channel=115
    -3, -2, 0, 0, 0, 4, 7, -4, 0,
    -- filter=191 channel=116
    -5, 10, -4, 3, 10, 10, -7, 4, 6,
    -- filter=191 channel=117
    1, 0, -3, -4, -3, -2, 5, -5, -5,
    -- filter=191 channel=118
    -5, 3, -2, -1, 0, -7, 1, -2, 5,
    -- filter=191 channel=119
    -4, 6, 4, 2, -3, 11, 2, 7, -1,
    -- filter=191 channel=120
    4, 5, -9, 12, 6, -5, -3, 6, -5,
    -- filter=191 channel=121
    0, 0, 1, -9, 9, 3, -7, -1, 7,
    -- filter=191 channel=122
    -16, -15, 28, -25, -2, 31, -28, -12, 17,
    -- filter=191 channel=123
    2, 2, 8, 7, -4, 3, 3, 3, 10,
    -- filter=191 channel=124
    1, 5, -6, 13, 6, -4, 6, 7, -3,
    -- filter=191 channel=125
    -9, 9, 15, -4, 14, 14, -8, 0, 15,
    -- filter=191 channel=126
    -8, 0, 0, -4, 3, -2, 2, 4, -2,
    -- filter=191 channel=127
    0, -3, 5, 1, -6, 3, 3, 2, 0,
    -- filter=192 channel=0
    -5, -3, 10, 2, 8, 9, 0, -8, 8,
    -- filter=192 channel=1
    1, 0, 1, 6, -2, 4, 2, -3, 4,
    -- filter=192 channel=2
    0, -5, 4, -5, 2, 6, 6, 0, -3,
    -- filter=192 channel=3
    6, 5, 1, 3, 6, 7, 10, 8, 15,
    -- filter=192 channel=4
    -7, 7, 1, 7, 6, 6, -2, -1, 7,
    -- filter=192 channel=5
    5, 0, 4, -4, -4, 3, -7, 3, 6,
    -- filter=192 channel=6
    -2, -6, 5, 1, 2, 8, 8, 5, 3,
    -- filter=192 channel=7
    4, 0, -1, 2, -6, -7, -3, -3, 1,
    -- filter=192 channel=8
    -6, -8, 4, -3, -1, -8, -5, 2, 4,
    -- filter=192 channel=9
    -5, 6, -4, -4, 6, -6, 0, -5, 1,
    -- filter=192 channel=10
    -5, 1, 1, -6, 5, -1, -3, -2, -12,
    -- filter=192 channel=11
    0, 2, -4, -3, 7, 6, 1, -6, -3,
    -- filter=192 channel=12
    -1, -4, -8, -2, -6, 0, 2, 4, 0,
    -- filter=192 channel=13
    4, -4, -3, 9, 12, 8, 5, -1, -9,
    -- filter=192 channel=14
    4, -2, 0, -4, -4, 4, -4, 1, -7,
    -- filter=192 channel=15
    -6, -10, -1, 5, 12, 11, -2, -7, -1,
    -- filter=192 channel=16
    8, -1, 3, 0, 7, -1, 5, 0, -4,
    -- filter=192 channel=17
    2, 7, -4, -2, -1, 3, -2, 0, -2,
    -- filter=192 channel=18
    -9, 0, -7, 11, 2, 6, 1, -3, -12,
    -- filter=192 channel=19
    -5, 5, 0, -6, 2, 7, 3, -3, 2,
    -- filter=192 channel=20
    1, 2, -2, 13, 15, 13, 1, 1, 2,
    -- filter=192 channel=21
    6, 10, 0, -3, -3, 4, 0, -5, -11,
    -- filter=192 channel=22
    1, 5, -5, 1, -1, 1, 7, 5, 1,
    -- filter=192 channel=23
    0, -14, 0, 15, 9, 5, -2, -4, -6,
    -- filter=192 channel=24
    5, 7, -3, -3, -5, -7, 5, -2, 1,
    -- filter=192 channel=25
    -6, 1, -4, -3, 9, 7, 1, -9, -16,
    -- filter=192 channel=26
    -6, 1, 3, 0, 6, -5, 0, 5, 5,
    -- filter=192 channel=27
    -4, -7, 3, 9, 9, 2, 0, -21, -20,
    -- filter=192 channel=28
    6, -6, 6, 0, -1, -6, -5, 3, -3,
    -- filter=192 channel=29
    -7, -3, -12, -3, 13, -2, -2, -7, -2,
    -- filter=192 channel=30
    1, 4, 10, 0, 1, 11, -5, -8, -12,
    -- filter=192 channel=31
    11, 0, 8, -2, 4, 5, -3, -8, -20,
    -- filter=192 channel=32
    4, -11, -10, 7, 12, 9, -4, -6, -6,
    -- filter=192 channel=33
    -4, 0, -7, -1, 1, 8, -4, 0, -5,
    -- filter=192 channel=34
    -5, -6, 8, 0, -4, 4, -9, -11, 1,
    -- filter=192 channel=35
    6, 0, 3, 0, 7, 7, -3, 4, -5,
    -- filter=192 channel=36
    -2, -3, 0, 6, 6, -8, -1, -7, -8,
    -- filter=192 channel=37
    3, -5, 3, 7, -6, -2, 2, 2, -1,
    -- filter=192 channel=38
    -5, -4, 1, 5, -2, 11, -4, 4, -10,
    -- filter=192 channel=39
    -6, 1, 0, -4, 8, 1, 5, -3, 4,
    -- filter=192 channel=40
    -1, 5, -6, 9, -1, 8, 9, 3, 3,
    -- filter=192 channel=41
    -6, 5, -13, -10, -12, -16, 0, -3, -4,
    -- filter=192 channel=42
    0, -2, -4, -5, 6, 3, -7, -9, -4,
    -- filter=192 channel=43
    -6, 0, -6, 1, 10, 6, 9, 10, 10,
    -- filter=192 channel=44
    2, 5, -1, 9, 1, 0, 0, -2, -1,
    -- filter=192 channel=45
    0, 4, 10, -3, 8, 5, -1, 1, 3,
    -- filter=192 channel=46
    0, -2, 1, -3, -3, 0, 3, 0, 5,
    -- filter=192 channel=47
    8, -2, 3, -4, -2, -4, 3, -1, -13,
    -- filter=192 channel=48
    0, -1, 0, 8, -3, 3, 0, -5, -15,
    -- filter=192 channel=49
    0, 0, -5, 4, 0, 3, -6, 0, 4,
    -- filter=192 channel=50
    10, -6, -1, -3, 0, 9, -3, -6, -15,
    -- filter=192 channel=51
    0, 0, -3, 5, -5, 7, -6, -5, 5,
    -- filter=192 channel=52
    2, -11, 1, 6, 4, 5, 1, -1, -2,
    -- filter=192 channel=53
    0, 0, 3, 0, -5, 3, -2, 0, -3,
    -- filter=192 channel=54
    2, 0, 0, 0, -4, 5, 5, 2, 2,
    -- filter=192 channel=55
    0, -2, -6, 0, 3, 6, -2, -9, -5,
    -- filter=192 channel=56
    5, 4, 0, 4, -7, 2, -4, 3, 5,
    -- filter=192 channel=57
    3, 1, -7, 5, -7, 3, 3, -2, 0,
    -- filter=192 channel=58
    4, 0, 1, 3, -5, 5, 5, -7, 9,
    -- filter=192 channel=59
    -5, 7, -1, 0, 2, 2, -8, 0, -14,
    -- filter=192 channel=60
    -7, -7, -6, 0, 1, -6, -1, -6, 7,
    -- filter=192 channel=61
    -2, 3, -2, -2, -2, -5, 6, -1, -2,
    -- filter=192 channel=62
    -2, 1, -2, -4, -5, -4, 7, 8, 7,
    -- filter=192 channel=63
    -7, 0, 4, 0, -1, 4, -5, -1, -2,
    -- filter=192 channel=64
    -3, 5, 7, 0, -4, -4, -6, 5, 5,
    -- filter=192 channel=65
    4, -7, -6, -2, 5, 2, -2, 6, -6,
    -- filter=192 channel=66
    -9, -1, -9, -9, -2, 0, 0, 3, -8,
    -- filter=192 channel=67
    2, -2, 7, -2, -5, 4, -3, 0, -4,
    -- filter=192 channel=68
    0, 5, 0, -6, 0, 2, -3, -1, -4,
    -- filter=192 channel=69
    6, 2, -4, 5, -8, -4, 3, 5, 0,
    -- filter=192 channel=70
    5, 1, 6, 2, 2, 6, 5, -2, -2,
    -- filter=192 channel=71
    0, 7, 4, 8, 10, 9, 0, 9, 10,
    -- filter=192 channel=72
    0, -1, -1, 5, 3, -5, -10, -12, -18,
    -- filter=192 channel=73
    -1, -4, -10, 3, 7, 6, -1, -3, -7,
    -- filter=192 channel=74
    0, -9, 7, 0, -7, 2, -1, -9, 0,
    -- filter=192 channel=75
    -1, -1, 3, 7, 3, 6, 5, -6, -3,
    -- filter=192 channel=76
    5, 1, -10, 10, 15, 14, 9, -1, 9,
    -- filter=192 channel=77
    6, -1, 7, 2, 5, 5, 0, -6, 5,
    -- filter=192 channel=78
    -1, 5, -1, -3, -6, -2, 4, -2, 1,
    -- filter=192 channel=79
    3, -2, -11, 11, 12, 4, 7, -5, -15,
    -- filter=192 channel=80
    1, -4, -2, 2, 1, 4, -1, -9, -18,
    -- filter=192 channel=81
    2, -2, 7, -7, 7, -4, -5, -6, -7,
    -- filter=192 channel=82
    -3, 0, -6, 0, -3, 8, -2, 4, -4,
    -- filter=192 channel=83
    5, 9, 4, 2, -3, -8, -4, 1, -4,
    -- filter=192 channel=84
    4, 0, 1, -3, 4, 0, -5, -6, -6,
    -- filter=192 channel=85
    3, 0, 6, 5, -3, -1, -6, 2, -5,
    -- filter=192 channel=86
    -4, -7, 2, -2, -8, -1, -8, -2, -6,
    -- filter=192 channel=87
    -8, 0, -4, 8, 1, 4, -2, -7, 5,
    -- filter=192 channel=88
    3, -3, 6, -1, 7, 3, 3, -6, 0,
    -- filter=192 channel=89
    5, -8, -10, 10, 9, 5, 2, -8, -18,
    -- filter=192 channel=90
    2, -1, 11, 5, 1, 2, 1, -4, 3,
    -- filter=192 channel=91
    1, -5, -3, 11, 10, 1, 2, -3, -4,
    -- filter=192 channel=92
    0, 0, 5, 0, -5, 8, -5, 0, 4,
    -- filter=192 channel=93
    7, -3, 7, 4, 4, -3, -8, -12, -10,
    -- filter=192 channel=94
    6, 1, -7, -1, 4, -2, 6, 6, 0,
    -- filter=192 channel=95
    3, -1, 0, -5, -1, -4, 1, 7, 4,
    -- filter=192 channel=96
    1, -3, 4, -5, 6, -6, 0, -2, 5,
    -- filter=192 channel=97
    1, -4, 2, 5, 10, 1, 0, 10, 6,
    -- filter=192 channel=98
    3, -6, -4, -1, 8, 8, -2, -2, -11,
    -- filter=192 channel=99
    5, -13, -8, -4, 3, -5, -6, -14, -12,
    -- filter=192 channel=100
    0, 2, -5, 1, -8, 3, -2, -8, -5,
    -- filter=192 channel=101
    -6, -2, -4, -5, 1, -4, 9, 0, 0,
    -- filter=192 channel=102
    6, 6, 0, -1, 0, -1, -6, -2, 2,
    -- filter=192 channel=103
    4, 6, 4, 2, 3, -3, -3, -6, -4,
    -- filter=192 channel=104
    8, 0, -5, 1, 5, 0, -9, -9, -17,
    -- filter=192 channel=105
    -3, -7, -8, 8, 10, 9, 0, -2, -3,
    -- filter=192 channel=106
    1, -2, 1, 5, 6, -2, 2, 4, 7,
    -- filter=192 channel=107
    5, -6, 0, 7, 5, 5, 0, 8, 5,
    -- filter=192 channel=108
    -1, -6, 5, 7, 1, -6, -5, 8, 3,
    -- filter=192 channel=109
    -6, -5, -1, -1, -2, 5, -1, -15, -14,
    -- filter=192 channel=110
    5, 3, 0, 2, 7, 1, -7, -3, -7,
    -- filter=192 channel=111
    0, -5, 6, 0, 3, -6, 7, -1, -4,
    -- filter=192 channel=112
    5, 0, 4, -5, 2, 0, -8, -10, -6,
    -- filter=192 channel=113
    2, 3, 0, -2, -1, 3, -5, -1, -10,
    -- filter=192 channel=114
    -5, -1, -2, 11, 1, 15, -1, -20, -15,
    -- filter=192 channel=115
    0, 6, 5, 0, -3, -7, 3, 7, 0,
    -- filter=192 channel=116
    8, 3, -8, 2, 0, -4, -8, -11, -15,
    -- filter=192 channel=117
    -3, -2, -1, 6, -5, 5, -3, -6, 4,
    -- filter=192 channel=118
    -1, -5, -2, 0, 0, -4, -3, -4, 7,
    -- filter=192 channel=119
    -3, -4, 5, 1, -8, -5, -11, -5, 3,
    -- filter=192 channel=120
    -5, -2, 5, 8, 5, -1, -9, -21, -18,
    -- filter=192 channel=121
    2, -5, -3, 0, -2, -4, -5, -2, 2,
    -- filter=192 channel=122
    3, 13, 17, 1, 4, -6, -5, -1, -14,
    -- filter=192 channel=123
    -5, -3, 1, 0, 2, -4, 1, -2, 6,
    -- filter=192 channel=124
    -1, -4, -5, 8, 6, 9, -3, -1, 1,
    -- filter=192 channel=125
    3, 4, -2, 7, 2, 0, -14, -10, -17,
    -- filter=192 channel=126
    -3, -11, -5, -5, 0, 8, 7, 2, 0,
    -- filter=192 channel=127
    6, 0, 4, -2, 0, -1, 1, -5, -7,
    -- filter=193 channel=0
    7, -3, -11, -4, 5, -11, -1, 5, 0,
    -- filter=193 channel=1
    -5, 0, -16, 2, 7, -5, 7, 17, 2,
    -- filter=193 channel=2
    -2, 0, -6, -6, 1, 6, -3, 0, 7,
    -- filter=193 channel=3
    -8, -13, -8, -5, 3, -5, -5, 2, 1,
    -- filter=193 channel=4
    -1, -4, -15, -7, -9, -2, 6, -7, 6,
    -- filter=193 channel=5
    10, 1, -16, 2, 6, -16, 0, 11, 0,
    -- filter=193 channel=6
    -4, -1, 0, -1, -5, 0, -8, -1, -5,
    -- filter=193 channel=7
    -2, 0, 1, -2, 1, 3, -7, 0, 1,
    -- filter=193 channel=8
    0, -4, 7, -4, 1, -5, 6, 0, 8,
    -- filter=193 channel=9
    -2, -1, 0, -3, -2, -3, -3, 1, -3,
    -- filter=193 channel=10
    -3, -4, 1, -4, -7, -1, 0, -7, -3,
    -- filter=193 channel=11
    -9, -4, 9, -13, -16, 1, 1, -5, -8,
    -- filter=193 channel=12
    1, -3, 1, -7, 0, 3, -2, 1, 1,
    -- filter=193 channel=13
    0, 5, 9, -4, 0, 13, -3, -7, -3,
    -- filter=193 channel=14
    -1, 0, -1, -2, 3, 3, -1, 0, 2,
    -- filter=193 channel=15
    0, 6, 4, -11, 1, 12, 3, 0, 7,
    -- filter=193 channel=16
    5, -1, -6, -3, 6, -3, 4, 2, -1,
    -- filter=193 channel=17
    5, 0, 2, -5, 6, 3, 6, 6, 2,
    -- filter=193 channel=18
    -1, 0, 1, -8, -4, 15, 1, 4, 6,
    -- filter=193 channel=19
    3, 6, -4, 6, -3, -7, 5, 0, -4,
    -- filter=193 channel=20
    -11, -3, 7, -12, -12, -4, -6, -15, -10,
    -- filter=193 channel=21
    -7, -1, -7, -3, -1, -9, -2, 1, 0,
    -- filter=193 channel=22
    4, 0, 5, -5, -2, 3, 0, 7, -1,
    -- filter=193 channel=23
    -10, 8, 11, -16, -1, 9, 0, -12, 14,
    -- filter=193 channel=24
    -4, -8, 6, -7, -4, -1, 5, 7, 0,
    -- filter=193 channel=25
    -7, 8, -4, -9, 0, -6, 0, 3, -1,
    -- filter=193 channel=26
    4, -7, -5, -3, 1, -9, 4, 5, 1,
    -- filter=193 channel=27
    -5, 4, 5, -1, 4, 8, 1, 0, 5,
    -- filter=193 channel=28
    2, -6, 3, 4, -5, -4, 3, -1, -5,
    -- filter=193 channel=29
    -13, -7, 8, -14, -12, 3, -1, -8, -7,
    -- filter=193 channel=30
    0, 0, -12, -3, 0, -4, 5, 0, -6,
    -- filter=193 channel=31
    -6, 10, 9, -12, 10, -5, -12, -10, 2,
    -- filter=193 channel=32
    -9, -3, 2, -2, 0, 11, 5, 0, -1,
    -- filter=193 channel=33
    -6, 11, -5, -6, 9, -1, 5, 8, 0,
    -- filter=193 channel=34
    7, 2, 11, 2, 13, -3, 8, 8, 4,
    -- filter=193 channel=35
    5, 6, 3, -4, 3, -6, 5, 2, -1,
    -- filter=193 channel=36
    -8, 2, 3, -3, -8, 2, 2, -5, -6,
    -- filter=193 channel=37
    -2, 5, -5, 4, 12, -10, 3, 20, 3,
    -- filter=193 channel=38
    3, -4, -3, 0, 0, -4, -3, -5, 4,
    -- filter=193 channel=39
    -7, 1, -1, -9, -2, -3, 0, -11, -2,
    -- filter=193 channel=40
    0, 7, 8, 5, 5, -4, 5, -8, 4,
    -- filter=193 channel=41
    -8, 7, 0, 3, 3, 11, 12, 8, -4,
    -- filter=193 channel=42
    0, 6, 4, -3, 7, 2, -3, -1, -3,
    -- filter=193 channel=43
    3, 0, 4, -4, 0, 7, 4, 2, 0,
    -- filter=193 channel=44
    0, 6, -2, -3, 2, -2, 4, 12, 0,
    -- filter=193 channel=45
    7, 0, -4, -3, 0, -3, -4, -3, -5,
    -- filter=193 channel=46
    1, 0, -7, 2, 2, -4, -3, 6, -6,
    -- filter=193 channel=47
    -3, 2, -8, 10, 3, -9, 1, 0, -3,
    -- filter=193 channel=48
    0, 6, -5, 3, 7, -9, 4, -6, 3,
    -- filter=193 channel=49
    0, -5, 2, -6, 4, 0, 0, -5, -4,
    -- filter=193 channel=50
    -2, 4, -1, 2, 9, 6, 4, 1, 0,
    -- filter=193 channel=51
    -4, 1, 2, -5, -2, 2, -7, 4, 7,
    -- filter=193 channel=52
    -2, -2, 9, -7, -4, -4, 1, -1, 8,
    -- filter=193 channel=53
    -4, 3, 3, -10, -11, 9, -2, -7, 0,
    -- filter=193 channel=54
    6, 4, -2, -3, 5, -4, -1, -6, -6,
    -- filter=193 channel=55
    -6, -3, 15, -17, -7, 8, -1, -14, 2,
    -- filter=193 channel=56
    5, -5, 5, -5, -4, 3, 1, -5, 0,
    -- filter=193 channel=57
    -4, -5, 7, 2, 3, 0, 3, -6, 0,
    -- filter=193 channel=58
    -3, -10, -11, -2, 2, -14, -4, 5, 0,
    -- filter=193 channel=59
    -7, 8, 6, 6, 6, 3, 1, 2, 1,
    -- filter=193 channel=60
    4, -1, 5, -6, 0, -2, -6, 3, 4,
    -- filter=193 channel=61
    0, 0, -7, 4, -4, -3, 7, -6, 5,
    -- filter=193 channel=62
    6, 2, 2, 2, 5, 6, -3, -6, 7,
    -- filter=193 channel=63
    -4, 0, -10, -2, -7, -14, -5, -6, -1,
    -- filter=193 channel=64
    -5, 4, -4, -4, -5, 7, -6, 2, 4,
    -- filter=193 channel=65
    -1, -6, 6, -4, 5, -3, 6, 6, -7,
    -- filter=193 channel=66
    -7, 0, -2, -5, 4, 8, 6, -4, -7,
    -- filter=193 channel=67
    0, 4, 6, -4, -5, 4, -4, 0, -1,
    -- filter=193 channel=68
    -7, -1, 1, -4, -5, -1, -6, 4, 0,
    -- filter=193 channel=69
    1, -6, -1, 0, 1, -4, 3, 2, -4,
    -- filter=193 channel=70
    8, 9, 0, 2, 9, 9, 4, 3, 9,
    -- filter=193 channel=71
    1, 5, -4, 0, 0, 3, 2, -1, -4,
    -- filter=193 channel=72
    -13, -1, 7, -11, -8, 9, -3, -15, -9,
    -- filter=193 channel=73
    -1, -2, 6, -2, -6, 0, -6, 2, 6,
    -- filter=193 channel=74
    0, 7, -5, -5, 5, -1, 5, 0, 0,
    -- filter=193 channel=75
    0, -4, -7, -2, 4, -14, 8, 13, -1,
    -- filter=193 channel=76
    2, 3, 2, -7, -3, 0, -5, -11, -1,
    -- filter=193 channel=77
    5, 3, 6, 1, -4, -2, -6, -6, 7,
    -- filter=193 channel=78
    -3, 0, -6, 3, 1, -11, 0, -4, -7,
    -- filter=193 channel=79
    -13, 10, 4, -8, 1, 17, 4, 1, 8,
    -- filter=193 channel=80
    -5, 3, -2, 0, -2, -2, 0, -8, -9,
    -- filter=193 channel=81
    -4, -3, -1, -1, -1, 6, -1, 3, -2,
    -- filter=193 channel=82
    7, -4, 1, -4, -2, -5, 1, -1, 5,
    -- filter=193 channel=83
    -6, 4, 0, 6, 0, -8, -3, -3, 0,
    -- filter=193 channel=84
    -8, 4, -5, -4, 5, 1, -5, -1, 5,
    -- filter=193 channel=85
    -2, 1, -3, 4, 0, -3, -6, -1, 0,
    -- filter=193 channel=86
    0, 0, 2, 0, 9, -4, -2, 0, 1,
    -- filter=193 channel=87
    3, -5, 5, -1, -3, 1, -6, -2, 6,
    -- filter=193 channel=88
    2, -1, 0, 1, -9, 1, -4, -11, 1,
    -- filter=193 channel=89
    -9, -2, 0, -1, -1, 3, 0, -10, -4,
    -- filter=193 channel=90
    2, -1, 5, -4, 0, -2, -4, -4, 5,
    -- filter=193 channel=91
    -4, -3, 0, -11, 5, 11, -6, -5, 3,
    -- filter=193 channel=92
    -1, 7, 3, -1, -2, 7, 1, 4, -5,
    -- filter=193 channel=93
    -5, 7, -4, 8, 2, -14, 0, 3, -1,
    -- filter=193 channel=94
    -4, -3, 3, 5, -1, -2, -6, -5, -4,
    -- filter=193 channel=95
    -3, 0, -5, 0, 2, 7, 5, 5, -5,
    -- filter=193 channel=96
    -5, -4, 7, 0, -4, 6, 1, -2, 5,
    -- filter=193 channel=97
    -4, -1, 1, -1, 2, -5, -3, 0, 0,
    -- filter=193 channel=98
    -7, -1, 5, -6, 6, 2, -9, -7, -2,
    -- filter=193 channel=99
    -1, 0, 1, -22, 0, 7, -3, -8, 3,
    -- filter=193 channel=100
    2, 0, 9, 4, 5, -3, 7, 6, 3,
    -- filter=193 channel=101
    0, -1, -7, -9, -2, -8, 6, -6, -4,
    -- filter=193 channel=102
    0, 4, -2, -6, 5, 3, 2, 1, 0,
    -- filter=193 channel=103
    8, 9, -3, 0, 4, -10, -7, -4, -2,
    -- filter=193 channel=104
    -4, 6, 3, 0, 1, -9, -7, -10, -11,
    -- filter=193 channel=105
    -4, -10, -1, 1, -5, 0, 3, -5, 0,
    -- filter=193 channel=106
    3, 2, 8, -6, -5, 5, 3, -5, 4,
    -- filter=193 channel=107
    4, -10, -2, 0, -7, 4, 5, -8, 3,
    -- filter=193 channel=108
    -2, 4, -3, -4, -7, -8, -6, 3, 0,
    -- filter=193 channel=109
    -9, 2, 6, 3, 4, 9, -1, 4, -4,
    -- filter=193 channel=110
    -6, 3, 8, -14, 0, -4, -4, -11, 1,
    -- filter=193 channel=111
    0, -2, 0, -1, -2, 1, -4, 0, -4,
    -- filter=193 channel=112
    7, 7, -5, -4, 7, -1, -3, 7, 7,
    -- filter=193 channel=113
    2, -1, 7, -1, 11, -2, 4, 8, 3,
    -- filter=193 channel=114
    0, 0, -6, -3, 1, 0, 5, 11, -7,
    -- filter=193 channel=115
    -1, -5, 2, 6, -7, 0, -3, -2, 5,
    -- filter=193 channel=116
    -13, -4, 5, -7, -9, 6, -5, -11, 3,
    -- filter=193 channel=117
    -2, 1, -6, -2, -5, -3, 0, -8, 6,
    -- filter=193 channel=118
    0, 1, 4, 0, 7, -5, -5, 5, 5,
    -- filter=193 channel=119
    6, 3, 2, 3, 5, 8, -3, 2, 6,
    -- filter=193 channel=120
    -12, -5, 9, -15, 4, -1, 2, -11, 4,
    -- filter=193 channel=121
    2, 8, 9, 2, -2, 3, 7, 4, -7,
    -- filter=193 channel=122
    0, 12, 1, 12, 13, -12, 4, -2, 1,
    -- filter=193 channel=123
    4, -3, 7, 0, 7, 4, -4, 7, -2,
    -- filter=193 channel=124
    3, 4, -5, -6, -11, -3, 0, -8, 3,
    -- filter=193 channel=125
    -4, 7, -3, -5, -1, 0, 0, -2, 2,
    -- filter=193 channel=126
    -5, 4, 6, 1, -10, -1, 3, -4, -9,
    -- filter=193 channel=127
    4, -4, 0, 5, 3, -6, 0, 8, 5,
    -- filter=194 channel=0
    0, 11, 10, -9, -8, -3, -17, -13, -8,
    -- filter=194 channel=1
    5, 5, 9, 1, -4, 2, -4, -10, -9,
    -- filter=194 channel=2
    4, 3, 0, 3, 4, -1, -3, 2, -5,
    -- filter=194 channel=3
    4, 4, 9, 5, -4, 6, 1, -1, -7,
    -- filter=194 channel=4
    2, 0, -8, 0, 2, 0, -3, -10, -6,
    -- filter=194 channel=5
    -5, 4, 2, -5, -1, -2, -10, -4, 4,
    -- filter=194 channel=6
    -1, -5, -7, -6, 1, -2, 7, 0, 1,
    -- filter=194 channel=7
    3, 0, -4, -5, 3, 5, 5, 2, 5,
    -- filter=194 channel=8
    0, -1, -2, 1, 4, 0, -7, -2, -6,
    -- filter=194 channel=9
    -1, -2, 3, -7, -3, -3, -8, -2, 6,
    -- filter=194 channel=10
    0, 8, -2, 8, 6, -4, -5, -3, 1,
    -- filter=194 channel=11
    6, -5, 0, 4, -7, -7, 6, 5, -3,
    -- filter=194 channel=12
    -7, 5, -3, 0, -3, -1, -2, -5, -4,
    -- filter=194 channel=13
    0, 5, -5, -3, -5, -8, 3, -7, 0,
    -- filter=194 channel=14
    5, -1, 2, 6, 4, 4, -7, 0, 5,
    -- filter=194 channel=15
    0, 4, -4, 1, -2, -3, -8, -2, -4,
    -- filter=194 channel=16
    -3, 0, 7, 0, 3, 7, 5, -2, 0,
    -- filter=194 channel=17
    2, -2, -2, 4, -3, 4, 6, -2, -6,
    -- filter=194 channel=18
    -2, -1, 5, -8, 0, -7, -12, -2, -4,
    -- filter=194 channel=19
    5, -3, -2, 1, -6, -2, 0, -5, -3,
    -- filter=194 channel=20
    2, 2, 0, 2, -2, 1, 10, 1, 9,
    -- filter=194 channel=21
    -4, -4, 1, 0, -2, -4, -5, 2, -2,
    -- filter=194 channel=22
    -1, -3, 9, 2, 2, 4, -7, 3, -6,
    -- filter=194 channel=23
    3, 0, 8, 6, -2, 10, -5, 1, 2,
    -- filter=194 channel=24
    -7, -2, 0, 0, 3, 6, -3, -2, 0,
    -- filter=194 channel=25
    -8, 3, 3, -9, -7, -1, -14, -3, 0,
    -- filter=194 channel=26
    -2, 3, 3, 0, 6, 3, 3, 6, 0,
    -- filter=194 channel=27
    5, 11, 7, 3, 1, 8, -16, -10, 2,
    -- filter=194 channel=28
    -4, 0, 6, 0, 2, 5, 6, 4, 3,
    -- filter=194 channel=29
    5, 0, -12, 6, -1, 1, 7, 4, -2,
    -- filter=194 channel=30
    3, -4, 0, 1, 0, 2, -13, 3, -7,
    -- filter=194 channel=31
    0, -5, -2, 9, -5, 9, 4, 10, 3,
    -- filter=194 channel=32
    0, 4, 5, -3, -3, -6, -11, -11, 2,
    -- filter=194 channel=33
    7, 4, 12, -8, -4, 0, -1, -7, -8,
    -- filter=194 channel=34
    -1, 0, 6, -5, -6, -1, -9, -1, 5,
    -- filter=194 channel=35
    -6, -6, 0, 2, 5, -4, -4, -2, 4,
    -- filter=194 channel=36
    1, -4, -1, 5, 7, -3, 1, 1, 0,
    -- filter=194 channel=37
    -6, 11, 9, -1, -4, 1, -16, -1, -10,
    -- filter=194 channel=38
    6, 9, 9, 6, 3, 0, -7, 2, 2,
    -- filter=194 channel=39
    1, 2, -6, 0, 0, -4, -3, 6, 0,
    -- filter=194 channel=40
    0, 1, -1, 3, 7, 4, 9, 0, -4,
    -- filter=194 channel=41
    -8, -5, -6, 3, -6, -2, 3, -7, -4,
    -- filter=194 channel=42
    0, -5, -3, 0, 5, 3, -5, -4, -5,
    -- filter=194 channel=43
    5, -2, -3, -2, 7, -5, -2, -2, -7,
    -- filter=194 channel=44
    4, -5, 8, 2, -6, -2, -9, -11, 1,
    -- filter=194 channel=45
    7, -3, 4, 0, 0, -4, 2, 1, 0,
    -- filter=194 channel=46
    7, -6, 0, 0, -6, 3, 0, 0, -4,
    -- filter=194 channel=47
    -5, 1, 1, 1, 6, -3, -6, 0, 1,
    -- filter=194 channel=48
    2, 0, 3, -9, 2, -3, -9, 2, 2,
    -- filter=194 channel=49
    -2, 1, -1, 2, -8, -4, -10, -10, -1,
    -- filter=194 channel=50
    3, 0, 1, 2, 2, 5, -4, -4, 7,
    -- filter=194 channel=51
    4, -1, -7, -1, -3, 1, 6, -5, 5,
    -- filter=194 channel=52
    6, -5, -4, -4, 5, -4, 0, 7, 7,
    -- filter=194 channel=53
    7, 3, -4, 3, -2, -4, -4, 1, 0,
    -- filter=194 channel=54
    7, 7, -2, -5, 5, 6, 3, 3, 1,
    -- filter=194 channel=55
    0, 9, -6, 5, -6, -4, 6, 3, 1,
    -- filter=194 channel=56
    -4, -4, 2, 4, -1, -2, 4, 4, -1,
    -- filter=194 channel=57
    -1, -7, 6, -1, 6, 4, 2, -8, 4,
    -- filter=194 channel=58
    -6, 9, 6, -3, 0, -2, -3, 0, -2,
    -- filter=194 channel=59
    5, 5, -2, 3, 0, -7, 2, -9, -5,
    -- filter=194 channel=60
    -1, -5, -2, -4, 7, -4, -1, -4, -5,
    -- filter=194 channel=61
    0, -5, -2, 4, -3, 4, 7, -4, -1,
    -- filter=194 channel=62
    4, -3, 0, -1, -5, 4, 4, 5, 5,
    -- filter=194 channel=63
    1, 0, -5, -6, 4, 5, -1, -7, -7,
    -- filter=194 channel=64
    3, -5, -2, 8, 2, 0, -3, -3, 2,
    -- filter=194 channel=65
    -6, 0, -3, -5, -3, -2, -3, 1, -4,
    -- filter=194 channel=66
    4, 4, -3, 2, -1, 0, -1, -6, -1,
    -- filter=194 channel=67
    -3, 0, 5, 3, -2, 0, -4, 2, 1,
    -- filter=194 channel=68
    -6, -2, -7, 7, -5, 5, -1, 2, 0,
    -- filter=194 channel=69
    1, 1, 4, -2, -5, 4, -1, 2, 5,
    -- filter=194 channel=70
    0, 9, 8, -4, 5, 7, -3, 3, -2,
    -- filter=194 channel=71
    2, 0, 9, 1, 6, -1, 2, 0, 2,
    -- filter=194 channel=72
    0, 2, -4, 2, 0, 6, 1, -3, -2,
    -- filter=194 channel=73
    2, -1, 0, 0, 1, 0, 3, -7, -2,
    -- filter=194 channel=74
    0, -3, 2, -2, 2, 2, -7, 3, -1,
    -- filter=194 channel=75
    6, 7, 12, 0, 4, 0, -10, -7, -4,
    -- filter=194 channel=76
    4, -5, -10, 11, -1, -8, 1, 6, -6,
    -- filter=194 channel=77
    -4, 1, 4, -1, 6, 7, -5, -6, -1,
    -- filter=194 channel=78
    4, -2, -1, -6, -1, 4, -5, 3, -2,
    -- filter=194 channel=79
    -3, 0, 7, -6, 3, 3, -7, -10, -1,
    -- filter=194 channel=80
    4, -4, -4, -1, -5, 6, -5, 1, 5,
    -- filter=194 channel=81
    -6, 5, 1, -6, -5, -4, -2, -6, -1,
    -- filter=194 channel=82
    0, 8, 7, 0, -4, 1, 8, 0, 7,
    -- filter=194 channel=83
    -3, 2, 1, -4, -2, 6, 0, -1, 4,
    -- filter=194 channel=84
    -4, 5, 3, -1, 0, 5, 0, -4, -4,
    -- filter=194 channel=85
    -4, 7, 0, -7, -4, 2, 1, 0, -2,
    -- filter=194 channel=86
    -3, 0, 7, -4, -7, -6, -5, 0, -3,
    -- filter=194 channel=87
    -5, 2, -8, 0, -3, -3, -2, 2, -2,
    -- filter=194 channel=88
    -5, 0, 4, 9, 2, 0, 3, 10, 0,
    -- filter=194 channel=89
    -2, 1, 0, 0, -2, -1, 2, -5, -10,
    -- filter=194 channel=90
    7, 1, -3, 9, 6, 10, 12, 10, 12,
    -- filter=194 channel=91
    2, 0, 0, -7, -1, 3, -5, 3, 0,
    -- filter=194 channel=92
    2, -1, 0, -3, -1, 7, -2, 3, -3,
    -- filter=194 channel=93
    -3, -4, -2, -2, -9, 3, -14, -10, -2,
    -- filter=194 channel=94
    -6, 0, -7, 7, 0, 0, 5, 0, 7,
    -- filter=194 channel=95
    1, -4, -5, -2, 4, 5, 0, -7, -6,
    -- filter=194 channel=96
    -2, 0, 6, 1, -5, -6, 3, 0, 0,
    -- filter=194 channel=97
    3, 8, 8, 0, 7, 5, 0, -4, -5,
    -- filter=194 channel=98
    -3, 11, 7, 2, -6, 4, -13, -11, -6,
    -- filter=194 channel=99
    -2, 1, 4, 2, 0, 3, -2, 0, 3,
    -- filter=194 channel=100
    -6, 2, -3, 6, 4, -2, 4, -1, 7,
    -- filter=194 channel=101
    0, 5, -4, 1, -6, 0, -4, 5, -8,
    -- filter=194 channel=102
    3, 3, 0, -2, -3, -2, 0, 4, 0,
    -- filter=194 channel=103
    -1, -2, -3, 3, 4, 5, -10, -5, -8,
    -- filter=194 channel=104
    5, 1, 0, 0, 0, 1, -8, 0, 0,
    -- filter=194 channel=105
    4, -8, -8, -1, 6, -7, 9, 8, 5,
    -- filter=194 channel=106
    4, 7, -3, 0, 0, -5, 4, 0, 5,
    -- filter=194 channel=107
    7, 0, 3, 6, -1, 2, -1, 9, -5,
    -- filter=194 channel=108
    1, 2, -4, 2, -4, 0, 0, 4, -1,
    -- filter=194 channel=109
    0, 0, -1, -3, -3, -3, -14, -7, 3,
    -- filter=194 channel=110
    -4, 7, 0, 9, 6, 3, -2, 8, 4,
    -- filter=194 channel=111
    -5, -7, -1, -6, 1, 5, 0, -4, 6,
    -- filter=194 channel=112
    -4, 3, 1, 2, 1, 0, -4, -3, -3,
    -- filter=194 channel=113
    -1, 4, 8, 8, -4, 0, 3, 6, -4,
    -- filter=194 channel=114
    -6, 1, 2, -10, -12, -4, -18, -8, 0,
    -- filter=194 channel=115
    1, -5, 4, -7, 0, -2, -1, -6, 5,
    -- filter=194 channel=116
    -8, -3, -4, -2, -1, 1, 0, 4, -2,
    -- filter=194 channel=117
    5, -2, 5, 4, -3, 3, 3, -4, 1,
    -- filter=194 channel=118
    -5, -2, 0, -6, -3, 4, 4, -2, 1,
    -- filter=194 channel=119
    0, 0, 4, 0, 0, 0, 2, 5, 11,
    -- filter=194 channel=120
    9, 9, 8, 7, -2, 2, -4, -3, 3,
    -- filter=194 channel=121
    -2, -1, 0, 0, 7, -3, 0, 0, -8,
    -- filter=194 channel=122
    5, -3, -2, 7, -3, -4, 0, 2, 4,
    -- filter=194 channel=123
    -1, 3, 2, 1, 0, -4, 0, 3, 1,
    -- filter=194 channel=124
    -2, -7, -7, -2, 5, 1, 8, 5, -2,
    -- filter=194 channel=125
    0, -7, -6, -7, -8, -4, -8, -3, 5,
    -- filter=194 channel=126
    4, 6, 2, -6, 0, -1, -4, -8, -6,
    -- filter=194 channel=127
    4, -1, 0, 3, -7, -4, 4, -3, 6,
    -- filter=195 channel=0
    6, 24, 20, -2, 26, 14, -9, -2, -11,
    -- filter=195 channel=1
    10, 22, 11, -2, 9, 11, -8, 4, 0,
    -- filter=195 channel=2
    -3, 2, 1, 0, -4, 4, 8, -3, -4,
    -- filter=195 channel=3
    -4, 0, 4, 1, 10, -5, -9, -4, -3,
    -- filter=195 channel=4
    7, -10, -7, 0, 7, 11, 5, 0, 6,
    -- filter=195 channel=5
    2, 22, 13, 4, 20, 4, 3, 9, -4,
    -- filter=195 channel=6
    5, 0, 1, 2, -1, 1, 5, -4, -6,
    -- filter=195 channel=7
    6, 5, 3, -4, 5, -2, 6, 1, -4,
    -- filter=195 channel=8
    1, 3, -3, -2, 3, 4, 3, 0, 2,
    -- filter=195 channel=9
    -5, -6, 2, -4, -10, -3, -5, -6, 4,
    -- filter=195 channel=10
    -6, 0, -7, 1, -9, -8, -3, 0, 3,
    -- filter=195 channel=11
    3, 2, 0, 4, 5, -2, -2, -5, 4,
    -- filter=195 channel=12
    -3, -3, -6, 1, 0, 0, 4, 6, 0,
    -- filter=195 channel=13
    -1, -5, -3, 6, -6, -6, 3, -5, 9,
    -- filter=195 channel=14
    -2, -3, 0, 6, 1, -4, -2, -3, -4,
    -- filter=195 channel=15
    6, 8, -2, -1, 2, 1, -3, 0, -3,
    -- filter=195 channel=16
    -4, -11, 2, -1, -9, -9, -5, -9, 4,
    -- filter=195 channel=17
    -1, 4, 0, 0, -1, 0, -2, 4, -4,
    -- filter=195 channel=18
    1, 8, 6, 1, 11, -3, -1, 7, 12,
    -- filter=195 channel=19
    -1, 0, 2, 3, -6, -5, 6, -1, -4,
    -- filter=195 channel=20
    -3, -1, -3, 6, 7, 1, -1, 4, 4,
    -- filter=195 channel=21
    -3, -7, -8, -5, -8, -8, -11, -10, -8,
    -- filter=195 channel=22
    8, 1, 7, -3, 13, -2, -8, 8, -1,
    -- filter=195 channel=23
    -6, 1, -2, 6, -9, -6, -6, -4, 4,
    -- filter=195 channel=24
    7, -2, 0, -4, 0, 2, 4, -1, 0,
    -- filter=195 channel=25
    -4, -8, -6, -1, -11, -2, 7, 2, 10,
    -- filter=195 channel=26
    3, 3, 0, -2, -4, -5, 2, 2, -3,
    -- filter=195 channel=27
    0, 0, -9, -11, 4, 4, 2, 10, 7,
    -- filter=195 channel=28
    0, -5, -2, 6, 4, -6, 5, -5, -7,
    -- filter=195 channel=29
    -4, 5, -7, -4, -1, -6, -7, 6, 8,
    -- filter=195 channel=30
    -4, 8, -4, -3, 5, 7, -5, -1, 1,
    -- filter=195 channel=31
    -4, -18, -12, -14, -17, -8, 4, 0, 1,
    -- filter=195 channel=32
    6, 3, -6, 7, 3, 0, -2, -2, 6,
    -- filter=195 channel=33
    -4, 10, 7, 0, 5, -9, -11, -7, 4,
    -- filter=195 channel=34
    7, 1, -7, 0, 6, 0, 8, 9, -6,
    -- filter=195 channel=35
    0, 1, 1, 4, -3, 4, 1, -6, -3,
    -- filter=195 channel=36
    7, -6, -7, 0, 0, -1, 1, -6, 0,
    -- filter=195 channel=37
    9, 18, 9, -7, 13, 0, -5, -3, -10,
    -- filter=195 channel=38
    -5, 4, -7, -7, 3, 1, -3, 3, 0,
    -- filter=195 channel=39
    3, -5, -1, 0, -7, -6, -1, -7, -3,
    -- filter=195 channel=40
    0, -7, 0, -8, -1, -1, 2, -8, 4,
    -- filter=195 channel=41
    0, -2, -6, 13, -8, -5, 2, -3, -7,
    -- filter=195 channel=42
    -8, -4, 7, -3, -1, -1, -7, 2, -7,
    -- filter=195 channel=43
    -1, 7, 6, 10, 5, 5, -11, -5, 2,
    -- filter=195 channel=44
    2, -5, -8, 0, -6, 2, -10, -7, 0,
    -- filter=195 channel=45
    4, 8, 3, -3, 9, -4, 4, 3, -6,
    -- filter=195 channel=46
    2, 8, 1, 4, 10, -4, -5, 7, -2,
    -- filter=195 channel=47
    -13, -3, -3, -9, -15, -8, -10, -12, 0,
    -- filter=195 channel=48
    1, -2, 0, -15, -4, 0, 0, 2, -3,
    -- filter=195 channel=49
    6, 5, -8, -5, 4, 7, -2, 0, 9,
    -- filter=195 channel=50
    -8, -7, 3, -8, -8, -3, -2, 0, 1,
    -- filter=195 channel=51
    6, 6, -7, 5, 1, 0, -1, -4, 0,
    -- filter=195 channel=52
    -1, 0, -8, 3, -2, -6, 9, 3, 3,
    -- filter=195 channel=53
    -6, -5, -6, -4, 7, -6, 2, 7, 3,
    -- filter=195 channel=54
    7, 2, 0, -2, -1, -1, 1, 6, 2,
    -- filter=195 channel=55
    2, 5, -11, 6, -2, -8, 4, 8, 13,
    -- filter=195 channel=56
    -3, -6, 0, 8, 5, -4, -1, 0, -8,
    -- filter=195 channel=57
    7, -4, -8, 1, 2, -2, 2, 0, 4,
    -- filter=195 channel=58
    7, 13, 15, 4, 13, 6, 1, 8, 0,
    -- filter=195 channel=59
    2, -1, -7, -3, -15, -6, 5, -10, -4,
    -- filter=195 channel=60
    -5, -5, -5, 7, -6, -2, 0, -4, 3,
    -- filter=195 channel=61
    5, 1, -9, 1, -3, -4, -1, 2, -6,
    -- filter=195 channel=62
    6, -6, -1, 3, 7, 1, -7, 1, 0,
    -- filter=195 channel=63
    0, 10, 10, 5, 5, 9, 5, 3, -3,
    -- filter=195 channel=64
    4, -2, -7, -6, -3, -2, 4, 0, -5,
    -- filter=195 channel=65
    -7, -1, 1, -3, -3, 5, -4, 4, 0,
    -- filter=195 channel=66
    7, -8, -9, 8, -9, 0, -2, -4, -6,
    -- filter=195 channel=67
    -2, -3, 4, 0, -4, -7, 2, 0, -5,
    -- filter=195 channel=68
    0, -4, -3, 0, 0, 4, 3, -1, 2,
    -- filter=195 channel=69
    4, -5, -5, 5, 2, -1, 4, 3, 7,
    -- filter=195 channel=70
    6, -4, -8, -7, -2, 5, -8, 9, 2,
    -- filter=195 channel=71
    -9, -9, -1, -6, -8, -4, 0, -4, -3,
    -- filter=195 channel=72
    0, -10, -7, -9, -7, -9, -4, 2, 8,
    -- filter=195 channel=73
    -2, 3, -5, 3, -7, -3, 7, 6, 1,
    -- filter=195 channel=74
    5, 1, -2, -3, -7, 2, 2, 0, -4,
    -- filter=195 channel=75
    3, 11, 17, -4, 15, -2, -2, 3, -9,
    -- filter=195 channel=76
    -5, 3, -10, 7, -3, -7, -1, -6, 2,
    -- filter=195 channel=77
    6, 4, -3, 2, -4, -5, 0, -2, 6,
    -- filter=195 channel=78
    -6, 3, -2, 5, 8, -2, 1, -6, 0,
    -- filter=195 channel=79
    11, 17, 1, -2, 15, 2, -13, 10, 12,
    -- filter=195 channel=80
    -10, -15, -1, -15, -15, 0, 2, -9, 3,
    -- filter=195 channel=81
    -3, 5, 4, -5, 1, -4, 0, -4, 2,
    -- filter=195 channel=82
    2, -1, 7, 1, 5, -7, 2, -7, 5,
    -- filter=195 channel=83
    -4, 3, 4, -7, -11, -4, 4, 6, -4,
    -- filter=195 channel=84
    -3, 4, -5, 1, 5, 0, 0, 0, 5,
    -- filter=195 channel=85
    2, 3, -3, 5, 5, 2, 4, -6, 4,
    -- filter=195 channel=86
    11, 3, 3, 7, 10, 7, -2, -1, 2,
    -- filter=195 channel=87
    4, -4, 0, 10, 4, 5, 3, -4, -2,
    -- filter=195 channel=88
    -5, -7, -5, 3, -5, -9, -2, 0, 3,
    -- filter=195 channel=89
    0, -8, 2, -8, -14, -3, 0, 1, -1,
    -- filter=195 channel=90
    2, -8, -8, -5, -14, -5, -1, -8, 3,
    -- filter=195 channel=91
    0, 4, -11, -4, 1, 7, 3, 7, 9,
    -- filter=195 channel=92
    1, -5, -7, -1, 0, -3, 6, 4, 5,
    -- filter=195 channel=93
    -8, 5, -3, -2, 6, -4, -9, 3, 5,
    -- filter=195 channel=94
    6, 0, -3, -5, -4, -6, 2, -5, -2,
    -- filter=195 channel=95
    -4, 7, -6, -6, -1, -3, 6, 0, 3,
    -- filter=195 channel=96
    4, -2, 6, 1, -7, 1, -5, -4, -1,
    -- filter=195 channel=97
    3, 0, 7, 3, -4, -3, 3, -7, -5,
    -- filter=195 channel=98
    -6, -3, 0, -10, -9, -6, 4, 5, 10,
    -- filter=195 channel=99
    -2, -12, -6, -4, -14, -5, 3, 0, 10,
    -- filter=195 channel=100
    5, 7, 3, 6, 9, -3, -1, -3, -1,
    -- filter=195 channel=101
    -3, -11, -2, -3, 3, 2, 3, 3, -3,
    -- filter=195 channel=102
    4, 2, 4, -2, -6, 7, -5, -5, 0,
    -- filter=195 channel=103
    -10, -7, -4, -2, -2, -5, -15, -4, -4,
    -- filter=195 channel=104
    -6, -10, 1, -6, -11, -7, -1, -2, -3,
    -- filter=195 channel=105
    8, 2, -4, 6, 5, -4, -5, 6, 4,
    -- filter=195 channel=106
    2, 0, -1, -6, -2, -3, -5, 2, -7,
    -- filter=195 channel=107
    7, 8, -5, -3, 13, 2, -12, 6, 2,
    -- filter=195 channel=108
    5, 7, 5, 4, 6, -2, -4, -4, -4,
    -- filter=195 channel=109
    4, 3, -3, 3, -2, 0, 1, 10, 14,
    -- filter=195 channel=110
    -5, 2, -6, 6, -1, -5, 7, -9, 7,
    -- filter=195 channel=111
    1, 4, -7, 7, 0, -7, 8, 7, 1,
    -- filter=195 channel=112
    0, 3, -4, -8, 7, 4, 6, -1, -3,
    -- filter=195 channel=113
    -6, 0, -1, 4, 0, -4, -5, -11, 3,
    -- filter=195 channel=114
    9, 22, 9, 7, 22, 4, -5, 16, 6,
    -- filter=195 channel=115
    3, 0, 0, -4, -5, -1, 3, -4, 7,
    -- filter=195 channel=116
    8, -5, -8, -11, -9, 2, 6, 5, 8,
    -- filter=195 channel=117
    -3, 0, -1, 1, -5, 2, -5, 4, 2,
    -- filter=195 channel=118
    -1, -3, -2, 4, -2, -8, -3, -3, -5,
    -- filter=195 channel=119
    2, -6, -1, 9, 4, -3, 8, 5, -8,
    -- filter=195 channel=120
    -2, 3, -5, -4, 0, -7, 4, 2, 7,
    -- filter=195 channel=121
    -4, -3, -2, 5, -9, 3, -3, -7, 2,
    -- filter=195 channel=122
    -24, -27, -14, -15, -29, -16, -14, -22, -4,
    -- filter=195 channel=123
    3, -5, -3, -2, 1, -4, 6, -4, -2,
    -- filter=195 channel=124
    0, 2, -4, 0, 8, -3, -10, -1, 2,
    -- filter=195 channel=125
    -6, -9, -3, -10, -6, 0, 0, 4, 8,
    -- filter=195 channel=126
    -6, 4, -5, 5, 1, 2, -9, -6, 7,
    -- filter=195 channel=127
    -6, 1, -4, 3, -4, -3, -5, -2, 5,
    -- filter=196 channel=0
    4, -9, 2, 9, -2, 2, 27, 13, 7,
    -- filter=196 channel=1
    -7, 7, 6, -3, -1, 12, -1, -6, 4,
    -- filter=196 channel=2
    3, 3, 0, -5, -8, -10, -3, -14, -6,
    -- filter=196 channel=3
    0, -26, -13, -22, -25, -2, -14, 1, 3,
    -- filter=196 channel=4
    -10, -18, -3, -22, -32, -12, -26, -29, -14,
    -- filter=196 channel=5
    -8, 0, 0, 0, -1, 1, 3, -1, 0,
    -- filter=196 channel=6
    6, 5, -5, 0, -10, -5, -2, -3, 0,
    -- filter=196 channel=7
    -4, 3, -2, 6, 5, 3, 4, 7, 0,
    -- filter=196 channel=8
    1, -7, 1, -15, -14, -7, -1, -4, 0,
    -- filter=196 channel=9
    6, 7, -1, 0, 15, 4, 4, 1, 0,
    -- filter=196 channel=10
    -2, 5, -7, 2, 0, 1, -15, -8, -5,
    -- filter=196 channel=11
    8, 6, 4, 7, 10, 2, 6, 14, -1,
    -- filter=196 channel=12
    -14, -16, 1, -2, -7, -10, -3, -17, -8,
    -- filter=196 channel=13
    -4, -6, -6, -9, -16, 6, -5, -10, 6,
    -- filter=196 channel=14
    3, -4, 6, -4, -3, 0, 4, 3, 2,
    -- filter=196 channel=15
    16, -3, -4, 4, 0, 0, 2, 4, 5,
    -- filter=196 channel=16
    -19, -6, -2, -7, 6, 8, -17, -3, -2,
    -- filter=196 channel=17
    6, -6, 1, -6, 0, 4, -6, -4, 6,
    -- filter=196 channel=18
    3, -8, 0, 8, -17, -3, 4, -1, 6,
    -- filter=196 channel=19
    5, -1, 6, 0, -7, 3, 3, -2, 0,
    -- filter=196 channel=20
    11, 5, 0, 6, 3, 6, 11, 8, 7,
    -- filter=196 channel=21
    -8, 19, 15, 4, 27, 9, -5, 0, -4,
    -- filter=196 channel=22
    4, -9, -4, 4, -11, -5, 0, 6, 1,
    -- filter=196 channel=23
    8, -4, 0, 8, -7, -5, 0, 12, 1,
    -- filter=196 channel=24
    7, -6, 0, 0, -1, -1, -4, -7, -1,
    -- filter=196 channel=25
    -7, 6, 0, -2, 2, -1, -8, -7, 0,
    -- filter=196 channel=26
    3, 4, 5, -8, 2, 4, -7, -12, -10,
    -- filter=196 channel=27
    11, 8, -2, 2, 8, -5, -7, 6, 2,
    -- filter=196 channel=28
    6, 6, 6, 2, -6, 6, 6, -5, -6,
    -- filter=196 channel=29
    4, 6, -11, 0, 0, -3, 0, 10, -6,
    -- filter=196 channel=30
    -4, 8, 0, 6, 9, 0, 4, -3, -1,
    -- filter=196 channel=31
    4, 12, 8, -3, 34, 10, -15, 8, -13,
    -- filter=196 channel=32
    9, 2, -10, -5, -15, -5, -1, -9, 0,
    -- filter=196 channel=33
    -4, 4, -2, 2, 7, -2, -2, 0, 0,
    -- filter=196 channel=34
    -5, -19, -12, -6, -22, -15, -19, -22, 1,
    -- filter=196 channel=35
    3, 0, -3, -5, 6, 0, -2, 7, 4,
    -- filter=196 channel=36
    7, 4, 1, 3, 4, -6, -2, -7, 0,
    -- filter=196 channel=37
    -4, 3, 1, 4, 1, 8, 7, -1, 6,
    -- filter=196 channel=38
    2, 11, 3, 3, 14, -3, 3, 7, 8,
    -- filter=196 channel=39
    9, -3, 1, 0, 5, 2, 0, 9, 4,
    -- filter=196 channel=40
    13, 1, 7, 7, 2, 0, 7, 13, 12,
    -- filter=196 channel=41
    -17, -22, 0, -27, -47, -6, -28, -51, -4,
    -- filter=196 channel=42
    2, 9, 3, 3, 10, 0, 9, 2, 5,
    -- filter=196 channel=43
    2, -9, -6, -4, -20, -15, 0, 6, 0,
    -- filter=196 channel=44
    0, 9, 2, -2, 14, 11, -4, -3, -5,
    -- filter=196 channel=45
    11, 6, 7, 14, 13, 10, 14, 10, 8,
    -- filter=196 channel=46
    1, 0, -6, -3, -5, 5, -1, 2, 3,
    -- filter=196 channel=47
    -10, 12, 7, -4, 23, 8, -15, 0, 0,
    -- filter=196 channel=48
    5, 15, 0, -3, 12, 9, -9, -4, -12,
    -- filter=196 channel=49
    9, 9, -5, -6, -9, -2, -2, 4, 0,
    -- filter=196 channel=50
    7, 15, -4, 13, 21, 0, 11, 11, 5,
    -- filter=196 channel=51
    5, 6, -2, 5, -5, 2, 4, 4, 6,
    -- filter=196 channel=52
    -3, -15, -4, -11, -16, -8, -10, -15, -3,
    -- filter=196 channel=53
    -6, -5, -6, 2, -7, 3, -7, -1, 6,
    -- filter=196 channel=54
    0, -2, -1, 0, -2, 6, 0, 7, 2,
    -- filter=196 channel=55
    13, -4, -5, 0, -5, -9, 7, 3, 4,
    -- filter=196 channel=56
    4, -6, -5, -7, -18, -5, -6, -14, -4,
    -- filter=196 channel=57
    -8, 2, 4, -4, -5, 1, -11, -13, -6,
    -- filter=196 channel=58
    -3, 0, -7, 5, -9, 2, 4, 0, 3,
    -- filter=196 channel=59
    -2, 4, 1, 2, 7, 8, -5, -3, 2,
    -- filter=196 channel=60
    1, 4, 6, -1, 2, -7, 7, -1, -6,
    -- filter=196 channel=61
    2, 1, -5, -7, 0, -1, -13, -10, -1,
    -- filter=196 channel=62
    5, 6, 3, 3, -7, -5, -2, -4, 2,
    -- filter=196 channel=63
    -4, -5, 5, -6, 0, 4, 0, -3, -2,
    -- filter=196 channel=64
    -5, 7, -1, 1, 0, -7, 4, 2, 3,
    -- filter=196 channel=65
    3, -3, -3, 1, 0, 0, -4, -2, -4,
    -- filter=196 channel=66
    -18, -16, -4, -5, -24, 3, -18, -23, -7,
    -- filter=196 channel=67
    7, -3, 4, 8, -7, -2, -3, 4, 4,
    -- filter=196 channel=68
    4, -4, -4, 1, -2, 4, -6, -7, -6,
    -- filter=196 channel=69
    -5, 1, 1, 0, -6, 8, -2, -7, -6,
    -- filter=196 channel=70
    5, -4, -13, 7, -2, -1, 6, 6, -3,
    -- filter=196 channel=71
    1, 1, 6, 0, 0, 9, -9, 0, -1,
    -- filter=196 channel=72
    5, 14, 0, 6, 30, -1, -5, 0, -3,
    -- filter=196 channel=73
    -2, -1, -1, -3, -5, -3, 3, -4, -4,
    -- filter=196 channel=74
    -1, 1, -4, 4, -3, -6, -7, 1, 3,
    -- filter=196 channel=75
    -9, 6, 0, 7, -10, 8, 9, 0, 2,
    -- filter=196 channel=76
    5, 4, 0, 2, 4, -2, 16, 16, 5,
    -- filter=196 channel=77
    4, 3, 0, -8, -7, -3, 3, -3, -4,
    -- filter=196 channel=78
    0, -2, 5, 5, -5, -6, 0, -8, -11,
    -- filter=196 channel=79
    0, -10, 0, 0, -11, -5, 0, 6, 6,
    -- filter=196 channel=80
    2, 20, 11, 6, 32, 13, -6, -3, -13,
    -- filter=196 channel=81
    -2, 2, -5, 0, -5, -6, -2, 6, -4,
    -- filter=196 channel=82
    1, 1, 0, 0, 6, 7, 7, 0, 6,
    -- filter=196 channel=83
    10, 14, 6, 3, 5, 0, 3, 6, 4,
    -- filter=196 channel=84
    8, -5, 2, -7, -5, -8, 0, -13, -7,
    -- filter=196 channel=85
    -2, 2, -6, 4, -2, -4, 1, 1, 2,
    -- filter=196 channel=86
    -3, -5, 2, -11, -6, -4, 1, -6, -1,
    -- filter=196 channel=87
    2, -7, 0, -6, -17, -7, -6, -14, -9,
    -- filter=196 channel=88
    3, 11, 0, -2, 5, -6, 5, 0, -6,
    -- filter=196 channel=89
    -3, 8, 3, -4, 2, 2, -4, 3, -3,
    -- filter=196 channel=90
    -5, 0, 0, 2, 8, -5, -14, -6, -6,
    -- filter=196 channel=91
    0, 13, 2, 1, 5, -4, 2, -5, 5,
    -- filter=196 channel=92
    -3, -3, -8, -5, -17, -11, -5, -6, -8,
    -- filter=196 channel=93
    -5, 14, 7, -10, 8, 6, -11, -8, -2,
    -- filter=196 channel=94
    -3, -7, 2, 0, 4, -2, 3, 3, 0,
    -- filter=196 channel=95
    -3, -1, -1, -12, -3, -6, -8, -7, -6,
    -- filter=196 channel=96
    4, 7, -5, 1, 9, 5, 6, -3, 0,
    -- filter=196 channel=97
    5, -9, -5, -1, 1, 7, 2, 0, 3,
    -- filter=196 channel=98
    -3, -1, -4, -4, 8, 0, -5, 0, -1,
    -- filter=196 channel=99
    7, 1, 0, 0, 12, -8, -17, -14, -2,
    -- filter=196 channel=100
    -2, -5, -5, 0, -7, -8, -5, -7, -14,
    -- filter=196 channel=101
    -10, -3, -4, -21, -11, -9, -19, -14, -11,
    -- filter=196 channel=102
    -2, 5, -3, -6, 0, 3, -5, 6, 1,
    -- filter=196 channel=103
    -3, 6, 4, 3, 28, 7, -4, -2, -5,
    -- filter=196 channel=104
    -1, 8, 8, 1, 30, 7, -13, 3, -13,
    -- filter=196 channel=105
    9, 2, 0, 0, -2, -7, 6, -1, 1,
    -- filter=196 channel=106
    10, 0, 1, 5, 6, 4, 10, 7, -4,
    -- filter=196 channel=107
    8, -7, -1, -1, -9, 5, 18, 9, 5,
    -- filter=196 channel=108
    -9, -9, -2, 0, -14, 3, 1, -3, -1,
    -- filter=196 channel=109
    -7, 1, -1, -8, -3, -1, -19, -3, -9,
    -- filter=196 channel=110
    0, 2, -2, -8, 0, 3, -4, -5, -2,
    -- filter=196 channel=111
    -4, 5, -1, 4, -7, 5, -4, 0, -2,
    -- filter=196 channel=112
    3, 4, -7, 5, 0, -7, 2, -1, 9,
    -- filter=196 channel=113
    -3, -3, 1, 1, 11, 5, 0, -5, -7,
    -- filter=196 channel=114
    14, -7, -6, 2, -13, -16, 17, -7, 0,
    -- filter=196 channel=115
    2, 3, 2, -5, -2, 2, 5, 3, 4,
    -- filter=196 channel=116
    -3, 13, 0, 2, 9, 1, -9, 2, -3,
    -- filter=196 channel=117
    -5, 2, 7, -1, 9, 5, -2, 7, 0,
    -- filter=196 channel=118
    3, 0, -5, 0, 4, 3, 0, 1, -1,
    -- filter=196 channel=119
    -5, -12, -2, -6, -28, -11, -20, -26, -6,
    -- filter=196 channel=120
    13, 13, 5, 4, 0, 7, 0, 9, -2,
    -- filter=196 channel=121
    -3, 2, -5, -8, -5, 5, -9, -15, -10,
    -- filter=196 channel=122
    -15, 24, 16, -4, 22, 23, -33, -10, -2,
    -- filter=196 channel=123
    0, -9, -9, -12, -5, 0, -13, -13, 0,
    -- filter=196 channel=124
    -2, -3, -2, -1, 2, -7, 6, 8, 6,
    -- filter=196 channel=125
    -5, 16, 6, -9, 12, 6, -16, -8, -6,
    -- filter=196 channel=126
    -5, 1, 6, -7, -15, 3, -3, -9, -4,
    -- filter=196 channel=127
    -2, 1, 0, -11, -12, 4, 1, -11, -2,
    -- filter=197 channel=0
    -5, 14, 9, 5, 16, 2, -3, 1, 0,
    -- filter=197 channel=1
    0, 1, 8, 5, 13, -2, 6, 5, -3,
    -- filter=197 channel=2
    0, 3, 0, 6, -5, 3, 1, 0, -1,
    -- filter=197 channel=3
    5, 2, 3, 4, 3, 8, 2, 6, 0,
    -- filter=197 channel=4
    -3, 0, 1, 5, 1, 8, 1, 10, 0,
    -- filter=197 channel=5
    -1, 6, 1, 1, 3, 2, 5, 7, 1,
    -- filter=197 channel=6
    -2, -7, 5, 4, 3, -5, -5, 2, -2,
    -- filter=197 channel=7
    0, 1, -1, 0, -3, 3, 4, 2, -5,
    -- filter=197 channel=8
    6, 4, -6, -1, 3, -1, 4, 0, -4,
    -- filter=197 channel=9
    7, 0, 1, -3, -2, 0, -3, 4, 7,
    -- filter=197 channel=10
    5, -7, 5, -1, 4, 5, -1, 1, -2,
    -- filter=197 channel=11
    5, -7, -3, 5, 5, -3, 4, 1, 3,
    -- filter=197 channel=12
    -4, 6, 1, -2, -5, 4, 0, 3, 1,
    -- filter=197 channel=13
    4, -8, -7, 0, 0, -6, 4, 0, -2,
    -- filter=197 channel=14
    -1, 0, 4, 2, -5, 0, -4, 6, 0,
    -- filter=197 channel=15
    2, -6, -1, -4, 2, 0, -5, -4, 4,
    -- filter=197 channel=16
    6, 0, 2, 2, 3, -7, 6, -4, 2,
    -- filter=197 channel=17
    3, -2, 2, 7, -1, 5, -6, -2, -3,
    -- filter=197 channel=18
    0, -3, 0, 7, 0, -8, 5, 0, 0,
    -- filter=197 channel=19
    6, -6, 0, 4, -6, -5, -7, -6, 5,
    -- filter=197 channel=20
    -6, -2, 4, 3, -7, 7, -1, 4, 5,
    -- filter=197 channel=21
    7, -5, 2, -6, -4, 3, 0, -4, 2,
    -- filter=197 channel=22
    -2, 5, 5, 6, 1, 1, -1, 4, -4,
    -- filter=197 channel=23
    -2, 0, -7, -3, -6, -1, 0, -9, -4,
    -- filter=197 channel=24
    -7, 5, -7, 3, 3, 0, 4, 3, 5,
    -- filter=197 channel=25
    0, -5, -6, -1, -1, -4, -1, 0, -3,
    -- filter=197 channel=26
    3, -3, 0, -3, -4, -4, -5, 0, -3,
    -- filter=197 channel=27
    7, 3, 3, 6, -8, 3, -3, -11, 7,
    -- filter=197 channel=28
    -4, 1, 4, 0, 5, 3, -3, -4, -4,
    -- filter=197 channel=29
    -1, -9, 4, -4, -8, -1, 1, -7, -4,
    -- filter=197 channel=30
    0, 6, 1, -7, 6, -1, 3, -2, 4,
    -- filter=197 channel=31
    2, 1, -2, 4, -12, 0, -8, -8, -3,
    -- filter=197 channel=32
    3, -6, 3, -3, -3, 5, 0, -10, 1,
    -- filter=197 channel=33
    4, -6, 4, 1, 5, 3, 0, -4, 4,
    -- filter=197 channel=34
    -2, -6, -8, 0, 1, 0, 5, 0, 5,
    -- filter=197 channel=35
    -6, -1, -6, -1, -4, -7, 1, -1, -5,
    -- filter=197 channel=36
    4, -5, -4, 4, -8, 1, -5, -3, 9,
    -- filter=197 channel=37
    6, 10, 3, -3, 4, 1, -2, 8, 5,
    -- filter=197 channel=38
    -5, -5, -6, -3, 2, 3, -2, -3, -6,
    -- filter=197 channel=39
    5, 1, -4, -4, -6, 0, -7, 6, 7,
    -- filter=197 channel=40
    0, -2, 7, 7, 1, 3, 6, 4, -6,
    -- filter=197 channel=41
    -3, -3, -12, 0, 6, -5, 0, -2, 0,
    -- filter=197 channel=42
    6, -4, 2, 6, 1, 6, -8, 2, 2,
    -- filter=197 channel=43
    -5, 5, 2, 3, -2, 5, 5, -5, 4,
    -- filter=197 channel=44
    2, -4, 1, 5, -4, -2, 2, -7, 6,
    -- filter=197 channel=45
    4, 3, 0, -5, 2, -1, 6, 7, 4,
    -- filter=197 channel=46
    0, 8, 0, -2, 7, 0, 1, 4, -5,
    -- filter=197 channel=47
    8, -3, 0, -5, -2, -4, -8, 0, 5,
    -- filter=197 channel=48
    8, -2, -5, -1, -4, -6, -8, 3, -4,
    -- filter=197 channel=49
    3, 4, 5, -5, -8, 1, 3, -5, -2,
    -- filter=197 channel=50
    0, 1, 6, -7, -8, 0, 0, 2, 4,
    -- filter=197 channel=51
    -4, 1, 6, 3, 2, 2, 6, 1, 0,
    -- filter=197 channel=52
    0, -6, 2, 5, -3, -3, 0, 2, 3,
    -- filter=197 channel=53
    1, 4, 0, 6, 5, 7, -1, -4, 5,
    -- filter=197 channel=54
    7, -1, 5, -1, 2, -7, -2, -5, -3,
    -- filter=197 channel=55
    5, 1, -6, 3, -9, -5, -4, -2, 6,
    -- filter=197 channel=56
    3, -2, -1, -1, -4, -4, 0, 4, 5,
    -- filter=197 channel=57
    0, -2, -2, -6, 0, -2, 3, 0, -3,
    -- filter=197 channel=58
    -7, -3, 2, 2, 12, 1, 4, -2, -7,
    -- filter=197 channel=59
    1, -3, -7, 3, -5, -7, -8, -5, 6,
    -- filter=197 channel=60
    0, 4, 5, 1, 0, 6, -1, 3, 4,
    -- filter=197 channel=61
    3, 2, 3, 5, 4, -2, -6, 5, 7,
    -- filter=197 channel=62
    6, 7, -6, 5, -2, 0, 5, 5, 1,
    -- filter=197 channel=63
    -8, 0, -4, 6, -3, -3, -2, -6, -3,
    -- filter=197 channel=64
    6, -3, -3, 1, -7, 3, 7, -2, -1,
    -- filter=197 channel=65
    -4, -2, 2, 4, -1, 0, 3, 3, 0,
    -- filter=197 channel=66
    -4, -2, 1, -1, 0, -2, 6, 0, 3,
    -- filter=197 channel=67
    -1, -7, 0, -3, -2, -7, -4, 2, -6,
    -- filter=197 channel=68
    0, -3, 3, 3, -2, 4, -5, -5, 2,
    -- filter=197 channel=69
    1, 3, -4, 2, 1, 0, 6, -3, -6,
    -- filter=197 channel=70
    8, -6, 2, 1, -9, -1, 1, -1, 2,
    -- filter=197 channel=71
    2, 0, -2, 0, 4, -6, 6, 5, 0,
    -- filter=197 channel=72
    2, 0, -3, -5, -6, 3, 1, -5, 0,
    -- filter=197 channel=73
    7, -3, -7, 4, -5, -2, 1, -2, 5,
    -- filter=197 channel=74
    1, -1, 0, 3, -5, 2, 0, -1, 0,
    -- filter=197 channel=75
    -4, 12, -3, -2, 15, -5, -5, 0, -6,
    -- filter=197 channel=76
    -5, -8, 2, 5, -5, 3, -7, -6, 4,
    -- filter=197 channel=77
    -1, 0, 2, 0, -4, -7, -2, 6, -7,
    -- filter=197 channel=78
    -6, 7, 3, -7, 4, 3, -2, -1, 4,
    -- filter=197 channel=79
    -3, -3, -3, 5, -7, -5, 0, 0, -2,
    -- filter=197 channel=80
    8, -5, -6, 4, -7, -10, -5, -2, 9,
    -- filter=197 channel=81
    0, -2, 3, -5, 4, -5, 4, -7, -2,
    -- filter=197 channel=82
    -2, 4, 0, 5, 2, -3, 2, -7, -6,
    -- filter=197 channel=83
    -1, 4, 2, 1, 5, 3, 6, 1, 6,
    -- filter=197 channel=84
    -2, 5, -2, 0, 1, -4, 3, 4, 2,
    -- filter=197 channel=85
    -1, -4, 6, 4, 3, -5, 4, 0, 4,
    -- filter=197 channel=86
    -5, 5, 4, 3, -2, 6, -8, -5, -3,
    -- filter=197 channel=87
    2, -2, -6, 3, -7, 2, -5, -4, -1,
    -- filter=197 channel=88
    -4, -3, -7, 6, -4, 2, 4, -2, -1,
    -- filter=197 channel=89
    1, 2, 3, 4, -10, -8, -8, -9, 5,
    -- filter=197 channel=90
    -6, -7, -2, -7, -4, 4, 3, 0, 7,
    -- filter=197 channel=91
    -4, -5, -1, -3, 0, 3, 1, 0, 5,
    -- filter=197 channel=92
    -2, -2, 1, -3, -6, 0, -2, 4, 2,
    -- filter=197 channel=93
    -5, -4, 0, -7, -6, -1, 2, 8, 2,
    -- filter=197 channel=94
    4, -1, 7, 0, -2, 6, 7, -5, 0,
    -- filter=197 channel=95
    4, -2, 0, -1, 0, 0, -1, 5, 4,
    -- filter=197 channel=96
    -7, 0, 2, -3, -1, -5, 0, 0, 0,
    -- filter=197 channel=97
    3, -1, 0, 4, 5, 0, 7, -1, -5,
    -- filter=197 channel=98
    0, -7, 1, 1, -5, -4, 1, -4, 1,
    -- filter=197 channel=99
    8, 2, -1, -5, -6, -3, -5, 0, 1,
    -- filter=197 channel=100
    0, 1, 6, -1, -4, -4, -3, 1, -8,
    -- filter=197 channel=101
    -5, -2, -1, -1, -3, 7, 6, 0, 9,
    -- filter=197 channel=102
    2, -1, -1, 0, 3, 3, 2, -7, 5,
    -- filter=197 channel=103
    7, 7, 3, 7, -4, 0, -6, -6, -7,
    -- filter=197 channel=104
    9, 3, 1, 0, -6, -1, 0, 5, 0,
    -- filter=197 channel=105
    -2, -4, -1, -5, -2, 0, 7, 7, 0,
    -- filter=197 channel=106
    0, 1, 4, 6, -7, -2, -5, -1, 2,
    -- filter=197 channel=107
    5, 1, 3, -6, 0, 6, 1, 3, -6,
    -- filter=197 channel=108
    6, 0, -1, -4, 3, 0, 4, 0, -2,
    -- filter=197 channel=109
    1, 0, -1, 4, -9, 3, -8, -10, -4,
    -- filter=197 channel=110
    -6, 0, 0, 4, -7, 5, -8, -8, 3,
    -- filter=197 channel=111
    0, -2, -8, 0, -3, -4, 5, -1, -3,
    -- filter=197 channel=112
    -3, 4, 6, -1, -6, -4, 4, 5, 4,
    -- filter=197 channel=113
    2, 0, 5, -1, -4, -8, 3, -5, 2,
    -- filter=197 channel=114
    -6, 11, -4, 9, 0, -4, 1, -3, 2,
    -- filter=197 channel=115
    0, 3, 5, -5, -4, 0, 4, 4, 1,
    -- filter=197 channel=116
    -3, 3, -3, -2, -2, -6, -6, 2, -1,
    -- filter=197 channel=117
    7, -2, 5, 1, 1, -7, 6, 0, 7,
    -- filter=197 channel=118
    2, 4, -7, 5, -2, 7, 6, -3, 4,
    -- filter=197 channel=119
    5, 3, -4, -7, 4, 4, -3, -4, 3,
    -- filter=197 channel=120
    1, 0, -3, 3, -11, -3, -4, -1, 8,
    -- filter=197 channel=121
    -1, 5, 0, -1, 3, 0, 2, 3, 2,
    -- filter=197 channel=122
    0, -6, -2, -5, -12, -5, 0, -4, 4,
    -- filter=197 channel=123
    -2, 6, 5, -2, -7, -1, 1, -7, 1,
    -- filter=197 channel=124
    -5, -2, 0, -7, -2, -6, 0, 7, 7,
    -- filter=197 channel=125
    7, -5, -2, -2, -12, -4, 4, -1, 2,
    -- filter=197 channel=126
    5, -4, -5, 0, 0, -3, -4, 1, 0,
    -- filter=197 channel=127
    -4, -1, -3, -5, 0, -4, -4, 2, -7,
    -- filter=198 channel=0
    0, 1, 3, 0, 0, -2, 4, 3, 5,
    -- filter=198 channel=1
    -4, -5, -6, -6, 0, 0, -6, 3, -1,
    -- filter=198 channel=2
    -5, -3, 2, 5, 7, 6, -7, 5, 6,
    -- filter=198 channel=3
    3, -6, -5, 6, -4, -6, -2, -2, 0,
    -- filter=198 channel=4
    6, -1, 6, 1, -2, -1, 4, 4, -4,
    -- filter=198 channel=5
    1, 6, -6, 6, 1, 1, 6, -4, 6,
    -- filter=198 channel=6
    -3, -3, -8, -6, 1, -5, 0, 2, 0,
    -- filter=198 channel=7
    0, -1, 0, 0, -5, 1, 3, 6, -4,
    -- filter=198 channel=8
    -2, 1, 0, 3, -1, -1, 6, -6, -5,
    -- filter=198 channel=9
    6, -5, 2, -7, 5, -5, 6, 5, -4,
    -- filter=198 channel=10
    1, 1, -2, 4, 3, 2, 2, -5, 0,
    -- filter=198 channel=11
    5, 4, 0, 3, -3, 0, -1, 6, 6,
    -- filter=198 channel=12
    2, 0, 2, 6, -4, -6, 7, 2, 0,
    -- filter=198 channel=13
    -3, 3, 5, -6, 0, 1, -8, 0, -7,
    -- filter=198 channel=14
    -2, 5, 0, 0, -1, 4, -6, -5, 1,
    -- filter=198 channel=15
    0, -6, -1, 1, 6, -8, 4, -3, -3,
    -- filter=198 channel=16
    1, -2, 4, 4, 2, 4, -1, -6, -2,
    -- filter=198 channel=17
    -5, 1, 0, 6, -5, 3, -1, 0, 4,
    -- filter=198 channel=18
    4, -3, -9, -6, 0, -3, 4, -7, -3,
    -- filter=198 channel=19
    1, 0, -4, 1, -2, 6, 3, 4, 0,
    -- filter=198 channel=20
    4, -2, -2, 4, -1, -8, -2, 3, 5,
    -- filter=198 channel=21
    -2, -3, -5, 2, 6, -1, 4, -7, -6,
    -- filter=198 channel=22
    6, 1, -1, 5, 1, -2, 2, 0, 6,
    -- filter=198 channel=23
    6, -4, 3, -3, -3, 1, 0, 4, -4,
    -- filter=198 channel=24
    0, 4, 0, 3, -3, -6, 0, -4, 0,
    -- filter=198 channel=25
    -5, 4, -4, 2, 0, 5, 3, -5, -1,
    -- filter=198 channel=26
    -6, 5, -3, -5, -5, -6, -3, 4, 6,
    -- filter=198 channel=27
    3, 4, 5, 1, 3, -4, -6, -8, -2,
    -- filter=198 channel=28
    -6, 4, 7, -4, 0, 6, -4, 0, 5,
    -- filter=198 channel=29
    -5, -7, -3, 4, -5, -1, -3, -2, 3,
    -- filter=198 channel=30
    -7, -7, 2, 4, 7, 5, -2, 0, -4,
    -- filter=198 channel=31
    -5, -1, -2, 7, 0, 6, -2, -1, -7,
    -- filter=198 channel=32
    -3, 1, -3, 0, 3, 0, -5, -1, -8,
    -- filter=198 channel=33
    0, -8, -1, -6, -1, -5, 1, 1, 1,
    -- filter=198 channel=34
    -1, 0, 0, -5, 3, 5, 0, 0, 6,
    -- filter=198 channel=35
    -2, -6, 6, -2, 3, 3, 4, -3, -5,
    -- filter=198 channel=36
    2, 3, 5, 7, -2, 2, 3, 5, 5,
    -- filter=198 channel=37
    -3, -6, -2, 5, 0, -5, 4, 7, 0,
    -- filter=198 channel=38
    -8, 0, -2, -6, 4, -2, -4, -6, 2,
    -- filter=198 channel=39
    -1, -6, -2, 8, 6, 1, 5, 0, 7,
    -- filter=198 channel=40
    2, 6, -3, 6, -2, -7, 2, -4, 5,
    -- filter=198 channel=41
    6, 2, 3, -7, 8, -5, -3, 6, -3,
    -- filter=198 channel=42
    -6, 0, 0, 1, 4, 5, 1, -3, 0,
    -- filter=198 channel=43
    6, 5, 1, 4, -4, -2, -6, 1, 2,
    -- filter=198 channel=44
    -4, -3, -6, 5, -5, -2, -5, -4, -7,
    -- filter=198 channel=45
    7, 0, -5, -5, 0, -4, -4, 7, 6,
    -- filter=198 channel=46
    -3, -3, 3, 1, -4, -5, 1, -6, -2,
    -- filter=198 channel=47
    0, -4, 4, 1, 7, -5, -2, 1, 2,
    -- filter=198 channel=48
    6, -5, -2, 0, -4, 3, -8, -6, -3,
    -- filter=198 channel=49
    -3, -5, 1, -4, -4, 5, -1, -1, -3,
    -- filter=198 channel=50
    -5, 1, -6, -1, 2, -5, 6, -1, -7,
    -- filter=198 channel=51
    -5, -3, 2, -6, 0, 5, 2, 3, -1,
    -- filter=198 channel=52
    -2, 1, -2, 5, 3, 5, 0, 4, 0,
    -- filter=198 channel=53
    7, -3, -2, 7, -6, 3, 0, -4, -1,
    -- filter=198 channel=54
    -6, 6, -2, -2, 6, -5, -3, 5, 0,
    -- filter=198 channel=55
    -5, 2, -3, 6, 6, -2, 5, -2, -3,
    -- filter=198 channel=56
    6, -5, -2, -2, 4, 2, 0, 0, 4,
    -- filter=198 channel=57
    -5, 6, -6, -3, -4, -5, 1, 1, -1,
    -- filter=198 channel=58
    -7, -3, -7, -5, -5, 4, 4, 2, 3,
    -- filter=198 channel=59
    0, -7, -6, -2, -2, -5, -9, 0, 0,
    -- filter=198 channel=60
    1, 1, 6, -3, 4, 5, -6, 6, 4,
    -- filter=198 channel=61
    0, 4, 6, -1, 6, -6, -4, 2, 5,
    -- filter=198 channel=62
    3, 3, -4, -2, -4, 5, 7, -1, 1,
    -- filter=198 channel=63
    2, 6, -1, 6, 0, 3, -1, 4, 0,
    -- filter=198 channel=64
    2, -5, 7, 5, 7, 3, -1, -2, 0,
    -- filter=198 channel=65
    6, -4, -7, 6, 6, 0, 1, 0, 0,
    -- filter=198 channel=66
    -3, -2, 2, -3, -1, -2, 3, -1, 0,
    -- filter=198 channel=67
    0, -4, 5, 4, -5, 5, 3, -3, -2,
    -- filter=198 channel=68
    -1, 4, -3, 1, -3, -6, 3, -3, 0,
    -- filter=198 channel=69
    -5, 6, 2, -1, 4, -4, 0, 4, 1,
    -- filter=198 channel=70
    0, 3, -5, 4, -1, -6, -7, -3, 2,
    -- filter=198 channel=71
    0, 4, 1, -5, 0, 5, -3, 2, 0,
    -- filter=198 channel=72
    4, 2, 6, -2, 2, 3, -1, 5, -4,
    -- filter=198 channel=73
    -2, 0, -3, 3, 6, 3, 4, -2, 5,
    -- filter=198 channel=74
    0, -7, -4, -3, 1, -4, 1, -1, -4,
    -- filter=198 channel=75
    1, 1, -2, -4, 4, -3, 6, 2, 1,
    -- filter=198 channel=76
    -1, 3, -5, 7, -5, -2, -5, 0, 0,
    -- filter=198 channel=77
    -3, 1, -3, 2, 1, -3, -7, 3, -3,
    -- filter=198 channel=78
    -5, -5, -7, 4, 4, 2, -5, -2, 6,
    -- filter=198 channel=79
    -1, -6, 0, 0, 1, 4, -8, 3, -6,
    -- filter=198 channel=80
    -8, 5, -2, -1, 4, 5, 0, -4, -2,
    -- filter=198 channel=81
    1, -2, -7, -2, 5, -6, -6, 2, 3,
    -- filter=198 channel=82
    -5, 2, -3, 3, 3, -6, 4, 3, 1,
    -- filter=198 channel=83
    2, -1, 1, 4, 0, 0, -5, 0, 3,
    -- filter=198 channel=84
    5, 6, 0, 2, -1, 2, 0, -7, 2,
    -- filter=198 channel=85
    2, -3, -1, 0, 0, 1, -2, 6, 2,
    -- filter=198 channel=86
    -2, -3, 5, -5, -5, -7, -5, 2, -3,
    -- filter=198 channel=87
    3, 0, 3, 6, -6, 6, 6, -5, 4,
    -- filter=198 channel=88
    5, -1, 6, -3, 1, 8, -5, 0, 4,
    -- filter=198 channel=89
    -9, 0, 4, -3, -1, -4, -7, -4, 2,
    -- filter=198 channel=90
    -4, 1, 1, 7, 4, -2, 5, 8, -1,
    -- filter=198 channel=91
    -3, -2, 1, 5, 4, 5, 0, -5, -6,
    -- filter=198 channel=92
    0, -3, 5, 0, -3, 0, 3, -3, 4,
    -- filter=198 channel=93
    4, 2, 2, 5, -7, 1, -4, -6, 3,
    -- filter=198 channel=94
    0, -6, -4, -2, 2, -6, 5, 1, 0,
    -- filter=198 channel=95
    -1, -7, -2, 1, -6, -6, 1, 6, 4,
    -- filter=198 channel=96
    0, 7, 1, -6, 1, 0, -2, 4, 6,
    -- filter=198 channel=97
    0, -6, 5, 1, -7, 0, 0, -1, 4,
    -- filter=198 channel=98
    -2, 3, 7, -7, -2, -2, -1, -7, -8,
    -- filter=198 channel=99
    0, 3, 5, 0, -3, 2, 0, -1, 6,
    -- filter=198 channel=100
    4, 1, -6, 1, 2, -6, -4, 1, 0,
    -- filter=198 channel=101
    0, 5, 6, 4, -6, 5, 0, 1, 0,
    -- filter=198 channel=102
    -6, 2, 1, 1, -6, 6, -1, 4, -5,
    -- filter=198 channel=103
    -4, 5, -3, 2, -6, 2, 3, -2, 6,
    -- filter=198 channel=104
    4, -3, -1, -2, 7, 0, -7, -5, -7,
    -- filter=198 channel=105
    -2, -4, -4, 3, 6, 4, -5, 7, -2,
    -- filter=198 channel=106
    0, 1, -1, -7, 7, 6, -3, 7, 0,
    -- filter=198 channel=107
    6, -6, -7, 4, 3, -1, 4, 1, 2,
    -- filter=198 channel=108
    -2, -5, 7, -6, 4, -5, -3, -2, -4,
    -- filter=198 channel=109
    -6, 2, -4, 0, 2, -4, -4, -2, 0,
    -- filter=198 channel=110
    0, -5, 7, -6, 0, 0, 1, 0, 5,
    -- filter=198 channel=111
    0, -1, -7, -2, -1, -2, 1, 0, -4,
    -- filter=198 channel=112
    1, -4, 0, 0, 0, 6, 5, -6, -5,
    -- filter=198 channel=113
    -1, 2, 1, -3, -6, 3, -2, 2, 3,
    -- filter=198 channel=114
    -4, -3, 0, 5, -2, 2, -9, -1, -1,
    -- filter=198 channel=115
    7, 0, 4, 1, -6, 4, 7, 3, 2,
    -- filter=198 channel=116
    -2, -2, 5, 5, -1, 4, 0, -6, -2,
    -- filter=198 channel=117
    -4, 5, -5, 0, -3, 3, -4, 5, -3,
    -- filter=198 channel=118
    1, 2, 4, -3, 0, -5, -5, -5, -3,
    -- filter=198 channel=119
    0, -4, 2, 2, 2, 2, 0, 6, -3,
    -- filter=198 channel=120
    2, -3, 2, 1, -2, -9, 2, 4, 1,
    -- filter=198 channel=121
    2, -6, 3, -3, 0, -4, 0, -4, -6,
    -- filter=198 channel=122
    -4, -2, 1, -1, 6, -1, 1, 0, 0,
    -- filter=198 channel=123
    0, 3, 3, 2, 4, 0, 4, 0, -5,
    -- filter=198 channel=124
    1, 4, 4, -6, 4, 6, 2, 3, 0,
    -- filter=198 channel=125
    4, 4, 2, -6, 0, 4, -3, -6, -7,
    -- filter=198 channel=126
    3, 0, -2, -8, 6, -6, 0, 0, -4,
    -- filter=198 channel=127
    -6, -1, 3, 0, 4, 2, 5, 1, 1,
    -- filter=199 channel=0
    -8, 11, -9, -9, 18, 10, -11, 5, 8,
    -- filter=199 channel=1
    4, 12, -3, -2, 15, 8, -14, 14, 1,
    -- filter=199 channel=2
    -3, 1, -7, -2, -4, -9, 0, 2, -2,
    -- filter=199 channel=3
    -7, -3, -8, -12, -8, 0, -1, 2, 11,
    -- filter=199 channel=4
    1, -2, 1, 1, 6, -5, 9, 10, 4,
    -- filter=199 channel=5
    -10, 7, -3, -6, 9, -2, -12, -2, -9,
    -- filter=199 channel=6
    3, -2, 3, -11, -11, -10, -5, 0, 2,
    -- filter=199 channel=7
    -6, 7, -2, 1, 1, -3, -4, 6, -5,
    -- filter=199 channel=8
    -6, -6, -5, 3, -5, 0, -2, 0, -1,
    -- filter=199 channel=9
    2, 5, 4, 0, 0, 0, 0, 2, 1,
    -- filter=199 channel=10
    0, -7, -13, -4, -15, -13, 5, 3, -8,
    -- filter=199 channel=11
    -1, -3, 3, -11, -15, -4, 3, -3, -6,
    -- filter=199 channel=12
    6, -6, -3, 2, 3, -8, -2, 1, -5,
    -- filter=199 channel=13
    0, -10, -4, -2, -1, -4, 14, 3, -2,
    -- filter=199 channel=14
    -1, -1, 1, -4, -1, 0, 4, -7, 3,
    -- filter=199 channel=15
    0, 2, 4, 3, 2, -8, -1, 3, -4,
    -- filter=199 channel=16
    1, -2, -3, 13, 2, 0, 6, 0, 0,
    -- filter=199 channel=17
    2, 4, 5, -3, 3, 0, -5, -6, -3,
    -- filter=199 channel=18
    0, 3, -5, -6, 3, 7, 8, 18, 8,
    -- filter=199 channel=19
    2, -4, 0, 7, -3, -5, 5, -5, 2,
    -- filter=199 channel=20
    -1, -11, 0, -15, -9, -12, -2, -1, 2,
    -- filter=199 channel=21
    13, -8, 1, 11, -1, 2, 2, 0, -11,
    -- filter=199 channel=22
    5, -6, -12, -7, -3, 2, 0, 2, 0,
    -- filter=199 channel=23
    -2, -12, -13, 4, -7, -25, 8, -1, -5,
    -- filter=199 channel=24
    2, -4, -1, 2, -3, 5, -6, -5, 0,
    -- filter=199 channel=25
    3, -3, -5, 12, 15, -4, 3, 7, 3,
    -- filter=199 channel=26
    8, 0, -10, -2, 6, 2, -4, -6, -4,
    -- filter=199 channel=27
    4, 3, -3, 15, 15, -12, 11, 26, 5,
    -- filter=199 channel=28
    -5, -6, -7, 3, 0, 7, 4, -2, -7,
    -- filter=199 channel=29
    -1, 0, 0, -11, -19, -7, 6, -2, -7,
    -- filter=199 channel=30
    6, 6, -4, -2, 5, 0, -9, 8, 5,
    -- filter=199 channel=31
    4, -12, -12, 7, -11, -18, 9, -7, -13,
    -- filter=199 channel=32
    -4, -5, -11, 0, 10, -3, 5, 13, 7,
    -- filter=199 channel=33
    -9, -7, -7, 5, 0, -2, -1, 16, 5,
    -- filter=199 channel=34
    0, -7, -14, -1, -10, -21, 0, 4, -15,
    -- filter=199 channel=35
    -3, 6, 7, -1, -1, -2, -3, -5, 6,
    -- filter=199 channel=36
    -3, -11, -5, 0, -13, -4, 13, -10, -12,
    -- filter=199 channel=37
    0, 17, -7, 1, 30, 14, -15, 13, 2,
    -- filter=199 channel=38
    1, 2, -8, 3, 3, -13, 8, 2, 2,
    -- filter=199 channel=39
    0, -6, 2, -9, -3, -3, 4, -6, -4,
    -- filter=199 channel=40
    1, 5, 0, -2, -9, -2, 5, 7, 6,
    -- filter=199 channel=41
    0, -14, 3, 8, -12, -12, 13, 0, 3,
    -- filter=199 channel=42
    1, 7, 9, -4, 12, 9, -4, -3, 2,
    -- filter=199 channel=43
    -1, 0, -6, -5, -5, -8, 0, 8, -3,
    -- filter=199 channel=44
    8, -1, -6, 7, 18, 0, 5, 4, 0,
    -- filter=199 channel=45
    0, 6, -2, 0, 2, 9, 1, -5, -1,
    -- filter=199 channel=46
    7, 0, 0, 8, 8, -2, -1, 8, 0,
    -- filter=199 channel=47
    13, 0, 2, 4, 4, 6, -2, 0, -4,
    -- filter=199 channel=48
    4, 8, -5, 8, 16, 10, 11, 17, 1,
    -- filter=199 channel=49
    4, -1, 0, -1, -3, -3, 5, 1, 13,
    -- filter=199 channel=50
    -3, 4, -3, 3, 2, 0, -2, 7, -1,
    -- filter=199 channel=51
    0, 5, -5, -3, -4, 0, -5, 5, -6,
    -- filter=199 channel=52
    5, -10, -2, 2, -6, -9, 6, 6, -9,
    -- filter=199 channel=53
    0, 2, 1, 3, -4, -3, -1, 1, -2,
    -- filter=199 channel=54
    4, 4, -6, 3, 5, 0, 6, -2, 3,
    -- filter=199 channel=55
    0, -13, -5, -6, -19, -20, 4, 1, 1,
    -- filter=199 channel=56
    -5, -10, -11, 0, -1, -5, 2, -4, -7,
    -- filter=199 channel=57
    3, 3, -7, -6, -3, 6, 2, 3, 5,
    -- filter=199 channel=58
    -10, -7, 1, -6, 4, 1, -6, -7, 5,
    -- filter=199 channel=59
    1, -7, -6, 17, 10, -5, 9, 10, 9,
    -- filter=199 channel=60
    6, -3, 5, -4, -1, -7, -6, 7, 2,
    -- filter=199 channel=61
    0, -2, -3, 0, -7, -3, 1, -7, -10,
    -- filter=199 channel=62
    -7, 0, 4, -5, 1, 0, -2, -5, 3,
    -- filter=199 channel=63
    -10, -3, -6, -13, -2, 4, -13, -5, -7,
    -- filter=199 channel=64
    -7, -11, 1, 6, -14, -4, -3, -6, 3,
    -- filter=199 channel=65
    -6, 3, -4, 6, -2, 0, -2, 0, 4,
    -- filter=199 channel=66
    -7, -10, -1, -1, -2, -7, 3, -3, -11,
    -- filter=199 channel=67
    0, 0, 4, -5, -5, -2, -5, -1, 3,
    -- filter=199 channel=68
    -4, -1, 3, 4, -4, 1, 0, 3, 9,
    -- filter=199 channel=69
    -3, -8, -6, 4, -8, 0, -8, 0, 4,
    -- filter=199 channel=70
    6, 2, -9, 9, 1, -8, 11, 10, -6,
    -- filter=199 channel=71
    -9, -9, 0, 0, 0, -7, -4, 6, 0,
    -- filter=199 channel=72
    0, -17, -4, 9, -15, -10, 1, -1, -13,
    -- filter=199 channel=73
    0, -4, -6, -1, 2, -2, 5, 0, 6,
    -- filter=199 channel=74
    2, -8, -9, 0, -4, -20, 5, 1, -18,
    -- filter=199 channel=75
    -4, -1, -1, -3, 17, 8, -9, 4, 11,
    -- filter=199 channel=76
    -7, 2, 3, -3, -12, -4, 3, -1, -7,
    -- filter=199 channel=77
    2, -6, -5, 4, -5, -3, -3, 1, -7,
    -- filter=199 channel=78
    -9, -5, -2, -9, 2, -10, -9, -3, -5,
    -- filter=199 channel=79
    0, 3, 2, 0, 8, 5, 0, 15, 6,
    -- filter=199 channel=80
    6, -2, -8, 1, -8, -10, 14, 2, 1,
    -- filter=199 channel=81
    2, -7, 0, -5, -3, -6, -7, 6, 2,
    -- filter=199 channel=82
    -3, 0, -5, -5, -6, -8, 1, 6, 4,
    -- filter=199 channel=83
    8, 3, 4, 2, 1, 1, 7, 2, 1,
    -- filter=199 channel=84
    6, -5, -3, 0, 0, -6, -2, 10, 5,
    -- filter=199 channel=85
    4, 1, 7, -4, 2, 0, -3, -6, -1,
    -- filter=199 channel=86
    0, -3, -5, -8, 7, -14, -1, -2, -2,
    -- filter=199 channel=87
    -7, -1, -2, -3, -12, -7, 4, -2, -2,
    -- filter=199 channel=88
    0, -1, -3, 9, -6, -12, 11, 0, -5,
    -- filter=199 channel=89
    -1, -1, 1, -3, -14, -5, 10, -4, -6,
    -- filter=199 channel=90
    5, -10, -7, 0, -10, -14, 13, -4, -15,
    -- filter=199 channel=91
    -3, -1, 0, 4, 10, -10, 9, 19, 2,
    -- filter=199 channel=92
    5, -5, -11, -4, 2, -4, 5, 0, -6,
    -- filter=199 channel=93
    9, 8, -1, 3, 10, 10, 6, 11, 7,
    -- filter=199 channel=94
    3, 3, -6, 0, 2, 4, -5, 4, 1,
    -- filter=199 channel=95
    -7, 1, 3, -7, -4, -9, 3, -4, -4,
    -- filter=199 channel=96
    7, 0, 4, 0, -3, 7, 0, -5, 11,
    -- filter=199 channel=97
    -9, -10, -6, -6, 3, -5, -3, 7, 0,
    -- filter=199 channel=98
    -4, 0, 0, 0, -1, -11, 6, 12, 3,
    -- filter=199 channel=99
    -7, -11, -11, -4, -16, -23, 7, -6, -16,
    -- filter=199 channel=100
    4, -8, -4, 0, -9, -7, -1, 6, 0,
    -- filter=199 channel=101
    -1, -7, -8, -3, 2, -8, 3, 10, -2,
    -- filter=199 channel=102
    3, -1, -3, 6, 7, -1, 7, -5, 1,
    -- filter=199 channel=103
    6, -7, 0, 2, 0, -8, -7, 0, -4,
    -- filter=199 channel=104
    2, -15, -7, 10, 0, -13, 2, -6, -11,
    -- filter=199 channel=105
    -9, 0, -7, -9, -6, -7, -1, 0, 0,
    -- filter=199 channel=106
    -4, -3, 8, -1, -10, 2, -1, 2, 0,
    -- filter=199 channel=107
    -11, -5, 1, -6, -9, 2, 2, -8, 3,
    -- filter=199 channel=108
    -8, -7, -5, -2, 0, -4, -7, 0, 2,
    -- filter=199 channel=109
    0, 3, -3, 13, 4, -14, 5, 24, -6,
    -- filter=199 channel=110
    -5, -12, -8, -6, -15, -16, -5, -1, -1,
    -- filter=199 channel=111
    -4, -9, -3, 4, 0, 3, 1, -3, -6,
    -- filter=199 channel=112
    -4, 7, -13, 6, 1, -6, -1, 5, -13,
    -- filter=199 channel=113
    -8, 1, -16, 8, -6, -8, -2, 1, -2,
    -- filter=199 channel=114
    -7, 3, -8, 1, 19, -1, -3, 15, 14,
    -- filter=199 channel=115
    3, 3, -3, 5, -7, 3, 2, -4, -1,
    -- filter=199 channel=116
    5, -2, -4, 8, -7, -2, 17, 4, 8,
    -- filter=199 channel=117
    3, 2, 0, 3, -2, -3, -3, -6, 4,
    -- filter=199 channel=118
    -6, -5, 3, 1, 6, 0, 5, -4, 0,
    -- filter=199 channel=119
    2, -2, -17, -4, 0, -19, 17, 0, -19,
    -- filter=199 channel=120
    -2, -4, -6, 1, -6, -14, 9, 13, -13,
    -- filter=199 channel=121
    -4, -10, -5, 9, -3, -13, 5, -5, 1,
    -- filter=199 channel=122
    17, 4, -9, 25, 7, -3, 12, 5, -2,
    -- filter=199 channel=123
    2, -3, -2, 7, -2, -9, 10, 0, -7,
    -- filter=199 channel=124
    4, -5, -6, -10, -2, 1, 5, -5, -1,
    -- filter=199 channel=125
    1, -9, -10, 12, -3, -14, 9, 0, -8,
    -- filter=199 channel=126
    0, -9, 1, -1, -6, -10, -4, -3, 4,
    -- filter=199 channel=127
    -3, -9, -8, -7, -4, 2, -4, 0, -4,
    -- filter=200 channel=0
    -10, -4, 8, 4, 0, 0, 3, 5, 8,
    -- filter=200 channel=1
    3, 4, 1, -1, 0, -3, 8, 0, 5,
    -- filter=200 channel=2
    -5, -2, 4, -1, -1, 3, -1, 3, 0,
    -- filter=200 channel=3
    0, -1, 1, -7, -10, 5, -3, -7, 9,
    -- filter=200 channel=4
    4, 2, -5, -12, -5, 3, -8, -3, 9,
    -- filter=200 channel=5
    -5, -8, -7, -3, -7, 0, 1, 8, -2,
    -- filter=200 channel=6
    -5, 6, -1, -5, 3, 2, -3, -7, 1,
    -- filter=200 channel=7
    2, -1, -1, 5, -5, 2, -4, -3, -5,
    -- filter=200 channel=8
    -5, -4, -2, 4, -4, 3, 6, 6, 1,
    -- filter=200 channel=9
    -2, 0, -5, 0, -8, 2, 0, 2, 6,
    -- filter=200 channel=10
    -3, 5, -9, -3, 2, -3, -4, 6, 1,
    -- filter=200 channel=11
    0, -1, 4, -3, -7, 5, -5, 2, -3,
    -- filter=200 channel=12
    -1, -3, 0, 0, 1, 6, 5, 0, 9,
    -- filter=200 channel=13
    4, 7, -7, 0, 5, 4, 0, 3, 0,
    -- filter=200 channel=14
    2, -4, 2, 0, 5, 0, 7, 7, -3,
    -- filter=200 channel=15
    5, -5, 7, 0, -8, -8, 1, -3, 0,
    -- filter=200 channel=16
    0, 2, -4, 2, -5, -3, -2, 7, 10,
    -- filter=200 channel=17
    7, 1, 4, -3, 0, 2, -2, 3, 0,
    -- filter=200 channel=18
    6, -4, 4, 3, -6, -1, -6, -9, 2,
    -- filter=200 channel=19
    3, 0, -2, -2, 4, 1, 5, -2, -1,
    -- filter=200 channel=20
    8, 14, 12, 10, -4, 9, -4, -8, -1,
    -- filter=200 channel=21
    -8, 0, -12, 5, 2, -1, 6, 13, 12,
    -- filter=200 channel=22
    3, 2, 5, 3, -3, 1, -7, -8, 2,
    -- filter=200 channel=23
    10, -1, -7, 0, -13, -5, -6, -3, -5,
    -- filter=200 channel=24
    -6, -6, -4, -7, 0, -4, 5, -6, 5,
    -- filter=200 channel=25
    -1, 3, -7, 6, -1, -1, 4, 8, 5,
    -- filter=200 channel=26
    1, -8, -2, -6, -3, 3, -8, -4, -2,
    -- filter=200 channel=27
    -1, -6, -2, -4, -8, -4, 0, -3, 8,
    -- filter=200 channel=28
    4, -2, -1, 3, 4, 7, -5, 6, 0,
    -- filter=200 channel=29
    4, 3, -1, -3, 2, 4, 3, -7, -7,
    -- filter=200 channel=30
    3, -9, -7, -3, 0, 3, 3, 8, 6,
    -- filter=200 channel=31
    -5, -11, -14, 7, -1, -7, 15, 18, 8,
    -- filter=200 channel=32
    10, 0, 3, 7, -7, -5, -3, 1, 5,
    -- filter=200 channel=33
    -6, 0, 0, 4, -2, -4, -7, 6, 1,
    -- filter=200 channel=34
    -2, -4, 8, -6, -4, -6, 6, 2, 3,
    -- filter=200 channel=35
    4, 2, 0, 3, -3, -3, -4, 7, -4,
    -- filter=200 channel=36
    3, -1, 5, 9, 5, -4, 7, 5, 5,
    -- filter=200 channel=37
    -1, -8, -3, -8, -3, 0, 3, 0, 6,
    -- filter=200 channel=38
    3, -8, 4, 6, -3, -8, 4, 7, 4,
    -- filter=200 channel=39
    0, 9, 2, -4, 5, 7, 6, -5, -1,
    -- filter=200 channel=40
    8, 3, -3, 0, 1, 1, 4, 1, -4,
    -- filter=200 channel=41
    5, 9, -1, 11, -2, 0, 2, -10, -2,
    -- filter=200 channel=42
    6, -8, -9, -6, 2, -5, 2, 3, -3,
    -- filter=200 channel=43
    -5, 0, 0, 0, -2, 2, 0, -3, -6,
    -- filter=200 channel=44
    0, -9, -8, -5, -1, -1, 2, 0, 10,
    -- filter=200 channel=45
    -2, -6, 1, -5, -4, 4, 4, 6, 1,
    -- filter=200 channel=46
    3, 2, 8, 0, 7, 0, -7, -1, 3,
    -- filter=200 channel=47
    -12, -8, -6, 4, -8, 0, 7, 11, 9,
    -- filter=200 channel=48
    -2, -6, -12, 6, -2, 0, 10, 8, 10,
    -- filter=200 channel=49
    9, -2, -1, -8, 0, -3, 0, -5, -4,
    -- filter=200 channel=50
    -6, -8, -1, 2, -1, -9, 7, -2, 8,
    -- filter=200 channel=51
    -2, 0, -1, 1, 4, -5, 6, -2, -4,
    -- filter=200 channel=52
    8, -5, -1, 7, 5, 1, -1, -8, 6,
    -- filter=200 channel=53
    -1, 6, 7, -2, 0, 3, -7, -9, 5,
    -- filter=200 channel=54
    -6, -1, 0, 0, -2, 5, -6, -4, -5,
    -- filter=200 channel=55
    6, 1, -5, 4, -5, -2, -7, -7, -5,
    -- filter=200 channel=56
    0, 2, -7, -4, 6, 2, -3, 5, -3,
    -- filter=200 channel=57
    -3, -1, 2, -7, 1, -3, -2, -3, -6,
    -- filter=200 channel=58
    0, -8, 6, -3, 5, -1, 3, 2, 7,
    -- filter=200 channel=59
    1, -7, -13, 6, -4, 4, 9, 1, 12,
    -- filter=200 channel=60
    -6, 1, 7, -7, 5, -3, -5, -2, -5,
    -- filter=200 channel=61
    0, 7, 3, -1, -2, -5, -4, -5, -2,
    -- filter=200 channel=62
    -5, -4, 2, 0, 0, 4, 0, 5, 6,
    -- filter=200 channel=63
    -6, -9, 2, -7, -7, -9, 4, -3, -8,
    -- filter=200 channel=64
    7, -3, -4, 0, 4, 0, 0, 0, 2,
    -- filter=200 channel=65
    6, 3, -1, -7, -4, -3, -3, 1, -1,
    -- filter=200 channel=66
    5, 1, 0, 9, 1, -2, -6, -8, 6,
    -- filter=200 channel=67
    6, -1, 4, 0, 1, 3, 4, -3, -1,
    -- filter=200 channel=68
    1, -3, -4, 2, 1, 5, 0, -2, 3,
    -- filter=200 channel=69
    4, -6, -4, 2, -1, 4, 6, -3, 0,
    -- filter=200 channel=70
    0, -6, -3, 5, -3, 6, 2, -5, 10,
    -- filter=200 channel=71
    6, -1, -3, 4, 0, 2, 4, -1, -4,
    -- filter=200 channel=72
    -4, -10, -11, 6, 3, -4, 5, 2, -3,
    -- filter=200 channel=73
    3, -6, -4, 2, 2, 4, -8, 0, -3,
    -- filter=200 channel=74
    5, -4, 1, -1, -8, -7, 0, 1, 3,
    -- filter=200 channel=75
    -6, -9, 6, -3, 2, 1, 5, 1, -1,
    -- filter=200 channel=76
    15, 9, 0, 11, 2, -1, -6, -9, -2,
    -- filter=200 channel=77
    -3, 2, 2, 1, 3, 5, 5, -7, 6,
    -- filter=200 channel=78
    2, 1, -3, 1, 0, -2, -5, 0, 1,
    -- filter=200 channel=79
    2, -6, -2, -2, -4, -7, -8, -8, 0,
    -- filter=200 channel=80
    -1, -12, -21, 3, -6, -11, 4, 13, 9,
    -- filter=200 channel=81
    3, 3, -5, -5, 0, 3, 7, -4, 4,
    -- filter=200 channel=82
    -5, -1, -2, 3, -5, 4, 6, -1, 5,
    -- filter=200 channel=83
    0, 1, 0, -6, 0, -6, 4, 11, 2,
    -- filter=200 channel=84
    1, 0, 2, -1, -7, 6, -3, -5, 9,
    -- filter=200 channel=85
    -4, -4, -4, 2, -5, 6, 3, -3, -5,
    -- filter=200 channel=86
    -7, 1, -4, 4, -8, 3, 6, -5, 6,
    -- filter=200 channel=87
    10, -2, 8, -4, -7, -5, 0, -11, -7,
    -- filter=200 channel=88
    5, 1, 1, 0, 0, 3, 6, 10, 3,
    -- filter=200 channel=89
    6, 1, -8, 9, -8, -8, 6, -3, 2,
    -- filter=200 channel=90
    1, 4, -5, 4, 2, 2, 5, 2, -5,
    -- filter=200 channel=91
    8, -7, -1, -8, 4, 1, -3, 1, 6,
    -- filter=200 channel=92
    -5, -7, 6, -7, -2, -1, -5, -7, -6,
    -- filter=200 channel=93
    -2, -6, -5, 3, 7, -4, 6, 7, 11,
    -- filter=200 channel=94
    2, 2, 3, 2, 6, 2, -4, 0, 5,
    -- filter=200 channel=95
    4, -4, 7, -7, -4, 7, 6, 4, -7,
    -- filter=200 channel=96
    -4, -5, 6, 7, -2, 5, 6, -7, 3,
    -- filter=200 channel=97
    -2, 2, -6, -5, -5, 4, 3, 1, -1,
    -- filter=200 channel=98
    -7, -8, -14, 0, -8, -2, 0, -2, 0,
    -- filter=200 channel=99
    3, 1, -9, 9, 0, -14, 4, 1, -6,
    -- filter=200 channel=100
    -4, -2, 1, -5, 1, 1, -1, -2, -1,
    -- filter=200 channel=101
    -4, 0, 5, -3, -5, -1, 1, -1, 0,
    -- filter=200 channel=102
    7, 5, 0, 0, 1, -3, 5, 2, 4,
    -- filter=200 channel=103
    -2, -5, -1, 1, -4, -12, 0, 11, 4,
    -- filter=200 channel=104
    -6, -3, -7, 7, 3, -7, 13, 16, 0,
    -- filter=200 channel=105
    1, 10, 3, 4, 4, -4, -6, -7, -3,
    -- filter=200 channel=106
    6, 2, 7, 8, 4, -5, -5, 2, -1,
    -- filter=200 channel=107
    0, 2, 0, 2, -8, 0, -8, -12, -7,
    -- filter=200 channel=108
    -4, 6, 2, 5, 5, 5, -6, -1, 7,
    -- filter=200 channel=109
    3, -5, -1, -4, 0, 4, -3, 0, 8,
    -- filter=200 channel=110
    -7, 1, 1, 6, -3, -12, 3, 4, -7,
    -- filter=200 channel=111
    0, 5, -3, 1, 3, 5, -1, 6, -5,
    -- filter=200 channel=112
    -7, 0, 5, -2, 1, 5, 0, 5, 1,
    -- filter=200 channel=113
    6, -5, -5, 6, 1, 0, -1, -2, 4,
    -- filter=200 channel=114
    7, -4, -4, -1, -12, -8, -4, -6, 2,
    -- filter=200 channel=115
    -3, -6, -2, -4, 5, 3, 5, 6, 4,
    -- filter=200 channel=116
    7, -7, -2, -2, -8, -5, 6, 1, 3,
    -- filter=200 channel=117
    -2, 6, -5, 0, 3, 1, -2, 0, 8,
    -- filter=200 channel=118
    0, 1, 0, -1, 1, -3, 0, -4, -3,
    -- filter=200 channel=119
    -6, -9, -2, 2, 0, 3, 0, -1, -5,
    -- filter=200 channel=120
    8, -11, -7, -10, -1, -7, -7, 2, 9,
    -- filter=200 channel=121
    1, -1, -2, 7, -7, 0, -3, 3, 4,
    -- filter=200 channel=122
    -8, -3, -9, 8, -3, 0, 11, 26, 19,
    -- filter=200 channel=123
    0, 6, -6, -4, -2, 5, 1, -8, -7,
    -- filter=200 channel=124
    0, 6, 8, -6, 0, 4, 5, -6, -4,
    -- filter=200 channel=125
    -4, 0, -2, 8, -5, -6, 11, -1, 6,
    -- filter=200 channel=126
    5, -4, -7, -1, -10, -6, -5, 0, -1,
    -- filter=200 channel=127
    -3, 6, 4, 5, -5, 0, 0, -5, 4,
    -- filter=201 channel=0
    -4, 2, -4, 6, 4, -2, -4, -6, 3,
    -- filter=201 channel=1
    -4, 4, 4, 2, 5, 7, -4, -2, -2,
    -- filter=201 channel=2
    -4, 3, 0, -5, 1, -6, 3, 7, -1,
    -- filter=201 channel=3
    2, -2, -3, -5, -6, 0, -5, 4, 6,
    -- filter=201 channel=4
    -7, -5, -1, -6, -6, 0, -4, 0, 5,
    -- filter=201 channel=5
    2, 7, 1, -1, -1, -6, 6, -2, 1,
    -- filter=201 channel=6
    -4, -2, 4, -4, 0, -3, -3, 3, 2,
    -- filter=201 channel=7
    -7, 6, 1, -3, 0, 3, 7, -6, 6,
    -- filter=201 channel=8
    7, -3, -3, 0, 5, 1, -6, 3, -5,
    -- filter=201 channel=9
    6, -1, -1, 1, 5, 3, -5, -2, -3,
    -- filter=201 channel=10
    -2, 0, 1, 2, 4, -2, 2, -2, -1,
    -- filter=201 channel=11
    2, 7, -4, -6, 0, 5, 4, 3, -3,
    -- filter=201 channel=12
    -1, 0, 5, -2, 6, -2, 0, 0, -5,
    -- filter=201 channel=13
    0, 0, -3, -1, 6, -1, 1, -2, -5,
    -- filter=201 channel=14
    -6, -1, -3, 0, 0, 5, 1, 7, 0,
    -- filter=201 channel=15
    4, -2, -4, -3, 3, -1, -3, 0, -2,
    -- filter=201 channel=16
    -7, -4, -1, -7, 1, -6, 2, 0, -2,
    -- filter=201 channel=17
    2, -5, 5, 6, 0, -4, -1, -6, -2,
    -- filter=201 channel=18
    5, 0, 6, 0, 1, -1, -5, 0, -1,
    -- filter=201 channel=19
    -6, 4, 7, 7, -7, -6, 5, -7, -7,
    -- filter=201 channel=20
    -4, -1, -5, -3, -6, 3, 0, -5, 1,
    -- filter=201 channel=21
    3, 0, 0, 4, 0, -7, 5, -1, -4,
    -- filter=201 channel=22
    0, 6, -2, 7, 3, -2, 2, -6, 7,
    -- filter=201 channel=23
    1, 0, -5, -3, 6, 6, -5, 7, -2,
    -- filter=201 channel=24
    1, -5, -1, 0, -3, -6, -6, 0, -6,
    -- filter=201 channel=25
    -6, -6, 2, 1, 7, -5, 3, 2, -7,
    -- filter=201 channel=26
    4, 1, 0, -1, 6, -2, 2, 5, 5,
    -- filter=201 channel=27
    6, 1, -4, 0, -7, -5, -7, 4, -6,
    -- filter=201 channel=28
    -3, 4, -4, -5, -6, 5, 5, -1, -7,
    -- filter=201 channel=29
    -2, 1, -5, 4, 7, -3, -2, -5, -3,
    -- filter=201 channel=30
    -2, -3, 1, 6, 6, 0, -5, 6, -2,
    -- filter=201 channel=31
    0, 4, -1, -1, -2, -2, -7, -1, 3,
    -- filter=201 channel=32
    3, -6, -6, -1, -4, -7, -3, -5, -3,
    -- filter=201 channel=33
    3, -5, -3, 5, -3, -4, -2, 0, -5,
    -- filter=201 channel=34
    6, 5, 7, 0, -2, -4, -4, -5, 5,
    -- filter=201 channel=35
    6, 1, 4, 0, 6, -5, 3, 1, 0,
    -- filter=201 channel=36
    -3, 0, -5, 0, -3, 2, 4, 2, -4,
    -- filter=201 channel=37
    5, 4, 5, 4, -3, 0, -7, -3, -5,
    -- filter=201 channel=38
    1, 2, 3, -4, 1, -4, -3, 2, -2,
    -- filter=201 channel=39
    5, -2, 0, -1, 0, -5, 0, -4, 1,
    -- filter=201 channel=40
    -7, 6, 4, 5, -1, 0, 0, 2, -3,
    -- filter=201 channel=41
    4, -5, -6, 5, -4, 2, 4, -6, -2,
    -- filter=201 channel=42
    -6, 7, 4, 1, 6, 0, 0, -7, 3,
    -- filter=201 channel=43
    -1, -1, -6, -3, 4, -5, 0, -3, 4,
    -- filter=201 channel=44
    2, -6, -7, 7, -1, 1, 1, 1, -5,
    -- filter=201 channel=45
    7, 5, -3, -3, 5, 4, -3, -2, 5,
    -- filter=201 channel=46
    -7, 3, 6, -6, -4, 2, 0, -5, 0,
    -- filter=201 channel=47
    -4, 3, -5, 4, -1, 3, -6, -2, 3,
    -- filter=201 channel=48
    -1, 2, -1, -6, 3, -2, -2, 4, 3,
    -- filter=201 channel=49
    -7, -2, 4, -5, -7, -1, -6, 0, -4,
    -- filter=201 channel=50
    -6, 5, 0, -5, 2, -5, -3, 4, -1,
    -- filter=201 channel=51
    5, -6, 5, 0, -3, 2, -7, 7, -4,
    -- filter=201 channel=52
    7, -3, -6, 2, 5, 4, -1, 5, -4,
    -- filter=201 channel=53
    -1, -3, -2, 6, 0, -4, 1, 0, 3,
    -- filter=201 channel=54
    2, 6, -3, 0, 5, -6, 1, 2, -5,
    -- filter=201 channel=55
    -7, -2, 5, 5, -1, 1, 3, -7, -6,
    -- filter=201 channel=56
    0, -7, 1, -3, 3, -6, 1, -1, 2,
    -- filter=201 channel=57
    0, -4, 1, 2, -5, 1, -4, -5, 6,
    -- filter=201 channel=58
    6, -6, 6, -3, -3, -6, -5, 0, 0,
    -- filter=201 channel=59
    4, -2, 0, -2, 3, 2, 6, -2, 0,
    -- filter=201 channel=60
    -3, 2, 0, -1, 0, -1, 1, -2, -3,
    -- filter=201 channel=61
    -3, -6, 0, 4, -7, -2, 7, -2, -2,
    -- filter=201 channel=62
    -1, 6, 0, -5, 2, -2, -1, 5, -6,
    -- filter=201 channel=63
    -1, -3, 0, 6, 0, -6, 5, -4, 6,
    -- filter=201 channel=64
    -4, -2, 4, -7, 7, -3, 0, -2, 6,
    -- filter=201 channel=65
    1, 0, -4, 2, -1, -6, -4, -1, 5,
    -- filter=201 channel=66
    4, -3, -1, -3, 3, 6, 6, -5, -5,
    -- filter=201 channel=67
    -5, -5, -1, 0, -2, 5, 6, -4, -7,
    -- filter=201 channel=68
    0, 0, -4, 2, -5, -5, 7, -6, 0,
    -- filter=201 channel=69
    0, -4, -5, -2, 0, -5, 5, 7, 6,
    -- filter=201 channel=70
    -4, -3, 4, -5, -2, 1, -1, 1, 0,
    -- filter=201 channel=71
    -1, 2, -7, 7, 2, 3, -5, -1, 6,
    -- filter=201 channel=72
    -2, -4, 2, 2, -3, 0, -6, 0, -6,
    -- filter=201 channel=73
    0, 4, 0, 4, -1, 2, 4, 2, 2,
    -- filter=201 channel=74
    -6, -1, -3, -6, 7, -5, -5, 2, -3,
    -- filter=201 channel=75
    5, -3, 4, 0, -1, -2, -3, 5, 6,
    -- filter=201 channel=76
    -1, 4, 0, 3, 3, 4, 0, 4, 1,
    -- filter=201 channel=77
    -6, 0, 1, 4, -1, 4, 1, 0, 6,
    -- filter=201 channel=78
    4, -4, 2, 7, 0, -3, -2, 1, -5,
    -- filter=201 channel=79
    4, -1, 3, -4, -5, -3, -2, -5, -2,
    -- filter=201 channel=80
    0, 2, 0, -2, -5, -5, 4, 4, -4,
    -- filter=201 channel=81
    0, 3, 0, 0, -3, -2, -5, -1, -4,
    -- filter=201 channel=82
    1, 0, -2, 0, -5, -6, -1, -6, 7,
    -- filter=201 channel=83
    4, -2, -1, 2, -4, 5, 0, -5, -1,
    -- filter=201 channel=84
    0, 3, -2, 2, 5, -7, 4, -2, 1,
    -- filter=201 channel=85
    0, 6, -6, 6, -3, 6, -6, -2, -3,
    -- filter=201 channel=86
    4, 2, 5, 3, 0, -1, -4, 0, -2,
    -- filter=201 channel=87
    -3, -4, 3, 1, -4, -1, 0, -5, -5,
    -- filter=201 channel=88
    -4, 4, 5, 7, -4, -2, 0, -6, -2,
    -- filter=201 channel=89
    -2, -6, 7, 6, 6, -7, 1, 0, 2,
    -- filter=201 channel=90
    -2, 0, -2, -4, 5, -6, 0, 4, 6,
    -- filter=201 channel=91
    -7, 5, 0, 0, 0, 2, 1, -1, -3,
    -- filter=201 channel=92
    3, 6, -1, -2, -5, 0, -3, 2, 7,
    -- filter=201 channel=93
    7, 6, 2, 1, -3, 1, 0, -7, -1,
    -- filter=201 channel=94
    -5, -2, 1, -3, 7, 3, -2, 4, -3,
    -- filter=201 channel=95
    6, 0, -3, 0, -3, -5, -5, -7, -1,
    -- filter=201 channel=96
    -2, 2, -1, 0, 6, -7, -4, 0, 0,
    -- filter=201 channel=97
    0, -4, -7, 3, 0, 3, 4, -2, -6,
    -- filter=201 channel=98
    0, -4, -5, 0, 3, 0, 6, -1, 0,
    -- filter=201 channel=99
    1, 0, -1, -5, -5, 3, -6, -6, 1,
    -- filter=201 channel=100
    2, 0, 4, 0, 0, 3, -6, -2, 6,
    -- filter=201 channel=101
    4, 3, -7, 2, 5, 1, 6, 7, -3,
    -- filter=201 channel=102
    3, 5, -6, -2, 3, 0, -2, -6, 4,
    -- filter=201 channel=103
    -3, 7, 2, -2, -2, -4, -5, 2, -2,
    -- filter=201 channel=104
    -5, 0, 6, -6, 6, -3, 0, -1, -1,
    -- filter=201 channel=105
    -5, -4, 6, 0, 6, 5, 0, -1, 4,
    -- filter=201 channel=106
    -2, 5, 1, 3, -1, 3, -5, -4, -1,
    -- filter=201 channel=107
    0, -1, 0, -1, -2, -6, 6, 0, 4,
    -- filter=201 channel=108
    -5, 0, -2, -4, -3, 7, -7, -4, -3,
    -- filter=201 channel=109
    5, 2, 2, -7, -3, -3, 2, 2, -1,
    -- filter=201 channel=110
    -6, -5, 0, 2, 0, -3, 1, 2, -6,
    -- filter=201 channel=111
    1, 6, 3, 6, 5, -6, -2, 0, -4,
    -- filter=201 channel=112
    6, 1, 0, -3, 1, -5, 0, 0, 0,
    -- filter=201 channel=113
    -4, 2, -6, 5, -2, -3, 1, 4, 5,
    -- filter=201 channel=114
    0, 6, -5, 3, -7, 6, -4, -2, -2,
    -- filter=201 channel=115
    -1, -2, 4, 4, 5, 3, 3, -6, 0,
    -- filter=201 channel=116
    2, -3, 1, 5, 0, -3, -3, 5, 3,
    -- filter=201 channel=117
    6, -6, 0, 4, 0, -7, 1, 3, 5,
    -- filter=201 channel=118
    -6, -4, -5, -2, 1, -4, 0, 7, 1,
    -- filter=201 channel=119
    -1, -2, 3, 3, -2, 3, 1, -5, -3,
    -- filter=201 channel=120
    2, 3, 7, 0, -4, 7, -7, 1, -6,
    -- filter=201 channel=121
    7, 2, 1, -5, -6, -5, 3, -2, 0,
    -- filter=201 channel=122
    0, -4, 1, -1, 3, -5, -2, -4, 0,
    -- filter=201 channel=123
    3, 3, 0, 1, -3, 0, -7, 6, 0,
    -- filter=201 channel=124
    6, 0, 5, 0, -3, -7, -7, -3, 1,
    -- filter=201 channel=125
    0, -2, 3, 6, -5, 1, 3, 0, -3,
    -- filter=201 channel=126
    -1, 3, -5, -6, -2, -5, -2, -3, 0,
    -- filter=201 channel=127
    0, 5, -5, 6, 5, 0, 4, 5, 5,
    -- filter=202 channel=0
    0, 7, -7, -6, -6, 3, 4, 3, -1,
    -- filter=202 channel=1
    1, 1, 0, -5, 2, -5, -6, 4, -4,
    -- filter=202 channel=2
    0, -2, 4, -4, 7, -6, -6, 3, 5,
    -- filter=202 channel=3
    0, 5, 5, 3, 1, 3, -2, 1, 4,
    -- filter=202 channel=4
    0, 0, 4, 3, -1, -4, 0, -2, -3,
    -- filter=202 channel=5
    -5, -1, 3, 2, 7, 0, 0, -5, -7,
    -- filter=202 channel=6
    1, 3, 7, -3, 7, 1, -5, 7, -4,
    -- filter=202 channel=7
    -7, 1, 4, -4, -6, -4, 3, 6, -1,
    -- filter=202 channel=8
    -4, -6, -5, 0, 0, 5, -4, -1, 0,
    -- filter=202 channel=9
    -6, -7, 4, 5, -2, 3, -5, 0, -1,
    -- filter=202 channel=10
    5, -4, 1, -1, 1, -6, 2, 1, -4,
    -- filter=202 channel=11
    -1, -3, 0, 6, 3, 6, -3, 5, -4,
    -- filter=202 channel=12
    4, 7, -5, -2, 2, -4, 0, 3, 7,
    -- filter=202 channel=13
    -5, 1, 0, 0, 3, 0, 0, 0, 6,
    -- filter=202 channel=14
    -3, 2, 5, -1, 4, -1, 6, -2, 0,
    -- filter=202 channel=15
    -3, -5, 1, 2, -1, -3, 0, 3, 2,
    -- filter=202 channel=16
    7, 3, -5, 2, 5, -1, -2, 3, 4,
    -- filter=202 channel=17
    -2, 4, -4, 4, -3, -1, -6, 6, -5,
    -- filter=202 channel=18
    -6, 0, -1, 2, 5, 5, 4, -6, -4,
    -- filter=202 channel=19
    7, -4, -2, 3, 2, 0, -2, 5, -7,
    -- filter=202 channel=20
    -3, -2, 5, -6, -4, -7, -5, -4, 1,
    -- filter=202 channel=21
    -4, -7, 2, 5, -3, 7, 0, 5, -1,
    -- filter=202 channel=22
    -1, -6, 5, -5, -1, -2, -6, 0, -4,
    -- filter=202 channel=23
    -1, -7, 0, 5, -3, -2, -4, -6, -3,
    -- filter=202 channel=24
    7, -4, 2, -1, 1, -2, -4, -3, 0,
    -- filter=202 channel=25
    3, 3, 2, -6, 6, -2, -1, 2, -1,
    -- filter=202 channel=26
    1, 1, 2, 6, 0, 1, 7, 2, 2,
    -- filter=202 channel=27
    -1, -1, -7, 1, -2, 4, -7, 0, -1,
    -- filter=202 channel=28
    -7, -6, 7, 3, -6, -3, 4, 0, 6,
    -- filter=202 channel=29
    6, -3, 0, 0, -3, 5, -1, -4, 4,
    -- filter=202 channel=30
    0, -7, -3, -4, 6, -4, 6, -3, -5,
    -- filter=202 channel=31
    4, -4, 3, -3, -4, -7, -5, -5, -4,
    -- filter=202 channel=32
    2, 0, 5, 1, 3, -2, -5, 1, -3,
    -- filter=202 channel=33
    0, 1, -5, 1, 3, 1, 6, 0, 6,
    -- filter=202 channel=34
    0, 4, -4, -2, 5, -6, 3, 0, -6,
    -- filter=202 channel=35
    -6, 1, 0, -4, 3, 3, -6, 3, 3,
    -- filter=202 channel=36
    1, 6, 5, -1, 4, -1, 0, 1, -1,
    -- filter=202 channel=37
    -7, 0, 1, 2, 6, -4, 5, -3, 5,
    -- filter=202 channel=38
    -6, 1, -3, 2, 4, 5, -4, -1, 5,
    -- filter=202 channel=39
    1, 0, -2, -5, -6, 4, 3, 4, -1,
    -- filter=202 channel=40
    3, 7, 3, 2, 5, 3, 3, -3, 4,
    -- filter=202 channel=41
    6, 0, 1, -6, 3, -6, -1, -3, 4,
    -- filter=202 channel=42
    -4, 7, -4, 1, 6, 1, 3, -6, 0,
    -- filter=202 channel=43
    -4, -7, 1, -2, -3, -5, 3, -6, 3,
    -- filter=202 channel=44
    -5, 0, 4, -5, 0, 0, 4, 2, 2,
    -- filter=202 channel=45
    -2, 2, -2, 3, -2, 4, 1, 3, -3,
    -- filter=202 channel=46
    7, 5, 6, 1, 4, 2, 7, 4, -2,
    -- filter=202 channel=47
    -7, 7, 5, -1, 5, -6, -1, 0, -6,
    -- filter=202 channel=48
    -2, -6, 0, 1, -1, -6, 6, -6, 1,
    -- filter=202 channel=49
    4, -5, -2, 6, -3, -4, 3, 0, 7,
    -- filter=202 channel=50
    -3, -7, 0, 0, -4, -1, -4, -7, 0,
    -- filter=202 channel=51
    0, 3, 1, -7, 1, -6, 6, 3, 2,
    -- filter=202 channel=52
    -7, 6, -6, -2, -2, -7, -7, 0, 0,
    -- filter=202 channel=53
    0, 6, -3, 4, 4, -4, -5, 5, -1,
    -- filter=202 channel=54
    3, 5, 1, -3, -3, -7, -1, -6, -7,
    -- filter=202 channel=55
    0, 2, 0, 0, 3, -6, -5, -1, -7,
    -- filter=202 channel=56
    2, 3, -5, 4, 6, 6, 5, -5, 0,
    -- filter=202 channel=57
    0, 3, 1, 0, 2, -6, 3, -1, 2,
    -- filter=202 channel=58
    -5, 0, 0, 0, -6, -6, 3, 6, 5,
    -- filter=202 channel=59
    -6, 0, 3, -1, 0, -4, -2, 6, 5,
    -- filter=202 channel=60
    -1, 6, 1, -6, -1, -3, -5, 1, 1,
    -- filter=202 channel=61
    4, -7, 0, 4, 0, 6, 4, -4, -1,
    -- filter=202 channel=62
    3, -1, -6, -7, 1, 7, -3, -1, -3,
    -- filter=202 channel=63
    2, -2, -1, 1, -5, -4, -7, -7, 1,
    -- filter=202 channel=64
    -2, -3, 0, 6, -3, -6, -3, 7, -3,
    -- filter=202 channel=65
    0, -6, 1, 1, 0, 4, -6, -2, 0,
    -- filter=202 channel=66
    6, -5, 5, -4, 4, -3, -1, -3, -5,
    -- filter=202 channel=67
    3, 5, -5, -6, 3, -4, 0, 0, -6,
    -- filter=202 channel=68
    -2, -7, 6, 2, 6, -7, 5, 2, 4,
    -- filter=202 channel=69
    -5, 4, 4, 2, 3, -5, 3, 1, 4,
    -- filter=202 channel=70
    -5, -7, 0, 1, -3, 2, 7, 5, -5,
    -- filter=202 channel=71
    4, 4, 6, -2, -7, -5, -4, -3, -6,
    -- filter=202 channel=72
    -5, 2, -6, -7, 7, 2, -3, 1, -5,
    -- filter=202 channel=73
    3, 0, -6, 2, -4, 6, -7, -6, -2,
    -- filter=202 channel=74
    -2, -4, -5, 0, -2, 3, -3, 7, 5,
    -- filter=202 channel=75
    3, -3, -7, 1, -3, -5, 0, -2, 0,
    -- filter=202 channel=76
    0, 5, -7, 6, 0, -4, 0, 1, -1,
    -- filter=202 channel=77
    -2, -6, 7, -2, -1, 6, 1, -5, -4,
    -- filter=202 channel=78
    1, -4, -1, -5, 1, -4, -4, 7, -2,
    -- filter=202 channel=79
    2, 4, -6, -3, 7, 4, 1, -6, 2,
    -- filter=202 channel=80
    6, -2, 5, 2, -6, -2, 7, 0, 0,
    -- filter=202 channel=81
    -7, 0, -7, 6, -6, -1, -5, 3, -6,
    -- filter=202 channel=82
    -3, 0, -4, 2, 0, 2, 5, -3, -6,
    -- filter=202 channel=83
    0, 7, -5, -6, 3, -3, -6, 5, -4,
    -- filter=202 channel=84
    -7, 5, 0, 0, 2, 0, -2, 1, 0,
    -- filter=202 channel=85
    -4, 4, -7, 0, -4, 0, -3, 3, 3,
    -- filter=202 channel=86
    3, -4, -1, 6, -5, 4, -2, -3, -1,
    -- filter=202 channel=87
    -4, 0, -5, -4, 5, -5, 6, 2, 0,
    -- filter=202 channel=88
    0, -2, -2, -6, 1, 6, 1, 0, -4,
    -- filter=202 channel=89
    -2, 0, 5, -5, -4, 5, -6, -3, 4,
    -- filter=202 channel=90
    -4, -6, 0, -5, 3, 3, -2, 0, 5,
    -- filter=202 channel=91
    2, -4, 5, 4, 0, -3, -3, -3, 0,
    -- filter=202 channel=92
    5, 5, 4, 3, -6, 3, -5, -4, -4,
    -- filter=202 channel=93
    -3, 1, -1, -3, -5, 0, 3, 0, -1,
    -- filter=202 channel=94
    -1, 6, 0, -1, 3, 0, -1, 6, 0,
    -- filter=202 channel=95
    7, -6, 6, 0, -7, 0, -4, -5, 6,
    -- filter=202 channel=96
    5, 0, -1, -6, -6, 2, 2, -4, -7,
    -- filter=202 channel=97
    -1, 4, 4, -4, 7, -5, 4, -3, 2,
    -- filter=202 channel=98
    0, -1, 5, -3, -3, 1, 2, -1, 6,
    -- filter=202 channel=99
    4, -2, 0, 3, -1, -5, -4, -1, -1,
    -- filter=202 channel=100
    0, 0, 3, -4, -4, -6, -4, -2, 2,
    -- filter=202 channel=101
    5, 4, 0, 3, -4, 6, -7, 4, -7,
    -- filter=202 channel=102
    0, 1, 1, -7, 2, 3, -4, 7, -1,
    -- filter=202 channel=103
    6, -5, -2, 0, -7, 3, 2, -1, 0,
    -- filter=202 channel=104
    6, 6, 5, -4, -6, 2, 0, 0, 2,
    -- filter=202 channel=105
    -5, 7, -7, 1, 2, 2, -1, 3, 4,
    -- filter=202 channel=106
    3, 0, -2, 3, 0, 2, 0, 4, -4,
    -- filter=202 channel=107
    -1, 2, 5, 0, 6, 4, -5, 6, 0,
    -- filter=202 channel=108
    -3, 1, 1, 5, -4, 3, -1, -1, 5,
    -- filter=202 channel=109
    1, -5, 0, 1, 0, 7, 5, -1, 5,
    -- filter=202 channel=110
    -2, 3, -6, 0, -5, 4, 0, -4, 5,
    -- filter=202 channel=111
    1, -2, -1, 6, -7, 0, -2, 0, 7,
    -- filter=202 channel=112
    6, 5, 1, 3, -6, 0, -4, 0, -4,
    -- filter=202 channel=113
    -6, -5, 0, 5, 2, 2, 1, 0, -6,
    -- filter=202 channel=114
    5, 0, 1, -7, 1, 0, 1, 1, -5,
    -- filter=202 channel=115
    -4, -4, -3, 1, -3, 4, -1, 6, 0,
    -- filter=202 channel=116
    2, -5, -4, 0, -3, 6, -6, -3, -5,
    -- filter=202 channel=117
    -3, 7, 2, -3, -3, 6, 4, 0, -3,
    -- filter=202 channel=118
    0, -2, 0, 3, 0, 3, 3, -5, 1,
    -- filter=202 channel=119
    2, 0, -1, 5, 5, -7, -3, -6, 7,
    -- filter=202 channel=120
    1, -4, -3, -2, 0, 0, 2, -4, -4,
    -- filter=202 channel=121
    -4, -5, 7, 1, 5, -7, -3, -2, 0,
    -- filter=202 channel=122
    1, -4, -1, -3, 5, 0, 1, -1, -7,
    -- filter=202 channel=123
    -1, -6, 1, -3, -3, 0, -2, -5, 2,
    -- filter=202 channel=124
    1, -2, 7, 5, 0, -7, 0, 3, -5,
    -- filter=202 channel=125
    -3, -7, 2, -7, 2, -7, 7, 3, -5,
    -- filter=202 channel=126
    -3, 6, -2, -7, -2, 0, 6, 5, 0,
    -- filter=202 channel=127
    0, -1, 5, 0, -6, -6, -1, 0, -4,
    -- filter=203 channel=0
    -5, -5, -3, -3, -3, 0, 7, -6, -7,
    -- filter=203 channel=1
    -3, -5, -9, -4, -3, 1, -4, 1, 7,
    -- filter=203 channel=2
    -4, -3, 6, -3, 4, -5, -9, -8, -3,
    -- filter=203 channel=3
    6, -8, 4, 3, -4, 1, 2, -4, -7,
    -- filter=203 channel=4
    3, 3, -3, -3, -1, -5, -5, -13, 2,
    -- filter=203 channel=5
    -3, -5, -1, 0, 2, -1, -4, 6, 3,
    -- filter=203 channel=6
    -7, 6, 1, 7, 6, -2, -6, 0, -4,
    -- filter=203 channel=7
    -5, 6, 3, -2, -6, 3, 5, -4, -4,
    -- filter=203 channel=8
    -7, -1, 0, 0, -4, -6, 3, -1, 4,
    -- filter=203 channel=9
    7, 4, 5, 1, -7, 6, 4, 8, -5,
    -- filter=203 channel=10
    1, -3, -4, 1, 11, -8, -4, 1, -7,
    -- filter=203 channel=11
    6, 0, 3, 0, 0, 6, 2, 6, 5,
    -- filter=203 channel=12
    5, 0, -1, -8, -2, -6, -6, 3, -2,
    -- filter=203 channel=13
    -2, 0, -6, -14, 14, 1, -9, 11, 1,
    -- filter=203 channel=14
    -6, -2, 0, 2, -6, -4, -2, -4, 3,
    -- filter=203 channel=15
    4, -4, -6, -5, 2, -7, -5, 1, -5,
    -- filter=203 channel=16
    -4, -1, -4, 1, -1, -7, 6, 7, 0,
    -- filter=203 channel=17
    -3, -1, -3, 1, 5, 2, 0, -6, 3,
    -- filter=203 channel=18
    6, 10, -8, -10, 20, -10, -10, 13, -3,
    -- filter=203 channel=19
    2, -7, -4, 1, 3, 3, -4, 0, 3,
    -- filter=203 channel=20
    5, -5, 6, -8, 6, -8, -10, 6, 0,
    -- filter=203 channel=21
    0, 2, 6, -6, -8, 3, 5, -4, 8,
    -- filter=203 channel=22
    4, 0, -1, 7, 6, -5, 1, 7, -4,
    -- filter=203 channel=23
    2, 0, -6, 10, 11, 0, -5, 17, -14,
    -- filter=203 channel=24
    5, -3, -4, -2, -2, 1, -3, -4, 4,
    -- filter=203 channel=25
    -1, 3, 1, -11, 6, -10, -14, 11, -2,
    -- filter=203 channel=26
    6, 0, 5, -4, 4, -3, -1, -4, 2,
    -- filter=203 channel=27
    6, -5, -2, -4, 13, -10, -19, 15, 4,
    -- filter=203 channel=28
    6, -4, 1, 6, -5, -5, 5, 4, 0,
    -- filter=203 channel=29
    1, 6, 6, -9, 5, 6, -3, 2, -7,
    -- filter=203 channel=30
    7, -2, -6, 3, -4, -5, -8, 5, 1,
    -- filter=203 channel=31
    -6, 0, 7, -8, 2, -7, -4, 7, 1,
    -- filter=203 channel=32
    2, -2, -2, -10, 16, 0, -17, 19, 2,
    -- filter=203 channel=33
    3, -2, 0, -7, 13, -7, -8, 9, -6,
    -- filter=203 channel=34
    -1, -9, -8, 18, -5, -6, 10, 1, -12,
    -- filter=203 channel=35
    4, 2, 0, 2, 0, 4, 4, 3, 4,
    -- filter=203 channel=36
    0, 2, 6, 0, -6, 5, 1, -7, -4,
    -- filter=203 channel=37
    -2, 1, 4, 0, -8, -4, 0, 4, -3,
    -- filter=203 channel=38
    5, 0, -4, -3, 5, -7, -11, 9, -6,
    -- filter=203 channel=39
    -5, 7, 4, 3, 6, -1, -8, -1, -5,
    -- filter=203 channel=40
    6, -5, -4, 6, 1, 4, 0, 3, -2,
    -- filter=203 channel=41
    4, 6, -9, 0, 15, -8, 7, 9, 0,
    -- filter=203 channel=42
    -5, 3, 7, -3, -2, -3, -1, -6, 1,
    -- filter=203 channel=43
    -8, 3, -5, 5, 3, -4, 3, -3, -10,
    -- filter=203 channel=44
    -3, -1, -2, -3, -4, 4, 5, -2, -4,
    -- filter=203 channel=45
    3, 5, -5, 2, 3, -3, -3, 3, -7,
    -- filter=203 channel=46
    -5, 1, -3, 0, 6, -3, 7, -6, -1,
    -- filter=203 channel=47
    5, 1, 5, 5, -6, -2, 1, -8, 2,
    -- filter=203 channel=48
    0, 0, 4, -8, -4, -6, -8, -3, 11,
    -- filter=203 channel=49
    -3, 9, 0, 0, 0, -1, -13, -3, 6,
    -- filter=203 channel=50
    1, 3, -6, -2, 4, -1, -8, 3, 3,
    -- filter=203 channel=51
    -1, 0, 0, -6, -2, -3, 0, 5, 3,
    -- filter=203 channel=52
    -2, -3, -3, 3, 3, 3, 4, 13, 1,
    -- filter=203 channel=53
    -3, 1, -5, 5, 2, 4, -3, 10, -5,
    -- filter=203 channel=54
    -6, -1, 0, 3, 2, -6, 5, 4, 0,
    -- filter=203 channel=55
    -1, 6, -4, 1, 16, -11, -15, 3, -9,
    -- filter=203 channel=56
    4, 2, 0, 5, 6, 1, -2, 2, -5,
    -- filter=203 channel=57
    -5, 1, 0, -5, 5, -7, -5, 1, -6,
    -- filter=203 channel=58
    7, -7, 7, 5, -5, 0, 7, 0, -1,
    -- filter=203 channel=59
    -6, 0, 8, -8, 9, -4, -14, 11, 1,
    -- filter=203 channel=60
    7, -1, 7, 4, -1, -5, 0, -1, -4,
    -- filter=203 channel=61
    0, 0, -6, -5, 0, -3, 3, 7, 6,
    -- filter=203 channel=62
    -4, 5, -5, 0, 0, -2, 2, 0, -6,
    -- filter=203 channel=63
    5, -1, 1, 0, 2, 2, 5, 0, 8,
    -- filter=203 channel=64
    4, 4, 6, 3, -1, 2, 8, -3, -6,
    -- filter=203 channel=65
    1, -3, 7, 6, 1, 6, -4, -7, -2,
    -- filter=203 channel=66
    5, 1, 2, -1, 6, 1, 2, 11, 3,
    -- filter=203 channel=67
    2, 5, -3, 1, -5, 3, 6, -6, -4,
    -- filter=203 channel=68
    0, -3, -4, -9, 0, -1, 4, 1, 7,
    -- filter=203 channel=69
    1, 0, 5, -4, 5, -1, -6, 0, -5,
    -- filter=203 channel=70
    3, -8, 1, 4, 1, -4, 0, 7, -3,
    -- filter=203 channel=71
    -1, -8, 5, -5, -1, -3, -1, -2, -5,
    -- filter=203 channel=72
    4, 4, 5, -10, 1, -1, -5, 0, 5,
    -- filter=203 channel=73
    3, -3, -7, -3, 5, -9, -3, 10, 7,
    -- filter=203 channel=74
    7, -5, -4, -5, 7, -8, -9, 12, -9,
    -- filter=203 channel=75
    6, 0, -1, 0, -1, 4, 0, -1, 1,
    -- filter=203 channel=76
    2, -2, 4, 0, 5, -1, -10, 4, -6,
    -- filter=203 channel=77
    -6, -1, -7, -4, 0, 1, -1, -2, 0,
    -- filter=203 channel=78
    -2, -2, -5, -1, -6, 0, 5, 2, -1,
    -- filter=203 channel=79
    -4, -1, 4, -12, 19, 0, -22, 17, -3,
    -- filter=203 channel=80
    2, 1, 6, -14, 4, -4, -17, 6, -2,
    -- filter=203 channel=81
    -6, 1, 6, 7, 0, 3, 6, 4, -7,
    -- filter=203 channel=82
    3, 4, 6, 7, 0, 1, 0, -1, -8,
    -- filter=203 channel=83
    0, 3, -6, 4, -7, 4, -2, -2, 11,
    -- filter=203 channel=84
    0, -2, -1, -10, 9, 0, 0, 1, 0,
    -- filter=203 channel=85
    5, -6, -2, -6, -4, 0, 5, 0, 4,
    -- filter=203 channel=86
    4, -3, -7, -6, -2, -2, 0, 5, -6,
    -- filter=203 channel=87
    0, 2, -1, 6, 0, 3, -4, 1, -10,
    -- filter=203 channel=88
    2, -2, -3, 0, -8, -3, 3, 6, -6,
    -- filter=203 channel=89
    0, 4, 4, -8, 14, 1, -11, 5, -4,
    -- filter=203 channel=90
    6, -5, -2, 0, -7, -2, 5, 5, -5,
    -- filter=203 channel=91
    7, 0, 0, -12, 11, -5, -17, 6, 4,
    -- filter=203 channel=92
    -2, 4, -4, 8, -7, 0, -2, 3, -8,
    -- filter=203 channel=93
    7, 2, 6, 2, 4, 1, 2, -4, 6,
    -- filter=203 channel=94
    -3, -6, -2, -6, 4, 0, 4, 0, -1,
    -- filter=203 channel=95
    5, -3, -5, 4, 4, 6, 0, 0, -5,
    -- filter=203 channel=96
    0, 0, 2, 1, 0, 0, 4, 3, 7,
    -- filter=203 channel=97
    1, 4, -2, -4, 0, 2, -6, -4, 2,
    -- filter=203 channel=98
    -5, 4, 0, -6, 15, -3, -6, 2, -7,
    -- filter=203 channel=99
    5, 0, -1, 1, 0, -13, -6, 12, -10,
    -- filter=203 channel=100
    8, -3, 2, 0, -5, -3, 6, 2, 0,
    -- filter=203 channel=101
    -4, -2, -2, -10, 4, -6, 0, -11, 3,
    -- filter=203 channel=102
    -5, 6, 0, -2, 5, 6, -7, -4, 7,
    -- filter=203 channel=103
    -4, 0, -1, 2, -3, -3, -7, -2, 1,
    -- filter=203 channel=104
    1, 4, -2, -11, 2, -3, -5, 0, 9,
    -- filter=203 channel=105
    -6, 2, -4, 0, 0, -2, -2, 5, 0,
    -- filter=203 channel=106
    -2, -6, -1, 5, 7, -3, -6, -9, 0,
    -- filter=203 channel=107
    0, -8, -6, 4, 2, -1, -5, 11, 3,
    -- filter=203 channel=108
    -7, -3, 1, 6, 4, -6, 5, -2, 6,
    -- filter=203 channel=109
    -2, 7, -1, 0, 19, -1, -17, 19, 0,
    -- filter=203 channel=110
    8, -6, -3, 1, 2, -6, -9, 4, 1,
    -- filter=203 channel=111
    -6, 6, -1, 4, 4, 6, 1, 2, 0,
    -- filter=203 channel=112
    -6, 1, -6, 0, 6, -2, 3, 6, 3,
    -- filter=203 channel=113
    1, -4, -4, 1, -4, -1, -9, 2, -7,
    -- filter=203 channel=114
    1, 6, -4, -15, 13, -5, -14, 12, 7,
    -- filter=203 channel=115
    2, -1, 3, 5, 8, -5, -6, -3, 3,
    -- filter=203 channel=116
    5, 10, 3, -9, 10, -4, -3, 10, 5,
    -- filter=203 channel=117
    0, 1, -2, 0, -2, -4, 0, 0, 5,
    -- filter=203 channel=118
    -6, -7, 3, 1, -4, -2, -1, 2, 0,
    -- filter=203 channel=119
    6, 3, 2, 13, -5, 0, 5, 6, -1,
    -- filter=203 channel=120
    2, -7, -6, -8, 9, -5, -10, 15, -9,
    -- filter=203 channel=121
    0, -2, 1, -4, 11, 2, -1, -1, -8,
    -- filter=203 channel=122
    -5, -4, 9, 0, -6, 4, 4, 1, 5,
    -- filter=203 channel=123
    6, -5, -6, 10, 3, -5, -1, 2, 3,
    -- filter=203 channel=124
    2, 4, -4, -6, 4, -5, -9, -1, -1,
    -- filter=203 channel=125
    -2, -1, 0, -6, 3, -8, -15, 10, 1,
    -- filter=203 channel=126
    -2, 7, 3, -8, 12, -5, -10, 1, -2,
    -- filter=203 channel=127
    -3, 0, 0, 4, -4, 3, -2, -2, 4,
    -- filter=204 channel=0
    3, -6, 6, 6, 0, 0, -2, -4, 0,
    -- filter=204 channel=1
    7, 0, 2, -2, 5, 2, 3, -1, -2,
    -- filter=204 channel=2
    1, -6, -1, -1, -4, 1, -4, 0, -6,
    -- filter=204 channel=3
    7, -1, -4, -4, -2, 0, 2, -5, -5,
    -- filter=204 channel=4
    2, 6, 2, -2, 4, 0, 3, 7, -1,
    -- filter=204 channel=5
    -7, 6, -6, 1, -7, 3, -3, 6, 4,
    -- filter=204 channel=6
    0, 0, 1, 0, 5, -2, -7, 4, 5,
    -- filter=204 channel=7
    1, -1, -4, 0, -2, 4, -5, 0, -1,
    -- filter=204 channel=8
    7, 4, 0, -2, -1, 1, -4, 1, 6,
    -- filter=204 channel=9
    5, -6, 5, -4, -6, 3, -4, -6, 1,
    -- filter=204 channel=10
    4, -4, -3, 0, 6, 0, 2, -1, 5,
    -- filter=204 channel=11
    2, -5, -3, -6, -2, -7, 2, -8, -2,
    -- filter=204 channel=12
    -5, -6, 0, 0, 0, -6, -1, 6, -1,
    -- filter=204 channel=13
    -5, -6, 2, 1, 7, -6, 1, -3, 3,
    -- filter=204 channel=14
    1, 0, 7, -5, -2, 1, -4, -2, 6,
    -- filter=204 channel=15
    -1, 5, -2, -5, 0, -1, 1, -4, 0,
    -- filter=204 channel=16
    5, 2, 4, -5, 0, -4, 6, 6, 5,
    -- filter=204 channel=17
    6, -6, -1, 0, -1, 5, 3, 6, -3,
    -- filter=204 channel=18
    -2, 2, 5, 3, 5, 0, -3, -2, 3,
    -- filter=204 channel=19
    7, 7, -6, 0, -3, 3, 0, 5, 5,
    -- filter=204 channel=20
    3, 6, -3, -6, 0, -5, 0, 2, -2,
    -- filter=204 channel=21
    -6, -3, -5, 4, -4, -5, -6, 3, 2,
    -- filter=204 channel=22
    -3, 3, 1, 6, -7, -3, -1, 3, 4,
    -- filter=204 channel=23
    -4, 6, -6, -2, 5, 2, -2, 0, -4,
    -- filter=204 channel=24
    -2, -3, 2, -7, 6, 1, -2, 2, 5,
    -- filter=204 channel=25
    2, 7, -7, 1, 1, -3, 0, -1, 1,
    -- filter=204 channel=26
    2, -5, 2, 5, 0, -3, -1, 0, -4,
    -- filter=204 channel=27
    -5, 1, 0, -7, -4, 1, -4, 6, 3,
    -- filter=204 channel=28
    -3, -1, -6, -3, -4, -2, 0, -4, 6,
    -- filter=204 channel=29
    1, -5, 0, 2, -4, 6, -8, -7, -1,
    -- filter=204 channel=30
    2, 6, 6, 4, 0, -5, -1, -5, -1,
    -- filter=204 channel=31
    0, 4, 5, -3, 0, -6, -5, 1, 7,
    -- filter=204 channel=32
    -2, 3, -6, -4, -4, 4, 1, 5, 3,
    -- filter=204 channel=33
    -6, -2, -2, 0, -3, -1, 5, 5, 1,
    -- filter=204 channel=34
    6, 1, 0, -2, 4, 5, 1, 3, 3,
    -- filter=204 channel=35
    0, 6, 4, -5, -3, -3, -4, -2, -2,
    -- filter=204 channel=36
    4, 3, -4, 6, -3, -7, -4, -1, -6,
    -- filter=204 channel=37
    -1, -4, -7, -2, -4, -2, -4, -7, -6,
    -- filter=204 channel=38
    0, 0, -7, -4, 0, 0, 6, -7, 6,
    -- filter=204 channel=39
    0, 4, -1, 1, -2, -6, 4, -4, -2,
    -- filter=204 channel=40
    -7, 7, -6, -2, 2, -2, 4, 2, -3,
    -- filter=204 channel=41
    -6, 2, 0, 6, 6, 4, -4, 0, 6,
    -- filter=204 channel=42
    -2, 3, 5, 4, -1, -5, -1, -3, -2,
    -- filter=204 channel=43
    -1, 5, 0, -5, -2, -6, -4, -1, -6,
    -- filter=204 channel=44
    -2, -6, 1, -6, -4, -2, -6, -3, -7,
    -- filter=204 channel=45
    0, 5, -3, -4, -3, 4, -7, 1, 3,
    -- filter=204 channel=46
    1, -7, 6, -2, 0, -2, 2, 5, 3,
    -- filter=204 channel=47
    2, -6, 5, -7, -5, -4, -3, 1, -5,
    -- filter=204 channel=48
    -3, 3, 7, -2, 1, 1, 2, -2, -5,
    -- filter=204 channel=49
    5, -3, -6, -4, 1, 5, 2, 0, 3,
    -- filter=204 channel=50
    0, 5, -5, 5, 5, 3, -2, -1, -7,
    -- filter=204 channel=51
    -4, -4, -5, 0, -2, 4, 0, -6, -4,
    -- filter=204 channel=52
    6, -4, -3, -7, 3, 5, 4, 0, 0,
    -- filter=204 channel=53
    7, 5, 0, -1, 3, 0, -2, -4, 4,
    -- filter=204 channel=54
    -5, -6, 5, 2, 0, 5, -2, 5, 0,
    -- filter=204 channel=55
    3, -3, 6, -1, -5, -1, -7, 5, -1,
    -- filter=204 channel=56
    -6, 1, -5, -1, 3, 0, 5, -4, -7,
    -- filter=204 channel=57
    -3, 5, 3, -5, -1, 4, 5, 5, 3,
    -- filter=204 channel=58
    1, 3, -4, 0, -3, -2, -1, 0, -2,
    -- filter=204 channel=59
    2, -6, -1, 5, -2, -2, 1, 2, -7,
    -- filter=204 channel=60
    6, 2, 5, 2, 5, 7, 5, -1, 0,
    -- filter=204 channel=61
    7, 5, -2, 1, -1, -5, 0, -4, 0,
    -- filter=204 channel=62
    -7, -4, -3, 1, 4, -1, 4, 5, 0,
    -- filter=204 channel=63
    6, 0, 6, 3, -7, -1, 3, 0, 6,
    -- filter=204 channel=64
    3, -7, 0, 6, -7, -3, -3, 5, 7,
    -- filter=204 channel=65
    0, 0, 5, -6, -2, 7, -3, 7, 5,
    -- filter=204 channel=66
    1, 4, -5, -2, -6, -4, -5, -4, -3,
    -- filter=204 channel=67
    1, 5, 0, 2, -3, -6, -2, -7, 5,
    -- filter=204 channel=68
    6, -3, 0, 7, -5, -6, -2, 0, 1,
    -- filter=204 channel=69
    0, 7, 3, 0, -6, 2, -5, -6, 0,
    -- filter=204 channel=70
    3, 0, 2, 5, -3, -7, 6, 2, -4,
    -- filter=204 channel=71
    -4, -5, -1, -3, -2, -4, 6, 5, -5,
    -- filter=204 channel=72
    2, -4, 0, 0, 3, 5, -6, 7, 6,
    -- filter=204 channel=73
    -6, 5, -5, 6, -8, -4, -3, -4, -1,
    -- filter=204 channel=74
    0, 2, 5, 1, 0, 1, 7, -4, 4,
    -- filter=204 channel=75
    2, 2, 4, 0, 2, 2, -5, 0, -4,
    -- filter=204 channel=76
    4, -4, 2, -1, -5, 1, -5, -6, -1,
    -- filter=204 channel=77
    3, -5, -6, -1, 0, -4, 3, -2, 2,
    -- filter=204 channel=78
    -7, -3, -1, 3, -5, 5, -5, 5, -2,
    -- filter=204 channel=79
    3, -8, -6, -5, 5, 3, 0, -2, -5,
    -- filter=204 channel=80
    -4, -4, -1, -2, 3, -1, 7, 3, -2,
    -- filter=204 channel=81
    2, 6, 3, 2, -7, 5, -5, -1, -2,
    -- filter=204 channel=82
    6, 6, 2, -7, -2, 2, 3, -7, 6,
    -- filter=204 channel=83
    -5, -4, -3, 1, -2, 3, 2, 4, -5,
    -- filter=204 channel=84
    0, 4, 4, -6, 6, -5, 6, 3, 5,
    -- filter=204 channel=85
    -1, -2, 0, 3, -1, 2, 4, -5, -4,
    -- filter=204 channel=86
    -2, -3, -4, -3, -2, -3, 0, 6, -1,
    -- filter=204 channel=87
    -5, 4, -6, 5, 0, -4, -7, 6, 4,
    -- filter=204 channel=88
    6, 0, 7, 1, -7, -6, -1, 5, -2,
    -- filter=204 channel=89
    2, 3, 5, 4, 4, -1, 6, -2, -5,
    -- filter=204 channel=90
    2, -5, 1, 6, -6, -2, 4, -7, -4,
    -- filter=204 channel=91
    -3, 1, 5, -7, 0, 5, 2, -6, 3,
    -- filter=204 channel=92
    4, -4, 0, 3, -7, 3, -3, 0, 3,
    -- filter=204 channel=93
    -3, -6, -1, -7, -6, -7, 0, -5, 0,
    -- filter=204 channel=94
    2, -5, -6, -2, -5, -2, 3, 0, -2,
    -- filter=204 channel=95
    0, 4, 5, 1, 0, 3, 0, -1, -2,
    -- filter=204 channel=96
    -5, 5, 7, -2, 7, 6, 2, 3, -5,
    -- filter=204 channel=97
    -4, 0, 5, -7, -6, -3, -4, 3, 0,
    -- filter=204 channel=98
    1, -7, -4, 1, -7, 4, -7, -4, 3,
    -- filter=204 channel=99
    2, 2, 0, 4, -4, 0, -2, 4, 6,
    -- filter=204 channel=100
    1, -6, -5, -1, -1, -6, 3, 5, 6,
    -- filter=204 channel=101
    5, 5, 7, -4, 4, -1, -3, -1, 1,
    -- filter=204 channel=102
    -1, 5, -1, -6, -6, 6, 6, -5, -5,
    -- filter=204 channel=103
    -7, 7, -1, 4, -7, -5, -7, -3, 3,
    -- filter=204 channel=104
    6, -7, 1, 6, -5, 5, 5, 0, 7,
    -- filter=204 channel=105
    5, -2, 0, -2, 2, 6, -4, -3, 6,
    -- filter=204 channel=106
    1, 7, -1, -1, 4, -3, -6, 1, -6,
    -- filter=204 channel=107
    1, -2, 4, -2, -4, 2, -5, 0, 6,
    -- filter=204 channel=108
    5, 4, 6, -5, -6, 4, -2, 0, -5,
    -- filter=204 channel=109
    -6, 3, 4, 4, 2, -5, 3, -6, 6,
    -- filter=204 channel=110
    -6, -4, -5, -3, 1, 0, -6, 1, -4,
    -- filter=204 channel=111
    -5, -3, 3, 4, -2, 3, 0, 2, 5,
    -- filter=204 channel=112
    -5, 0, -7, 6, -1, 2, 1, 2, 7,
    -- filter=204 channel=113
    6, 0, -7, -4, -7, 1, -4, 4, 0,
    -- filter=204 channel=114
    -5, 0, -3, -7, 0, 1, 1, -5, -7,
    -- filter=204 channel=115
    1, 2, -5, -2, 0, -1, 1, 7, -5,
    -- filter=204 channel=116
    -7, -7, -4, -5, -6, 1, 2, 5, 6,
    -- filter=204 channel=117
    6, -4, -5, 3, 0, 6, -5, 7, -7,
    -- filter=204 channel=118
    -4, 0, -2, -4, 3, 2, 4, 5, 6,
    -- filter=204 channel=119
    -6, 0, 1, 6, -4, -3, 6, -7, 3,
    -- filter=204 channel=120
    1, 1, -5, 1, -6, -7, -4, 5, 0,
    -- filter=204 channel=121
    -6, 2, -2, 0, 4, 0, -6, 5, 6,
    -- filter=204 channel=122
    -2, 1, 2, 3, -1, -4, -2, 1, 0,
    -- filter=204 channel=123
    -6, 7, -3, 7, 2, -3, 0, -4, -5,
    -- filter=204 channel=124
    -5, 0, -4, -4, 3, -3, 3, 5, 0,
    -- filter=204 channel=125
    2, -6, 6, -7, 2, -7, 3, 4, -4,
    -- filter=204 channel=126
    0, -5, 2, 2, 1, 0, 1, -3, 2,
    -- filter=204 channel=127
    0, 3, 5, 3, 1, 0, -1, 6, -5,
    -- filter=205 channel=0
    -18, -1, -1, -5, 0, 4, 0, 11, 14,
    -- filter=205 channel=1
    -15, -5, 5, -7, 11, 10, 0, 5, 0,
    -- filter=205 channel=2
    -3, 4, -8, -5, 5, 4, 4, -4, -7,
    -- filter=205 channel=3
    -9, 0, 9, -3, -2, 9, -1, 8, 7,
    -- filter=205 channel=4
    4, -6, -2, -12, -4, 0, -11, -6, 0,
    -- filter=205 channel=5
    -17, -9, -4, -2, 5, 18, 6, 14, 12,
    -- filter=205 channel=6
    10, 8, -3, 6, -6, -5, 1, -5, -5,
    -- filter=205 channel=7
    -2, -7, 0, 1, 0, 7, -4, -6, 1,
    -- filter=205 channel=8
    2, 0, 0, -5, -2, 1, -7, -2, -7,
    -- filter=205 channel=9
    6, 0, -5, 2, 8, 4, -3, 9, 7,
    -- filter=205 channel=10
    9, 7, -5, 9, 3, -1, 1, 0, -12,
    -- filter=205 channel=11
    13, 5, 10, 8, -9, -9, -1, -4, 2,
    -- filter=205 channel=12
    -6, 2, 1, -8, 6, -9, 4, -4, -1,
    -- filter=205 channel=13
    -3, 8, 0, 6, 3, -12, 3, -4, -10,
    -- filter=205 channel=14
    0, 2, -5, -3, 5, 5, -7, 6, 3,
    -- filter=205 channel=15
    11, 10, 2, 4, 0, -13, 4, -12, -2,
    -- filter=205 channel=16
    -10, 0, -8, -1, 1, -2, 0, 11, 9,
    -- filter=205 channel=17
    -6, 6, 2, 5, -3, 0, 2, 0, 1,
    -- filter=205 channel=18
    11, 11, 6, 2, 0, -10, 0, -11, -7,
    -- filter=205 channel=19
    -4, 2, -3, -1, 2, 2, 2, 0, -2,
    -- filter=205 channel=20
    18, 17, 14, 10, -11, -8, 2, -15, 2,
    -- filter=205 channel=21
    -3, 6, 0, 9, 14, -3, -1, 8, 5,
    -- filter=205 channel=22
    -8, -7, 2, 3, 1, -1, -5, -8, -2,
    -- filter=205 channel=23
    15, 15, -12, 8, -17, -14, -5, -10, -12,
    -- filter=205 channel=24
    3, 0, -5, -7, 6, 0, 0, -5, 7,
    -- filter=205 channel=25
    1, 9, -10, 5, 12, -9, 6, -3, -5,
    -- filter=205 channel=26
    -5, 2, -3, 4, -2, -2, -5, 7, -3,
    -- filter=205 channel=27
    13, 7, -4, 12, -10, -6, -3, -9, -9,
    -- filter=205 channel=28
    -2, -3, 3, 2, -6, 1, -1, 3, 1,
    -- filter=205 channel=29
    12, 14, 12, 12, -6, -10, 8, -11, 4,
    -- filter=205 channel=30
    -3, -9, -4, 1, 1, -1, -4, 7, 0,
    -- filter=205 channel=31
    12, 9, -12, 18, 3, -1, 5, -9, 5,
    -- filter=205 channel=32
    -2, 3, -1, 10, 0, -10, 4, -9, -11,
    -- filter=205 channel=33
    -9, 2, -3, 5, 9, -1, 1, 4, 0,
    -- filter=205 channel=34
    -6, -16, -14, -9, -7, -8, -12, -3, -8,
    -- filter=205 channel=35
    4, 1, 2, -6, 7, -7, -3, 2, -6,
    -- filter=205 channel=36
    9, 3, -8, 2, -1, 0, -8, -7, 2,
    -- filter=205 channel=37
    -22, -14, -11, -4, -3, 4, -3, 2, 2,
    -- filter=205 channel=38
    -2, 10, 5, 7, 1, -2, -1, 3, -6,
    -- filter=205 channel=39
    0, 10, 0, -2, 2, -3, -2, -2, 5,
    -- filter=205 channel=40
    0, -2, 0, -2, 1, -5, -7, -7, 1,
    -- filter=205 channel=41
    -2, -2, 10, -15, 0, -17, -8, -8, -19,
    -- filter=205 channel=42
    2, -7, -1, -5, 5, 10, 3, 2, -1,
    -- filter=205 channel=43
    -5, -1, -3, -1, 2, -3, 1, 2, -5,
    -- filter=205 channel=44
    -9, -3, -6, -1, 0, 6, 5, -1, 8,
    -- filter=205 channel=45
    1, -1, 6, -4, 1, 8, 0, 0, 0,
    -- filter=205 channel=46
    -5, 4, 6, -2, -4, -6, 4, 0, -7,
    -- filter=205 channel=47
    -4, 0, -5, -5, 12, 3, 1, 4, 7,
    -- filter=205 channel=48
    2, -2, -13, 3, 6, -3, -4, 3, 5,
    -- filter=205 channel=49
    4, 8, 5, -5, -10, -7, 3, -1, -1,
    -- filter=205 channel=50
    11, -2, -7, 14, -2, -8, 4, 0, 0,
    -- filter=205 channel=51
    3, 7, 6, -2, 5, 0, -5, -6, -5,
    -- filter=205 channel=52
    -2, -5, -2, -4, -3, -8, -8, 0, 1,
    -- filter=205 channel=53
    1, 0, -5, 6, 2, -1, 1, -9, 5,
    -- filter=205 channel=54
    6, -3, 0, -5, 5, -4, -2, 6, -2,
    -- filter=205 channel=55
    11, 16, 4, 9, -8, -20, 6, -14, -6,
    -- filter=205 channel=56
    -1, -5, -2, 1, -3, 0, 3, -5, -7,
    -- filter=205 channel=57
    -6, 0, -1, -5, 3, -5, -7, 1, -3,
    -- filter=205 channel=58
    -12, -8, 1, -3, 8, 1, -2, 4, 6,
    -- filter=205 channel=59
    -6, 10, 1, 15, 4, -3, -3, -2, -14,
    -- filter=205 channel=60
    -7, -3, -3, 1, 6, 0, 3, 4, 0,
    -- filter=205 channel=61
    6, 7, -3, -5, -3, 5, 4, -3, 2,
    -- filter=205 channel=62
    -5, 0, -3, 3, -1, 0, -6, -5, 4,
    -- filter=205 channel=63
    0, -3, 5, 2, -2, 4, -2, 10, 0,
    -- filter=205 channel=64
    9, -2, -1, 3, 3, 0, -3, -7, -2,
    -- filter=205 channel=65
    -5, 0, 1, 2, 0, 7, 4, -7, 1,
    -- filter=205 channel=66
    -5, 1, -8, -10, -3, -13, -1, -2, -5,
    -- filter=205 channel=67
    0, 4, 2, 3, -4, -3, -4, 6, 0,
    -- filter=205 channel=68
    2, 3, -3, -4, -8, 0, -1, 4, -2,
    -- filter=205 channel=69
    -2, 0, -6, 2, 4, -6, 0, -5, 0,
    -- filter=205 channel=70
    -1, 5, -14, 6, -4, -1, -3, -5, -10,
    -- filter=205 channel=71
    6, 4, -6, 5, 4, -5, 3, 0, -4,
    -- filter=205 channel=72
    3, 14, -2, 19, 12, -5, -4, -8, -6,
    -- filter=205 channel=73
    10, 0, -7, 11, -6, -5, -5, -8, -10,
    -- filter=205 channel=74
    2, 1, -4, -2, -10, -11, 1, -12, -4,
    -- filter=205 channel=75
    -13, -9, 8, -14, 3, 16, 9, 18, 6,
    -- filter=205 channel=76
    6, 3, 6, 5, -7, -9, 0, -2, -4,
    -- filter=205 channel=77
    -5, -4, 4, -1, -4, 0, -3, 0, -1,
    -- filter=205 channel=78
    -3, -1, 3, 0, 0, 0, 5, 0, 7,
    -- filter=205 channel=79
    2, 11, -3, 10, 1, -17, 1, 0, -6,
    -- filter=205 channel=80
    7, 11, 1, 22, 8, -10, 9, 3, -8,
    -- filter=205 channel=81
    7, 3, -1, -1, 0, -3, 0, 1, -5,
    -- filter=205 channel=82
    6, 0, -5, 1, -4, -3, -2, 1, 0,
    -- filter=205 channel=83
    5, 0, 3, -4, 6, 1, -3, 0, 4,
    -- filter=205 channel=84
    5, -4, -2, 6, -9, 0, -2, -3, -4,
    -- filter=205 channel=85
    -3, 0, 0, -2, -4, 5, 5, 3, 0,
    -- filter=205 channel=86
    -11, -4, 0, -12, 2, -4, -7, -5, 7,
    -- filter=205 channel=87
    -1, 3, -1, -9, -2, 0, -7, -11, -10,
    -- filter=205 channel=88
    5, -1, 3, 1, -4, 0, -9, -3, 0,
    -- filter=205 channel=89
    5, 15, -1, 16, 11, -19, -2, -13, -16,
    -- filter=205 channel=90
    1, 2, -3, -4, -6, -1, -9, -4, -5,
    -- filter=205 channel=91
    11, 7, -9, 9, -10, -5, -8, 0, 2,
    -- filter=205 channel=92
    3, 0, 1, -10, -4, 0, -6, 1, -3,
    -- filter=205 channel=93
    -16, -8, -5, 2, -4, 9, 0, 7, 7,
    -- filter=205 channel=94
    2, -7, 7, -4, -1, -4, -4, 6, 2,
    -- filter=205 channel=95
    -1, 4, 7, 5, -6, 0, -1, 0, 3,
    -- filter=205 channel=96
    0, 3, 8, 0, 5, -6, 4, 2, -4,
    -- filter=205 channel=97
    -8, 7, 2, 0, 10, 7, 3, 7, -3,
    -- filter=205 channel=98
    5, 12, 0, 9, 5, -15, -1, 6, 0,
    -- filter=205 channel=99
    17, 13, -5, 11, 4, -14, -1, -17, 0,
    -- filter=205 channel=100
    3, -2, 3, 2, -5, -1, -1, -4, 4,
    -- filter=205 channel=101
    0, 5, 4, 1, -2, -2, 1, 0, -6,
    -- filter=205 channel=102
    -5, 0, 0, 3, 2, -6, 0, 0, -2,
    -- filter=205 channel=103
    -4, -1, -3, 0, 7, 9, 3, 6, 12,
    -- filter=205 channel=104
    6, 9, -5, 12, 3, 3, -6, 1, -1,
    -- filter=205 channel=105
    6, 0, 5, 6, -4, -1, 2, -6, 3,
    -- filter=205 channel=106
    -2, -4, 7, 1, -9, -5, 4, -5, -3,
    -- filter=205 channel=107
    2, 10, 5, 1, -12, 0, 2, -13, -5,
    -- filter=205 channel=108
    -7, -1, 5, 0, -2, 7, -7, 0, 6,
    -- filter=205 channel=109
    0, 3, -14, 5, -5, -14, -5, -12, -2,
    -- filter=205 channel=110
    7, -2, 1, 3, 0, 0, 1, 0, 0,
    -- filter=205 channel=111
    4, 5, -5, 0, -5, -6, -2, -3, -5,
    -- filter=205 channel=112
    4, -1, -10, 6, -5, 5, 7, 0, -2,
    -- filter=205 channel=113
    4, -1, -8, 9, 4, -1, 5, -1, -9,
    -- filter=205 channel=114
    -4, 3, -6, 1, -7, -3, -4, -8, 3,
    -- filter=205 channel=115
    -2, 1, 5, -7, -2, -1, -4, 1, 4,
    -- filter=205 channel=116
    14, 0, -2, 13, -1, -15, -5, -11, -9,
    -- filter=205 channel=117
    3, 6, 0, 4, -3, 0, 3, 0, -6,
    -- filter=205 channel=118
    2, 5, 6, 4, 7, 7, -1, -1, 3,
    -- filter=205 channel=119
    7, -11, -7, -9, -16, -8, -11, -8, -1,
    -- filter=205 channel=120
    26, 13, -2, 12, -20, -1, -6, -7, -9,
    -- filter=205 channel=121
    -1, -2, -1, -4, 2, -12, -5, -6, -4,
    -- filter=205 channel=122
    -13, -10, -8, 3, 14, 3, -2, 9, 5,
    -- filter=205 channel=123
    -6, -7, -12, -5, -6, -9, -1, -7, 3,
    -- filter=205 channel=124
    5, 0, 6, -4, -8, -4, 2, 4, -4,
    -- filter=205 channel=125
    16, 11, 0, 3, -1, -15, 2, -6, -6,
    -- filter=205 channel=126
    3, 10, 8, 13, 13, -9, 4, -5, -7,
    -- filter=205 channel=127
    -8, -2, -4, -5, 0, -4, -7, 2, 0,
    -- filter=206 channel=0
    -8, 23, 25, -7, 38, 46, -20, 17, 19,
    -- filter=206 channel=1
    -7, 14, 12, 0, 35, 26, -20, 3, 1,
    -- filter=206 channel=2
    1, -3, -4, 1, -9, 0, 5, -8, 3,
    -- filter=206 channel=3
    2, 1, 2, -8, 6, 2, -3, -2, -3,
    -- filter=206 channel=4
    -6, -1, 6, -7, -1, 0, -10, -4, -4,
    -- filter=206 channel=5
    -15, 5, 9, -1, 23, 16, -12, -2, -4,
    -- filter=206 channel=6
    -7, 0, 1, -6, 9, 15, -4, 6, -4,
    -- filter=206 channel=7
    1, 6, -6, 6, 4, 2, 4, -1, -1,
    -- filter=206 channel=8
    3, -4, -6, -2, -6, -4, -3, -9, 1,
    -- filter=206 channel=9
    7, 0, 5, 5, 1, 3, 2, -7, 0,
    -- filter=206 channel=10
    7, -6, -14, 9, -8, -13, 2, -15, -12,
    -- filter=206 channel=11
    1, -10, 4, -1, -1, 8, 6, -1, 1,
    -- filter=206 channel=12
    -7, -10, 6, -2, -4, 7, -6, -9, -4,
    -- filter=206 channel=13
    2, -6, -7, 3, -5, -7, -4, 0, 2,
    -- filter=206 channel=14
    -6, 1, 0, -4, 1, 0, 0, -4, 5,
    -- filter=206 channel=15
    -4, 3, 6, 1, 14, 14, 1, 7, 8,
    -- filter=206 channel=16
    0, 0, -6, 5, 0, -2, -4, -13, -6,
    -- filter=206 channel=17
    -4, 6, -6, 1, 6, -6, 6, -3, -2,
    -- filter=206 channel=18
    -14, 0, 3, 0, 21, 17, -12, 14, -2,
    -- filter=206 channel=19
    -5, 6, 4, 0, 0, 2, -5, 1, 1,
    -- filter=206 channel=20
    -7, -7, 5, -7, -7, 1, 4, 0, 4,
    -- filter=206 channel=21
    2, -6, 0, -4, -19, -17, -1, -4, -10,
    -- filter=206 channel=22
    -8, 10, 2, -1, 21, 8, -7, 10, -1,
    -- filter=206 channel=23
    0, -14, -7, 2, -6, 4, 10, -7, -4,
    -- filter=206 channel=24
    -3, -1, 4, -1, 2, -5, -3, -3, 1,
    -- filter=206 channel=25
    7, -1, 3, 8, -7, -1, 4, 0, 0,
    -- filter=206 channel=26
    -3, 0, -3, 1, 0, -1, -1, -9, 6,
    -- filter=206 channel=27
    4, 7, -7, 4, 6, 1, 4, 3, 11,
    -- filter=206 channel=28
    -4, -3, -5, -6, 5, -1, -4, 6, 1,
    -- filter=206 channel=29
    0, -12, -2, 4, -8, 7, 3, 5, -8,
    -- filter=206 channel=30
    2, 3, 10, 0, 1, 15, -3, 7, 14,
    -- filter=206 channel=31
    16, -16, -9, 8, -32, -12, 15, -17, 5,
    -- filter=206 channel=32
    1, -4, 2, -9, 15, 6, -3, -4, 4,
    -- filter=206 channel=33
    -4, 3, 6, 3, 13, 11, -6, 0, 4,
    -- filter=206 channel=34
    -12, -6, -7, 0, -15, 4, -6, -8, -2,
    -- filter=206 channel=35
    -1, -6, 5, -6, 0, -1, -2, 0, 0,
    -- filter=206 channel=36
    2, -15, -13, 3, -16, -7, 4, -6, -11,
    -- filter=206 channel=37
    -13, 18, 14, -3, 29, 30, -20, 3, 5,
    -- filter=206 channel=38
    3, -3, -1, 4, -9, 0, -2, 2, 5,
    -- filter=206 channel=39
    3, -3, 2, -5, 1, -6, 1, -3, 0,
    -- filter=206 channel=40
    6, 0, -4, 10, -2, 9, 2, 8, 1,
    -- filter=206 channel=41
    -10, -20, 1, -6, -14, 2, -14, -8, -4,
    -- filter=206 channel=42
    0, 3, 5, 2, 4, 2, -1, -2, 0,
    -- filter=206 channel=43
    -7, 4, 7, 0, 10, 7, -9, 0, -6,
    -- filter=206 channel=44
    0, 9, 10, 1, 2, 13, -4, 4, 5,
    -- filter=206 channel=45
    -3, 9, 5, 4, 5, 2, -1, 12, 8,
    -- filter=206 channel=46
    5, 3, 0, 2, 1, 2, 5, -2, -5,
    -- filter=206 channel=47
    0, -2, -4, -7, -4, 0, 3, -8, 3,
    -- filter=206 channel=48
    -1, 6, -6, -3, -3, -2, -6, 3, 5,
    -- filter=206 channel=49
    4, 7, 0, 6, 11, 5, 1, 2, -5,
    -- filter=206 channel=50
    11, 0, 0, -1, 5, 0, 5, 1, 6,
    -- filter=206 channel=51
    -6, 2, -2, 5, 1, -1, -5, 3, 0,
    -- filter=206 channel=52
    -7, -11, 2, -2, -3, -4, -4, -10, -3,
    -- filter=206 channel=53
    -4, 1, 0, 2, 1, 6, 5, -4, 3,
    -- filter=206 channel=54
    -4, -4, 7, 2, 1, -5, -4, 4, -1,
    -- filter=206 channel=55
    4, -7, -7, 1, -4, -12, 0, 4, -4,
    -- filter=206 channel=56
    -10, 2, -4, -6, -7, -6, 2, 3, 3,
    -- filter=206 channel=57
    -8, -5, -5, -8, -6, 2, -1, 3, -4,
    -- filter=206 channel=58
    -11, 8, 9, -5, 12, 19, -10, 0, 0,
    -- filter=206 channel=59
    2, -4, -9, 4, -3, -9, 5, 3, 5,
    -- filter=206 channel=60
    -2, -5, 1, 7, 6, -6, 3, 3, -1,
    -- filter=206 channel=61
    2, -10, -2, 6, -10, -4, 0, 0, -10,
    -- filter=206 channel=62
    0, -5, 2, -1, 3, -2, -4, -5, -7,
    -- filter=206 channel=63
    -4, 1, 7, -6, 0, 11, 2, -2, 2,
    -- filter=206 channel=64
    3, 1, -2, 5, -12, -3, 8, 4, -1,
    -- filter=206 channel=65
    7, 2, -3, 4, -2, 6, -3, 4, -3,
    -- filter=206 channel=66
    -6, -16, -5, -5, -14, -1, -2, -11, 0,
    -- filter=206 channel=67
    -1, 8, 0, -7, 6, 3, -5, -6, 1,
    -- filter=206 channel=68
    6, -8, -6, 6, 1, 3, 4, -5, -7,
    -- filter=206 channel=69
    -2, -7, 7, -5, 0, 0, -2, -3, -3,
    -- filter=206 channel=70
    1, 4, 11, 0, 14, 7, -4, 2, 1,
    -- filter=206 channel=71
    5, -9, -9, 1, -5, -9, 5, 3, 1,
    -- filter=206 channel=72
    14, -11, -8, 14, -18, -17, 3, -6, 3,
    -- filter=206 channel=73
    2, 1, -4, 4, -1, -3, -1, 0, 0,
    -- filter=206 channel=74
    -3, -16, 1, -4, -2, 0, 0, -6, -3,
    -- filter=206 channel=75
    -10, 12, 6, -1, 25, 26, -18, 0, 5,
    -- filter=206 channel=76
    -4, 0, -2, 0, 2, -10, 8, 8, -10,
    -- filter=206 channel=77
    -3, 2, -4, -3, -7, 2, 0, 6, -4,
    -- filter=206 channel=78
    -7, 0, 2, -9, -6, -2, 0, -2, -3,
    -- filter=206 channel=79
    -3, 6, 1, 6, 24, 24, -7, 9, 7,
    -- filter=206 channel=80
    0, -17, -7, -1, -17, -19, 5, -11, 0,
    -- filter=206 channel=81
    -4, -3, 0, 2, -3, -2, 5, -1, 0,
    -- filter=206 channel=82
    -1, -1, 1, 0, -2, 3, 1, -3, 1,
    -- filter=206 channel=83
    4, -3, -6, 9, -4, -5, 0, 0, -1,
    -- filter=206 channel=84
    1, -4, 3, -7, 7, 12, -4, -7, 9,
    -- filter=206 channel=85
    -1, 2, -1, 5, 5, 6, -6, -5, 1,
    -- filter=206 channel=86
    -3, -5, 4, 2, -5, 1, -4, -13, -2,
    -- filter=206 channel=87
    -1, -11, 3, -6, -4, 7, -6, -2, 1,
    -- filter=206 channel=88
    2, -13, 2, 1, -8, -18, 4, -10, -8,
    -- filter=206 channel=89
    7, -5, -13, 5, -6, -8, 0, -7, -7,
    -- filter=206 channel=90
    -1, -15, -5, 6, -16, -9, 6, 0, -7,
    -- filter=206 channel=91
    0, 1, 5, 5, 10, 3, 5, 0, 4,
    -- filter=206 channel=92
    -1, -4, -2, -4, -5, 0, -2, 0, -3,
    -- filter=206 channel=93
    1, 0, 12, -4, 9, 7, -15, -3, 1,
    -- filter=206 channel=94
    -3, 5, 6, 7, 4, 6, -3, -2, -7,
    -- filter=206 channel=95
    -4, 2, -7, 4, 0, 3, -2, -8, 1,
    -- filter=206 channel=96
    2, 9, -2, 5, 0, 0, 0, -1, 1,
    -- filter=206 channel=97
    1, -5, -3, 2, 0, 8, 0, 2, -5,
    -- filter=206 channel=98
    2, -12, -9, 2, -12, 1, 0, -7, -12,
    -- filter=206 channel=99
    4, -31, -2, 6, -33, -17, 15, -23, -4,
    -- filter=206 channel=100
    0, 3, -4, -3, -4, -6, 3, 5, -11,
    -- filter=206 channel=101
    8, -11, 2, -5, 3, -11, -3, -6, -3,
    -- filter=206 channel=102
    7, 3, -2, 1, 1, 3, -4, 0, -1,
    -- filter=206 channel=103
    1, 2, -6, -4, 2, 6, -9, -5, 0,
    -- filter=206 channel=104
    8, -12, -11, 0, -22, -25, 4, -8, -3,
    -- filter=206 channel=105
    -1, -2, 4, 3, 3, 2, 7, -2, 3,
    -- filter=206 channel=106
    4, -7, 0, 2, -1, 4, 6, 1, 2,
    -- filter=206 channel=107
    -3, 9, 13, 4, 20, 22, -1, 1, 12,
    -- filter=206 channel=108
    -11, -4, 6, -9, 10, 1, -2, 7, 0,
    -- filter=206 channel=109
    -1, 0, -14, 2, 8, 0, -2, -2, -8,
    -- filter=206 channel=110
    6, -16, -8, -1, -18, -7, 5, -3, -3,
    -- filter=206 channel=111
    0, 1, -5, -3, 3, 4, 2, 2, -8,
    -- filter=206 channel=112
    7, 7, -1, 0, 11, -1, 0, 0, 2,
    -- filter=206 channel=113
    8, 0, -10, -1, -9, -6, 2, 1, -2,
    -- filter=206 channel=114
    -11, 21, 19, -15, 44, 46, -24, 11, 18,
    -- filter=206 channel=115
    2, -6, -2, 6, -3, -6, 4, -1, -7,
    -- filter=206 channel=116
    3, -4, -4, 4, -14, -9, 2, -2, -5,
    -- filter=206 channel=117
    0, -2, -8, -1, -1, -2, 7, 0, -7,
    -- filter=206 channel=118
    -4, 4, 3, -1, 2, 0, -1, -2, -7,
    -- filter=206 channel=119
    -7, -4, -7, -1, -4, 5, -5, -11, -4,
    -- filter=206 channel=120
    -5, -12, 0, 0, -3, 11, 5, -3, 1,
    -- filter=206 channel=121
    -8, -2, -10, 1, -4, -9, -2, -6, -10,
    -- filter=206 channel=122
    2, -5, -5, 4, -17, -21, 9, -16, -4,
    -- filter=206 channel=123
    -9, -9, -1, 4, -9, -6, 1, 2, -4,
    -- filter=206 channel=124
    -4, -3, 0, 5, 4, 2, 4, -5, -2,
    -- filter=206 channel=125
    4, -21, -14, 8, -24, -17, 8, -14, 2,
    -- filter=206 channel=126
    -2, -1, 5, -9, 3, 10, -7, 0, 2,
    -- filter=206 channel=127
    -1, 0, -6, 3, 3, -8, -2, 0, -6,
    -- filter=207 channel=0
    -3, 2, -5, -7, 7, -4, 4, 4, -3,
    -- filter=207 channel=1
    1, 0, 7, -1, 2, 5, -2, 0, 7,
    -- filter=207 channel=2
    -1, -7, 0, -5, 0, -6, -7, 7, 7,
    -- filter=207 channel=3
    -5, 0, -7, -5, -7, 0, 0, 6, 2,
    -- filter=207 channel=4
    6, 0, -7, 1, -4, -3, 7, -2, 0,
    -- filter=207 channel=5
    6, 4, -1, 0, -5, -2, 5, 7, 5,
    -- filter=207 channel=6
    -2, 4, 4, -4, -3, -4, -2, 3, -6,
    -- filter=207 channel=7
    0, -4, 1, 1, 6, -4, 1, -7, 2,
    -- filter=207 channel=8
    -4, -1, 5, 3, -4, -6, -1, -2, -4,
    -- filter=207 channel=9
    -4, -5, -6, 4, 5, -1, 1, 7, 5,
    -- filter=207 channel=10
    -1, -5, 5, 4, -3, -6, -2, 6, 5,
    -- filter=207 channel=11
    -3, -2, -2, 1, 2, -6, -5, 3, -5,
    -- filter=207 channel=12
    3, -6, 6, -3, -2, -5, 5, 5, 0,
    -- filter=207 channel=13
    -1, 0, -7, 2, 1, -4, 3, 4, -4,
    -- filter=207 channel=14
    4, 5, 2, 0, 6, 0, -1, 6, 7,
    -- filter=207 channel=15
    -4, -6, 1, 6, 0, 5, -5, -4, -7,
    -- filter=207 channel=16
    -2, 5, 6, -1, -5, -3, 1, -4, 2,
    -- filter=207 channel=17
    -5, 5, 5, -2, 1, 6, -6, -5, 6,
    -- filter=207 channel=18
    0, 5, 0, -3, -1, -4, 0, -3, -1,
    -- filter=207 channel=19
    6, 1, -7, 2, 2, 2, -3, -6, -6,
    -- filter=207 channel=20
    -5, 1, 0, 2, 2, -5, -7, -4, -3,
    -- filter=207 channel=21
    -1, 6, -5, 3, 1, 5, -2, -1, 3,
    -- filter=207 channel=22
    -4, 7, 4, -6, 4, -5, 7, -5, 4,
    -- filter=207 channel=23
    -2, -7, -3, -3, -7, 2, -2, -7, -6,
    -- filter=207 channel=24
    7, -7, 6, 0, 0, 3, 4, -2, 6,
    -- filter=207 channel=25
    -1, 4, 0, 4, 5, 2, -5, 0, 2,
    -- filter=207 channel=26
    2, 3, 2, -1, -5, -3, -5, -5, -1,
    -- filter=207 channel=27
    -1, 2, -6, -1, 0, 6, -3, -5, 0,
    -- filter=207 channel=28
    1, -4, 5, 6, -5, 7, -4, 1, -2,
    -- filter=207 channel=29
    0, 0, 5, -4, 4, 1, 6, 1, -1,
    -- filter=207 channel=30
    0, 5, -4, 3, 2, -1, 3, 1, -4,
    -- filter=207 channel=31
    0, 0, -5, -1, -6, -7, 0, 3, -2,
    -- filter=207 channel=32
    4, 1, 5, -7, -2, 4, -2, 4, 0,
    -- filter=207 channel=33
    5, -2, -2, 7, 6, -5, 3, -7, 1,
    -- filter=207 channel=34
    0, 0, 5, 3, -5, 2, -7, 2, -3,
    -- filter=207 channel=35
    0, -3, -4, -3, -2, -5, -3, -5, 0,
    -- filter=207 channel=36
    -6, -4, 2, -3, -7, 0, -7, 0, 6,
    -- filter=207 channel=37
    -4, 2, -6, -1, 6, -3, -2, 0, -5,
    -- filter=207 channel=38
    -7, 7, -5, -1, 2, 1, -3, -6, -6,
    -- filter=207 channel=39
    -4, 5, -3, -2, -1, 1, 2, -6, 1,
    -- filter=207 channel=40
    -6, -7, 5, 0, 1, 5, -1, -7, -4,
    -- filter=207 channel=41
    0, -5, -4, 5, 4, 0, -3, -4, -6,
    -- filter=207 channel=42
    0, -3, 7, -7, -6, 1, -5, 4, -2,
    -- filter=207 channel=43
    4, 0, -3, 0, -1, 3, 1, 1, -2,
    -- filter=207 channel=44
    -7, 1, -6, -5, -1, 2, 0, 0, -6,
    -- filter=207 channel=45
    -3, 6, -2, -1, -3, 3, 5, 0, 7,
    -- filter=207 channel=46
    4, -1, 0, 1, 0, 1, -4, -3, -2,
    -- filter=207 channel=47
    -5, -3, 5, -1, 3, -3, 6, 0, -3,
    -- filter=207 channel=48
    -1, -2, 7, 2, -3, -2, 4, 4, 0,
    -- filter=207 channel=49
    4, 4, 4, -1, 4, 0, -3, 0, -2,
    -- filter=207 channel=50
    -2, -3, 2, 5, 2, 2, -1, 0, 7,
    -- filter=207 channel=51
    0, 1, 3, -5, -4, 1, 2, -1, -3,
    -- filter=207 channel=52
    -6, 5, -6, -5, 1, 0, 0, -6, 4,
    -- filter=207 channel=53
    -5, -6, 1, 6, 5, 0, -1, -6, 5,
    -- filter=207 channel=54
    -4, 6, -3, 6, -7, 7, 2, 0, -1,
    -- filter=207 channel=55
    2, -2, -1, 4, -3, 6, 1, 5, -4,
    -- filter=207 channel=56
    3, 6, -2, -2, -2, -6, -6, 6, 5,
    -- filter=207 channel=57
    5, -5, 4, 0, 7, -1, 6, -1, -2,
    -- filter=207 channel=58
    7, 6, -1, -1, 7, 2, -4, 3, -2,
    -- filter=207 channel=59
    3, 1, 2, 1, 4, -2, 6, -7, 4,
    -- filter=207 channel=60
    -2, 2, -2, 6, -5, 5, 4, 5, 4,
    -- filter=207 channel=61
    -1, -3, -2, 3, 0, 2, 7, 6, -4,
    -- filter=207 channel=62
    -1, -5, 2, 2, -6, 1, -2, -4, -5,
    -- filter=207 channel=63
    -6, 0, -7, -2, -4, 1, -6, 4, 4,
    -- filter=207 channel=64
    3, 4, 0, -3, 6, -6, 0, 3, 6,
    -- filter=207 channel=65
    -2, 6, -1, -2, 2, -3, 1, -5, 5,
    -- filter=207 channel=66
    2, 0, 3, 5, 2, 1, 6, -3, -4,
    -- filter=207 channel=67
    3, 0, 0, 2, 3, 6, 1, -5, -6,
    -- filter=207 channel=68
    6, -6, 6, 2, -1, -5, -4, 5, 5,
    -- filter=207 channel=69
    4, 5, -6, -6, -7, 0, 3, 1, 2,
    -- filter=207 channel=70
    0, 2, -7, -7, -4, -6, 0, 0, -3,
    -- filter=207 channel=71
    -5, -6, -6, -5, -6, -4, -6, -2, -6,
    -- filter=207 channel=72
    2, -1, -6, 1, -5, -7, -2, 2, 3,
    -- filter=207 channel=73
    1, -6, -1, 3, -7, -6, -3, -1, -4,
    -- filter=207 channel=74
    4, -5, -6, -7, 0, 4, -3, -4, 3,
    -- filter=207 channel=75
    4, 0, 0, -2, 0, 0, 3, 2, 2,
    -- filter=207 channel=76
    4, 0, 4, 0, 0, -2, -1, 4, 0,
    -- filter=207 channel=77
    4, -1, 0, 0, -7, -3, -1, -2, -4,
    -- filter=207 channel=78
    -7, -4, -3, 5, -1, -1, 5, 5, -4,
    -- filter=207 channel=79
    4, -1, 3, -2, -7, -6, -4, -6, 2,
    -- filter=207 channel=80
    -3, 0, 0, 3, -2, -4, 5, -2, -6,
    -- filter=207 channel=81
    7, 4, -2, 2, 4, 0, -4, -5, -3,
    -- filter=207 channel=82
    -4, 4, -4, 0, 0, 4, -6, 0, -3,
    -- filter=207 channel=83
    -7, 2, 2, 1, 1, -2, 1, -1, 4,
    -- filter=207 channel=84
    4, -1, 5, 1, 5, 3, 0, -4, 6,
    -- filter=207 channel=85
    7, -4, 2, 2, 0, -4, 7, 6, -5,
    -- filter=207 channel=86
    0, -3, -5, 0, 1, 4, 4, 7, 6,
    -- filter=207 channel=87
    -5, 7, -4, -6, 0, 4, 1, 0, 6,
    -- filter=207 channel=88
    3, 2, 4, -3, 0, 3, 6, -4, -3,
    -- filter=207 channel=89
    5, -5, 4, -4, 2, 2, 4, -7, -1,
    -- filter=207 channel=90
    -7, 3, -1, -6, -7, 6, 0, -3, 4,
    -- filter=207 channel=91
    4, -5, 0, -2, -4, -6, 5, -3, 2,
    -- filter=207 channel=92
    3, 0, 5, 0, 6, 0, 0, -3, 7,
    -- filter=207 channel=93
    -4, -5, 1, -7, 4, -3, 4, -6, 0,
    -- filter=207 channel=94
    -6, -4, 0, -6, -2, -4, 5, -3, -2,
    -- filter=207 channel=95
    -5, -7, -6, -2, -3, -7, 6, -2, 2,
    -- filter=207 channel=96
    5, 5, 2, -7, -6, 0, -7, 7, -2,
    -- filter=207 channel=97
    -1, 7, -4, 1, -4, 0, 0, 5, -5,
    -- filter=207 channel=98
    3, 0, -5, -4, -3, 4, -1, -7, 7,
    -- filter=207 channel=99
    6, -7, 3, 0, 4, 4, 3, -7, -5,
    -- filter=207 channel=100
    6, -5, 4, 0, -1, 2, 1, 7, -3,
    -- filter=207 channel=101
    -4, -3, -7, 7, 0, 2, 3, -1, -4,
    -- filter=207 channel=102
    -5, 5, -3, -6, 3, 7, 0, -3, 2,
    -- filter=207 channel=103
    -5, -4, -2, -3, -5, 7, -3, -7, -1,
    -- filter=207 channel=104
    0, -3, 3, -3, 6, -4, 0, 5, 3,
    -- filter=207 channel=105
    1, 6, 0, 6, 5, -3, 1, -2, -5,
    -- filter=207 channel=106
    4, 1, 3, 3, 4, 6, -1, -1, 3,
    -- filter=207 channel=107
    1, -5, -4, -7, -6, 0, -3, 6, 0,
    -- filter=207 channel=108
    -1, 5, -7, -6, -7, 1, -4, -1, 1,
    -- filter=207 channel=109
    -2, -2, -1, -2, -2, -6, -2, 4, 5,
    -- filter=207 channel=110
    2, 2, -3, -3, -2, 5, -6, -2, -2,
    -- filter=207 channel=111
    3, -1, 5, -1, 2, -6, -4, -5, 5,
    -- filter=207 channel=112
    -2, 3, 1, 5, 6, 3, 5, -5, -1,
    -- filter=207 channel=113
    0, 0, 2, -1, 0, -6, -7, -2, -6,
    -- filter=207 channel=114
    6, 4, -5, -6, -5, -3, 4, -6, -4,
    -- filter=207 channel=115
    -5, -3, 6, -1, -4, -1, 6, 3, -1,
    -- filter=207 channel=116
    7, -4, 5, 3, -2, 4, -1, -2, -1,
    -- filter=207 channel=117
    0, -1, 5, -2, 6, 0, -5, -4, -1,
    -- filter=207 channel=118
    -1, -1, 0, 0, -7, -5, -6, 6, 0,
    -- filter=207 channel=119
    4, 0, 5, 4, -6, -6, 0, 1, 6,
    -- filter=207 channel=120
    1, 2, 0, 6, 4, -4, 3, -4, 7,
    -- filter=207 channel=121
    5, 1, 0, -3, 2, 3, 5, 4, -3,
    -- filter=207 channel=122
    -3, 5, 5, -3, 1, 0, -7, 4, -5,
    -- filter=207 channel=123
    4, -7, 0, 0, 6, -6, 3, 0, -2,
    -- filter=207 channel=124
    4, 0, -1, -1, -2, 7, -5, -6, 0,
    -- filter=207 channel=125
    -5, -3, -5, 0, 2, -4, 1, 5, -1,
    -- filter=207 channel=126
    0, 7, 6, 0, 0, -7, 7, -5, 5,
    -- filter=207 channel=127
    0, 5, -6, 2, 3, 7, 1, 0, -6,
    -- filter=208 channel=0
    -1, 2, -7, -1, -7, -11, 0, -4, -7,
    -- filter=208 channel=1
    -1, -2, -5, 7, -7, -9, 1, -8, 4,
    -- filter=208 channel=2
    2, -7, -8, 3, 1, 3, -1, -1, 3,
    -- filter=208 channel=3
    -7, 8, -1, 4, 3, -6, 2, -3, -5,
    -- filter=208 channel=4
    4, -11, -6, -3, -7, -8, 5, 6, 7,
    -- filter=208 channel=5
    -5, -3, 3, 2, -6, 1, -5, -6, -4,
    -- filter=208 channel=6
    1, 5, 2, 7, 0, 0, 0, 3, 7,
    -- filter=208 channel=7
    4, -3, -6, 1, -5, 5, 0, 7, 5,
    -- filter=208 channel=8
    1, 0, 0, 3, 2, 5, 5, 6, -6,
    -- filter=208 channel=9
    -6, 0, 4, -4, 3, 0, -2, 3, 1,
    -- filter=208 channel=10
    4, 3, 0, 8, -4, -2, 8, -9, 1,
    -- filter=208 channel=11
    0, 5, 0, -3, 0, 0, 0, 9, 9,
    -- filter=208 channel=12
    10, -9, 2, -2, 1, 2, 1, 0, -7,
    -- filter=208 channel=13
    10, -8, -8, 2, -2, -8, 1, -1, -5,
    -- filter=208 channel=14
    4, 3, -1, 0, -5, 7, 0, -5, 1,
    -- filter=208 channel=15
    -5, 0, 4, 3, -4, -7, 0, -1, -3,
    -- filter=208 channel=16
    -2, -4, -2, 4, 3, 1, 4, -8, 7,
    -- filter=208 channel=17
    1, 0, 4, 1, 2, -3, -4, -5, -2,
    -- filter=208 channel=18
    -1, -3, -7, -2, -5, -3, 8, -6, -6,
    -- filter=208 channel=19
    7, 5, 5, -6, 6, 5, 5, 4, 5,
    -- filter=208 channel=20
    5, 6, 10, -5, 5, 5, 6, 4, 4,
    -- filter=208 channel=21
    11, -7, -2, 7, 4, 7, 3, -9, 10,
    -- filter=208 channel=22
    1, 0, 5, -5, -6, 0, -1, -5, 1,
    -- filter=208 channel=23
    2, -8, 1, -4, -9, -3, -3, -7, -6,
    -- filter=208 channel=24
    -5, -3, -3, 7, -7, 0, 6, 5, 0,
    -- filter=208 channel=25
    -2, -13, -10, 8, -11, -6, 5, -6, -6,
    -- filter=208 channel=26
    -4, -2, -2, 2, -1, 0, -1, -3, 1,
    -- filter=208 channel=27
    -3, -2, -6, -4, -17, -14, 4, -15, -7,
    -- filter=208 channel=28
    4, 7, -2, 2, 5, -1, 2, 0, 4,
    -- filter=208 channel=29
    -2, 1, 10, -1, 10, 3, 3, 2, 7,
    -- filter=208 channel=30
    -7, 0, -2, 0, -6, -6, 0, 2, 0,
    -- filter=208 channel=31
    8, -9, 6, 0, -3, -4, 6, 1, -5,
    -- filter=208 channel=32
    -3, -8, 2, 3, -8, -1, 6, -7, -3,
    -- filter=208 channel=33
    -3, -8, 5, 0, -14, -3, -4, -11, 0,
    -- filter=208 channel=34
    -6, 5, -2, 4, -7, -8, 8, -9, 0,
    -- filter=208 channel=35
    1, 7, 1, 0, -4, 1, -1, 6, 5,
    -- filter=208 channel=36
    0, -1, 3, 2, -3, 10, 0, 0, 7,
    -- filter=208 channel=37
    0, -3, 0, 6, -9, 0, 7, 2, -1,
    -- filter=208 channel=38
    5, 2, -1, -2, -4, -4, -1, -2, 0,
    -- filter=208 channel=39
    6, 0, 6, -2, 4, 7, -4, 6, 3,
    -- filter=208 channel=40
    0, 7, 4, 7, 6, -1, 0, 6, 4,
    -- filter=208 channel=41
    12, 3, -3, 15, 9, -10, 17, 6, -8,
    -- filter=208 channel=42
    5, 2, -2, 2, -4, -5, -1, 4, 4,
    -- filter=208 channel=43
    -7, 2, -2, 3, 2, 0, 3, -4, 5,
    -- filter=208 channel=44
    0, 0, 0, 4, -10, 0, -2, 3, -2,
    -- filter=208 channel=45
    5, 7, 6, -4, 7, 3, 7, -2, 11,
    -- filter=208 channel=46
    5, 5, -2, -3, 7, 0, 2, 4, 4,
    -- filter=208 channel=47
    8, 0, -2, 1, -11, 3, 4, -2, 0,
    -- filter=208 channel=48
    0, 1, -8, -3, -1, 2, -3, 0, -3,
    -- filter=208 channel=49
    2, -7, -1, -6, -4, 0, -1, 2, -4,
    -- filter=208 channel=50
    -5, -4, -6, -5, 0, -3, -6, 0, -7,
    -- filter=208 channel=51
    -1, 7, 7, 2, 0, 4, 4, 7, 2,
    -- filter=208 channel=52
    -3, 1, -7, 0, 1, -6, 3, -8, -7,
    -- filter=208 channel=53
    -5, -2, 5, -1, 1, -2, -3, -2, -4,
    -- filter=208 channel=54
    -6, -3, 3, -5, 1, -1, -2, -2, -1,
    -- filter=208 channel=55
    -2, -5, 0, -6, -4, -7, -1, -1, -7,
    -- filter=208 channel=56
    4, 0, -1, 4, -6, 0, -3, 0, -8,
    -- filter=208 channel=57
    2, -8, 3, 4, -6, -3, 7, -4, -1,
    -- filter=208 channel=58
    -4, -7, -1, 6, 3, 0, -2, -5, 6,
    -- filter=208 channel=59
    -3, 1, -5, 7, -9, -4, -2, -1, -10,
    -- filter=208 channel=60
    2, 5, -6, 7, -1, 1, 2, -1, -6,
    -- filter=208 channel=61
    0, 2, 2, 8, -7, 0, 1, 6, -4,
    -- filter=208 channel=62
    2, -2, -1, -5, 0, 5, 3, -5, 3,
    -- filter=208 channel=63
    7, 0, -2, 4, -4, 9, 5, -4, 8,
    -- filter=208 channel=64
    8, 0, -1, 7, 0, 7, 2, -5, -4,
    -- filter=208 channel=65
    -2, -6, 7, 6, 5, 3, 3, 4, -5,
    -- filter=208 channel=66
    0, -8, 0, 7, -3, 0, -2, -8, -1,
    -- filter=208 channel=67
    6, 3, 2, 4, 3, 6, 2, 4, -5,
    -- filter=208 channel=68
    6, 1, 7, -2, 1, 4, -5, 8, -2,
    -- filter=208 channel=69
    7, -5, -3, 6, 5, 4, 3, 1, 2,
    -- filter=208 channel=70
    -4, -1, -3, -9, -10, -8, -5, -14, -12,
    -- filter=208 channel=71
    6, 0, 6, -3, -2, 3, 0, -7, 3,
    -- filter=208 channel=72
    5, 2, 2, -2, -5, -5, 0, -10, 4,
    -- filter=208 channel=73
    5, -8, 2, 2, -10, -10, 1, -3, 0,
    -- filter=208 channel=74
    -5, -2, 0, 0, -9, -3, -2, 0, -4,
    -- filter=208 channel=75
    6, 5, 6, 1, -12, -9, 0, 1, 0,
    -- filter=208 channel=76
    9, 6, 12, 0, 0, -3, 9, 11, -2,
    -- filter=208 channel=77
    8, -1, -7, -3, -3, -4, -2, 6, 0,
    -- filter=208 channel=78
    -5, -1, 5, -1, -5, 5, -1, 1, -2,
    -- filter=208 channel=79
    2, -4, -12, 0, -3, -14, 8, 2, -3,
    -- filter=208 channel=80
    0, 0, -8, -1, -15, -3, 10, -14, -2,
    -- filter=208 channel=81
    -2, 0, 1, 6, 7, 3, 4, 6, 6,
    -- filter=208 channel=82
    -1, 3, -2, 4, -1, 1, 4, -1, 4,
    -- filter=208 channel=83
    -5, 4, -4, -5, 1, -6, 5, -6, 8,
    -- filter=208 channel=84
    -2, -2, -5, -4, -3, -1, 2, 3, -1,
    -- filter=208 channel=85
    3, 5, 5, 0, 3, 2, -3, -3, 5,
    -- filter=208 channel=86
    3, -8, 5, 0, -8, 1, 3, 1, -2,
    -- filter=208 channel=87
    -6, 0, -2, 7, 1, -5, -6, 2, 3,
    -- filter=208 channel=88
    -2, 6, 7, 6, 3, 8, 0, 7, 10,
    -- filter=208 channel=89
    0, 2, 3, 2, -3, -1, 1, -9, -3,
    -- filter=208 channel=90
    -2, -1, 6, -4, 2, 10, 6, 1, 5,
    -- filter=208 channel=91
    2, -4, -3, 1, -11, 0, -2, -9, 4,
    -- filter=208 channel=92
    5, 1, -4, -4, -3, -3, 3, -3, -1,
    -- filter=208 channel=93
    1, -5, 1, 0, -1, 3, 8, 1, 4,
    -- filter=208 channel=94
    1, 0, 6, 7, -2, 5, 7, 5, -4,
    -- filter=208 channel=95
    5, 0, 2, 7, 5, 2, 1, 0, 2,
    -- filter=208 channel=96
    5, -5, 4, 7, -6, -4, 2, 3, 0,
    -- filter=208 channel=97
    -1, -3, 0, -5, -2, -1, -7, -7, 0,
    -- filter=208 channel=98
    9, -1, -6, -3, -12, -7, 7, 0, -1,
    -- filter=208 channel=99
    8, -8, -2, -6, -4, 0, 3, -5, 3,
    -- filter=208 channel=100
    0, 3, 2, 0, 2, -6, -6, 2, -5,
    -- filter=208 channel=101
    -6, 2, 3, 0, -7, 2, 0, 4, -3,
    -- filter=208 channel=102
    7, 0, 6, 0, 3, -6, 1, -6, 5,
    -- filter=208 channel=103
    -3, 2, 4, 2, -6, 6, 7, -2, 0,
    -- filter=208 channel=104
    4, -6, 6, 8, -4, -6, -1, 0, -1,
    -- filter=208 channel=105
    5, 9, 0, 1, 4, 7, 5, 12, 5,
    -- filter=208 channel=106
    6, 11, 2, 3, 5, -5, 8, 3, -5,
    -- filter=208 channel=107
    6, 5, -3, -8, 7, 3, -3, 3, 0,
    -- filter=208 channel=108
    0, 7, -7, 5, 1, -2, 0, 5, 0,
    -- filter=208 channel=109
    1, -12, -10, 2, -11, -4, -2, -2, -5,
    -- filter=208 channel=110
    4, 4, 1, -5, 2, -5, 4, -4, 4,
    -- filter=208 channel=111
    8, 5, 7, 9, -1, 0, 7, 3, -2,
    -- filter=208 channel=112
    -3, -3, 6, 4, 3, 1, 3, -3, -7,
    -- filter=208 channel=113
    6, -5, 1, 6, -12, -2, 0, -4, -11,
    -- filter=208 channel=114
    5, -5, -11, 4, -6, -13, 7, -5, -5,
    -- filter=208 channel=115
    0, 1, -2, 2, -6, -6, -1, 4, 3,
    -- filter=208 channel=116
    1, -13, 0, 5, 0, -8, -3, -6, 2,
    -- filter=208 channel=117
    0, 0, -3, 3, 3, 2, -1, -7, 2,
    -- filter=208 channel=118
    0, -3, 5, -6, -3, -1, -6, 0, -6,
    -- filter=208 channel=119
    5, -3, -9, -4, -6, 0, -2, -6, 0,
    -- filter=208 channel=120
    -6, -7, -7, -2, -9, -6, 0, -9, 6,
    -- filter=208 channel=121
    3, -2, -7, 6, -5, -1, 6, -1, -1,
    -- filter=208 channel=122
    15, 0, -3, 14, 0, 2, 15, -4, 0,
    -- filter=208 channel=123
    6, 5, -6, -2, -6, -3, -6, -4, -1,
    -- filter=208 channel=124
    -1, 7, 3, -4, 0, 6, -4, 4, 7,
    -- filter=208 channel=125
    -1, -9, -9, 1, -14, 0, 10, -5, -7,
    -- filter=208 channel=126
    9, -5, -1, 5, 1, -7, -3, 0, -11,
    -- filter=208 channel=127
    4, -5, -3, -1, -3, -3, 0, -4, 3,
    -- filter=209 channel=0
    8, -2, -19, -3, -25, -8, 5, -20, -16,
    -- filter=209 channel=1
    0, -4, -10, -16, -27, -21, -6, -18, -9,
    -- filter=209 channel=2
    9, -2, -4, -2, 3, -2, -6, -3, -4,
    -- filter=209 channel=3
    7, -2, -4, -4, 1, 0, 0, -2, -5,
    -- filter=209 channel=4
    3, 3, 0, -21, -7, -16, -16, -7, -3,
    -- filter=209 channel=5
    -5, -7, -6, -1, -18, -4, 0, -3, -13,
    -- filter=209 channel=6
    2, -6, -7, 2, -7, 6, 0, -7, -3,
    -- filter=209 channel=7
    -2, 6, -6, -4, 0, 6, -3, 1, 4,
    -- filter=209 channel=8
    4, -8, 2, -2, -9, 0, -4, -12, 0,
    -- filter=209 channel=9
    -3, 2, 2, -4, 6, 3, 8, -2, 3,
    -- filter=209 channel=10
    -5, 3, -4, 2, 10, -1, -6, 6, -1,
    -- filter=209 channel=11
    -12, -5, -5, 7, 15, 0, 2, 1, 7,
    -- filter=209 channel=12
    -1, 0, -2, 3, 0, -9, -6, -11, -5,
    -- filter=209 channel=13
    -4, 8, 3, 2, 8, 7, -11, -9, 0,
    -- filter=209 channel=14
    0, 4, -2, -5, 2, 1, 1, 2, -7,
    -- filter=209 channel=15
    8, 6, -4, 10, 10, -1, -10, 2, -3,
    -- filter=209 channel=16
    -5, 0, 3, -14, -9, 3, -9, 3, 3,
    -- filter=209 channel=17
    0, -2, 1, 0, 0, 7, 6, 5, 5,
    -- filter=209 channel=18
    5, 4, -10, 5, 18, 7, -9, -4, -10,
    -- filter=209 channel=19
    0, 0, 6, -2, -1, -5, 4, -1, -1,
    -- filter=209 channel=20
    -11, -11, 3, 1, 17, 9, 0, 17, 6,
    -- filter=209 channel=21
    -11, 3, 7, 4, -7, 6, 7, 12, 3,
    -- filter=209 channel=22
    -4, -10, -5, 0, -4, -1, -2, -9, -7,
    -- filter=209 channel=23
    2, -4, -12, 12, 19, -2, 5, 11, -27,
    -- filter=209 channel=24
    6, 6, -5, -3, 1, 6, 0, 1, 0,
    -- filter=209 channel=25
    9, 7, -8, -8, 2, -5, -18, -7, -2,
    -- filter=209 channel=26
    8, 1, 0, -1, 4, 6, -2, 2, 8,
    -- filter=209 channel=27
    23, 19, -11, 9, 4, -11, -13, 0, -23,
    -- filter=209 channel=28
    -4, 4, 0, -2, -6, 2, 1, -6, 3,
    -- filter=209 channel=29
    -6, 1, -1, 5, 26, 1, -11, 6, 7,
    -- filter=209 channel=30
    10, 12, -7, -7, 1, -15, -3, -8, -3,
    -- filter=209 channel=31
    10, 17, -8, 15, 10, -15, 17, 14, -12,
    -- filter=209 channel=32
    10, 3, -5, -3, 11, -2, -10, -9, -19,
    -- filter=209 channel=33
    15, -1, -4, 11, 10, -1, -11, -4, -12,
    -- filter=209 channel=34
    -11, -9, -4, 2, -23, -26, -11, -17, -13,
    -- filter=209 channel=35
    -4, -1, 3, 6, -1, -2, 0, 3, 0,
    -- filter=209 channel=36
    -4, -1, 7, -7, 7, -7, -9, -7, 5,
    -- filter=209 channel=37
    -5, -11, -9, -6, -23, -12, -15, -25, -6,
    -- filter=209 channel=38
    5, 2, -3, -1, 14, 0, -6, 3, -1,
    -- filter=209 channel=39
    2, 5, 7, 0, 9, 0, -9, 8, 9,
    -- filter=209 channel=40
    -9, 2, 6, 5, 1, 7, 7, 2, 6,
    -- filter=209 channel=41
    -4, -7, 2, -9, -9, 4, -21, -19, -3,
    -- filter=209 channel=42
    -2, 10, -5, 0, -1, 2, 6, 0, -1,
    -- filter=209 channel=43
    2, -3, -8, 1, 0, -2, -6, -5, 0,
    -- filter=209 channel=44
    5, -3, -8, 0, -9, -14, 3, -6, -12,
    -- filter=209 channel=45
    0, 5, 6, 5, -2, 4, 1, 0, -3,
    -- filter=209 channel=46
    -3, -5, -6, -8, 2, -8, 3, -6, 4,
    -- filter=209 channel=47
    -4, -10, 3, -10, -7, -2, -9, -6, 7,
    -- filter=209 channel=48
    14, 9, -1, -7, -2, -12, 0, -12, -10,
    -- filter=209 channel=49
    3, 11, -1, 5, 3, -5, -10, -11, -11,
    -- filter=209 channel=50
    9, 10, -4, 15, 13, -2, 9, 5, -10,
    -- filter=209 channel=51
    -3, -1, -5, -4, -1, -4, -2, 3, -4,
    -- filter=209 channel=52
    -7, -10, -14, 2, -2, -2, -1, -4, -5,
    -- filter=209 channel=53
    -5, 4, 5, -4, 11, 7, 3, 0, -5,
    -- filter=209 channel=54
    5, -6, 1, -5, -4, -6, -3, -6, -5,
    -- filter=209 channel=55
    3, 7, -5, 5, 27, 0, -5, 6, -12,
    -- filter=209 channel=56
    1, -5, -9, 1, -4, -4, -9, -8, -12,
    -- filter=209 channel=57
    -2, -4, 2, -1, 3, -5, -10, -8, -7,
    -- filter=209 channel=58
    -6, -5, 2, 2, -4, -5, 0, 0, 5,
    -- filter=209 channel=59
    6, 12, -1, 6, 9, 0, -6, -7, 2,
    -- filter=209 channel=60
    5, -5, 1, -5, 3, 4, -6, -3, -5,
    -- filter=209 channel=61
    -1, -8, -5, -2, 1, -7, 3, 2, 0,
    -- filter=209 channel=62
    0, -1, -6, 1, -4, 0, -1, 8, 1,
    -- filter=209 channel=63
    0, -1, -3, -4, 4, 6, 7, -4, -2,
    -- filter=209 channel=64
    -9, -3, -5, 1, 4, 7, 0, -5, -4,
    -- filter=209 channel=65
    1, -6, 4, 0, -3, 0, -3, -1, -6,
    -- filter=209 channel=66
    -9, -3, -2, -9, -9, 2, -8, -11, -7,
    -- filter=209 channel=67
    0, -2, 5, -4, 2, -5, -1, 4, 1,
    -- filter=209 channel=68
    -5, 9, 7, -4, -5, 4, -4, 5, 4,
    -- filter=209 channel=69
    -7, 1, -1, -1, -8, -6, 4, -1, 0,
    -- filter=209 channel=70
    18, 0, -4, 5, -3, -20, 3, -5, -24,
    -- filter=209 channel=71
    4, 3, 0, -1, 1, 4, 5, 4, -1,
    -- filter=209 channel=72
    12, 6, 4, 12, 21, 0, 1, 6, 4,
    -- filter=209 channel=73
    6, 11, 1, -2, 13, -9, -13, -3, -15,
    -- filter=209 channel=74
    5, 0, -13, 6, 1, -21, -2, 0, -23,
    -- filter=209 channel=75
    4, -13, -2, -4, -26, -9, -10, -5, -9,
    -- filter=209 channel=76
    -13, -6, 3, -4, 11, 18, -7, 13, 11,
    -- filter=209 channel=77
    -1, -2, -4, -1, -4, 0, 3, 0, -2,
    -- filter=209 channel=78
    -2, -6, -7, -4, -7, 1, 4, -3, -4,
    -- filter=209 channel=79
    8, 10, -6, 2, 19, -2, -18, -6, -21,
    -- filter=209 channel=80
    12, 23, -1, -3, 8, -2, 0, 12, 8,
    -- filter=209 channel=81
    7, 5, 3, -3, 5, 6, 5, 1, 1,
    -- filter=209 channel=82
    -6, -2, 1, -1, -4, 4, 8, 3, 1,
    -- filter=209 channel=83
    -1, 12, 0, 4, 8, 0, -3, 0, -5,
    -- filter=209 channel=84
    3, -1, -7, -3, 0, -11, -17, -3, -9,
    -- filter=209 channel=85
    4, 1, 0, 2, 1, 4, -4, -4, 0,
    -- filter=209 channel=86
    -6, -10, -9, 0, -7, -6, -5, -4, -12,
    -- filter=209 channel=87
    -2, -15, -2, -6, 0, 2, -6, -3, -3,
    -- filter=209 channel=88
    1, 2, 4, 1, -2, -8, 1, 0, -5,
    -- filter=209 channel=89
    11, 14, -3, 9, 26, 10, -1, 2, -13,
    -- filter=209 channel=90
    -4, -1, -2, -4, -1, -5, 1, 7, 3,
    -- filter=209 channel=91
    9, 8, -12, 6, 16, -11, -19, 1, -12,
    -- filter=209 channel=92
    -6, 0, -3, 0, -6, 1, 5, -11, -2,
    -- filter=209 channel=93
    1, -6, -1, -8, -21, -12, -4, -11, 0,
    -- filter=209 channel=94
    -1, 5, -5, -6, -5, 7, 0, -5, -6,
    -- filter=209 channel=95
    -6, 3, 6, -2, 4, 4, -3, 6, 0,
    -- filter=209 channel=96
    2, -3, -4, 4, 3, -3, 1, 5, 6,
    -- filter=209 channel=97
    6, 5, -5, 4, 0, 3, -1, 9, -2,
    -- filter=209 channel=98
    12, 20, 1, 8, 19, -9, -11, -4, -9,
    -- filter=209 channel=99
    5, 8, -8, 11, 19, -17, 2, 10, -20,
    -- filter=209 channel=100
    -6, -5, -4, -4, 4, 2, 2, 3, 0,
    -- filter=209 channel=101
    7, -1, 7, -11, 0, -11, -5, -8, -5,
    -- filter=209 channel=102
    -1, -3, -7, 0, -4, -1, 1, 1, -2,
    -- filter=209 channel=103
    0, -1, -3, -9, -14, -7, -4, -2, 0,
    -- filter=209 channel=104
    2, 13, 8, 9, 9, -5, -3, 9, -4,
    -- filter=209 channel=105
    -15, -9, 3, -6, 5, 4, -8, 6, 4,
    -- filter=209 channel=106
    -4, -7, 4, 1, 9, 5, 2, 7, 5,
    -- filter=209 channel=107
    -4, -4, 0, 5, 2, -7, -8, 7, -3,
    -- filter=209 channel=108
    1, -6, 4, -4, -6, 5, 1, -1, -3,
    -- filter=209 channel=109
    15, 4, -7, 0, 12, -11, -12, -7, -20,
    -- filter=209 channel=110
    5, 0, 0, 1, 4, 1, -3, 8, -4,
    -- filter=209 channel=111
    -2, 1, 5, -5, 0, -4, -9, 3, -1,
    -- filter=209 channel=112
    8, 0, 1, -1, -7, -6, -3, -6, -14,
    -- filter=209 channel=113
    4, 1, -1, 9, 3, 8, -3, 2, -9,
    -- filter=209 channel=114
    5, 5, -4, 0, -4, -17, -12, -9, -21,
    -- filter=209 channel=115
    3, -3, 6, 6, -2, 1, 5, -1, 1,
    -- filter=209 channel=116
    6, 11, 10, 0, 16, -12, -11, 0, -9,
    -- filter=209 channel=117
    4, 0, 2, -1, 4, -2, 6, 3, 7,
    -- filter=209 channel=118
    -7, 7, -1, -7, -5, 5, 5, 2, 4,
    -- filter=209 channel=119
    -6, -15, -5, 0, -11, -7, -10, -15, -14,
    -- filter=209 channel=120
    16, 15, -3, 18, 13, -16, -7, 2, -24,
    -- filter=209 channel=121
    -4, 4, 0, -7, 0, 0, -1, 4, -6,
    -- filter=209 channel=122
    -15, 0, -11, -11, -16, -3, -6, 5, -1,
    -- filter=209 channel=123
    -9, -9, -11, -7, -1, -2, -5, -1, -10,
    -- filter=209 channel=124
    -1, 1, 0, 5, 5, 0, -10, 3, 5,
    -- filter=209 channel=125
    2, 15, 2, 7, 19, -8, 0, -1, -3,
    -- filter=209 channel=126
    -3, -6, -2, 7, 12, 13, -6, 8, 5,
    -- filter=209 channel=127
    -8, -7, 4, 1, 0, -1, 2, -8, -4,
    -- filter=210 channel=0
    4, -3, 2, -4, 0, 5, 2, 2, -6,
    -- filter=210 channel=1
    -6, -7, -6, -5, -6, -1, 5, -4, 0,
    -- filter=210 channel=2
    3, 3, -7, 4, 3, -3, 6, 1, 7,
    -- filter=210 channel=3
    0, -4, -2, 0, -5, 4, 1, -2, 0,
    -- filter=210 channel=4
    1, 4, 1, 3, -7, -3, -7, -5, 1,
    -- filter=210 channel=5
    -5, -4, -5, 3, 3, -2, -1, 0, 5,
    -- filter=210 channel=6
    1, 1, -7, -7, 4, -5, 4, -5, 6,
    -- filter=210 channel=7
    -2, -1, -4, -7, 5, -2, -6, 6, -6,
    -- filter=210 channel=8
    6, -4, -1, -4, -1, -1, 4, -1, -6,
    -- filter=210 channel=9
    -1, 0, -2, -2, 3, 5, 5, 6, -5,
    -- filter=210 channel=10
    7, -2, 0, 4, 1, -3, 0, 5, -7,
    -- filter=210 channel=11
    6, -2, 1, -5, -3, 3, -4, 2, -5,
    -- filter=210 channel=12
    2, 0, 2, -5, -5, -6, 0, 6, 7,
    -- filter=210 channel=13
    4, 3, 6, -3, 0, -1, 6, 3, -1,
    -- filter=210 channel=14
    1, 4, -4, -4, -2, -2, -3, -2, -4,
    -- filter=210 channel=15
    6, -4, 3, -5, -7, 3, 3, -3, -3,
    -- filter=210 channel=16
    -1, 5, 2, -2, 2, 1, 2, -7, -2,
    -- filter=210 channel=17
    -7, 4, 7, -2, -5, 1, -5, 0, -1,
    -- filter=210 channel=18
    0, 0, -5, 0, -1, -6, -2, 6, -3,
    -- filter=210 channel=19
    -3, 4, 0, 5, 0, -2, -6, -3, -2,
    -- filter=210 channel=20
    -6, -4, 1, 4, -6, 0, -5, -6, 0,
    -- filter=210 channel=21
    1, 6, -1, 1, -1, -3, -2, 4, -3,
    -- filter=210 channel=22
    -1, 6, -1, 0, 7, 0, -1, -3, 7,
    -- filter=210 channel=23
    -6, -4, -1, 4, 0, -4, 1, 0, 3,
    -- filter=210 channel=24
    -6, 5, 1, -3, -1, 0, 5, 5, 6,
    -- filter=210 channel=25
    -3, -2, -1, 0, 1, -4, -4, 0, -3,
    -- filter=210 channel=26
    0, 0, 5, 2, -1, -4, -1, 2, -1,
    -- filter=210 channel=27
    -5, 0, 5, 0, 1, -7, -4, -1, 5,
    -- filter=210 channel=28
    -3, 2, 6, 0, 0, 0, 4, -5, -3,
    -- filter=210 channel=29
    -2, -7, 4, -4, -2, -7, -2, 6, -5,
    -- filter=210 channel=30
    -3, 3, -7, 2, -7, 0, 4, -1, -4,
    -- filter=210 channel=31
    -3, 5, 0, 4, 0, -4, 0, -1, 2,
    -- filter=210 channel=32
    0, 0, -1, -3, -2, -5, 0, -5, 1,
    -- filter=210 channel=33
    0, -3, -6, -1, 4, -2, 4, -2, -1,
    -- filter=210 channel=34
    0, 2, 5, 0, -7, -7, 7, 0, -7,
    -- filter=210 channel=35
    0, -4, -5, -3, -4, -5, 1, 6, 5,
    -- filter=210 channel=36
    -4, -7, -2, 0, -5, -5, 0, -5, 2,
    -- filter=210 channel=37
    0, 0, 5, 4, 7, 0, -4, -2, -4,
    -- filter=210 channel=38
    0, 0, 0, -1, 0, -7, 3, -6, 2,
    -- filter=210 channel=39
    -4, -2, 6, 4, -3, 0, -5, -5, 2,
    -- filter=210 channel=40
    3, 2, -4, 5, 4, -4, -2, -5, 3,
    -- filter=210 channel=41
    7, -7, 5, -1, 3, -2, 6, -7, -5,
    -- filter=210 channel=42
    -5, -1, -7, -2, -4, 1, -1, 4, 0,
    -- filter=210 channel=43
    2, -3, 0, -4, 2, 5, 1, 6, -5,
    -- filter=210 channel=44
    -2, 6, -1, 1, -6, -4, 4, -7, 0,
    -- filter=210 channel=45
    6, -1, 2, -5, 3, 3, 0, -1, 5,
    -- filter=210 channel=46
    3, -4, -3, -3, 2, -3, -7, 6, 3,
    -- filter=210 channel=47
    -6, -6, 5, 3, 6, 3, -1, 4, 2,
    -- filter=210 channel=48
    -5, -7, 5, 3, 3, -5, -6, -3, -2,
    -- filter=210 channel=49
    -5, 0, -6, 2, -1, 6, -6, 2, -6,
    -- filter=210 channel=50
    -7, 5, -6, -7, 3, 4, 1, 0, 1,
    -- filter=210 channel=51
    -3, 0, 2, -4, 6, 0, 4, -1, 5,
    -- filter=210 channel=52
    2, 7, -4, 0, -3, 0, 4, 5, 5,
    -- filter=210 channel=53
    4, 6, 2, 5, -1, 0, 5, -3, 0,
    -- filter=210 channel=54
    2, -5, -5, -1, 4, 5, 2, -2, -6,
    -- filter=210 channel=55
    1, 0, -6, 5, -6, 3, 4, 0, -7,
    -- filter=210 channel=56
    4, 0, 0, -1, 3, 2, -1, -6, -2,
    -- filter=210 channel=57
    -3, 2, -6, 1, -2, 0, -6, -6, 7,
    -- filter=210 channel=58
    -5, -5, 0, 2, 6, 0, -7, 0, 0,
    -- filter=210 channel=59
    3, 4, -6, -3, -7, 4, 1, -2, 0,
    -- filter=210 channel=60
    3, -4, -2, -2, 3, -4, -7, 4, 0,
    -- filter=210 channel=61
    -7, 4, 6, 3, 2, -2, 1, 2, 4,
    -- filter=210 channel=62
    -1, -6, 3, 7, 1, -3, 3, 2, 0,
    -- filter=210 channel=63
    1, 0, -3, 0, 4, 3, 0, 3, 2,
    -- filter=210 channel=64
    3, 2, 4, 1, 2, 1, -6, 0, 5,
    -- filter=210 channel=65
    -6, -7, -1, 1, 1, 3, 7, -2, -5,
    -- filter=210 channel=66
    -3, -1, 5, -1, 1, -1, 6, -1, -2,
    -- filter=210 channel=67
    3, 7, -7, -3, -2, 0, -4, -6, -3,
    -- filter=210 channel=68
    2, 0, 1, -5, 0, 7, 0, 1, 0,
    -- filter=210 channel=69
    -5, -3, 6, 5, -4, 1, 3, -7, 6,
    -- filter=210 channel=70
    3, -1, -2, 0, 0, -1, -7, -3, -5,
    -- filter=210 channel=71
    -1, 0, -3, 4, 4, 1, 1, -5, 0,
    -- filter=210 channel=72
    5, -7, 2, -5, -4, -3, -6, 4, 0,
    -- filter=210 channel=73
    0, 1, 0, 1, 3, 1, -4, 5, -5,
    -- filter=210 channel=74
    2, 5, -1, -7, -3, 4, -4, -4, 0,
    -- filter=210 channel=75
    -6, -2, 5, 6, 0, 1, -2, -1, -5,
    -- filter=210 channel=76
    -1, -3, -5, 4, 1, -2, -4, 6, 7,
    -- filter=210 channel=77
    -2, -1, 1, 0, 5, 6, 2, -3, -5,
    -- filter=210 channel=78
    -2, -4, -7, 0, 1, 7, -1, 0, 2,
    -- filter=210 channel=79
    3, 7, 6, 5, -1, 6, 2, -1, 0,
    -- filter=210 channel=80
    -3, 4, -3, -6, 6, 5, -2, -8, -3,
    -- filter=210 channel=81
    4, 2, 6, -6, -5, -5, 4, 4, 0,
    -- filter=210 channel=82
    0, -2, -2, -2, 0, 3, 3, -3, 0,
    -- filter=210 channel=83
    3, 0, -4, 4, 0, 3, -4, -1, 3,
    -- filter=210 channel=84
    2, -5, -3, -3, -6, 3, -6, -2, -2,
    -- filter=210 channel=85
    7, 3, 0, 0, -7, 0, 0, -2, 1,
    -- filter=210 channel=86
    1, 0, 7, 5, 4, 0, 5, 6, 4,
    -- filter=210 channel=87
    1, -7, 1, -2, -2, 0, -2, 3, -6,
    -- filter=210 channel=88
    0, 3, 3, 5, 0, 5, -6, 2, -7,
    -- filter=210 channel=89
    -5, -2, 7, 4, -4, 5, -3, 5, 5,
    -- filter=210 channel=90
    6, 3, 2, 4, -4, 3, -3, -2, -5,
    -- filter=210 channel=91
    -1, -7, -3, 1, -2, 2, 0, -7, -2,
    -- filter=210 channel=92
    0, 3, 2, -6, -6, 6, 6, -1, -5,
    -- filter=210 channel=93
    -6, -3, -1, -1, 7, 4, 3, -1, 3,
    -- filter=210 channel=94
    -6, 3, 2, 2, 0, 1, -4, -4, -5,
    -- filter=210 channel=95
    -7, 2, -2, -4, 0, 6, 0, -1, -2,
    -- filter=210 channel=96
    1, 4, -4, 5, 7, -6, -3, -4, 1,
    -- filter=210 channel=97
    5, 3, 0, 5, -6, 0, 5, 0, 6,
    -- filter=210 channel=98
    -2, 0, -4, 0, -3, 0, -2, 2, 0,
    -- filter=210 channel=99
    -5, 0, 5, -6, -7, -2, 4, 6, -5,
    -- filter=210 channel=100
    0, -4, 5, -5, -5, 1, -6, 3, 0,
    -- filter=210 channel=101
    -6, 3, 7, 4, 6, -1, -3, -6, 5,
    -- filter=210 channel=102
    4, 1, 4, -5, 1, 4, 1, -5, -4,
    -- filter=210 channel=103
    4, 1, 2, 3, 0, 2, -3, -6, -6,
    -- filter=210 channel=104
    4, 1, 3, -4, -3, -4, 6, -2, 4,
    -- filter=210 channel=105
    -2, -4, 2, 4, 4, 3, -1, 2, -5,
    -- filter=210 channel=106
    -5, 0, 0, 2, -2, 0, -2, 2, 1,
    -- filter=210 channel=107
    -6, 0, -3, -2, -6, -7, 1, -2, 5,
    -- filter=210 channel=108
    0, -1, 0, 0, 5, 0, 1, 6, 0,
    -- filter=210 channel=109
    -2, -4, 2, -1, 0, -2, 7, -7, 5,
    -- filter=210 channel=110
    -5, -1, 1, -6, 5, -5, 6, -7, -1,
    -- filter=210 channel=111
    1, 0, -5, 0, 0, 2, 4, -1, -2,
    -- filter=210 channel=112
    4, -2, 6, -6, 2, 7, -5, -4, 3,
    -- filter=210 channel=113
    3, 0, -6, 6, -4, -4, 2, -3, -4,
    -- filter=210 channel=114
    -6, 1, 0, -3, -5, -2, 3, -1, 3,
    -- filter=210 channel=115
    0, 3, 1, 7, 3, -5, 3, -3, -3,
    -- filter=210 channel=116
    0, 0, 1, -7, 4, -7, -6, 1, 4,
    -- filter=210 channel=117
    3, 1, 3, -1, 6, 4, -3, 5, 4,
    -- filter=210 channel=118
    1, -2, 3, 5, 0, -5, 6, 7, 1,
    -- filter=210 channel=119
    6, 5, -7, 3, -2, 7, -1, 4, 2,
    -- filter=210 channel=120
    -4, -1, -5, -4, 0, -7, 1, 0, -5,
    -- filter=210 channel=121
    -3, 1, 2, -2, -3, 3, 0, 5, -2,
    -- filter=210 channel=122
    -3, -7, 0, -4, 5, 3, 5, 4, -6,
    -- filter=210 channel=123
    -6, 0, -3, -6, -3, -3, 4, -3, -2,
    -- filter=210 channel=124
    -5, 1, -3, -5, -6, -1, 2, 6, -3,
    -- filter=210 channel=125
    -5, -2, -1, 1, -7, 3, -2, 0, 6,
    -- filter=210 channel=126
    -5, 0, -6, -2, -2, -3, 3, 0, 4,
    -- filter=210 channel=127
    -5, -6, -1, -5, -1, -4, -3, 5, 6,
    -- filter=211 channel=0
    0, -2, -1, 4, 3, -19, -10, 6, -9,
    -- filter=211 channel=1
    3, -2, 5, 9, 15, -17, -3, 1, 8,
    -- filter=211 channel=2
    2, 1, -8, -7, 5, -6, 3, 0, 0,
    -- filter=211 channel=3
    1, -3, 16, -8, -22, 2, -4, 5, -6,
    -- filter=211 channel=4
    6, -10, -1, -7, 17, -13, 2, -3, 10,
    -- filter=211 channel=5
    6, 2, 2, 10, -6, -3, -2, 6, -3,
    -- filter=211 channel=6
    -1, 5, 0, 5, -2, 0, 4, -5, 6,
    -- filter=211 channel=7
    7, -5, -7, -4, 1, 7, 4, 0, -5,
    -- filter=211 channel=8
    0, 0, 1, -2, -10, 8, -2, -7, 1,
    -- filter=211 channel=9
    6, 0, 10, 7, -12, 0, 1, 8, -5,
    -- filter=211 channel=10
    -4, -4, 9, 3, -2, 4, 4, 13, 0,
    -- filter=211 channel=11
    4, 5, -11, -1, 4, -2, -1, 10, -2,
    -- filter=211 channel=12
    5, 0, 9, -5, 8, -5, -1, 17, 3,
    -- filter=211 channel=13
    12, -8, 7, -10, 15, -12, -6, 10, -1,
    -- filter=211 channel=14
    -2, -2, 3, -5, 6, -7, -6, 0, 0,
    -- filter=211 channel=15
    4, 2, 0, 1, 5, -3, -7, 11, 0,
    -- filter=211 channel=16
    7, -1, 16, 2, -1, 2, 4, 11, -10,
    -- filter=211 channel=17
    2, -4, 4, 1, -3, 6, -2, -2, 0,
    -- filter=211 channel=18
    4, 2, -6, -3, 9, -21, -9, 7, 7,
    -- filter=211 channel=19
    0, 5, 0, -5, -6, -3, 0, 0, 7,
    -- filter=211 channel=20
    -2, -3, -10, -1, 0, -5, -3, 5, 2,
    -- filter=211 channel=21
    0, 0, 9, 4, -6, -8, -5, 2, -6,
    -- filter=211 channel=22
    0, -2, 13, 10, 0, 4, 0, 7, -10,
    -- filter=211 channel=23
    -23, -13, 32, 11, -25, 7, -7, 34, -25,
    -- filter=211 channel=24
    -6, -5, 1, 1, -6, 5, -6, 3, 1,
    -- filter=211 channel=25
    1, -13, 16, -7, 13, -10, -14, 21, 5,
    -- filter=211 channel=26
    -3, -3, 3, 5, 5, -6, -3, 3, -3,
    -- filter=211 channel=27
    0, -27, 19, 16, -10, -14, -22, 21, -18,
    -- filter=211 channel=28
    1, 0, -2, 5, 4, 1, 7, 3, -3,
    -- filter=211 channel=29
    -1, -2, -10, 1, 11, -2, -3, 5, 1,
    -- filter=211 channel=30
    3, -10, 4, 0, -8, -7, -7, 9, -1,
    -- filter=211 channel=31
    -13, -16, 29, 16, -25, -1, -3, 18, -33,
    -- filter=211 channel=32
    -1, -5, 17, 7, 4, -18, -9, 27, 2,
    -- filter=211 channel=33
    -6, -15, 25, 14, -7, -5, -9, 20, -22,
    -- filter=211 channel=34
    -12, 10, 25, 12, -15, 25, -5, 13, -2,
    -- filter=211 channel=35
    2, 3, 5, -6, 7, -4, -6, 6, -3,
    -- filter=211 channel=36
    -2, 3, -7, -8, 2, -5, 0, 9, 12,
    -- filter=211 channel=37
    2, -6, 6, 9, 9, -15, -9, 7, -1,
    -- filter=211 channel=38
    -9, -8, 19, 6, -7, 2, -1, 7, -14,
    -- filter=211 channel=39
    -5, 3, 0, 1, 4, -10, -4, 2, -2,
    -- filter=211 channel=40
    -1, 0, 2, -7, 1, -7, -5, 8, -12,
    -- filter=211 channel=41
    13, 5, 2, -18, 47, -20, 6, -7, 30,
    -- filter=211 channel=42
    0, -4, 5, 7, 1, -9, -5, 0, -4,
    -- filter=211 channel=43
    -9, 4, 3, -2, -17, 7, 3, 11, -5,
    -- filter=211 channel=44
    -5, -5, 13, 11, 0, 0, -1, -1, -5,
    -- filter=211 channel=45
    -7, -9, -3, 5, -7, -10, 1, 4, -9,
    -- filter=211 channel=46
    -4, 3, 0, 2, 1, 8, 6, 1, 0,
    -- filter=211 channel=47
    0, -1, 16, 0, -8, -4, -2, 12, -4,
    -- filter=211 channel=48
    1, -11, 12, 4, -1, -21, -3, 2, -2,
    -- filter=211 channel=49
    5, -12, 3, 0, 4, -9, -7, 0, -1,
    -- filter=211 channel=50
    3, -19, 15, 0, -10, -10, -5, 4, -6,
    -- filter=211 channel=51
    0, -6, -1, 1, 0, 3, -3, 1, 2,
    -- filter=211 channel=52
    -2, -2, 16, 2, 0, 12, 4, 9, -4,
    -- filter=211 channel=53
    1, -4, 6, 3, -5, -6, 5, 12, 2,
    -- filter=211 channel=54
    4, -1, -4, 6, -5, 0, 1, 5, 3,
    -- filter=211 channel=55
    -4, 1, -1, -1, 0, -9, -8, 19, -7,
    -- filter=211 channel=56
    -6, 0, -2, 8, -5, -1, 4, 9, 5,
    -- filter=211 channel=57
    8, 0, -3, 1, 14, 3, 7, -5, 12,
    -- filter=211 channel=58
    7, 3, -7, 12, -2, -2, 1, 7, 7,
    -- filter=211 channel=59
    2, -12, 14, -8, 15, -23, 0, 13, 0,
    -- filter=211 channel=60
    -6, -3, 7, -4, 2, -4, -1, -5, 6,
    -- filter=211 channel=61
    3, -5, 10, -1, -1, 6, -3, 7, 4,
    -- filter=211 channel=62
    3, -6, 2, 0, 2, 3, -2, 3, 0,
    -- filter=211 channel=63
    4, -4, -5, 8, 1, 1, 1, -1, 5,
    -- filter=211 channel=64
    7, 3, -9, -5, 0, -4, 4, 6, -5,
    -- filter=211 channel=65
    6, 4, 2, 0, 0, 0, -3, -6, -2,
    -- filter=211 channel=66
    4, 0, 14, -5, 29, -1, 0, 10, 3,
    -- filter=211 channel=67
    1, -6, -4, 1, 2, -5, 0, 0, -7,
    -- filter=211 channel=68
    7, 5, -7, -3, 12, -4, -7, -4, 2,
    -- filter=211 channel=69
    7, -6, 8, 5, -1, -6, -6, 0, -5,
    -- filter=211 channel=70
    0, -3, 19, 9, -16, 0, -2, 14, -17,
    -- filter=211 channel=71
    -2, -5, 5, -7, -4, 5, 6, 5, -3,
    -- filter=211 channel=72
    8, -17, 7, 6, 3, -16, -1, 14, -15,
    -- filter=211 channel=73
    1, 5, 3, -9, 4, -7, -8, -1, 0,
    -- filter=211 channel=74
    -4, -12, 25, 7, -13, 0, -2, 13, -12,
    -- filter=211 channel=75
    -3, -3, 12, 12, -10, -12, -3, 21, -9,
    -- filter=211 channel=76
    0, 0, -5, -2, 13, -5, -9, 0, -1,
    -- filter=211 channel=77
    -3, -4, -3, -3, 3, 8, 2, 3, -4,
    -- filter=211 channel=78
    -6, -3, 9, -1, -6, 8, 2, -6, 4,
    -- filter=211 channel=79
    3, -13, 20, -7, 3, -23, -14, 31, -9,
    -- filter=211 channel=80
    2, -22, 21, -3, 2, -18, 3, 21, -13,
    -- filter=211 channel=81
    1, 3, 5, 5, -2, 0, -5, -4, 2,
    -- filter=211 channel=82
    -3, 2, 0, 0, -5, 6, -2, 4, -6,
    -- filter=211 channel=83
    -4, -5, -6, 7, -2, -6, 5, -7, -7,
    -- filter=211 channel=84
    4, -2, 0, -7, 9, -7, -5, 15, 2,
    -- filter=211 channel=85
    5, -1, 1, 0, -6, -1, -5, 4, -2,
    -- filter=211 channel=86
    -1, 1, 10, 3, 2, 5, -9, 21, -6,
    -- filter=211 channel=87
    4, 7, 2, 6, -5, 0, -8, 16, 10,
    -- filter=211 channel=88
    0, -4, -4, -3, -8, 8, 7, 3, 5,
    -- filter=211 channel=89
    0, -6, 11, -1, 8, -13, -1, 2, -7,
    -- filter=211 channel=90
    -1, 4, 9, 6, -19, 14, 5, 13, -9,
    -- filter=211 channel=91
    4, -17, 6, 5, 5, -11, -9, 20, -3,
    -- filter=211 channel=92
    1, 5, 10, -2, -2, 18, 9, 1, -2,
    -- filter=211 channel=93
    0, -11, -1, 4, 2, -16, -4, -3, 7,
    -- filter=211 channel=94
    2, 7, 3, -5, 7, -6, 6, 1, 0,
    -- filter=211 channel=95
    2, 1, -3, -5, -7, -3, 1, 0, -5,
    -- filter=211 channel=96
    -5, -9, -1, 0, 9, -3, -3, 0, 7,
    -- filter=211 channel=97
    -5, -5, 5, 3, -9, 0, 4, 6, -13,
    -- filter=211 channel=98
    3, -21, 10, 4, -1, -17, -5, 15, -11,
    -- filter=211 channel=99
    -6, -3, 17, 3, -16, 4, 4, 21, -19,
    -- filter=211 channel=100
    -2, 5, -6, 2, 0, 9, 3, -7, 14,
    -- filter=211 channel=101
    1, -1, 7, -8, 8, -1, 0, -10, 8,
    -- filter=211 channel=102
    5, 1, 4, 4, 6, 6, 4, 6, -3,
    -- filter=211 channel=103
    2, -5, 9, 10, -15, -5, 4, 12, -21,
    -- filter=211 channel=104
    4, -18, 16, 1, -4, -20, -5, 5, -7,
    -- filter=211 channel=105
    6, 1, -6, 0, 10, -8, -7, 0, -2,
    -- filter=211 channel=106
    4, -1, 0, -1, 2, 1, 0, -12, 10,
    -- filter=211 channel=107
    -6, -1, -2, -3, 2, -3, 0, 1, 2,
    -- filter=211 channel=108
    8, 0, -2, -6, 4, 0, 1, 0, 2,
    -- filter=211 channel=109
    7, -22, 19, 5, 6, -10, -13, 22, 1,
    -- filter=211 channel=110
    -8, 0, 16, 2, -1, 4, -1, 16, -10,
    -- filter=211 channel=111
    1, 6, -2, -2, 1, -6, -6, 4, 2,
    -- filter=211 channel=112
    -9, -14, 14, 11, -16, -1, -2, 10, -13,
    -- filter=211 channel=113
    -14, -2, 13, 3, -19, 10, -1, 6, -16,
    -- filter=211 channel=114
    -3, -10, 0, 3, 19, -28, -11, 16, 0,
    -- filter=211 channel=115
    -4, -4, -6, -1, -3, 4, 4, 7, 0,
    -- filter=211 channel=116
    12, -13, -1, -3, 19, -11, -7, 5, 4,
    -- filter=211 channel=117
    1, 0, 2, -10, 8, -14, 3, 0, 7,
    -- filter=211 channel=118
    1, -6, 0, -6, -4, 4, -1, -4, 6,
    -- filter=211 channel=119
    1, 20, 10, 0, -5, 20, 4, 2, 5,
    -- filter=211 channel=120
    -5, -13, 15, 8, -26, -5, -8, 14, -22,
    -- filter=211 channel=121
    5, 3, 1, 3, 7, -6, -3, 11, 0,
    -- filter=211 channel=122
    -2, -9, 19, 11, -1, 4, 7, 13, -15,
    -- filter=211 channel=123
    0, 12, 11, 12, -1, 14, -1, 8, -2,
    -- filter=211 channel=124
    -3, 6, -8, 3, 6, 2, -6, 0, -5,
    -- filter=211 channel=125
    7, -18, 19, 3, -2, -22, -1, 20, -7,
    -- filter=211 channel=126
    5, 0, -7, -5, 11, -14, -4, -5, 0,
    -- filter=211 channel=127
    -5, 6, 0, -2, 4, -6, 3, 3, 11,
    -- filter=212 channel=0
    3, 1, 8, 0, -8, 2, 9, -1, 1,
    -- filter=212 channel=1
    -2, -10, 11, -4, -7, 10, -1, 16, 1,
    -- filter=212 channel=2
    -2, -6, 0, -1, 1, -7, 0, -6, -3,
    -- filter=212 channel=3
    7, 14, 1, 5, 0, -16, 7, -8, -1,
    -- filter=212 channel=4
    7, 5, -6, -2, 0, -21, -1, -5, -23,
    -- filter=212 channel=5
    -2, -10, 0, 1, -12, 5, 5, -3, -3,
    -- filter=212 channel=6
    1, 3, 4, 3, 8, -5, 5, -2, -3,
    -- filter=212 channel=7
    0, 0, -1, -4, 4, -3, -6, 7, 3,
    -- filter=212 channel=8
    -8, 0, 1, -10, 3, 12, 7, -4, 4,
    -- filter=212 channel=9
    3, -9, -5, -4, -7, 6, 0, -5, 4,
    -- filter=212 channel=10
    -11, 1, 1, 0, -7, 11, 0, -4, -5,
    -- filter=212 channel=11
    0, 0, -3, -2, 5, -6, 10, -6, -8,
    -- filter=212 channel=12
    1, 7, 9, -3, 6, 22, -1, 18, 18,
    -- filter=212 channel=13
    4, 2, 4, 4, -3, 13, -4, 13, -4,
    -- filter=212 channel=14
    -3, 6, 0, -1, -4, -3, -4, 5, 1,
    -- filter=212 channel=15
    -7, -9, 2, 7, 0, -1, -2, -6, -9,
    -- filter=212 channel=16
    -4, 5, 11, -6, -5, 13, 3, -10, 13,
    -- filter=212 channel=17
    -2, -6, -2, -3, 1, 2, 0, 0, 0,
    -- filter=212 channel=18
    0, -12, 3, 9, -10, -5, -4, 2, -16,
    -- filter=212 channel=19
    0, 6, 6, 5, 6, 1, -7, 2, 1,
    -- filter=212 channel=20
    0, 6, -9, 9, 5, 4, 3, 0, 8,
    -- filter=212 channel=21
    0, -2, 9, -3, -18, 19, -1, -18, -3,
    -- filter=212 channel=22
    4, -1, 2, -3, -9, 10, 6, -6, 8,
    -- filter=212 channel=23
    -7, 0, 10, 1, -19, 19, -5, -25, 11,
    -- filter=212 channel=24
    6, 1, 5, -5, -5, 7, 0, 0, -5,
    -- filter=212 channel=25
    -10, -2, 16, -7, -10, 19, -4, -5, 10,
    -- filter=212 channel=26
    0, 2, 0, -7, -5, 4, -6, 4, 6,
    -- filter=212 channel=27
    -11, -5, 16, 10, -32, 18, 5, -29, 5,
    -- filter=212 channel=28
    -7, 0, -4, -2, -3, -3, -7, -6, -7,
    -- filter=212 channel=29
    0, -5, -8, 8, -2, -10, -1, 0, 1,
    -- filter=212 channel=30
    7, 3, -4, 2, -10, 8, 5, -4, 3,
    -- filter=212 channel=31
    -3, -7, 20, 0, -31, 20, -9, -37, 9,
    -- filter=212 channel=32
    -6, -12, 0, 7, -15, 5, 8, -3, 3,
    -- filter=212 channel=33
    1, -7, 7, 0, -13, 6, 1, -14, 2,
    -- filter=212 channel=34
    -13, 6, 17, -13, 3, 35, -11, -12, 33,
    -- filter=212 channel=35
    3, 0, -4, -5, 0, -1, -6, -5, 6,
    -- filter=212 channel=36
    0, 1, 1, -10, 3, 12, -10, -4, 10,
    -- filter=212 channel=37
    9, -7, 9, 0, -5, 5, 6, 6, 4,
    -- filter=212 channel=38
    -4, -9, 4, 3, -8, 10, 0, -15, 9,
    -- filter=212 channel=39
    8, 1, 2, -3, 0, -9, 5, 9, 1,
    -- filter=212 channel=40
    0, -5, -3, -3, -2, 2, 5, 1, -4,
    -- filter=212 channel=41
    -7, 9, 8, -14, 10, 21, -13, 24, 11,
    -- filter=212 channel=42
    9, -7, 0, 0, -3, -14, 0, 0, -10,
    -- filter=212 channel=43
    2, 3, -2, -4, 8, -7, 2, -6, 6,
    -- filter=212 channel=44
    8, -3, 15, 2, -4, 15, -1, -1, 4,
    -- filter=212 channel=45
    1, -3, -5, 0, -5, -6, -2, 0, -2,
    -- filter=212 channel=46
    -4, -2, -4, -8, 6, -3, 5, 0, -1,
    -- filter=212 channel=47
    -1, 0, 6, -1, -6, 5, 4, -14, 9,
    -- filter=212 channel=48
    -3, 0, 3, -4, -10, 14, -1, -15, 3,
    -- filter=212 channel=49
    2, -9, -8, 1, -3, -15, 8, -7, -19,
    -- filter=212 channel=50
    -3, 0, 15, -5, -10, 12, 4, -9, 2,
    -- filter=212 channel=51
    -4, 2, -2, -7, 0, 0, 0, 3, 0,
    -- filter=212 channel=52
    -6, 3, 7, 0, 4, 15, -2, -3, 13,
    -- filter=212 channel=53
    -1, -1, 3, -4, -7, -6, 1, 5, -2,
    -- filter=212 channel=54
    -4, 5, 5, -6, 7, -1, -5, -2, 0,
    -- filter=212 channel=55
    -13, -6, 6, -4, 0, 8, -7, 0, 2,
    -- filter=212 channel=56
    -2, 6, 7, -5, -4, 15, -2, -2, 17,
    -- filter=212 channel=57
    -5, 8, 5, 1, 9, 8, -5, 8, -4,
    -- filter=212 channel=58
    3, -6, 1, 1, 4, -3, 1, 7, -6,
    -- filter=212 channel=59
    -6, -3, 9, 1, -16, 17, -8, -11, -6,
    -- filter=212 channel=60
    2, -1, 4, -5, 6, 3, -7, -4, -3,
    -- filter=212 channel=61
    4, -5, 3, -9, 6, 6, -3, -3, 1,
    -- filter=212 channel=62
    -6, -5, -3, 5, 0, 0, -6, 5, -6,
    -- filter=212 channel=63
    -8, -2, -5, 1, 4, 3, 2, 5, -1,
    -- filter=212 channel=64
    0, 7, -1, -7, -2, 8, -5, 3, -3,
    -- filter=212 channel=65
    0, 4, 0, -2, 6, -4, 5, 2, -3,
    -- filter=212 channel=66
    -3, -1, 8, -13, 15, 30, -10, 26, 14,
    -- filter=212 channel=67
    -4, -3, 0, -8, 0, -5, 2, 6, 2,
    -- filter=212 channel=68
    6, 7, -3, -2, -2, -8, 6, 9, 3,
    -- filter=212 channel=69
    3, -7, -1, 6, 0, 5, 3, 6, 5,
    -- filter=212 channel=70
    -1, -7, 15, 4, -10, 9, 7, -11, 6,
    -- filter=212 channel=71
    0, 2, 8, 4, 2, 1, -6, -10, -1,
    -- filter=212 channel=72
    -8, 1, 16, -10, -20, 10, -4, -20, 2,
    -- filter=212 channel=73
    5, 0, 1, -6, 0, -7, -2, 2, 1,
    -- filter=212 channel=74
    0, 0, 20, -2, -10, 36, -6, -20, 16,
    -- filter=212 channel=75
    -2, -8, 0, 4, -8, -10, 5, 2, 1,
    -- filter=212 channel=76
    -5, -6, 3, 7, 1, -1, 1, 9, -1,
    -- filter=212 channel=77
    -2, -1, -1, 6, -5, 1, -4, 0, 6,
    -- filter=212 channel=78
    0, -2, -2, -5, -1, 5, -5, -7, 6,
    -- filter=212 channel=79
    -8, 0, 12, 13, -16, -4, 1, -5, -6,
    -- filter=212 channel=80
    -5, -12, 21, 0, -22, 17, -1, -13, 0,
    -- filter=212 channel=81
    5, -6, -2, 0, 5, -4, 0, 0, -4,
    -- filter=212 channel=82
    2, -4, -1, -1, 4, -6, 0, 4, 3,
    -- filter=212 channel=83
    -7, -6, -6, 0, -6, 6, 2, -9, -8,
    -- filter=212 channel=84
    -1, 2, 4, 0, 0, 0, -1, -7, 0,
    -- filter=212 channel=85
    -3, 4, -3, 6, 0, 4, -6, 0, 2,
    -- filter=212 channel=86
    -5, -7, 2, 5, -8, 16, -3, -2, 14,
    -- filter=212 channel=87
    4, -8, 4, 0, 4, 10, -4, 0, 17,
    -- filter=212 channel=88
    -7, -2, 12, -9, 2, 18, -5, -13, 9,
    -- filter=212 channel=89
    -8, -10, 14, 1, -7, 10, -11, 2, -2,
    -- filter=212 channel=90
    -11, 6, 16, -3, -4, 20, -16, -8, 10,
    -- filter=212 channel=91
    -3, -11, -3, 4, -9, 0, 1, -19, -2,
    -- filter=212 channel=92
    -1, 3, 11, -12, -1, 13, 3, 2, 17,
    -- filter=212 channel=93
    5, 2, 5, 10, -8, 10, 12, -6, 0,
    -- filter=212 channel=94
    -4, 3, 1, 2, -6, 6, 4, 1, 2,
    -- filter=212 channel=95
    2, 3, -2, 0, 4, -3, 4, -5, 2,
    -- filter=212 channel=96
    3, -3, 5, -2, -2, -9, -4, 6, -11,
    -- filter=212 channel=97
    -6, -1, 3, 1, -5, -7, -6, -11, 4,
    -- filter=212 channel=98
    -7, -5, 12, 2, -23, 3, -3, -17, 3,
    -- filter=212 channel=99
    -14, 2, 10, -6, -21, 36, -11, -29, 20,
    -- filter=212 channel=100
    -5, -4, 3, 2, 5, 12, -7, 0, 10,
    -- filter=212 channel=101
    8, 6, 3, 0, 0, -8, 2, 2, -17,
    -- filter=212 channel=102
    -6, 1, 0, -4, -2, 0, -6, 6, 4,
    -- filter=212 channel=103
    -3, 4, 9, 7, -16, 7, -1, -19, 2,
    -- filter=212 channel=104
    -5, -12, 5, -7, -9, 11, -8, -16, 3,
    -- filter=212 channel=105
    7, -4, -3, 7, 5, -4, 0, 10, 9,
    -- filter=212 channel=106
    6, -6, -6, 1, 7, -10, 1, 3, 4,
    -- filter=212 channel=107
    8, 0, 2, -2, 5, 1, 7, -3, 9,
    -- filter=212 channel=108
    -10, -3, 0, 0, 4, -8, -3, 9, 0,
    -- filter=212 channel=109
    -11, -11, 0, 4, -18, 17, 2, -22, -1,
    -- filter=212 channel=110
    0, -2, 11, -8, 0, 10, -5, -11, 7,
    -- filter=212 channel=111
    1, 6, -1, 3, 7, 8, 0, 5, -4,
    -- filter=212 channel=112
    0, -12, 9, -1, -16, 20, 5, -15, 3,
    -- filter=212 channel=113
    -13, -5, 13, -2, -10, 16, 6, -11, 12,
    -- filter=212 channel=114
    7, -2, 0, 2, -13, -6, 15, -2, -6,
    -- filter=212 channel=115
    6, -3, -5, 6, -1, 2, 4, 3, 1,
    -- filter=212 channel=116
    2, -2, 1, -8, -16, -3, 0, -1, -9,
    -- filter=212 channel=117
    3, -1, 3, -1, -2, 0, -7, 0, -7,
    -- filter=212 channel=118
    7, 5, 4, 0, 7, -3, -6, 4, 2,
    -- filter=212 channel=119
    -6, 6, 11, -11, 7, 31, -10, -4, 34,
    -- filter=212 channel=120
    0, -2, 5, 2, -20, 16, 10, -32, 18,
    -- filter=212 channel=121
    -11, 5, -2, -9, -3, 10, 0, 0, 0,
    -- filter=212 channel=122
    0, 6, 24, -3, -10, 33, -1, -23, 16,
    -- filter=212 channel=123
    -4, -2, 7, -6, 8, 16, -5, -4, 13,
    -- filter=212 channel=124
    10, -3, -6, 2, -4, 4, 3, 6, 0,
    -- filter=212 channel=125
    -1, -7, 15, -9, -20, 24, 0, -22, -1,
    -- filter=212 channel=126
    0, 0, 4, -5, -1, 0, -1, 8, -2,
    -- filter=212 channel=127
    -2, -4, -4, -6, 7, -2, -10, 1, 0,
    -- filter=213 channel=0
    7, 3, -13, 18, 0, -16, 12, 7, -4,
    -- filter=213 channel=1
    4, 5, -2, 15, 11, -9, 2, 13, 1,
    -- filter=213 channel=2
    -6, 2, 1, -4, -9, -5, 5, -1, -3,
    -- filter=213 channel=3
    -3, -6, -3, 0, -1, -15, 0, -3, -8,
    -- filter=213 channel=4
    -3, -5, -6, 6, -10, -14, 8, 10, -10,
    -- filter=213 channel=5
    -2, 1, 10, 6, -1, 7, 4, 0, 3,
    -- filter=213 channel=6
    1, -6, 0, 7, -9, -10, 5, -4, -12,
    -- filter=213 channel=7
    -4, 2, -1, 4, -3, -2, 1, 0, 3,
    -- filter=213 channel=8
    -3, -9, 0, -2, -1, -4, 8, -1, 5,
    -- filter=213 channel=9
    -6, 0, 0, -8, -7, -1, 4, 5, 6,
    -- filter=213 channel=10
    -9, 0, 4, -1, 0, 4, -12, 2, 5,
    -- filter=213 channel=11
    -1, -1, -2, 8, -8, -8, -4, -4, 1,
    -- filter=213 channel=12
    2, 7, 3, -6, 4, 6, 1, -2, -2,
    -- filter=213 channel=13
    5, 3, 4, -8, 4, -18, -1, 5, -4,
    -- filter=213 channel=14
    -5, 1, -2, -6, -5, 2, 2, 5, -5,
    -- filter=213 channel=15
    11, 4, -12, 0, -7, -21, -1, -6, -18,
    -- filter=213 channel=16
    -15, -6, 19, -9, -4, 21, -10, 9, 8,
    -- filter=213 channel=17
    6, -3, -2, -4, -5, 2, 0, 0, 3,
    -- filter=213 channel=18
    12, 0, -27, 1, 2, -28, 0, 0, -22,
    -- filter=213 channel=19
    -3, -5, 3, -1, 6, -7, 3, 4, 4,
    -- filter=213 channel=20
    0, 3, -15, 1, -1, -15, 2, -6, -17,
    -- filter=213 channel=21
    -15, -4, 15, -24, 12, 31, -5, 7, 21,
    -- filter=213 channel=22
    4, 0, -13, 9, -2, -9, 4, -7, -10,
    -- filter=213 channel=23
    11, -3, -4, 6, -12, -23, 3, -15, -15,
    -- filter=213 channel=24
    -7, 0, 0, 3, -4, 0, -7, 0, 2,
    -- filter=213 channel=25
    4, 6, 3, -6, 8, -16, -1, 4, 7,
    -- filter=213 channel=26
    -12, -10, 1, -9, -6, 5, -2, 5, 15,
    -- filter=213 channel=27
    14, -7, -16, 3, -9, -38, 16, 2, -6,
    -- filter=213 channel=28
    3, 4, -5, 0, 5, -5, -6, 3, 3,
    -- filter=213 channel=29
    3, -6, -10, 8, -4, -14, -2, 4, -12,
    -- filter=213 channel=30
    -6, 1, -7, 0, -7, -12, 6, 4, -2,
    -- filter=213 channel=31
    -12, -5, 17, -22, -14, 17, -5, -8, 5,
    -- filter=213 channel=32
    13, 7, -12, 3, -9, -29, 14, 0, -12,
    -- filter=213 channel=33
    9, 11, -6, 2, -7, -25, 9, -4, -18,
    -- filter=213 channel=34
    2, -3, 1, 0, -9, -6, 12, -12, -1,
    -- filter=213 channel=35
    4, -2, -5, -1, 6, 4, -2, 2, -6,
    -- filter=213 channel=36
    -8, -11, 10, -10, 5, 10, -12, 5, 3,
    -- filter=213 channel=37
    -8, 7, 2, 14, 0, 3, -2, 6, 1,
    -- filter=213 channel=38
    0, 3, 5, 3, -10, -4, 5, -6, 2,
    -- filter=213 channel=39
    3, -1, -10, -2, 5, -8, 2, -4, -10,
    -- filter=213 channel=40
    1, 0, -11, 1, -4, -4, 7, 0, -12,
    -- filter=213 channel=41
    4, -7, 14, -2, 5, 2, -11, -2, 4,
    -- filter=213 channel=42
    -2, -6, -7, 0, 0, -9, -3, 2, -1,
    -- filter=213 channel=43
    9, -6, -16, 11, -6, -20, -1, -1, -12,
    -- filter=213 channel=44
    -4, -1, 11, -9, 6, 1, 1, 8, 13,
    -- filter=213 channel=45
    -5, 1, -3, 1, -1, 0, 6, 4, -5,
    -- filter=213 channel=46
    -1, 4, 0, 0, 0, 2, -1, 0, -4,
    -- filter=213 channel=47
    -18, -7, 15, -22, 6, 20, -2, 6, 23,
    -- filter=213 channel=48
    0, 0, -3, -7, -2, -2, -4, 11, 3,
    -- filter=213 channel=49
    10, 4, -18, 11, -7, -13, 4, -7, -14,
    -- filter=213 channel=50
    -4, 2, 1, -1, 3, -1, 2, -4, 1,
    -- filter=213 channel=51
    2, 6, 5, 6, -5, -1, -1, 6, -6,
    -- filter=213 channel=52
    6, 0, 3, -1, -11, -11, -3, -8, -6,
    -- filter=213 channel=53
    -2, -2, -1, 4, -7, -1, 2, 1, -2,
    -- filter=213 channel=54
    4, 4, -5, -2, 0, -2, -1, -2, 1,
    -- filter=213 channel=55
    6, -2, -13, 7, -1, -22, 9, -1, -13,
    -- filter=213 channel=56
    5, -9, -1, -3, -2, 4, 7, 4, 3,
    -- filter=213 channel=57
    1, -4, 0, -7, 0, -3, -3, -2, -7,
    -- filter=213 channel=58
    -8, -3, 7, 0, 9, 5, -7, 1, 7,
    -- filter=213 channel=59
    4, 4, -4, -9, -1, 4, -3, 3, 6,
    -- filter=213 channel=60
    0, -1, 7, 4, -7, -1, 5, 4, -1,
    -- filter=213 channel=61
    1, 2, 8, 1, 4, 6, 5, -2, 2,
    -- filter=213 channel=62
    -5, 3, 0, -7, 0, 5, -5, 1, 0,
    -- filter=213 channel=63
    -5, 4, 6, -10, 0, 14, -2, -2, 12,
    -- filter=213 channel=64
    -6, 3, 0, 3, 3, 2, 2, -3, -3,
    -- filter=213 channel=65
    6, 1, -1, -4, -2, 0, 6, 0, -3,
    -- filter=213 channel=66
    0, 1, 0, -2, 0, 7, 2, 9, 4,
    -- filter=213 channel=67
    4, 0, 3, -5, 3, -5, -4, -2, 0,
    -- filter=213 channel=68
    -5, -6, 2, -2, -2, 0, 1, 6, 4,
    -- filter=213 channel=69
    3, 0, 8, 4, 6, 3, 0, -5, 5,
    -- filter=213 channel=70
    3, -5, -6, 11, -8, -11, 13, -9, -18,
    -- filter=213 channel=71
    -3, -2, 5, 0, 0, 5, 1, 0, -1,
    -- filter=213 channel=72
    -6, -4, 4, -13, -3, 14, -11, 5, 14,
    -- filter=213 channel=73
    11, -1, -16, 0, -4, -17, 0, -2, 0,
    -- filter=213 channel=74
    7, -10, 0, 2, -13, -8, 2, 0, 0,
    -- filter=213 channel=75
    6, 12, 5, 5, 14, -6, 0, 0, -4,
    -- filter=213 channel=76
    11, -5, -16, 3, -8, -18, 10, -8, -6,
    -- filter=213 channel=77
    6, -3, 3, 0, -5, -3, 5, -2, 0,
    -- filter=213 channel=78
    -2, 3, -1, -11, -5, 9, -10, -6, 0,
    -- filter=213 channel=79
    14, 8, -30, 13, -8, -37, 6, -10, -25,
    -- filter=213 channel=80
    -22, 2, 6, -14, 0, 16, -5, 9, 20,
    -- filter=213 channel=81
    2, -5, 1, -2, -7, 1, 3, 6, -2,
    -- filter=213 channel=82
    0, 1, 5, -2, -8, -7, -3, 4, -7,
    -- filter=213 channel=83
    0, -1, 3, -2, 5, -2, -5, 6, 5,
    -- filter=213 channel=84
    2, -7, -3, 1, -8, -23, 0, -2, -12,
    -- filter=213 channel=85
    0, 6, 7, 2, -5, 4, 2, -3, 0,
    -- filter=213 channel=86
    -6, -11, -6, 4, 0, 0, -3, -8, -4,
    -- filter=213 channel=87
    1, -5, -9, 2, -10, -4, 0, 0, -8,
    -- filter=213 channel=88
    -2, 3, 5, -10, 4, 11, -6, 0, 18,
    -- filter=213 channel=89
    -6, 1, 0, -1, 0, -17, 1, 8, 4,
    -- filter=213 channel=90
    -9, -8, 8, -6, -7, 11, -2, 1, 13,
    -- filter=213 channel=91
    6, -1, -16, 5, -8, -17, 1, -5, -4,
    -- filter=213 channel=92
    5, 4, 1, 6, 0, 3, 6, -6, -2,
    -- filter=213 channel=93
    -9, 1, 14, 0, 8, 15, -5, 13, 13,
    -- filter=213 channel=94
    -2, 1, -2, 5, 4, 0, 0, -5, 1,
    -- filter=213 channel=95
    5, 2, -2, -8, -5, 2, -4, 2, -3,
    -- filter=213 channel=96
    -5, -3, -6, 0, 5, 3, 0, 6, 6,
    -- filter=213 channel=97
    -1, 2, 0, 0, 3, 4, 2, 0, -7,
    -- filter=213 channel=98
    0, 6, 0, -4, 0, -17, -1, 4, -2,
    -- filter=213 channel=99
    -2, 0, 0, -7, -8, 6, -6, -4, 14,
    -- filter=213 channel=100
    -8, -5, 4, -5, -5, -3, -5, -4, -6,
    -- filter=213 channel=101
    -3, -6, -4, -6, -3, -4, 5, 8, -1,
    -- filter=213 channel=102
    -6, 2, -7, -4, 0, -1, -5, 2, 0,
    -- filter=213 channel=103
    -15, 0, 13, -4, 11, 29, -6, 0, 7,
    -- filter=213 channel=104
    -16, 1, 14, -10, -4, 23, -18, 1, 13,
    -- filter=213 channel=105
    0, 4, 0, -2, 6, -11, -4, 3, -6,
    -- filter=213 channel=106
    0, 2, -2, -3, 4, 1, -5, 0, 0,
    -- filter=213 channel=107
    13, 2, -10, 4, -12, -28, 3, -15, -16,
    -- filter=213 channel=108
    -2, -3, 7, 6, -1, -6, 3, 0, 0,
    -- filter=213 channel=109
    11, -10, -7, 0, -2, -19, 8, -1, 0,
    -- filter=213 channel=110
    -3, -2, 11, -14, -9, 4, -4, 0, 1,
    -- filter=213 channel=111
    5, 3, 4, 0, -1, 1, -6, 2, 8,
    -- filter=213 channel=112
    -2, -4, 1, 7, -7, -1, 6, 1, 4,
    -- filter=213 channel=113
    -6, 8, -3, -4, -5, -2, 1, -5, 3,
    -- filter=213 channel=114
    17, 9, -33, 18, -4, -44, 17, -1, -21,
    -- filter=213 channel=115
    -5, 1, -4, -5, -3, -3, 4, 0, 2,
    -- filter=213 channel=116
    1, 0, -11, -9, 5, -15, -4, 3, -3,
    -- filter=213 channel=117
    0, 5, 5, -10, 7, -2, 0, 8, 2,
    -- filter=213 channel=118
    1, -4, -4, 1, -1, -4, 6, 2, 7,
    -- filter=213 channel=119
    -2, -6, 0, -2, -10, 2, -3, 0, 3,
    -- filter=213 channel=120
    15, -10, -13, 11, -10, -18, 14, -14, 2,
    -- filter=213 channel=121
    1, 1, 0, -2, 1, 2, -6, 6, 4,
    -- filter=213 channel=122
    -19, -5, 35, -26, 12, 43, -23, 13, 39,
    -- filter=213 channel=123
    0, 8, 10, 2, 0, 5, -6, -4, -2,
    -- filter=213 channel=124
    -3, -6, -12, -1, 0, -3, 6, -2, 0,
    -- filter=213 channel=125
    -2, -8, -2, -6, -8, -3, -6, -1, 5,
    -- filter=213 channel=126
    1, 10, 2, -5, 6, -1, 2, 12, -8,
    -- filter=213 channel=127
    -7, 2, -3, -1, 5, 0, 0, 7, -1,
    -- filter=214 channel=0
    3, 3, -5, 2, -8, -9, 6, -2, -7,
    -- filter=214 channel=1
    9, 0, 0, 1, -6, -12, 2, 2, 0,
    -- filter=214 channel=2
    -2, -6, -2, 0, 0, -5, -3, -3, -4,
    -- filter=214 channel=3
    1, 0, 9, -5, -2, 4, -2, 0, 5,
    -- filter=214 channel=4
    -5, -4, 5, -4, -1, -10, -2, -7, -10,
    -- filter=214 channel=5
    -1, 0, 8, 1, 2, 7, 3, 2, -3,
    -- filter=214 channel=6
    -4, -4, -7, -4, -8, -2, 0, 0, 3,
    -- filter=214 channel=7
    -6, -1, 2, -1, 5, 2, -1, 7, -3,
    -- filter=214 channel=8
    2, -9, -6, -7, -3, -6, -7, -7, -8,
    -- filter=214 channel=9
    3, 7, 1, 5, -6, -5, 0, 0, -8,
    -- filter=214 channel=10
    10, 8, -3, -1, 5, -5, -2, 0, -8,
    -- filter=214 channel=11
    -7, 4, -7, -1, -3, 7, 3, 6, -3,
    -- filter=214 channel=12
    -2, 3, -6, 2, -11, -4, 0, -3, -4,
    -- filter=214 channel=13
    1, -3, 1, 1, -14, -9, 1, -12, -2,
    -- filter=214 channel=14
    1, 4, 6, 4, 7, -6, 0, 5, -3,
    -- filter=214 channel=15
    -1, 2, -5, -2, -12, 0, -4, -2, -8,
    -- filter=214 channel=16
    4, 10, 12, 12, 9, 7, 3, 10, -2,
    -- filter=214 channel=17
    0, 7, 4, 2, 3, 0, 0, 0, -3,
    -- filter=214 channel=18
    -1, -10, 0, -11, -10, -20, -15, -17, -17,
    -- filter=214 channel=19
    0, 5, 2, -5, -4, -5, 3, 0, -2,
    -- filter=214 channel=20
    0, -6, 0, 5, -4, -1, -1, 1, 3,
    -- filter=214 channel=21
    11, 8, 9, 18, 11, 9, 11, 6, 7,
    -- filter=214 channel=22
    1, -4, 1, -5, -7, -6, -8, 1, -7,
    -- filter=214 channel=23
    -6, 6, -2, -1, -13, 0, -15, -18, -15,
    -- filter=214 channel=24
    3, -4, -3, 1, -4, -2, 0, 4, 3,
    -- filter=214 channel=25
    2, -8, -10, 1, -6, -5, -1, -9, -11,
    -- filter=214 channel=26
    5, -1, 3, 10, 4, 3, 0, 2, 3,
    -- filter=214 channel=27
    2, -2, -6, -13, -17, -18, -18, -23, -15,
    -- filter=214 channel=28
    -4, 1, 2, 4, -2, 5, -3, -7, -7,
    -- filter=214 channel=29
    -9, 4, -4, 3, 0, -3, -8, 0, 1,
    -- filter=214 channel=30
    1, 2, 0, -8, -2, -2, 1, -9, -3,
    -- filter=214 channel=31
    10, 9, 11, 10, 3, 10, 1, -12, -2,
    -- filter=214 channel=32
    -3, -8, -1, -14, -9, -19, -3, -13, -6,
    -- filter=214 channel=33
    1, 6, 3, -6, -18, -7, -7, -16, -9,
    -- filter=214 channel=34
    -4, 2, -1, 0, -13, -10, 1, -1, -1,
    -- filter=214 channel=35
    -6, -7, 4, 2, -3, 0, 6, 5, -3,
    -- filter=214 channel=36
    10, 3, -3, -1, 2, 8, 0, 1, 10,
    -- filter=214 channel=37
    9, 0, -2, 9, 0, 0, -4, 3, -4,
    -- filter=214 channel=38
    4, -5, -1, -4, -8, -5, -3, -9, -10,
    -- filter=214 channel=39
    6, 2, -3, -7, 2, 4, -1, 4, -2,
    -- filter=214 channel=40
    4, 9, 1, -4, 0, -2, 0, 3, -4,
    -- filter=214 channel=41
    1, 5, -10, 2, -8, -16, -6, -3, -7,
    -- filter=214 channel=42
    -2, 4, -5, 5, -6, -8, 0, -8, 0,
    -- filter=214 channel=43
    -6, 3, -2, -8, 0, 0, 5, 0, 0,
    -- filter=214 channel=44
    8, -5, 10, -3, -6, -1, 4, -10, -9,
    -- filter=214 channel=45
    -3, 1, -2, 0, 3, -3, -4, -4, -5,
    -- filter=214 channel=46
    -4, 0, 1, -4, 5, -7, 5, 2, -5,
    -- filter=214 channel=47
    4, 11, 9, 14, 1, 8, 12, -6, 5,
    -- filter=214 channel=48
    5, 2, 0, 3, -7, -2, -5, -11, -12,
    -- filter=214 channel=49
    -5, -4, 3, 0, -2, -2, 2, -8, 0,
    -- filter=214 channel=50
    6, -8, -7, 2, -10, -1, -4, -9, -2,
    -- filter=214 channel=51
    4, -5, 7, 2, -6, 4, -1, 5, 1,
    -- filter=214 channel=52
    7, -5, 0, 3, -6, -5, 2, 3, -6,
    -- filter=214 channel=53
    -8, 0, -4, -5, -4, -4, -8, 4, -4,
    -- filter=214 channel=54
    0, -4, -2, -5, 7, -4, 0, 6, 3,
    -- filter=214 channel=55
    -8, -6, -1, -6, -13, -10, -4, -16, -7,
    -- filter=214 channel=56
    0, 2, 1, 4, -7, 4, 1, -3, -2,
    -- filter=214 channel=57
    0, 7, -5, 0, 3, 0, -3, 2, 5,
    -- filter=214 channel=58
    0, 6, 4, -1, -3, 3, 0, 4, -1,
    -- filter=214 channel=59
    0, 3, 0, -5, -3, -13, 2, -10, -8,
    -- filter=214 channel=60
    0, 1, -2, 0, -2, -5, -4, 3, -4,
    -- filter=214 channel=61
    7, 0, 1, 3, 5, -4, -2, -7, -1,
    -- filter=214 channel=62
    4, -3, -2, 3, 0, 5, -1, -6, 6,
    -- filter=214 channel=63
    -2, 8, 0, 4, 7, 10, 7, 4, 1,
    -- filter=214 channel=64
    0, 3, -2, 2, 5, 3, 6, -2, 5,
    -- filter=214 channel=65
    3, -2, 0, -2, -2, 0, -1, 3, -3,
    -- filter=214 channel=66
    -4, -9, -3, 3, 0, 0, 2, -7, 3,
    -- filter=214 channel=67
    0, -7, -6, -2, -5, 7, -3, -3, 4,
    -- filter=214 channel=68
    5, -3, -2, 6, -4, 3, 0, -6, 0,
    -- filter=214 channel=69
    -4, 5, 0, -5, -4, 4, -4, 3, 2,
    -- filter=214 channel=70
    5, -9, -2, -1, -7, -8, -15, -11, -5,
    -- filter=214 channel=71
    0, 5, -1, -1, 2, 8, 8, 3, -2,
    -- filter=214 channel=72
    1, 7, 4, -1, 5, 0, -9, -6, 0,
    -- filter=214 channel=73
    -5, -5, -1, -6, -1, -10, -12, -5, -5,
    -- filter=214 channel=74
    -2, -6, -9, 2, -13, -5, -7, -12, 0,
    -- filter=214 channel=75
    3, 6, 9, 6, -3, 0, 1, -2, -9,
    -- filter=214 channel=76
    3, 0, 3, -3, 2, 7, 6, -4, 2,
    -- filter=214 channel=77
    5, -5, -5, 6, -2, -6, 4, 3, -3,
    -- filter=214 channel=78
    -5, 1, 8, -3, 3, 9, -4, 3, 3,
    -- filter=214 channel=79
    -2, -8, -10, -12, -20, -9, -10, -6, -22,
    -- filter=214 channel=80
    11, 6, 10, 7, -4, -4, -5, -7, -10,
    -- filter=214 channel=81
    7, 4, 4, -2, -3, -4, -5, 0, -3,
    -- filter=214 channel=82
    6, 5, -3, -5, -5, -4, -1, 0, -2,
    -- filter=214 channel=83
    -3, -5, 4, 6, -4, -1, -9, 2, -2,
    -- filter=214 channel=84
    -6, -10, -7, -9, -13, -4, -9, -3, -7,
    -- filter=214 channel=85
    -4, 2, 1, 6, -5, 3, 1, -6, 3,
    -- filter=214 channel=86
    8, -6, -6, -6, -6, 0, -4, -3, -6,
    -- filter=214 channel=87
    -6, -10, 2, 1, 2, -3, -5, 1, 5,
    -- filter=214 channel=88
    10, 4, 5, 5, 7, 0, 2, 2, 4,
    -- filter=214 channel=89
    -3, -4, 2, -3, -12, -9, -9, -14, -17,
    -- filter=214 channel=90
    2, 0, 7, 12, 4, 7, 3, -3, 8,
    -- filter=214 channel=91
    -4, -13, -5, -2, -13, -5, -10, -6, -9,
    -- filter=214 channel=92
    7, 0, 3, 0, 0, -8, 3, -4, -1,
    -- filter=214 channel=93
    2, -7, 6, 8, 1, -1, -3, 1, -8,
    -- filter=214 channel=94
    1, 1, -1, -4, 6, 0, -5, 3, 0,
    -- filter=214 channel=95
    2, -4, -5, -6, 4, -2, 5, -1, -6,
    -- filter=214 channel=96
    3, 4, 3, 6, -4, 1, -1, 1, 2,
    -- filter=214 channel=97
    1, 9, 14, 7, 9, 7, 4, 7, 5,
    -- filter=214 channel=98
    0, 4, -7, -5, -9, -5, 0, -10, -13,
    -- filter=214 channel=99
    2, 2, 4, -4, -6, -5, -9, -4, 0,
    -- filter=214 channel=100
    0, -6, -8, 2, 3, 0, -1, -6, 0,
    -- filter=214 channel=101
    3, -3, -4, -2, -6, -5, -7, -4, -8,
    -- filter=214 channel=102
    -3, -6, 7, 4, -4, 2, 4, 3, 1,
    -- filter=214 channel=103
    3, 2, 5, 11, -2, 13, 0, 0, 0,
    -- filter=214 channel=104
    5, 5, 5, 10, -2, 1, 0, 1, -2,
    -- filter=214 channel=105
    -2, -5, -4, 1, -1, 6, 4, -5, 4,
    -- filter=214 channel=106
    -2, 2, 2, 9, 6, 0, 1, 7, -1,
    -- filter=214 channel=107
    1, 2, -4, 0, -5, -9, 1, 4, 0,
    -- filter=214 channel=108
    -2, 6, -5, -6, 0, 6, -2, -4, 2,
    -- filter=214 channel=109
    -8, -13, 0, -13, -21, -11, -17, -10, -14,
    -- filter=214 channel=110
    7, 8, 7, 4, 6, 3, 6, 0, 2,
    -- filter=214 channel=111
    6, 0, -6, -4, 3, 2, -5, 5, 0,
    -- filter=214 channel=112
    -3, 0, 3, -3, -3, 1, 1, -5, -5,
    -- filter=214 channel=113
    9, 6, 0, 2, -10, 0, 1, 0, -6,
    -- filter=214 channel=114
    -6, -14, -9, -1, -15, -21, -1, -17, -10,
    -- filter=214 channel=115
    3, -3, 1, 3, -5, 7, 1, 1, 4,
    -- filter=214 channel=116
    4, 0, -9, 0, -7, -13, -4, -8, -11,
    -- filter=214 channel=117
    -2, -3, -6, 2, -8, -8, 5, 1, -8,
    -- filter=214 channel=118
    1, -4, 6, 0, 6, 3, 0, 3, -4,
    -- filter=214 channel=119
    -8, -1, -6, -3, -8, -3, -11, -6, 0,
    -- filter=214 channel=120
    0, -11, -10, -10, -14, -10, -8, -8, -11,
    -- filter=214 channel=121
    7, -2, 7, 4, -1, 0, 4, -10, -10,
    -- filter=214 channel=122
    20, 8, 24, 22, 15, 10, 12, -2, 11,
    -- filter=214 channel=123
    -1, -1, -1, 4, -7, -3, 5, -3, 0,
    -- filter=214 channel=124
    -7, 1, -1, -3, 1, 3, -2, -3, -8,
    -- filter=214 channel=125
    6, -7, 0, 3, -4, -9, -8, -16, -10,
    -- filter=214 channel=126
    -2, 8, -1, 5, -10, -12, -1, 3, -13,
    -- filter=214 channel=127
    1, 3, -1, 0, 0, -6, -2, 0, 0,
    -- filter=215 channel=0
    5, 0, -1, -7, -8, 2, -4, -9, -6,
    -- filter=215 channel=1
    2, 6, 1, -4, -6, 4, -9, 0, -1,
    -- filter=215 channel=2
    -4, 2, 1, -4, 4, -6, 6, 1, 6,
    -- filter=215 channel=3
    1, -3, -1, 0, 3, 1, 6, 1, -3,
    -- filter=215 channel=4
    2, 1, 2, -2, 1, -2, -4, 7, 2,
    -- filter=215 channel=5
    9, 2, 0, -1, 2, -5, 3, -2, -5,
    -- filter=215 channel=6
    7, 1, 6, -6, -3, 7, -1, 2, -3,
    -- filter=215 channel=7
    2, 3, 6, -1, 0, -6, 7, 0, 4,
    -- filter=215 channel=8
    -4, 0, -5, 6, 4, -1, 6, 5, 0,
    -- filter=215 channel=9
    -3, -7, -2, -3, -3, 1, -1, 0, 0,
    -- filter=215 channel=10
    8, -3, 2, 4, -3, -4, -8, -1, -7,
    -- filter=215 channel=11
    6, -6, 8, 0, 7, 0, -1, 1, 2,
    -- filter=215 channel=12
    -2, -4, 5, -1, 6, 6, -6, 5, -1,
    -- filter=215 channel=13
    3, -7, 6, -6, 0, -2, -8, 4, 6,
    -- filter=215 channel=14
    1, 4, 4, -1, 5, 0, -6, -5, 6,
    -- filter=215 channel=15
    7, 4, 1, 5, -9, 6, -10, 1, 0,
    -- filter=215 channel=16
    6, 6, 5, 4, 2, 0, -4, 4, 3,
    -- filter=215 channel=17
    6, -3, -2, 7, 1, 7, 1, -7, -7,
    -- filter=215 channel=18
    5, -4, 3, -4, -3, 7, -4, -3, 1,
    -- filter=215 channel=19
    0, 4, 0, 6, -5, -6, 2, 5, 2,
    -- filter=215 channel=20
    -5, -6, 2, 5, 0, -2, 2, 1, 5,
    -- filter=215 channel=21
    4, 6, -3, 6, 1, -3, -1, 2, 4,
    -- filter=215 channel=22
    1, -4, 4, -7, 0, 7, 4, 7, 4,
    -- filter=215 channel=23
    3, 4, 3, 2, 4, -1, 0, 0, 5,
    -- filter=215 channel=24
    3, 1, -5, -3, -3, 6, 5, 0, -6,
    -- filter=215 channel=25
    4, -5, -6, 0, -3, -7, 0, 4, 1,
    -- filter=215 channel=26
    1, 3, -3, 2, 7, -3, -1, 1, -3,
    -- filter=215 channel=27
    3, 2, 7, -11, 0, 1, -11, -9, 2,
    -- filter=215 channel=28
    0, 0, -5, 4, -2, 0, 6, 6, -4,
    -- filter=215 channel=29
    -5, -6, 0, -4, 0, 0, -2, 4, 0,
    -- filter=215 channel=30
    0, -7, -4, 0, -5, 2, -3, 0, -1,
    -- filter=215 channel=31
    -2, -4, -8, -6, 2, 1, 2, 4, -7,
    -- filter=215 channel=32
    4, 0, 7, -1, -9, 1, -11, 0, 8,
    -- filter=215 channel=33
    6, -7, 8, -5, -11, 2, -7, -3, -6,
    -- filter=215 channel=34
    -2, 5, -2, -5, 6, 3, 6, 11, -4,
    -- filter=215 channel=35
    -1, 3, -4, 3, -1, 5, -5, 0, -1,
    -- filter=215 channel=36
    0, -5, 2, 1, 7, -6, 0, 2, -2,
    -- filter=215 channel=37
    3, -3, 0, 3, -5, -5, -6, 1, 0,
    -- filter=215 channel=38
    4, 4, -6, 1, 3, 3, -4, 0, 1,
    -- filter=215 channel=39
    1, 1, -2, -3, -5, -6, -3, -7, -2,
    -- filter=215 channel=40
    -4, 7, 5, -4, -3, 3, 0, -3, 1,
    -- filter=215 channel=41
    8, 7, -5, 12, 0, 7, -7, 4, -2,
    -- filter=215 channel=42
    1, 1, 0, -1, -7, -1, -6, 4, 4,
    -- filter=215 channel=43
    2, -4, 4, 0, 0, 7, -1, -2, -3,
    -- filter=215 channel=44
    -6, -4, -5, 0, 6, -1, -6, 6, -8,
    -- filter=215 channel=45
    7, 1, 0, -4, 6, -3, 4, -6, -4,
    -- filter=215 channel=46
    -3, 3, 1, 0, -6, 7, -7, -4, 0,
    -- filter=215 channel=47
    6, 0, -4, -5, 5, -2, -2, 7, 4,
    -- filter=215 channel=48
    6, -9, -6, 0, -7, -2, -5, -7, -1,
    -- filter=215 channel=49
    -1, -8, 2, -3, -3, 6, -3, -5, 0,
    -- filter=215 channel=50
    -6, -6, 5, -2, -5, -1, 3, -6, -8,
    -- filter=215 channel=51
    3, 4, -2, 0, 7, -5, 5, -2, -5,
    -- filter=215 channel=52
    -4, 0, 0, 3, -3, 6, 5, -3, 0,
    -- filter=215 channel=53
    1, 4, 3, 5, 2, 8, 3, -3, 0,
    -- filter=215 channel=54
    4, 5, 0, 0, 2, 3, -6, -7, -3,
    -- filter=215 channel=55
    0, 0, -3, 0, -5, 6, -2, -7, -3,
    -- filter=215 channel=56
    -3, 0, 0, 4, 6, 4, 1, -4, 3,
    -- filter=215 channel=57
    4, -3, -4, -1, 4, 5, -5, 6, 6,
    -- filter=215 channel=58
    0, 8, 5, 3, 0, -7, 0, -1, 3,
    -- filter=215 channel=59
    3, 1, 0, -2, 0, -2, -9, 6, 0,
    -- filter=215 channel=60
    1, -1, -4, 4, -3, -1, 1, -2, 1,
    -- filter=215 channel=61
    -3, 0, -3, -3, 9, -4, -2, 3, 4,
    -- filter=215 channel=62
    5, 6, -6, -6, -3, 1, 4, 0, -2,
    -- filter=215 channel=63
    -1, 7, -2, 6, 0, -4, -4, 0, -1,
    -- filter=215 channel=64
    -1, 3, -5, -2, 6, 7, 2, -2, 6,
    -- filter=215 channel=65
    0, 3, -3, 0, 4, -2, 3, -4, -3,
    -- filter=215 channel=66
    -5, -4, -1, 2, 0, 0, 0, -5, 2,
    -- filter=215 channel=67
    3, -6, 1, 4, -5, 3, 2, 0, -7,
    -- filter=215 channel=68
    3, 4, 4, 4, -6, 0, -6, 1, -1,
    -- filter=215 channel=69
    3, -5, -5, 7, -3, 4, -6, -5, 3,
    -- filter=215 channel=70
    5, 6, 7, -4, 1, -4, 0, 0, 3,
    -- filter=215 channel=71
    6, 1, 3, 7, -1, -8, 5, 0, -6,
    -- filter=215 channel=72
    -1, -7, -1, 7, 4, -2, -4, -1, -3,
    -- filter=215 channel=73
    6, 2, -4, 0, 1, 4, -6, 6, 4,
    -- filter=215 channel=74
    -5, 0, 1, 3, 5, -2, 4, 7, 6,
    -- filter=215 channel=75
    11, 6, -1, 10, -6, 3, -10, 0, -5,
    -- filter=215 channel=76
    -2, -1, -1, 3, -4, 0, 2, 1, 7,
    -- filter=215 channel=77
    5, 3, 0, 7, 7, -4, 0, 4, 1,
    -- filter=215 channel=78
    4, -4, 4, -5, 7, -1, 6, -1, 6,
    -- filter=215 channel=79
    13, -3, 9, 2, -11, 10, -12, -9, 1,
    -- filter=215 channel=80
    -3, -4, 1, -3, -4, 5, -6, -2, -5,
    -- filter=215 channel=81
    0, -4, -7, -5, 4, 7, 2, 2, -2,
    -- filter=215 channel=82
    2, -5, 3, -2, 6, -3, 3, -6, -4,
    -- filter=215 channel=83
    -7, -3, 1, 1, -1, 6, 0, 6, 4,
    -- filter=215 channel=84
    8, -4, 3, -2, 4, 6, -6, 1, 0,
    -- filter=215 channel=85
    5, -3, 5, -2, 1, 6, 0, 0, 0,
    -- filter=215 channel=86
    7, 6, 0, 4, -3, 3, 3, 0, 1,
    -- filter=215 channel=87
    8, -1, 2, 3, 7, 2, -3, -2, -6,
    -- filter=215 channel=88
    3, 5, -5, 4, 9, -1, 1, 6, 2,
    -- filter=215 channel=89
    7, -2, 0, 6, -4, -5, -9, -7, 5,
    -- filter=215 channel=90
    0, 0, -4, -3, 6, -5, 2, 5, 4,
    -- filter=215 channel=91
    -2, -1, 0, -9, -5, -4, -7, -7, 4,
    -- filter=215 channel=92
    -4, 7, -6, -5, -1, -3, -3, 1, 5,
    -- filter=215 channel=93
    3, 7, -6, 3, 3, 3, 0, -3, -10,
    -- filter=215 channel=94
    0, 6, -7, 6, -5, -5, 4, -2, 0,
    -- filter=215 channel=95
    2, 5, 0, -1, -5, 2, -4, 6, -2,
    -- filter=215 channel=96
    5, -5, 3, 6, 0, 5, 1, 0, 1,
    -- filter=215 channel=97
    -5, 6, -6, 3, 4, 1, -2, -5, 1,
    -- filter=215 channel=98
    -5, 0, 7, -5, -6, -2, -11, -4, 3,
    -- filter=215 channel=99
    4, 4, 1, -1, 3, -5, 2, 7, -3,
    -- filter=215 channel=100
    4, 7, -4, -3, 1, -4, 0, -6, 7,
    -- filter=215 channel=101
    2, -2, -1, 0, -5, -7, 1, -4, -2,
    -- filter=215 channel=102
    2, 4, 3, 4, -4, -1, -3, -1, 4,
    -- filter=215 channel=103
    4, 1, 5, 0, 4, -9, 0, 1, -4,
    -- filter=215 channel=104
    -2, -6, 0, 0, 5, 1, -7, 9, 0,
    -- filter=215 channel=105
    7, -1, -4, 0, -1, -2, 0, 5, 1,
    -- filter=215 channel=106
    -1, 4, -3, 5, 3, -1, -4, -6, 1,
    -- filter=215 channel=107
    4, 1, 8, -2, 0, 1, -6, -5, -5,
    -- filter=215 channel=108
    2, -4, 7, 3, 4, -3, -2, -7, 1,
    -- filter=215 channel=109
    4, -5, 3, 0, -5, 7, -4, -8, -2,
    -- filter=215 channel=110
    8, 3, -4, 8, 5, 1, -1, 2, 1,
    -- filter=215 channel=111
    3, -5, 4, 0, -7, -6, 2, 4, 0,
    -- filter=215 channel=112
    4, 6, 0, 0, 3, 5, 1, 5, 4,
    -- filter=215 channel=113
    -2, -3, -6, 1, -1, 6, -4, -1, 0,
    -- filter=215 channel=114
    12, -8, -1, -2, -11, 6, -12, -7, -5,
    -- filter=215 channel=115
    5, 3, 1, 0, 1, 1, 3, -1, 3,
    -- filter=215 channel=116
    0, 2, -2, -5, -1, 2, 0, -8, 4,
    -- filter=215 channel=117
    -4, -2, -3, -4, 5, 5, -1, 1, -3,
    -- filter=215 channel=118
    5, 1, 1, 5, -6, 7, -4, -1, 2,
    -- filter=215 channel=119
    -1, 12, 7, -8, 0, 5, -1, 11, 2,
    -- filter=215 channel=120
    -5, -7, -1, -4, -5, -2, 3, 8, -7,
    -- filter=215 channel=121
    -2, 8, -2, -3, 2, 2, 2, -4, -2,
    -- filter=215 channel=122
    -6, 0, -6, -4, 1, 2, 0, 3, 3,
    -- filter=215 channel=123
    3, 3, 0, 7, -2, 1, 4, -1, -5,
    -- filter=215 channel=124
    1, 2, -5, 6, 1, 0, -5, -6, 5,
    -- filter=215 channel=125
    0, -11, 3, -9, 0, 1, 2, -2, -5,
    -- filter=215 channel=126
    3, -5, -5, 12, -4, 7, -3, -4, 3,
    -- filter=215 channel=127
    2, 1, -4, -5, -6, 4, -3, -4, 1,
    -- filter=216 channel=0
    -4, -7, 1, -9, -2, 0, -10, -4, 0,
    -- filter=216 channel=1
    -12, -9, -8, -10, -20, 1, -13, -15, -2,
    -- filter=216 channel=2
    1, 4, 4, -3, 6, -3, -4, 4, 3,
    -- filter=216 channel=3
    0, -3, -9, 2, -6, -7, 0, -6, -2,
    -- filter=216 channel=4
    3, -2, -15, -2, -7, 0, 2, -8, 1,
    -- filter=216 channel=5
    -11, -5, 6, -17, -13, -3, -3, -4, 8,
    -- filter=216 channel=6
    4, -5, -5, 6, 2, -6, 5, -2, -3,
    -- filter=216 channel=7
    3, 4, -1, -3, 1, -5, -3, 0, -2,
    -- filter=216 channel=8
    -6, 4, -3, 1, 0, 4, -7, -4, -1,
    -- filter=216 channel=9
    -4, -3, 1, 0, -2, 5, 5, 0, 11,
    -- filter=216 channel=10
    -7, -9, 6, 2, -6, 6, -8, -9, 3,
    -- filter=216 channel=11
    6, -2, -2, 0, -3, 3, 7, -6, -1,
    -- filter=216 channel=12
    0, 1, -1, 3, -7, -7, -2, -8, -1,
    -- filter=216 channel=13
    -3, -5, 0, -6, -11, -5, 0, -8, 7,
    -- filter=216 channel=14
    0, 3, 4, 2, -7, -2, -6, 3, 7,
    -- filter=216 channel=15
    -6, 0, -1, 0, 3, 3, -6, -4, 0,
    -- filter=216 channel=16
    -2, 0, 0, -6, -11, 6, -9, 0, 2,
    -- filter=216 channel=17
    -2, 0, -2, -4, 3, -3, 1, -2, -5,
    -- filter=216 channel=18
    -4, -2, 4, 1, -6, 0, -4, -17, 9,
    -- filter=216 channel=19
    2, 5, -5, -6, -5, 0, -2, 3, 0,
    -- filter=216 channel=20
    -4, -9, -1, 3, 7, -9, 1, 0, 0,
    -- filter=216 channel=21
    -17, -7, 7, -8, -5, 11, -14, 4, 6,
    -- filter=216 channel=22
    5, 0, -5, -1, -2, -3, -5, 5, 1,
    -- filter=216 channel=23
    0, 10, 14, -5, 4, 0, -6, 13, 9,
    -- filter=216 channel=24
    -4, -5, 1, -1, 0, 2, 5, 6, -6,
    -- filter=216 channel=25
    -12, -5, 18, -14, -5, 6, -15, -8, 21,
    -- filter=216 channel=26
    -11, 0, 8, -13, -8, -2, -9, -11, -1,
    -- filter=216 channel=27
    -8, 12, 22, -14, 2, 12, -17, -2, 28,
    -- filter=216 channel=28
    4, 3, 1, 0, 0, 3, 6, -3, 7,
    -- filter=216 channel=29
    0, 2, -4, 3, 3, 0, 9, 3, -3,
    -- filter=216 channel=30
    5, 2, 5, -3, -9, -3, -8, -2, 1,
    -- filter=216 channel=31
    -18, 1, 22, -15, 11, 21, -8, 15, 27,
    -- filter=216 channel=32
    -5, 3, -2, -2, 0, 3, -4, -8, 5,
    -- filter=216 channel=33
    -9, -3, 10, -4, -1, 10, -10, -8, 5,
    -- filter=216 channel=34
    2, -1, 0, -9, -3, 1, -2, 0, 12,
    -- filter=216 channel=35
    -4, -3, 6, 2, 5, 5, -3, 7, -5,
    -- filter=216 channel=36
    0, -8, 4, -5, -7, 0, -3, -9, -3,
    -- filter=216 channel=37
    -5, -4, -8, -17, -17, -10, -9, -14, -3,
    -- filter=216 channel=38
    -1, 8, 5, -2, -3, 0, -10, -2, 4,
    -- filter=216 channel=39
    -4, -4, -8, -1, 0, 3, 1, -4, -5,
    -- filter=216 channel=40
    -4, -9, -4, -2, -1, 1, 5, -4, -7,
    -- filter=216 channel=41
    -4, -9, 6, -7, -21, 2, -14, -12, 0,
    -- filter=216 channel=42
    0, 7, 8, 0, -3, 0, 0, -4, 6,
    -- filter=216 channel=43
    0, -6, -4, 2, 2, -9, 5, 0, -1,
    -- filter=216 channel=44
    -6, -1, 0, -22, -11, 10, -13, 2, 2,
    -- filter=216 channel=45
    5, -4, -7, -2, 0, -7, 2, 5, -5,
    -- filter=216 channel=46
    -7, 0, 3, -6, 5, 0, -2, 2, -4,
    -- filter=216 channel=47
    -17, -4, 13, -14, -12, 8, -17, -2, 9,
    -- filter=216 channel=48
    0, -5, 15, -19, -1, 18, -6, 3, 22,
    -- filter=216 channel=49
    7, 5, 3, -4, -6, -3, -3, -3, 0,
    -- filter=216 channel=50
    -5, 8, 9, -1, 11, 12, -6, 7, 16,
    -- filter=216 channel=51
    4, -7, 5, 4, 3, 7, 3, 1, 5,
    -- filter=216 channel=52
    -6, -1, -4, -4, -1, 0, -7, -5, 1,
    -- filter=216 channel=53
    1, -4, -4, 6, 0, 4, 3, -6, 1,
    -- filter=216 channel=54
    0, -1, 3, 1, -5, 1, -5, -6, 7,
    -- filter=216 channel=55
    -6, -1, 1, -3, 5, 6, -7, -5, 0,
    -- filter=216 channel=56
    -6, 3, -4, 0, -6, 10, 5, -2, 5,
    -- filter=216 channel=57
    5, -3, -1, 0, -9, 4, -8, -9, 2,
    -- filter=216 channel=58
    -5, -5, -8, -4, -8, -1, -7, -2, -1,
    -- filter=216 channel=59
    -2, -5, 17, -18, -1, 13, -14, -10, 18,
    -- filter=216 channel=60
    3, -2, -3, -5, -1, 4, 2, -3, 4,
    -- filter=216 channel=61
    -2, 1, -3, 5, 6, -4, -6, -2, -5,
    -- filter=216 channel=62
    2, 5, 1, 3, 6, 1, -7, -7, -3,
    -- filter=216 channel=63
    1, -5, 0, 0, -11, 2, -1, -8, 0,
    -- filter=216 channel=64
    2, 3, 2, 4, 4, 0, -1, 0, 0,
    -- filter=216 channel=65
    5, 2, 0, -3, -7, -4, 3, -6, 0,
    -- filter=216 channel=66
    -6, -1, 0, -10, -14, 0, -2, -3, 3,
    -- filter=216 channel=67
    4, 3, -6, -2, -4, -4, 0, -5, -4,
    -- filter=216 channel=68
    -6, -1, -1, 5, -4, 0, 1, -1, -2,
    -- filter=216 channel=69
    6, -3, 1, 1, 2, 1, 0, 0, 8,
    -- filter=216 channel=70
    -6, 9, 2, -4, 6, 0, 0, 8, 9,
    -- filter=216 channel=71
    3, -7, -7, 5, 0, 0, -2, -4, 0,
    -- filter=216 channel=72
    -7, -1, 19, -14, -3, 19, -4, -5, 14,
    -- filter=216 channel=73
    3, 2, -1, -1, -4, 2, -7, 6, 7,
    -- filter=216 channel=74
    -5, 3, 9, -13, 13, 13, -9, 1, 6,
    -- filter=216 channel=75
    -6, -8, -6, -11, -12, -2, -4, -9, -2,
    -- filter=216 channel=76
    6, -13, -8, 6, -5, -16, -1, -2, -15,
    -- filter=216 channel=77
    -8, 5, -2, 5, 0, -5, -4, 3, 2,
    -- filter=216 channel=78
    -9, -5, 8, 0, 1, 4, 2, 5, 1,
    -- filter=216 channel=79
    0, -10, 3, -14, -6, -7, -1, -19, -3,
    -- filter=216 channel=80
    -5, 2, 24, -13, -2, 27, -12, 0, 24,
    -- filter=216 channel=81
    4, 1, 6, -4, 7, -3, 5, -7, 0,
    -- filter=216 channel=82
    3, -6, -3, 2, -5, -5, -7, 1, -6,
    -- filter=216 channel=83
    -1, 10, 0, -8, 2, 15, -10, 4, 7,
    -- filter=216 channel=84
    -2, 4, -5, -4, -3, 6, -5, -6, -3,
    -- filter=216 channel=85
    -7, -2, 5, 6, 5, -6, -4, -5, 0,
    -- filter=216 channel=86
    4, -3, -6, -5, -11, 2, -8, -4, 0,
    -- filter=216 channel=87
    1, -1, -7, 0, -6, -7, -1, 0, 2,
    -- filter=216 channel=88
    -9, 2, -1, 3, -2, 6, 1, -1, -5,
    -- filter=216 channel=89
    -13, 0, 9, -6, -4, 9, -5, -3, 4,
    -- filter=216 channel=90
    1, -6, -2, 1, 0, 0, -8, 2, 1,
    -- filter=216 channel=91
    1, 9, 9, -14, 3, -1, -11, 0, 14,
    -- filter=216 channel=92
    0, 0, -5, 0, 0, 0, -1, -3, 0,
    -- filter=216 channel=93
    -3, -5, 7, -17, -8, 0, -10, -3, 9,
    -- filter=216 channel=94
    4, 1, -4, 1, 4, 4, -4, 1, 0,
    -- filter=216 channel=95
    -6, 0, 2, -4, -2, -1, -2, -7, 0,
    -- filter=216 channel=96
    -1, -3, 2, -6, -7, -4, -1, 0, 1,
    -- filter=216 channel=97
    1, 0, -2, 0, 8, -2, 4, -1, -6,
    -- filter=216 channel=98
    -12, 7, 19, -9, -5, 23, -5, -7, 25,
    -- filter=216 channel=99
    -10, 14, 6, -10, 7, 21, -13, 14, 19,
    -- filter=216 channel=100
    2, -6, -5, 0, -4, -3, -3, 6, 6,
    -- filter=216 channel=101
    -1, 5, -6, -6, -3, -6, -3, 1, -10,
    -- filter=216 channel=102
    2, 4, -4, -6, -4, 3, -5, 5, 7,
    -- filter=216 channel=103
    -14, -4, 14, -7, 0, 6, -16, 3, 4,
    -- filter=216 channel=104
    -15, 1, 15, -12, 4, 22, -11, 5, 11,
    -- filter=216 channel=105
    -3, -1, -6, 10, -7, -7, 9, 0, -12,
    -- filter=216 channel=106
    -4, -8, 0, 0, -6, -1, 6, -1, -9,
    -- filter=216 channel=107
    -3, -5, -5, -1, 3, -3, 1, 1, -3,
    -- filter=216 channel=108
    -9, -3, 5, -4, -1, 4, 3, -8, -1,
    -- filter=216 channel=109
    -10, 6, 22, -7, -3, 9, -8, -2, 27,
    -- filter=216 channel=110
    -5, 5, 5, 2, 2, 7, 0, -2, 7,
    -- filter=216 channel=111
    -7, 5, -6, 3, -8, 5, 4, -8, -4,
    -- filter=216 channel=112
    0, -2, 3, 0, 7, 2, -6, 0, 9,
    -- filter=216 channel=113
    -6, 1, 6, -4, 8, 11, -12, 2, 7,
    -- filter=216 channel=114
    0, -1, -6, -12, -19, -10, -5, -3, 8,
    -- filter=216 channel=115
    3, -1, -4, -6, -1, -2, 4, 6, 5,
    -- filter=216 channel=116
    4, 9, 17, -5, -7, 10, -14, 2, 15,
    -- filter=216 channel=117
    -3, -3, -6, 0, -1, -3, -4, 1, -2,
    -- filter=216 channel=118
    7, -4, 0, -2, 5, 6, 0, 1, -1,
    -- filter=216 channel=119
    -7, 2, 12, -6, 0, 4, 0, 10, 2,
    -- filter=216 channel=120
    -6, 20, 15, -5, 14, 17, -14, 12, 26,
    -- filter=216 channel=121
    1, -2, 4, -10, -5, 0, -5, -3, -2,
    -- filter=216 channel=122
    -25, -16, 1, -24, -17, 17, -21, -3, 22,
    -- filter=216 channel=123
    0, 0, -4, -2, 7, 3, 4, 5, 7,
    -- filter=216 channel=124
    -1, -3, -7, -1, 0, -6, 8, 1, 5,
    -- filter=216 channel=125
    -13, 3, 15, -19, 7, 11, -18, 3, 23,
    -- filter=216 channel=126
    -2, -4, 0, -1, -4, -3, -1, -14, 7,
    -- filter=216 channel=127
    1, 0, 3, -3, -6, 5, -8, 1, -1,
    -- filter=217 channel=0
    4, -10, 6, -9, 2, 9, 8, -6, -3,
    -- filter=217 channel=1
    -2, -6, 1, 0, 16, 11, 7, -9, -9,
    -- filter=217 channel=2
    2, 5, 6, 7, 6, -8, -2, 5, 8,
    -- filter=217 channel=3
    21, 4, -7, 6, 32, 19, 4, 6, 0,
    -- filter=217 channel=4
    -11, 26, 0, 44, 25, -6, -10, 17, 25,
    -- filter=217 channel=5
    -10, -8, -1, 0, 9, 0, 2, 0, 2,
    -- filter=217 channel=6
    -6, -10, 0, 7, 2, 0, 4, -2, 4,
    -- filter=217 channel=7
    2, 7, -1, 3, 0, 0, 3, -4, 0,
    -- filter=217 channel=8
    1, 16, 6, 14, 2, -1, -6, -5, 6,
    -- filter=217 channel=9
    -11, -7, 0, 3, 15, 3, -3, -7, -4,
    -- filter=217 channel=10
    9, -13, -14, 1, 15, 18, 0, -8, -7,
    -- filter=217 channel=11
    -4, -5, 4, 5, 12, 4, -1, -4, 2,
    -- filter=217 channel=12
    6, -3, 1, -7, 13, -6, 2, -4, -6,
    -- filter=217 channel=13
    6, -16, -10, -3, 31, 16, 0, -11, -10,
    -- filter=217 channel=14
    3, -3, 6, -3, -1, 5, -3, 0, -2,
    -- filter=217 channel=15
    -9, -14, -4, -2, 14, 12, 8, -10, -9,
    -- filter=217 channel=16
    -1, -12, -3, 5, 3, 9, 3, 6, -6,
    -- filter=217 channel=17
    3, -4, 1, -7, 5, 6, 0, 3, -3,
    -- filter=217 channel=18
    -23, -24, 1, -1, 32, 7, 10, -12, -19,
    -- filter=217 channel=19
    -4, 3, -2, 4, 5, 6, 5, 0, -2,
    -- filter=217 channel=20
    -9, 2, 3, 12, 20, 11, -6, 0, 1,
    -- filter=217 channel=21
    -9, -7, 2, -3, 3, 0, -5, 0, 1,
    -- filter=217 channel=22
    -4, -4, 4, 3, -6, 1, 2, 0, 0,
    -- filter=217 channel=23
    -11, -23, -14, 8, 28, 18, 1, -14, -27,
    -- filter=217 channel=24
    3, 5, 4, -4, -3, 4, 1, -8, 5,
    -- filter=217 channel=25
    -20, -26, -4, 22, 39, 1, -7, -12, -12,
    -- filter=217 channel=26
    -13, -5, 3, 5, 6, -13, 0, 0, -6,
    -- filter=217 channel=27
    -40, -26, 8, 42, 45, 10, -9, -41, -10,
    -- filter=217 channel=28
    -5, -6, -4, 5, 6, 5, 1, -3, 4,
    -- filter=217 channel=29
    -8, -5, 6, 4, 12, 2, 2, -9, -4,
    -- filter=217 channel=30
    -23, -11, 6, 19, 21, 4, -9, -16, -1,
    -- filter=217 channel=31
    -17, -15, -1, 8, 32, 10, -9, -15, -10,
    -- filter=217 channel=32
    -21, -18, 2, 12, 39, 11, 0, -24, -6,
    -- filter=217 channel=33
    -6, -25, -17, -3, 28, 23, 15, -2, -20,
    -- filter=217 channel=34
    -2, -8, -15, 2, -14, -5, -4, -3, 1,
    -- filter=217 channel=35
    7, 2, 7, 0, -4, -7, 7, -2, -6,
    -- filter=217 channel=36
    0, 5, 0, 9, 9, -5, -16, -6, 5,
    -- filter=217 channel=37
    -17, -8, 8, 10, 18, -3, -6, -6, 4,
    -- filter=217 channel=38
    -11, -11, -2, -2, 17, 13, 6, -5, -5,
    -- filter=217 channel=39
    -7, -5, 4, 9, 12, 7, 5, -10, -6,
    -- filter=217 channel=40
    -2, -4, 2, 2, 0, -2, -1, 1, 1,
    -- filter=217 channel=41
    9, -11, -15, -34, -14, 4, -7, 3, -17,
    -- filter=217 channel=42
    -5, 2, 7, 4, 11, -2, 0, 0, -3,
    -- filter=217 channel=43
    3, -12, -7, -3, 12, 3, 13, -2, -15,
    -- filter=217 channel=44
    -7, -6, 12, 16, 12, 0, -4, -7, -5,
    -- filter=217 channel=45
    -6, -1, -5, -5, -2, 3, 0, -1, 6,
    -- filter=217 channel=46
    -2, -3, 0, 0, -1, -1, 7, -1, 2,
    -- filter=217 channel=47
    -11, -8, -5, -2, 18, 12, 6, -4, -7,
    -- filter=217 channel=48
    -32, -13, 10, 32, 39, 5, -9, -23, 1,
    -- filter=217 channel=49
    -15, -5, 4, 28, 18, -4, -5, -12, 7,
    -- filter=217 channel=50
    -10, -5, 10, 6, 13, 7, -7, -12, -13,
    -- filter=217 channel=51
    -1, -5, 4, 7, -7, -5, -1, -2, 1,
    -- filter=217 channel=52
    -7, 5, 1, 15, -1, -6, 1, 0, 2,
    -- filter=217 channel=53
    -7, -5, 1, 11, 12, 9, 0, 3, -1,
    -- filter=217 channel=54
    2, -5, 0, -1, 4, -3, -4, 5, -3,
    -- filter=217 channel=55
    -4, -15, 8, 0, 16, 16, 4, -15, -16,
    -- filter=217 channel=56
    -5, 13, -7, 1, 0, 3, -8, 0, 6,
    -- filter=217 channel=57
    -1, -4, 3, -7, 3, -7, 6, -5, -2,
    -- filter=217 channel=58
    5, 0, 0, 4, -10, 5, 2, 5, 2,
    -- filter=217 channel=59
    -17, -13, -2, 0, 20, 13, 6, -2, -4,
    -- filter=217 channel=60
    6, 7, -2, 0, -1, -5, -4, 3, 1,
    -- filter=217 channel=61
    -1, 0, 0, 6, 5, -6, -12, -2, -4,
    -- filter=217 channel=62
    8, -1, 0, -4, 0, 1, -3, 0, -3,
    -- filter=217 channel=63
    0, -4, -1, -11, -5, 0, -1, 2, -11,
    -- filter=217 channel=64
    7, 6, -5, -5, 0, 5, -3, -3, 7,
    -- filter=217 channel=65
    7, 0, 3, 7, 7, -5, -1, 3, 3,
    -- filter=217 channel=66
    10, -5, -9, -15, 0, 3, 8, -7, -1,
    -- filter=217 channel=67
    2, 2, 3, 8, -7, 3, 7, 1, -4,
    -- filter=217 channel=68
    -8, 2, -2, 5, 2, 0, -6, -6, 3,
    -- filter=217 channel=69
    4, -2, -4, 1, 0, 4, 0, 0, -3,
    -- filter=217 channel=70
    -2, -7, 6, 17, 14, 7, 4, -11, 0,
    -- filter=217 channel=71
    3, 7, -18, -8, 7, 4, 3, 10, 2,
    -- filter=217 channel=72
    -8, -17, 2, 10, 13, 3, 0, -16, -5,
    -- filter=217 channel=73
    -21, -12, 3, 13, 21, -2, 6, -17, 5,
    -- filter=217 channel=74
    -20, 0, 5, 17, 3, -13, -11, -13, -4,
    -- filter=217 channel=75
    0, -18, -22, -20, 18, 23, 2, 7, -14,
    -- filter=217 channel=76
    -1, -6, -7, -2, 16, 15, -1, -4, -6,
    -- filter=217 channel=77
    -1, -7, -7, 6, 5, 0, -4, -6, 2,
    -- filter=217 channel=78
    2, -13, -7, 5, 2, 5, 5, -1, -9,
    -- filter=217 channel=79
    -17, -28, -7, 5, 41, 22, 5, -24, -25,
    -- filter=217 channel=80
    -5, -19, 5, 4, 31, 9, 0, -19, -8,
    -- filter=217 channel=81
    -1, -2, 0, -3, -6, -7, 1, 4, 5,
    -- filter=217 channel=82
    8, 1, -10, -5, -2, 0, -3, -3, 3,
    -- filter=217 channel=83
    -4, 4, 7, 5, 2, 3, -8, -1, -6,
    -- filter=217 channel=84
    -23, 2, 1, 16, 12, 2, -12, -8, 8,
    -- filter=217 channel=85
    0, -5, 6, -7, -5, 1, 7, 4, 0,
    -- filter=217 channel=86
    -6, -6, 5, 4, -5, -10, -2, 0, 0,
    -- filter=217 channel=87
    0, 10, -1, 10, 6, 1, 4, 2, 0,
    -- filter=217 channel=88
    -3, 7, 9, 6, 1, -5, -9, -15, 2,
    -- filter=217 channel=89
    -8, -27, 4, 3, 40, 18, 2, -20, -19,
    -- filter=217 channel=90
    0, 10, 3, -3, -3, -2, 0, 3, -5,
    -- filter=217 channel=91
    -19, -1, 6, 35, 24, 2, -7, -25, -3,
    -- filter=217 channel=92
    6, 0, -6, 2, -7, 3, 5, 5, -3,
    -- filter=217 channel=93
    -23, -8, 5, 25, 21, -1, -5, -18, -9,
    -- filter=217 channel=94
    -4, 5, -3, 0, 4, 2, 4, -4, 0,
    -- filter=217 channel=95
    12, -4, -8, 8, 0, 4, 1, 5, -2,
    -- filter=217 channel=96
    0, -3, 0, 1, -3, -4, 2, 3, 4,
    -- filter=217 channel=97
    19, 0, -9, -1, -1, 4, 3, 19, 1,
    -- filter=217 channel=98
    -16, -25, -1, 19, 44, 14, 12, -26, -11,
    -- filter=217 channel=99
    -13, -5, 5, 10, 28, 3, -15, -26, -7,
    -- filter=217 channel=100
    -6, -5, 0, 1, -6, 6, 0, 2, -7,
    -- filter=217 channel=101
    -7, 12, 4, 31, 21, -1, -9, 13, 21,
    -- filter=217 channel=102
    0, -2, 6, -1, 1, 6, 3, 0, -4,
    -- filter=217 channel=103
    -2, -13, -12, -8, 16, 17, 10, 7, 4,
    -- filter=217 channel=104
    -6, -8, 10, 7, 14, 0, -7, -6, 2,
    -- filter=217 channel=105
    -5, -6, 0, -4, 6, 3, 4, -6, -6,
    -- filter=217 channel=106
    0, -4, 1, 4, -1, -1, 8, 3, -4,
    -- filter=217 channel=107
    -13, -9, -1, 10, 13, 7, -3, 0, -1,
    -- filter=217 channel=108
    7, 0, -3, -6, 0, 0, 2, 2, 0,
    -- filter=217 channel=109
    -28, -12, 4, 21, 34, 1, -2, -28, -11,
    -- filter=217 channel=110
    2, 0, -2, 0, 6, 3, 6, 1, -7,
    -- filter=217 channel=111
    -1, -6, -4, -9, -8, -6, 2, -6, -6,
    -- filter=217 channel=112
    -10, -1, -4, 17, 5, -8, -6, -8, 1,
    -- filter=217 channel=113
    0, -8, -13, -6, 13, 16, 11, -2, -12,
    -- filter=217 channel=114
    -38, -25, 9, 29, 37, 3, 0, -24, -8,
    -- filter=217 channel=115
    -4, 4, -2, -5, -1, 4, 0, -3, 0,
    -- filter=217 channel=116
    -28, -12, 12, 25, 35, 2, -6, -21, 0,
    -- filter=217 channel=117
    -9, -7, -5, 0, 14, 4, -6, 0, 4,
    -- filter=217 channel=118
    -6, -3, 0, -4, -8, 4, 2, -3, -5,
    -- filter=217 channel=119
    0, 12, -4, 9, -5, -2, -10, 1, 0,
    -- filter=217 channel=120
    -42, 0, 19, 42, 33, -11, -20, -37, -1,
    -- filter=217 channel=121
    12, -9, -9, 0, 2, 18, 14, -3, -10,
    -- filter=217 channel=122
    -5, 0, -7, 4, 23, 4, -13, 0, 0,
    -- filter=217 channel=123
    -3, 4, -10, 4, -6, -4, -3, 0, 0,
    -- filter=217 channel=124
    0, -2, -2, 7, 5, 3, 0, -1, 4,
    -- filter=217 channel=125
    -19, -17, 6, 14, 26, 6, -4, -22, -6,
    -- filter=217 channel=126
    12, -11, -8, -10, 10, 22, 15, 9, -13,
    -- filter=217 channel=127
    6, -1, 3, -3, 2, 3, 1, -7, -8,
    -- filter=218 channel=0
    2, 7, -1, 1, -2, 8, -5, -2, 7,
    -- filter=218 channel=1
    0, 8, 5, 1, 5, 7, 1, 2, 5,
    -- filter=218 channel=2
    6, -4, 6, 1, 3, -3, 3, -6, -7,
    -- filter=218 channel=3
    -5, 8, 1, -6, -5, 4, 6, -1, 4,
    -- filter=218 channel=4
    2, 0, 0, 2, 1, -5, 1, -2, 3,
    -- filter=218 channel=5
    6, 6, 4, -3, -3, 4, 0, -1, 0,
    -- filter=218 channel=6
    7, -2, 5, 1, 1, -4, 7, 1, -1,
    -- filter=218 channel=7
    1, -3, -2, 6, 5, 4, 5, 5, 2,
    -- filter=218 channel=8
    -1, -7, -4, 4, -6, 5, 6, -2, -6,
    -- filter=218 channel=9
    1, -6, -4, -5, 6, 1, -1, 5, 0,
    -- filter=218 channel=10
    -2, -5, 4, -5, 0, 1, 3, 6, -3,
    -- filter=218 channel=11
    0, 1, -4, 1, 4, 0, -6, 3, 4,
    -- filter=218 channel=12
    4, 2, 1, 0, 4, 4, -5, -7, -7,
    -- filter=218 channel=13
    -5, 1, -5, -6, 6, 0, 0, 6, -4,
    -- filter=218 channel=14
    0, 2, 2, -4, -3, 4, -3, -2, -6,
    -- filter=218 channel=15
    1, -7, 3, -2, -2, 6, 0, 4, 5,
    -- filter=218 channel=16
    -3, 3, -4, -4, 6, 1, -2, -6, -6,
    -- filter=218 channel=17
    -1, 7, -4, -2, 6, -2, 7, -2, -6,
    -- filter=218 channel=18
    1, 2, 0, -4, 3, 0, 2, -4, -2,
    -- filter=218 channel=19
    -4, 2, -5, -3, 1, 6, -7, 4, -4,
    -- filter=218 channel=20
    4, 2, -1, -5, -6, -3, -5, -4, -4,
    -- filter=218 channel=21
    -1, 1, 0, 0, -1, -7, -4, -6, 2,
    -- filter=218 channel=22
    3, -2, -4, 6, 3, -4, -1, -5, -1,
    -- filter=218 channel=23
    0, -6, 2, 0, -3, 0, 6, -2, 2,
    -- filter=218 channel=24
    2, -4, 0, 1, -7, 2, -4, -1, -4,
    -- filter=218 channel=25
    1, 3, -8, -6, 0, 1, -3, -4, -7,
    -- filter=218 channel=26
    -1, -1, 5, -4, 6, 2, -6, 4, 6,
    -- filter=218 channel=27
    -7, -10, 2, -7, -7, -8, -7, -6, -6,
    -- filter=218 channel=28
    -6, -5, 0, -4, 0, -3, 5, 4, 1,
    -- filter=218 channel=29
    -5, 6, 0, 2, -2, -1, -3, 0, 3,
    -- filter=218 channel=30
    0, -3, -7, 1, 1, -3, 1, -7, 3,
    -- filter=218 channel=31
    -3, -1, -1, -5, 2, -5, -1, 6, -7,
    -- filter=218 channel=32
    3, -3, 1, -8, 0, -7, -4, -5, -7,
    -- filter=218 channel=33
    6, 5, -6, -7, 0, -2, 2, -3, 1,
    -- filter=218 channel=34
    6, 4, 0, 4, -2, 0, 5, 6, 2,
    -- filter=218 channel=35
    -2, 0, -1, 2, 5, 0, -3, -3, -7,
    -- filter=218 channel=36
    2, 0, 1, 4, 2, 5, -6, -5, -1,
    -- filter=218 channel=37
    4, 1, -3, -4, -1, 0, 0, -4, -7,
    -- filter=218 channel=38
    2, -3, 0, -3, -5, 0, -1, 4, 2,
    -- filter=218 channel=39
    3, -1, -2, 6, -3, -5, 3, 5, 5,
    -- filter=218 channel=40
    -5, 7, -5, -6, 6, 2, -2, 4, 2,
    -- filter=218 channel=41
    8, 4, 1, 4, 3, -7, -4, 4, 0,
    -- filter=218 channel=42
    -3, -1, 4, -6, 4, 4, -2, -2, -3,
    -- filter=218 channel=43
    8, 3, 8, 3, -3, -1, -5, 1, 6,
    -- filter=218 channel=44
    -4, 3, -2, -5, 3, -6, 2, -2, 6,
    -- filter=218 channel=45
    3, -4, -5, 2, -5, 0, 5, -2, 0,
    -- filter=218 channel=46
    0, 5, -6, -3, 5, -2, 3, 3, 1,
    -- filter=218 channel=47
    4, -2, 3, 3, -3, 6, 4, 6, 2,
    -- filter=218 channel=48
    -3, -5, 1, 0, -7, 2, -5, 3, 2,
    -- filter=218 channel=49
    2, 6, 2, 0, -1, -5, 4, 1, -6,
    -- filter=218 channel=50
    0, 1, -3, -3, -6, 2, -3, -2, -3,
    -- filter=218 channel=51
    -5, 0, 0, 5, -5, -5, 0, -4, -5,
    -- filter=218 channel=52
    7, -1, -1, 4, 0, 4, -3, -4, 4,
    -- filter=218 channel=53
    1, -1, 0, 3, -7, -2, -1, -4, 3,
    -- filter=218 channel=54
    3, -2, 0, -4, 6, 0, 3, -1, 4,
    -- filter=218 channel=55
    6, 4, 0, -2, 0, -7, -1, 2, 0,
    -- filter=218 channel=56
    1, -6, -6, -6, -2, 4, 4, 5, 5,
    -- filter=218 channel=57
    4, -1, 3, -6, -6, 0, -6, 4, -7,
    -- filter=218 channel=58
    4, -2, -2, 0, -2, 3, -5, -3, 5,
    -- filter=218 channel=59
    -2, -6, -5, -6, -6, -1, 4, 1, 0,
    -- filter=218 channel=60
    0, 7, -5, -3, 5, 2, 0, 6, -4,
    -- filter=218 channel=61
    5, 7, 4, -1, -2, -1, 4, 2, 4,
    -- filter=218 channel=62
    7, -6, -3, -6, -6, 6, 3, 0, 2,
    -- filter=218 channel=63
    1, -5, 0, 5, 2, -4, 3, 7, 1,
    -- filter=218 channel=64
    -1, 3, 1, 6, 1, 1, 1, -4, 1,
    -- filter=218 channel=65
    1, 2, 1, -5, -2, 4, 3, -2, 4,
    -- filter=218 channel=66
    6, -2, -6, 4, 5, -3, 7, -3, 1,
    -- filter=218 channel=67
    0, -2, 4, 5, 4, 4, 4, 1, 0,
    -- filter=218 channel=68
    5, 1, -4, 5, 1, -3, 5, 4, -6,
    -- filter=218 channel=69
    -5, -6, 4, 0, -2, -1, -4, 4, 0,
    -- filter=218 channel=70
    2, -2, 1, -2, -3, -7, 0, 4, 6,
    -- filter=218 channel=71
    4, 0, 4, -2, -2, 1, -4, 7, -4,
    -- filter=218 channel=72
    0, 5, -6, 2, -5, -3, 1, 3, 4,
    -- filter=218 channel=73
    6, 2, 3, -4, -2, 1, -6, -1, 0,
    -- filter=218 channel=74
    0, 2, -1, 2, 5, 1, 2, -5, -1,
    -- filter=218 channel=75
    7, 8, -5, 0, 1, 5, 4, -3, 4,
    -- filter=218 channel=76
    -1, -5, -4, 4, -4, -7, 1, 6, 1,
    -- filter=218 channel=77
    5, 0, 0, -6, -3, 5, 0, 2, 0,
    -- filter=218 channel=78
    7, 4, -5, -5, 5, -6, -7, -5, -4,
    -- filter=218 channel=79
    -6, 0, -1, -5, -6, -8, 1, 0, 0,
    -- filter=218 channel=80
    -6, -8, -5, -5, 3, 0, -7, 0, -3,
    -- filter=218 channel=81
    3, -3, 0, -5, -1, -2, 5, -2, 0,
    -- filter=218 channel=82
    -5, -3, -2, 2, 0, 3, 2, 7, 5,
    -- filter=218 channel=83
    4, 2, 0, 0, -2, -6, 0, -7, -3,
    -- filter=218 channel=84
    -7, 1, -4, 7, -1, -5, 1, -3, -5,
    -- filter=218 channel=85
    -3, 1, 0, -4, 6, 3, -1, 5, 6,
    -- filter=218 channel=86
    -5, 0, -6, 2, 4, -5, 7, -5, 3,
    -- filter=218 channel=87
    6, 4, 7, -1, 0, 1, -2, -6, -6,
    -- filter=218 channel=88
    -5, -3, 2, 1, 6, 7, 7, 0, 2,
    -- filter=218 channel=89
    0, -4, 0, 1, -5, -5, -8, 3, -5,
    -- filter=218 channel=90
    -5, -2, -5, 2, -5, 1, -2, 0, 1,
    -- filter=218 channel=91
    6, -8, 3, 0, -7, 3, 1, -8, -8,
    -- filter=218 channel=92
    7, -6, 0, 1, -5, 0, 0, -2, -5,
    -- filter=218 channel=93
    -1, -6, -1, -3, -1, 5, 4, -6, -6,
    -- filter=218 channel=94
    2, 5, 1, -2, -5, 1, 0, -3, 3,
    -- filter=218 channel=95
    -1, -4, -3, -5, -5, 0, 0, 0, 2,
    -- filter=218 channel=96
    2, -3, -1, 3, 2, -3, -7, 1, 1,
    -- filter=218 channel=97
    -2, 4, 4, -6, 4, 1, -6, 2, 1,
    -- filter=218 channel=98
    2, -5, 4, 1, -3, -4, -1, -1, 0,
    -- filter=218 channel=99
    -5, -6, 1, 5, 3, 2, 5, -6, 0,
    -- filter=218 channel=100
    4, 3, -4, -2, -4, -7, 2, 0, 5,
    -- filter=218 channel=101
    1, 1, 1, 0, -1, -5, 0, 6, -7,
    -- filter=218 channel=102
    0, 1, -4, 5, -1, -2, 4, 6, -4,
    -- filter=218 channel=103
    6, -4, 3, -3, 3, -4, -6, -2, 0,
    -- filter=218 channel=104
    4, -3, 1, -4, 1, -4, 5, -4, 3,
    -- filter=218 channel=105
    4, 3, 5, -2, -6, -3, -6, 4, 5,
    -- filter=218 channel=106
    3, 4, -3, -4, 7, 0, -6, 0, -4,
    -- filter=218 channel=107
    -3, 5, -3, 3, 0, -6, -3, -5, 3,
    -- filter=218 channel=108
    0, 2, -4, -3, 2, -1, 0, 5, 2,
    -- filter=218 channel=109
    -1, -4, 0, 0, -3, -6, -4, 1, -1,
    -- filter=218 channel=110
    4, 1, -7, 0, 0, -1, 0, 2, 5,
    -- filter=218 channel=111
    7, 1, -5, 1, 5, -7, 0, 1, 5,
    -- filter=218 channel=112
    6, -7, -6, -2, 0, 4, -2, -5, 2,
    -- filter=218 channel=113
    0, 0, -4, -1, 0, -4, 3, 1, 4,
    -- filter=218 channel=114
    0, 0, -1, 6, 0, 4, -7, 3, 6,
    -- filter=218 channel=115
    -5, 0, -1, 1, -3, -6, 4, 2, 5,
    -- filter=218 channel=116
    -6, 7, -6, 0, -2, -6, -1, 2, 1,
    -- filter=218 channel=117
    2, -3, -2, -5, 7, 2, 2, -2, 0,
    -- filter=218 channel=118
    6, 4, -6, -1, 2, 4, 1, 5, 0,
    -- filter=218 channel=119
    0, -6, -2, 6, -7, -6, -7, 4, 0,
    -- filter=218 channel=120
    1, 1, 5, -2, -2, 5, 0, 1, 4,
    -- filter=218 channel=121
    4, 2, -4, 0, -5, -8, -5, 0, 0,
    -- filter=218 channel=122
    8, -4, -6, 4, -4, 0, -4, 3, 0,
    -- filter=218 channel=123
    -5, 1, 4, -1, 4, 3, 4, -6, 0,
    -- filter=218 channel=124
    -1, 2, 4, 4, 6, 0, -4, 2, 4,
    -- filter=218 channel=125
    4, -3, 3, -2, 4, -7, 2, -5, 1,
    -- filter=218 channel=126
    0, -5, 1, -6, 3, 0, 0, 4, -6,
    -- filter=218 channel=127
    6, 1, 3, 5, -3, 7, -1, 2, -5,
    -- filter=219 channel=0
    3, 5, -4, -8, 3, 8, -3, 9, 5,
    -- filter=219 channel=1
    -6, -9, -9, 2, 0, -10, -4, 1, 0,
    -- filter=219 channel=2
    -5, -3, 7, -6, -5, -4, -4, -3, 6,
    -- filter=219 channel=3
    8, 28, 21, -11, 1, 10, -7, 0, 0,
    -- filter=219 channel=4
    6, 9, 12, -7, -4, 6, -7, -8, 6,
    -- filter=219 channel=5
    -4, 6, 3, -7, 10, 5, -9, 6, 0,
    -- filter=219 channel=6
    -2, 5, -2, 5, 2, 5, 8, -5, 8,
    -- filter=219 channel=7
    2, 5, -2, 6, 6, -6, 0, 7, -3,
    -- filter=219 channel=8
    7, -2, -5, -2, -3, 6, -6, -6, -2,
    -- filter=219 channel=9
    -3, -4, 5, -3, -7, 3, 6, -4, 0,
    -- filter=219 channel=10
    1, 11, 12, 0, 0, -3, 4, 0, -5,
    -- filter=219 channel=11
    3, 0, 12, -4, -5, -11, 0, -2, 3,
    -- filter=219 channel=12
    -2, 5, 0, 2, -8, 0, 0, 0, -1,
    -- filter=219 channel=13
    0, 10, 16, -2, -15, -17, -3, -11, -14,
    -- filter=219 channel=14
    0, -5, 6, -1, 3, -4, -3, 2, -5,
    -- filter=219 channel=15
    8, 13, 11, -3, -16, -10, 4, -14, -18,
    -- filter=219 channel=16
    -6, 0, -2, -4, 6, 6, 4, 2, -2,
    -- filter=219 channel=17
    0, -3, -6, -2, 2, 6, 2, 3, -6,
    -- filter=219 channel=18
    -1, 13, 20, 4, -15, -11, 4, -7, -12,
    -- filter=219 channel=19
    -2, 4, 1, -2, 6, 4, -6, 1, 5,
    -- filter=219 channel=20
    3, 16, 21, -11, -14, -1, 0, 0, -3,
    -- filter=219 channel=21
    -3, -11, -11, -1, 3, 7, 3, -2, 9,
    -- filter=219 channel=22
    5, 4, 7, 4, -1, -8, 7, 0, -6,
    -- filter=219 channel=23
    13, 21, 19, -12, -29, -5, 4, -22, -2,
    -- filter=219 channel=24
    -2, 2, -4, 2, 2, -6, 2, 1, -1,
    -- filter=219 channel=25
    0, 3, 10, 5, -5, -8, 7, 4, -10,
    -- filter=219 channel=26
    2, 1, -9, 0, 9, -1, -7, 4, 3,
    -- filter=219 channel=27
    0, 13, 7, -5, -23, -12, 3, -6, -11,
    -- filter=219 channel=28
    -7, 7, 0, -4, 0, -6, -6, -7, 3,
    -- filter=219 channel=29
    3, 13, 10, -3, -4, -10, 8, 1, -5,
    -- filter=219 channel=30
    -10, -2, 7, 5, -10, -8, -8, -4, -3,
    -- filter=219 channel=31
    1, 9, 8, 4, -1, 11, -2, 0, -5,
    -- filter=219 channel=32
    -1, 9, 22, 2, -13, -15, 7, -5, -8,
    -- filter=219 channel=33
    5, 6, 17, -2, -11, -6, -4, -13, -4,
    -- filter=219 channel=34
    0, 9, 9, 6, 0, 8, 4, 1, 6,
    -- filter=219 channel=35
    -7, -2, 0, 3, -1, -2, 1, 6, -6,
    -- filter=219 channel=36
    -6, -4, -2, 4, -4, -1, -6, -5, 10,
    -- filter=219 channel=37
    -13, -1, -3, -1, -3, 7, -8, 4, 0,
    -- filter=219 channel=38
    -4, 13, 7, -4, -6, -4, 0, 0, -1,
    -- filter=219 channel=39
    -2, 3, 2, -1, 0, -6, 3, -2, 0,
    -- filter=219 channel=40
    -4, 7, 2, -4, -3, 0, 1, -3, -6,
    -- filter=219 channel=41
    6, 5, 7, 6, 6, -17, 5, 8, -12,
    -- filter=219 channel=42
    4, 0, -5, -5, 1, 2, 0, -1, 7,
    -- filter=219 channel=43
    9, 14, 17, 0, 0, -1, 1, -4, -9,
    -- filter=219 channel=44
    -7, 2, 0, 5, 0, 6, -5, -2, 0,
    -- filter=219 channel=45
    -4, 5, 5, -6, -5, 7, -5, 8, 2,
    -- filter=219 channel=46
    -5, 7, -5, 3, -1, 1, 5, 6, -8,
    -- filter=219 channel=47
    -7, -9, -8, 3, 10, 7, -6, 2, 5,
    -- filter=219 channel=48
    0, 0, -7, 1, -1, -13, 0, 1, 0,
    -- filter=219 channel=49
    -5, -1, 3, -5, -8, -14, -5, -8, -1,
    -- filter=219 channel=50
    -1, -2, 8, -1, -2, -10, 5, 1, 0,
    -- filter=219 channel=51
    -4, 5, -6, 0, -1, 0, 0, -6, -6,
    -- filter=219 channel=52
    5, 9, 10, -9, -5, -4, -5, -4, -3,
    -- filter=219 channel=53
    6, 9, 5, -8, 0, 3, -1, -5, -6,
    -- filter=219 channel=54
    6, -6, -4, -3, -4, -3, 0, -5, -6,
    -- filter=219 channel=55
    2, 13, 23, -9, -19, -19, 6, -18, -3,
    -- filter=219 channel=56
    6, 8, 4, -7, -5, 0, 3, 0, 1,
    -- filter=219 channel=57
    -1, -4, -1, 3, 1, 3, 6, -1, 1,
    -- filter=219 channel=58
    0, 1, 1, -1, 3, 3, -5, 12, 0,
    -- filter=219 channel=59
    -5, -1, 2, 0, 2, -11, 0, -5, -9,
    -- filter=219 channel=60
    -3, 1, -3, -2, 1, -3, 5, -6, 0,
    -- filter=219 channel=61
    0, -5, -6, -3, -9, -1, -4, -6, -5,
    -- filter=219 channel=62
    7, -2, 5, 0, 7, 7, 4, -8, -6,
    -- filter=219 channel=63
    -7, -8, -2, 8, 13, 10, 1, 9, 2,
    -- filter=219 channel=64
    -1, -2, 7, -4, 0, -6, 2, 5, 6,
    -- filter=219 channel=65
    4, -2, 4, -3, 1, -6, -6, 2, 0,
    -- filter=219 channel=66
    7, 0, 2, 3, -6, 0, 4, -1, -1,
    -- filter=219 channel=67
    0, -4, -3, 3, 4, 5, 5, -2, -6,
    -- filter=219 channel=68
    -5, 2, 1, 6, -8, 2, 2, -8, 7,
    -- filter=219 channel=69
    6, -4, 1, 4, 6, -1, 9, -3, 4,
    -- filter=219 channel=70
    -1, 14, 11, -11, -13, -6, -3, -13, -17,
    -- filter=219 channel=71
    11, 11, 7, -2, -2, 0, 0, 3, -4,
    -- filter=219 channel=72
    -2, 6, 0, -5, -9, -6, 6, -10, -1,
    -- filter=219 channel=73
    1, 2, 7, 3, -17, -10, -5, 0, -7,
    -- filter=219 channel=74
    -2, 0, -1, 2, -11, 2, -2, -9, 3,
    -- filter=219 channel=75
    4, 7, 0, 4, 16, -3, -7, 6, -10,
    -- filter=219 channel=76
    1, 5, 18, 3, -14, -5, 11, -9, -6,
    -- filter=219 channel=77
    -2, -6, 2, -2, 7, 2, 5, 1, 3,
    -- filter=219 channel=78
    5, -3, -5, -3, 11, 0, 3, 2, -1,
    -- filter=219 channel=79
    2, 19, 27, 2, -29, -24, 15, -8, -12,
    -- filter=219 channel=80
    -4, -9, -1, 11, 0, -4, 1, 7, -5,
    -- filter=219 channel=81
    -3, 7, -7, 1, 0, -1, 4, -1, 3,
    -- filter=219 channel=82
    -1, 5, 7, -8, 3, -3, 0, 1, 0,
    -- filter=219 channel=83
    0, 1, 5, -1, -8, 2, 1, 7, -2,
    -- filter=219 channel=84
    2, 5, 10, -3, -12, -12, 1, 2, 3,
    -- filter=219 channel=85
    0, -6, 1, -1, -6, 1, 4, 5, 7,
    -- filter=219 channel=86
    -8, -4, 5, -7, 1, 4, -1, -5, 1,
    -- filter=219 channel=87
    -2, 11, 3, -1, -9, 3, 7, 1, 6,
    -- filter=219 channel=88
    4, -3, -10, 6, 4, 1, -2, -4, 0,
    -- filter=219 channel=89
    -2, 4, 21, 0, -5, -11, 1, -7, -13,
    -- filter=219 channel=90
    8, 8, -1, 3, 0, 12, -11, -3, 0,
    -- filter=219 channel=91
    0, 2, 5, -8, -25, -10, -8, -6, -11,
    -- filter=219 channel=92
    6, 1, 3, -9, 5, 0, 0, 2, 1,
    -- filter=219 channel=93
    -3, -13, -13, 5, -2, 8, -1, 11, 7,
    -- filter=219 channel=94
    5, 5, -3, -6, 0, -4, -3, -2, -5,
    -- filter=219 channel=95
    3, -2, 6, 0, 5, 0, 0, 1, -2,
    -- filter=219 channel=96
    0, 0, 0, 4, -5, 0, -1, -4, 0,
    -- filter=219 channel=97
    5, 6, 5, 1, 4, 5, 4, -4, -7,
    -- filter=219 channel=98
    -3, 4, 9, -1, -4, -10, 6, 3, 2,
    -- filter=219 channel=99
    8, 14, 2, -2, -10, 4, 4, -7, -4,
    -- filter=219 channel=100
    8, -3, -4, 0, 6, 0, -1, 1, 3,
    -- filter=219 channel=101
    6, 6, 10, -3, -2, 5, 2, -7, -4,
    -- filter=219 channel=102
    2, 1, 0, -6, 4, 0, -4, 6, 4,
    -- filter=219 channel=103
    3, 4, 0, 9, 8, 6, -7, 3, 2,
    -- filter=219 channel=104
    2, -5, 0, 4, -4, 1, -3, 5, 4,
    -- filter=219 channel=105
    0, 14, 11, 2, -9, 6, 8, -5, -5,
    -- filter=219 channel=106
    -2, 0, 2, 4, -8, 4, 1, 2, 4,
    -- filter=219 channel=107
    6, 6, 8, -5, -4, -3, -6, -8, 3,
    -- filter=219 channel=108
    1, 7, -3, 11, 10, 2, 6, 10, -1,
    -- filter=219 channel=109
    0, 2, 9, -2, -12, -21, 4, -10, -7,
    -- filter=219 channel=110
    -1, 12, 4, 4, -8, 13, -7, -8, 6,
    -- filter=219 channel=111
    -3, 1, 6, 2, -4, 2, 0, 9, 4,
    -- filter=219 channel=112
    4, 3, 9, -4, -10, -6, -6, -2, -3,
    -- filter=219 channel=113
    5, 12, 0, -7, 1, 7, -1, -3, -7,
    -- filter=219 channel=114
    -4, 9, 13, 7, -6, -21, 10, -1, -9,
    -- filter=219 channel=115
    4, 0, 6, -6, -5, 3, -4, -5, 5,
    -- filter=219 channel=116
    -4, 6, 11, 2, -12, -19, 3, -6, -6,
    -- filter=219 channel=117
    5, -3, -2, -6, -9, -9, -2, -3, 3,
    -- filter=219 channel=118
    0, 3, -4, 7, -5, -6, -2, 4, 7,
    -- filter=219 channel=119
    10, 1, 5, 0, 5, -1, -9, 6, 1,
    -- filter=219 channel=120
    11, 10, 18, 0, -24, -14, -1, -9, 1,
    -- filter=219 channel=121
    0, -1, -2, -5, 3, 2, -4, 4, 2,
    -- filter=219 channel=122
    -9, -18, -10, 12, 7, 14, -2, 9, 0,
    -- filter=219 channel=123
    5, 2, -3, 6, -1, -3, -2, 5, 2,
    -- filter=219 channel=124
    -2, -2, 9, 3, 0, 3, 9, -5, 1,
    -- filter=219 channel=125
    -3, 7, 8, 1, -1, -11, -5, 2, -7,
    -- filter=219 channel=126
    8, 13, 11, -3, 9, -5, 7, -7, 0,
    -- filter=219 channel=127
    -5, 0, -5, -4, 6, -3, 9, -1, -4,
    -- filter=220 channel=0
    5, 0, -6, 9, 2, -3, -2, 2, -7,
    -- filter=220 channel=1
    5, -3, -6, 14, -1, 0, 10, 1, -7,
    -- filter=220 channel=2
    4, -8, -5, -8, 1, 4, -4, -1, -2,
    -- filter=220 channel=3
    13, 0, 3, -12, -2, 9, -6, -2, 3,
    -- filter=220 channel=4
    -7, -9, -1, -10, -5, 4, -2, -10, -6,
    -- filter=220 channel=5
    9, -5, -18, 13, 4, -15, 12, 6, -8,
    -- filter=220 channel=6
    -1, 9, 0, -12, -9, -6, 2, -3, -7,
    -- filter=220 channel=7
    1, 4, 5, -2, 2, 6, 1, -4, 0,
    -- filter=220 channel=8
    -3, 3, -4, -3, -7, -5, 2, -2, -6,
    -- filter=220 channel=9
    6, 5, -4, 0, -4, 1, 0, -5, 2,
    -- filter=220 channel=10
    1, 7, 4, -5, -5, -4, 5, -4, 8,
    -- filter=220 channel=11
    0, 13, 5, -2, -11, -4, -5, -2, 0,
    -- filter=220 channel=12
    -5, -6, -6, -7, -2, 0, 2, -7, 5,
    -- filter=220 channel=13
    4, 9, 9, -12, -9, 6, -10, -13, -4,
    -- filter=220 channel=14
    -2, -5, -2, -5, 2, 1, -1, 1, 4,
    -- filter=220 channel=15
    17, 13, 15, -18, -9, 4, -4, -15, 0,
    -- filter=220 channel=16
    -7, -10, -17, 4, 8, -6, 8, 12, 0,
    -- filter=220 channel=17
    2, -3, -5, 0, 6, 0, -4, -3, 0,
    -- filter=220 channel=18
    10, 10, 18, -6, -16, 4, -7, -8, 2,
    -- filter=220 channel=19
    3, 0, -7, -5, -2, -6, -6, -4, 2,
    -- filter=220 channel=20
    0, 8, 10, -14, -7, -1, -2, -2, 2,
    -- filter=220 channel=21
    5, 0, -15, 8, 14, -5, 11, 5, -3,
    -- filter=220 channel=22
    0, 6, 2, -1, 3, -1, 1, 3, -9,
    -- filter=220 channel=23
    16, 22, 16, -14, -8, 0, -9, -17, -7,
    -- filter=220 channel=24
    -5, 3, -1, 0, 7, -1, -1, 0, -4,
    -- filter=220 channel=25
    9, 3, -3, -6, -5, 2, 11, 0, -6,
    -- filter=220 channel=26
    2, -8, -8, 0, 1, -14, 0, 0, -9,
    -- filter=220 channel=27
    15, 14, 0, -1, 0, -4, 4, 0, -8,
    -- filter=220 channel=28
    -5, -6, 7, -2, 1, 0, 1, -4, 5,
    -- filter=220 channel=29
    4, 10, 10, -6, -13, 1, -8, -5, 3,
    -- filter=220 channel=30
    -1, -2, -5, 0, -4, -11, 10, 7, -4,
    -- filter=220 channel=31
    13, 14, -3, 2, 6, -1, 10, 9, -2,
    -- filter=220 channel=32
    10, 14, 17, -13, -4, -4, 0, -14, -9,
    -- filter=220 channel=33
    6, 8, 0, -6, 5, -3, -4, -2, 0,
    -- filter=220 channel=34
    4, 5, -2, -4, -4, 0, -10, 3, -10,
    -- filter=220 channel=35
    5, -4, 6, 3, -5, 5, -2, -6, 7,
    -- filter=220 channel=36
    -13, -1, -5, -11, -9, 0, 1, -5, 4,
    -- filter=220 channel=37
    -5, -12, -10, 11, 0, -8, 3, 5, -6,
    -- filter=220 channel=38
    14, 8, -3, 3, 8, -3, 5, 4, -4,
    -- filter=220 channel=39
    -3, 4, 5, -9, -4, -1, 1, -4, 5,
    -- filter=220 channel=40
    0, 2, 0, -10, -5, 7, -3, -4, -2,
    -- filter=220 channel=41
    -1, 0, 6, 4, -16, 1, -1, -9, 8,
    -- filter=220 channel=42
    2, -1, -10, 0, 8, -6, 10, 8, 0,
    -- filter=220 channel=43
    5, 5, 9, -4, -14, -4, -6, -3, -2,
    -- filter=220 channel=44
    3, -8, -5, 6, 0, 0, 7, 6, -10,
    -- filter=220 channel=45
    0, 0, 5, 2, 1, 3, 3, 2, -4,
    -- filter=220 channel=46
    6, 4, -4, 6, -7, -5, -3, -3, 6,
    -- filter=220 channel=47
    3, -6, -22, 11, 16, -6, 14, 8, -5,
    -- filter=220 channel=48
    2, -3, -9, -3, -1, -9, 0, 4, 0,
    -- filter=220 channel=49
    6, -2, 1, -5, -12, 8, -7, -12, -5,
    -- filter=220 channel=50
    9, 8, 6, 0, 6, -3, 4, -3, -2,
    -- filter=220 channel=51
    0, -7, 5, -1, 0, -1, 0, 5, 5,
    -- filter=220 channel=52
    8, 5, 8, -1, -7, -6, -1, -10, -6,
    -- filter=220 channel=53
    -2, 0, 2, 0, -8, -2, -8, -9, -6,
    -- filter=220 channel=54
    -2, 4, 2, 2, 0, -5, -3, 3, -1,
    -- filter=220 channel=55
    11, 20, 14, -10, -6, -1, -9, -17, -7,
    -- filter=220 channel=56
    -2, 2, -7, -10, -10, 0, -4, -5, 3,
    -- filter=220 channel=57
    -8, -6, -4, -1, 3, 1, 0, 0, -5,
    -- filter=220 channel=58
    -3, -2, -12, 0, -2, -12, 6, 10, -1,
    -- filter=220 channel=59
    12, 0, -2, 0, 1, 0, 1, 4, 0,
    -- filter=220 channel=60
    1, -5, 2, -5, -6, -7, -4, -2, -4,
    -- filter=220 channel=61
    4, 0, -4, -3, 0, -5, -5, 1, 1,
    -- filter=220 channel=62
    -5, -2, 0, -2, -6, -1, 5, 6, 4,
    -- filter=220 channel=63
    0, -7, -8, 5, 8, -7, 8, 3, 2,
    -- filter=220 channel=64
    -2, -2, 6, -9, 0, 0, 1, -1, 4,
    -- filter=220 channel=65
    0, -1, 6, 2, -5, 3, -5, 0, -1,
    -- filter=220 channel=66
    -4, -2, -5, -3, -12, -7, -8, 0, -3,
    -- filter=220 channel=67
    -4, 1, -1, 1, 0, -5, -2, -8, -4,
    -- filter=220 channel=68
    0, 5, 3, -4, 0, -3, 0, 3, 4,
    -- filter=220 channel=69
    4, 2, -2, 0, 0, -5, -6, 2, 3,
    -- filter=220 channel=70
    16, 5, 5, -10, -3, 7, -2, -11, 1,
    -- filter=220 channel=71
    0, 3, 3, 0, -1, -5, -1, -2, 8,
    -- filter=220 channel=72
    0, 11, -4, 1, -2, 0, 8, 6, 3,
    -- filter=220 channel=73
    -1, 0, 3, -13, -14, 3, 0, -3, 2,
    -- filter=220 channel=74
    -2, 1, -3, -9, -7, -2, -7, 2, -5,
    -- filter=220 channel=75
    13, 8, -2, 10, 0, 3, 3, -1, -1,
    -- filter=220 channel=76
    9, 15, 17, -8, -15, -3, -7, -7, -5,
    -- filter=220 channel=77
    0, 3, 0, -3, -7, 2, 5, 6, -1,
    -- filter=220 channel=78
    7, 1, -5, 10, 7, -8, 4, -3, 5,
    -- filter=220 channel=79
    10, 15, 19, -8, -19, 5, -4, -7, -6,
    -- filter=220 channel=80
    5, 12, -3, 10, 1, 0, 8, 12, 3,
    -- filter=220 channel=81
    0, 7, 0, -2, 6, 7, -4, 5, 2,
    -- filter=220 channel=82
    -3, -3, 1, 5, -3, 5, -3, -1, 6,
    -- filter=220 channel=83
    -1, -3, -8, 6, -2, -4, -3, 3, -3,
    -- filter=220 channel=84
    -1, 9, 4, -14, -10, -8, 2, -1, 0,
    -- filter=220 channel=85
    3, 6, -2, 0, -6, -6, -1, 6, 0,
    -- filter=220 channel=86
    4, -3, -5, 1, 0, -1, -1, -3, -5,
    -- filter=220 channel=87
    -6, -2, 11, -6, -4, -9, -8, -13, 1,
    -- filter=220 channel=88
    -10, -8, -11, -10, -6, 0, 1, 3, -6,
    -- filter=220 channel=89
    20, 9, 7, -12, -9, 6, -10, 1, 0,
    -- filter=220 channel=90
    -7, -4, -9, 1, 5, 2, -9, 3, 5,
    -- filter=220 channel=91
    -6, 14, 12, -12, -7, 1, -5, -10, 2,
    -- filter=220 channel=92
    3, 0, -3, 4, -4, 2, 0, 2, -1,
    -- filter=220 channel=93
    -11, -7, -23, 4, 1, -5, 9, 12, -9,
    -- filter=220 channel=94
    5, 2, -3, 6, 2, -2, 7, 2, -1,
    -- filter=220 channel=95
    -1, -5, 1, -7, -8, 4, -9, 3, -5,
    -- filter=220 channel=96
    3, 0, -2, 0, 3, 0, -3, -2, 2,
    -- filter=220 channel=97
    11, 0, -2, 7, 2, 4, 0, 4, -3,
    -- filter=220 channel=98
    18, 9, 6, 3, -3, -5, 0, 3, -3,
    -- filter=220 channel=99
    10, 8, 12, -5, -7, -7, -7, -7, -2,
    -- filter=220 channel=100
    -6, 5, -1, -6, -6, 3, -7, -6, -1,
    -- filter=220 channel=101
    -7, -9, -6, -13, -3, -4, -14, -5, 2,
    -- filter=220 channel=102
    -6, -3, -3, 2, -2, -6, -7, 2, -4,
    -- filter=220 channel=103
    11, -8, -14, 20, 21, -10, 1, 16, -2,
    -- filter=220 channel=104
    0, 5, 0, 11, 0, -6, 12, 3, 1,
    -- filter=220 channel=105
    8, -1, 0, -12, -4, -8, -10, -10, -5,
    -- filter=220 channel=106
    0, 6, 6, -6, 0, 3, -7, -6, 3,
    -- filter=220 channel=107
    5, 10, 5, -14, -15, 3, -9, -7, -4,
    -- filter=220 channel=108
    3, 5, 3, 3, -4, -5, -3, -3, 5,
    -- filter=220 channel=109
    12, 13, 1, -8, -13, -1, -2, 0, -12,
    -- filter=220 channel=110
    9, 13, 7, -2, -4, 3, 0, 2, 1,
    -- filter=220 channel=111
    -1, 3, 0, 6, -8, 5, -2, 0, -3,
    -- filter=220 channel=112
    12, 6, 1, 0, 0, -6, 1, 0, 3,
    -- filter=220 channel=113
    4, 12, 2, 1, -3, 0, 4, 2, -2,
    -- filter=220 channel=114
    12, 7, 6, -12, -7, -9, 5, -7, -6,
    -- filter=220 channel=115
    -2, 0, -3, -2, -1, -6, -7, 5, 2,
    -- filter=220 channel=116
    1, 8, 4, -3, -5, -2, 9, 1, -10,
    -- filter=220 channel=117
    0, -5, 0, 0, 1, 3, 2, -3, -1,
    -- filter=220 channel=118
    1, 0, 2, -2, 2, 1, 1, 0, 4,
    -- filter=220 channel=119
    -6, -8, 0, -8, -14, -7, -5, -10, -5,
    -- filter=220 channel=120
    5, 4, 5, -14, -18, -1, -4, 0, -18,
    -- filter=220 channel=121
    0, -3, -3, 0, -5, -1, 0, -8, -2,
    -- filter=220 channel=122
    -2, -13, -24, 16, 19, -19, 14, 20, -6,
    -- filter=220 channel=123
    -2, -4, -2, 1, -2, -7, -3, -4, -3,
    -- filter=220 channel=124
    -4, 3, 1, -2, -2, 1, 2, -10, -4,
    -- filter=220 channel=125
    5, 8, -4, -1, -7, -1, -1, 5, 4,
    -- filter=220 channel=126
    4, 3, 2, 3, 0, 3, 2, -5, 5,
    -- filter=220 channel=127
    3, 0, 6, -6, -3, 0, -5, -7, -2,
    -- filter=221 channel=0
    -8, 9, -8, -6, 19, -14, 2, 15, -5,
    -- filter=221 channel=1
    2, 11, -12, -7, 12, 0, -10, 8, -12,
    -- filter=221 channel=2
    4, 6, -2, -1, -6, -6, -2, -5, 1,
    -- filter=221 channel=3
    -3, -4, 0, 0, -12, -14, -17, -3, -20,
    -- filter=221 channel=4
    6, -6, -4, -11, -5, -10, -8, -9, -4,
    -- filter=221 channel=5
    -2, 0, -7, 4, 0, 0, -5, -5, -5,
    -- filter=221 channel=6
    1, -4, -2, -8, 7, 6, 0, -1, 0,
    -- filter=221 channel=7
    -1, 0, 0, -2, 1, 2, 3, 1, 4,
    -- filter=221 channel=8
    -6, 8, 2, 3, 2, 13, 5, -2, -1,
    -- filter=221 channel=9
    -4, 1, 3, -3, 6, 0, 0, -7, -5,
    -- filter=221 channel=10
    -3, -5, 5, -1, 10, -8, -1, 4, 0,
    -- filter=221 channel=11
    -1, -5, -10, 0, -6, -3, -2, -8, 0,
    -- filter=221 channel=12
    0, 16, 0, -2, 12, 8, -1, 14, 4,
    -- filter=221 channel=13
    -7, 10, -7, -10, 18, -14, 0, 11, -7,
    -- filter=221 channel=14
    5, 6, 6, -7, -3, 2, 6, -1, -6,
    -- filter=221 channel=15
    -2, -2, 0, -2, 2, -16, -7, 3, -11,
    -- filter=221 channel=16
    -1, 9, 5, 4, -1, -5, 0, -3, -13,
    -- filter=221 channel=17
    -5, 5, 2, -1, -4, 1, 3, -5, -3,
    -- filter=221 channel=18
    -10, 7, -14, -6, 20, -6, 0, 8, -13,
    -- filter=221 channel=19
    7, 1, -1, -4, 1, -5, -3, 4, -5,
    -- filter=221 channel=20
    -7, -1, -3, -8, -2, -4, -6, 3, -8,
    -- filter=221 channel=21
    -7, 0, -4, 6, -2, -13, -3, -4, -2,
    -- filter=221 channel=22
    6, 3, 0, -1, 1, -8, 4, -3, 8,
    -- filter=221 channel=23
    -1, 2, -4, 5, 12, -10, 1, -4, 0,
    -- filter=221 channel=24
    6, 0, 3, 0, 7, -4, 2, -5, -3,
    -- filter=221 channel=25
    -6, 14, -12, -1, 14, -6, 1, 15, -8,
    -- filter=221 channel=26
    0, 6, -1, 6, 0, 2, 2, -3, -7,
    -- filter=221 channel=27
    4, 20, -14, 0, 19, -17, 9, 2, -7,
    -- filter=221 channel=28
    6, 0, 6, -6, -6, 1, 3, 7, -1,
    -- filter=221 channel=29
    -8, 5, -15, -8, -4, -10, -6, 0, -2,
    -- filter=221 channel=30
    3, 8, -6, -6, 8, -12, 4, -1, -13,
    -- filter=221 channel=31
    -6, 8, 0, 8, 1, -9, 8, -6, -9,
    -- filter=221 channel=32
    -12, 13, -17, -8, 19, -8, -11, 13, -17,
    -- filter=221 channel=33
    -3, 14, -5, -6, 11, -12, -3, 7, -15,
    -- filter=221 channel=34
    6, 0, 13, 7, 20, 24, -2, 9, 24,
    -- filter=221 channel=35
    6, 0, -5, 0, -6, -6, -5, -2, 3,
    -- filter=221 channel=36
    1, -4, -10, 3, 6, -11, 6, -2, -7,
    -- filter=221 channel=37
    -2, 14, 1, 2, 12, -8, -4, 6, -2,
    -- filter=221 channel=38
    -6, 3, 3, 0, 2, -9, -1, 2, -11,
    -- filter=221 channel=39
    0, -2, -6, -1, -2, -3, -1, -6, 0,
    -- filter=221 channel=40
    -3, -4, -2, -4, -5, -2, -3, -5, -5,
    -- filter=221 channel=41
    -12, -4, 20, -8, 15, 25, -7, 0, 10,
    -- filter=221 channel=42
    2, 4, -6, -2, -4, -5, -5, 4, -9,
    -- filter=221 channel=43
    -2, 4, 2, -9, -1, -11, -4, 0, -10,
    -- filter=221 channel=44
    5, 8, 1, 6, 0, -7, 4, 2, -2,
    -- filter=221 channel=45
    8, 5, -10, 3, -6, -2, 3, 4, -7,
    -- filter=221 channel=46
    -7, -7, 2, -4, -4, 8, 1, -1, 7,
    -- filter=221 channel=47
    1, 0, -8, 9, 9, -9, 5, 1, -11,
    -- filter=221 channel=48
    -3, 15, -6, -6, 8, -10, 0, 4, -11,
    -- filter=221 channel=49
    4, 3, -10, 3, 4, -11, 4, -3, -3,
    -- filter=221 channel=50
    4, -2, -6, 3, 10, -13, 3, 0, -2,
    -- filter=221 channel=51
    -5, -2, 3, -7, -2, 7, -3, 5, 4,
    -- filter=221 channel=52
    -4, 6, -4, 7, 16, 6, 4, 0, 3,
    -- filter=221 channel=53
    0, 6, 2, -7, 0, -10, 6, 5, -2,
    -- filter=221 channel=54
    4, 1, -7, 0, 2, -6, 3, 0, -4,
    -- filter=221 channel=55
    -9, 10, -2, -2, 17, -18, 3, 2, -14,
    -- filter=221 channel=56
    -3, 0, 13, 5, 4, 7, -1, 5, 5,
    -- filter=221 channel=57
    2, 0, 0, 1, -3, -3, -2, 0, 1,
    -- filter=221 channel=58
    10, 4, -5, -6, -5, 5, 3, -8, 1,
    -- filter=221 channel=59
    -12, 6, -5, 0, 17, -4, 2, 12, -17,
    -- filter=221 channel=60
    6, -6, 0, 6, 1, -4, 4, 0, -6,
    -- filter=221 channel=61
    0, 6, -2, 3, 11, 0, 6, -1, 3,
    -- filter=221 channel=62
    3, -6, 3, 5, 5, 0, -3, 4, 5,
    -- filter=221 channel=63
    4, 0, 3, 3, -6, -4, 6, -4, -1,
    -- filter=221 channel=64
    3, -6, 4, 5, -8, 0, 4, -6, -6,
    -- filter=221 channel=65
    -4, 6, 0, 5, 1, 5, 5, 6, 4,
    -- filter=221 channel=66
    -5, 14, -3, 6, 26, 8, 4, 13, -6,
    -- filter=221 channel=67
    -3, 7, 3, -3, -6, -2, -3, 0, 0,
    -- filter=221 channel=68
    -1, -5, -3, -3, 3, -6, 2, -4, -3,
    -- filter=221 channel=69
    -8, 6, 4, -4, 0, 3, 3, 1, 1,
    -- filter=221 channel=70
    -10, 9, -11, 2, 14, -10, -6, 9, 2,
    -- filter=221 channel=71
    -5, -11, 0, 0, -10, 0, -9, -6, -12,
    -- filter=221 channel=72
    -5, 1, -5, -4, 4, -7, -2, 7, -12,
    -- filter=221 channel=73
    -3, 3, -10, 4, 10, -13, 0, 10, 0,
    -- filter=221 channel=74
    6, 0, 0, 4, 16, -2, 5, 2, 7,
    -- filter=221 channel=75
    0, 5, -1, -7, 5, 2, -8, 2, -4,
    -- filter=221 channel=76
    -2, 4, -3, -11, 4, -6, 0, 3, -13,
    -- filter=221 channel=77
    4, 0, 5, -5, 4, -1, -5, 7, 6,
    -- filter=221 channel=78
    0, 6, -1, 0, -3, 2, 5, -3, 5,
    -- filter=221 channel=79
    -13, 20, -14, -7, 32, -11, -11, 10, -16,
    -- filter=221 channel=80
    -2, 12, -7, -5, 18, -10, -5, 2, -11,
    -- filter=221 channel=81
    -5, 6, -3, 3, -1, 2, 1, -1, 5,
    -- filter=221 channel=82
    -1, -7, 0, -2, -3, -7, -3, -1, -7,
    -- filter=221 channel=83
    4, 1, -3, 7, -5, -10, -1, -6, -5,
    -- filter=221 channel=84
    -1, 12, -9, -4, 18, -6, 3, 2, 3,
    -- filter=221 channel=85
    -5, -4, 5, 0, 4, 0, 0, -2, -2,
    -- filter=221 channel=86
    -3, 6, -6, -3, 9, -1, -1, 8, -2,
    -- filter=221 channel=87
    3, 5, -2, -7, 9, 4, 5, -4, 9,
    -- filter=221 channel=88
    3, -5, 6, 8, -4, -6, -6, 2, 5,
    -- filter=221 channel=89
    -13, 5, -8, -9, 15, -16, -9, 13, -15,
    -- filter=221 channel=90
    2, -5, 9, 3, -1, 6, -2, -1, 0,
    -- filter=221 channel=91
    4, 4, -10, 3, 8, -17, 4, 4, -11,
    -- filter=221 channel=92
    5, -5, 4, 0, -5, 0, -5, 5, 7,
    -- filter=221 channel=93
    9, 9, -3, 5, 0, -13, 4, 0, -14,
    -- filter=221 channel=94
    7, -4, 3, -3, 7, -7, -3, -5, -3,
    -- filter=221 channel=95
    1, -5, 3, 7, 6, -3, 0, 7, 5,
    -- filter=221 channel=96
    4, 4, -7, -6, 6, -5, 0, -2, 0,
    -- filter=221 channel=97
    -3, 0, 0, 5, -10, -4, -4, -8, -9,
    -- filter=221 channel=98
    -3, 10, -5, 0, 20, -14, 1, 15, -10,
    -- filter=221 channel=99
    4, 2, 2, 6, 13, -10, 0, 6, -5,
    -- filter=221 channel=100
    -4, 6, 9, 8, 8, 16, -3, 0, 12,
    -- filter=221 channel=101
    -5, -4, -11, 5, -12, -8, -8, -2, -14,
    -- filter=221 channel=102
    4, -4, 5, -4, -4, 3, 6, 1, 1,
    -- filter=221 channel=103
    -4, 4, -10, 5, -3, -11, 1, 6, -19,
    -- filter=221 channel=104
    2, 4, 0, 3, 6, -16, 7, 2, -13,
    -- filter=221 channel=105
    -3, 5, 2, -6, 5, 1, -3, -2, 0,
    -- filter=221 channel=106
    -1, -6, 0, -9, -4, 6, 0, 0, 8,
    -- filter=221 channel=107
    -6, -1, -10, -5, 2, -13, -2, 0, -6,
    -- filter=221 channel=108
    5, -1, 7, 1, -6, 10, 3, -8, -3,
    -- filter=221 channel=109
    0, 10, -11, -1, 29, -14, 8, 2, -13,
    -- filter=221 channel=110
    2, 0, -5, 7, 1, -7, -2, 0, -3,
    -- filter=221 channel=111
    -1, -5, 7, -2, 3, -2, -4, -4, -6,
    -- filter=221 channel=112
    -2, 6, -2, -1, 14, -9, -3, -2, 2,
    -- filter=221 channel=113
    -6, 5, -6, 4, 15, -6, -1, 0, -8,
    -- filter=221 channel=114
    -12, 26, -16, -14, 30, -14, -10, 17, -5,
    -- filter=221 channel=115
    -2, 5, 7, -2, 8, -3, -1, 5, 5,
    -- filter=221 channel=116
    -10, 15, -10, -2, 9, -16, -9, 2, -5,
    -- filter=221 channel=117
    1, -2, 2, -8, -3, -4, -6, 6, 2,
    -- filter=221 channel=118
    -1, 4, 0, -2, -3, 4, -6, -6, 4,
    -- filter=221 channel=119
    -2, 6, 18, 3, 7, 30, 6, 8, 25,
    -- filter=221 channel=120
    5, 11, -3, 9, 8, -10, 0, 4, 0,
    -- filter=221 channel=121
    -11, -1, 1, -1, 13, 8, -3, 0, -5,
    -- filter=221 channel=122
    9, -4, 0, 12, 3, -11, 10, 0, -7,
    -- filter=221 channel=123
    -4, -5, 0, -3, 7, 15, -3, 4, 5,
    -- filter=221 channel=124
    -4, 1, -8, 0, 3, 0, 4, -6, 2,
    -- filter=221 channel=125
    4, 9, 0, 5, 10, -13, 4, 7, -16,
    -- filter=221 channel=126
    -7, -3, 3, -3, 14, -1, -3, 7, -1,
    -- filter=221 channel=127
    1, 2, 6, 7, 7, 3, -2, -4, -3,
    -- filter=222 channel=0
    7, -5, 4, -5, -1, 0, -8, 0, 2,
    -- filter=222 channel=1
    6, 7, 4, -5, 11, 10, 0, 4, 0,
    -- filter=222 channel=2
    -3, -3, 4, -1, 6, -3, -2, 2, -2,
    -- filter=222 channel=3
    1, -7, 0, 1, 0, 3, -8, -3, 0,
    -- filter=222 channel=4
    4, 12, -6, 0, 2, 0, 0, 2, 0,
    -- filter=222 channel=5
    -7, -4, 2, 5, 9, -7, 0, 0, -10,
    -- filter=222 channel=6
    5, 2, -4, 7, -2, 2, -6, -1, -4,
    -- filter=222 channel=7
    -1, 0, 0, 3, 0, 2, -1, -2, 3,
    -- filter=222 channel=8
    4, 3, -2, 4, 1, 4, 2, -7, 0,
    -- filter=222 channel=9
    -9, 6, -5, -7, 0, -1, -2, 0, -1,
    -- filter=222 channel=10
    -1, -2, 8, -7, 9, -2, 4, 6, 0,
    -- filter=222 channel=11
    -4, -7, -5, -4, -7, -9, -1, -8, 0,
    -- filter=222 channel=12
    2, 3, -4, -3, -4, -2, 7, 2, 8,
    -- filter=222 channel=13
    -1, 0, -3, -3, 5, 10, -2, 0, 0,
    -- filter=222 channel=14
    3, 1, 0, 3, -4, 2, -5, 0, 0,
    -- filter=222 channel=15
    -10, -5, 0, -8, 4, -12, -7, -6, 0,
    -- filter=222 channel=16
    -4, 2, 0, 4, 11, 9, 0, 6, 0,
    -- filter=222 channel=17
    4, -3, -4, 3, -5, 0, -1, 2, -5,
    -- filter=222 channel=18
    0, -11, 2, 0, -4, -4, -1, 6, -9,
    -- filter=222 channel=19
    -4, -2, 7, 1, 0, 0, 6, 7, 0,
    -- filter=222 channel=20
    0, 4, -6, 1, 1, -11, -6, -11, -2,
    -- filter=222 channel=21
    -4, -7, 5, -8, 12, 10, -2, 5, -2,
    -- filter=222 channel=22
    2, -4, 5, -3, -3, -7, -4, 0, -7,
    -- filter=222 channel=23
    -9, -2, -3, -6, 5, -18, 7, -8, -16,
    -- filter=222 channel=24
    5, 0, 3, 0, -6, -1, -6, 2, 6,
    -- filter=222 channel=25
    -3, 5, 7, -6, 11, 6, 7, 10, -6,
    -- filter=222 channel=26
    -4, 0, 0, 3, -2, 0, 4, -2, -2,
    -- filter=222 channel=27
    -13, 7, -8, -9, 16, -5, 9, 6, -13,
    -- filter=222 channel=28
    -2, -6, -4, 1, -3, -1, -3, -3, 1,
    -- filter=222 channel=29
    -5, 0, -4, -3, -6, 1, -4, -7, -4,
    -- filter=222 channel=30
    -9, -1, -4, 4, 3, 2, 6, -1, -3,
    -- filter=222 channel=31
    -10, -7, 7, -10, 9, -3, 6, 4, -15,
    -- filter=222 channel=32
    -9, -5, 0, -2, 2, -7, -2, 2, -4,
    -- filter=222 channel=33
    -3, 0, -2, -5, 2, -4, -2, 6, 2,
    -- filter=222 channel=34
    -4, -1, -9, -1, -1, -8, -1, -4, 0,
    -- filter=222 channel=35
    3, 5, -7, 2, 1, 2, 5, 3, 1,
    -- filter=222 channel=36
    -2, 1, 4, 3, 8, 2, 3, -9, 4,
    -- filter=222 channel=37
    5, 8, 10, 0, 4, 6, 3, 2, -6,
    -- filter=222 channel=38
    -12, 1, 5, 1, 2, -3, -2, 4, 0,
    -- filter=222 channel=39
    -6, 0, -2, -3, 1, -7, -2, -1, -6,
    -- filter=222 channel=40
    -6, 3, -6, -2, 5, 5, 6, -4, 0,
    -- filter=222 channel=41
    5, 1, -7, -5, 5, 10, -4, 9, 2,
    -- filter=222 channel=42
    0, -4, 1, 0, -3, 3, -8, -4, 0,
    -- filter=222 channel=43
    0, 6, 2, 0, -3, -8, 2, 7, 4,
    -- filter=222 channel=44
    -2, -2, 3, 1, 6, -1, -4, 9, 2,
    -- filter=222 channel=45
    1, 2, 1, -1, -4, -6, -6, 0, 0,
    -- filter=222 channel=46
    0, -5, 0, 0, -5, 7, -2, -3, 3,
    -- filter=222 channel=47
    -13, -5, 13, -2, 9, 12, 0, 6, 3,
    -- filter=222 channel=48
    -6, 8, 8, -5, 3, 6, 2, 5, -10,
    -- filter=222 channel=49
    0, 8, 0, 6, 0, 0, -6, -4, 2,
    -- filter=222 channel=50
    -13, -1, -8, -1, -3, 0, -2, -5, -1,
    -- filter=222 channel=51
    1, -5, 7, 1, -4, 1, -1, 0, 1,
    -- filter=222 channel=52
    -5, 7, -1, 6, 9, -9, 1, -3, 0,
    -- filter=222 channel=53
    1, 0, 3, 2, -5, 0, -5, -8, 1,
    -- filter=222 channel=54
    3, 7, -3, 0, 1, 5, -4, 7, 6,
    -- filter=222 channel=55
    -14, -10, -2, 2, -6, -2, 4, 5, -1,
    -- filter=222 channel=56
    0, 1, -2, 6, 0, 1, 3, 5, -5,
    -- filter=222 channel=57
    0, 0, 4, -3, 6, 1, 4, 0, 4,
    -- filter=222 channel=58
    -3, -3, 2, 0, 3, 9, 3, -2, 7,
    -- filter=222 channel=59
    -17, -5, -2, -4, 6, 0, -3, -1, -5,
    -- filter=222 channel=60
    1, 4, 5, -3, 3, -2, 6, 4, 5,
    -- filter=222 channel=61
    2, -2, -4, 0, 8, -5, 4, -1, -5,
    -- filter=222 channel=62
    0, 0, 5, 2, -6, -2, -6, -5, 0,
    -- filter=222 channel=63
    2, -6, 3, -7, 4, -3, 4, 1, -7,
    -- filter=222 channel=64
    0, -2, 4, 7, -7, 2, 7, 3, -4,
    -- filter=222 channel=65
    -4, 4, 5, -3, -3, -3, 1, 0, -1,
    -- filter=222 channel=66
    0, -3, 4, 3, 3, 10, -6, -2, 4,
    -- filter=222 channel=67
    1, -2, 1, -1, 3, 3, 6, 3, 3,
    -- filter=222 channel=68
    3, -6, 5, -3, 2, 2, 0, 0, 6,
    -- filter=222 channel=69
    6, 4, -2, 0, 0, -5, -7, -6, 3,
    -- filter=222 channel=70
    -9, -5, -1, 1, 7, -7, 0, -4, 0,
    -- filter=222 channel=71
    2, -2, -4, -6, 3, 2, 2, 3, 5,
    -- filter=222 channel=72
    -17, -3, -3, -11, 7, 5, -4, 0, -10,
    -- filter=222 channel=73
    -9, 6, -5, 5, 6, 0, 3, 0, 0,
    -- filter=222 channel=74
    0, 4, -7, 7, 10, -13, 0, -2, -7,
    -- filter=222 channel=75
    -8, -4, 4, -5, 6, 8, -5, 8, 7,
    -- filter=222 channel=76
    -1, 1, 0, 2, 0, -8, -3, -4, 4,
    -- filter=222 channel=77
    -5, 2, 0, 3, 0, -5, -1, -6, 0,
    -- filter=222 channel=78
    -6, 0, 7, 6, 8, 3, -4, -4, -6,
    -- filter=222 channel=79
    -11, -14, 0, -11, 5, 0, -1, 4, 4,
    -- filter=222 channel=80
    -19, -1, 10, -17, 14, 2, 0, 6, -9,
    -- filter=222 channel=81
    -1, 3, 0, -4, 0, 0, 0, 5, 0,
    -- filter=222 channel=82
    6, -6, 2, -5, 0, 0, -5, -2, -1,
    -- filter=222 channel=83
    1, 0, -7, -3, -3, 0, 1, 0, -7,
    -- filter=222 channel=84
    0, -1, 0, -4, 9, 0, 0, -5, -9,
    -- filter=222 channel=85
    2, 4, 4, -5, -7, 6, 3, -3, -2,
    -- filter=222 channel=86
    3, 5, -7, 6, -1, -3, 0, 6, -1,
    -- filter=222 channel=87
    -4, 3, 4, 2, 2, -4, 8, -7, -6,
    -- filter=222 channel=88
    -8, 2, 0, 0, -3, 4, -2, 1, -10,
    -- filter=222 channel=89
    -10, -8, 7, -3, -3, 1, 6, 1, -7,
    -- filter=222 channel=90
    0, -2, -4, -3, -3, -8, 7, 3, -5,
    -- filter=222 channel=91
    0, 8, -6, 1, 1, 0, -2, -4, -10,
    -- filter=222 channel=92
    0, -5, -5, 2, 1, 0, -6, 2, 6,
    -- filter=222 channel=93
    -7, 9, -1, 3, 16, 0, 7, 7, -1,
    -- filter=222 channel=94
    -1, -7, 7, 0, 2, -2, 7, 1, 6,
    -- filter=222 channel=95
    1, 3, 8, 2, 5, 1, 5, 0, 0,
    -- filter=222 channel=96
    0, 4, 1, 3, -7, 3, 3, -1, -2,
    -- filter=222 channel=97
    4, -3, 5, -1, 2, -4, -1, -5, 1,
    -- filter=222 channel=98
    -7, 0, 6, -14, 11, -4, 5, 0, -5,
    -- filter=222 channel=99
    -21, 8, -4, -2, -2, -11, 14, -10, -9,
    -- filter=222 channel=100
    9, 0, -6, 3, -7, 3, -3, 3, -4,
    -- filter=222 channel=101
    -2, 8, 2, -2, 2, 3, -5, -2, 0,
    -- filter=222 channel=102
    -1, -1, -1, -5, 1, 3, 3, -1, 5,
    -- filter=222 channel=103
    -19, -6, 1, -10, 4, 0, -5, 8, -8,
    -- filter=222 channel=104
    -12, 6, 3, -7, 10, 0, 5, 5, -10,
    -- filter=222 channel=105
    3, -3, -8, 0, -1, -2, -5, 1, -5,
    -- filter=222 channel=106
    -3, 5, -3, 2, -5, -5, 4, -4, 0,
    -- filter=222 channel=107
    7, 4, 1, 3, 4, -10, 3, 0, -5,
    -- filter=222 channel=108
    3, -8, 1, -7, -4, -3, -4, -2, 6,
    -- filter=222 channel=109
    -16, 4, -5, 1, 14, -2, 9, 6, -10,
    -- filter=222 channel=110
    -9, -1, -6, -10, -1, 5, 1, 2, -2,
    -- filter=222 channel=111
    0, -7, 6, -1, -3, 1, 2, 6, -6,
    -- filter=222 channel=112
    -11, 2, 2, 7, 10, -6, -5, 6, -9,
    -- filter=222 channel=113
    -10, -1, -4, -1, 0, -1, -7, 0, -7,
    -- filter=222 channel=114
    -2, -3, -2, 0, 2, -8, 2, -1, 0,
    -- filter=222 channel=115
    0, -1, -4, 2, 2, -4, 1, -2, 0,
    -- filter=222 channel=116
    -1, -3, 0, 0, -1, 0, 10, -1, -12,
    -- filter=222 channel=117
    -1, -5, -2, -4, -5, 7, 1, -3, -6,
    -- filter=222 channel=118
    -2, -3, -3, 2, 2, 2, -1, 0, 3,
    -- filter=222 channel=119
    7, 4, -5, 13, 0, -8, 6, 2, -3,
    -- filter=222 channel=120
    -12, 1, -6, 7, 9, -5, 9, -1, -8,
    -- filter=222 channel=121
    5, -3, 4, -2, 0, 5, -3, 0, 3,
    -- filter=222 channel=122
    -20, -1, 15, -11, 19, 9, 4, 3, -5,
    -- filter=222 channel=123
    4, -2, 1, 9, 6, 2, -2, 1, 0,
    -- filter=222 channel=124
    -5, 4, 4, 4, 5, -3, 2, 1, 2,
    -- filter=222 channel=125
    -8, -4, 7, -4, 5, -5, 9, 2, -9,
    -- filter=222 channel=126
    -5, -4, 4, -5, 7, 10, -9, 0, 3,
    -- filter=222 channel=127
    0, -1, -6, 0, 4, -5, 0, -3, 4,
    -- filter=223 channel=0
    3, -1, 0, -6, 4, -1, -4, -5, 0,
    -- filter=223 channel=1
    -6, -2, -6, -7, 2, 1, -3, 0, -5,
    -- filter=223 channel=2
    5, -6, 6, -2, -3, -4, 1, -7, 1,
    -- filter=223 channel=3
    4, 2, 5, -6, -3, 4, 7, -2, -2,
    -- filter=223 channel=4
    0, 0, 1, 6, 7, -3, -4, 2, 2,
    -- filter=223 channel=5
    -5, -1, -5, 1, -7, 3, -3, 1, 5,
    -- filter=223 channel=6
    -3, -2, -7, 6, 2, 4, 1, 1, 2,
    -- filter=223 channel=7
    5, 6, 2, -7, -3, -6, 4, 7, 5,
    -- filter=223 channel=8
    -1, -1, -2, 0, -5, 0, 0, 5, 7,
    -- filter=223 channel=9
    1, -1, -2, 3, 3, 0, 3, 4, -1,
    -- filter=223 channel=10
    7, 2, -6, 5, 2, -4, 2, -5, 5,
    -- filter=223 channel=11
    -5, -6, 1, 2, -6, -4, -1, 1, -3,
    -- filter=223 channel=12
    7, -7, 7, 3, 7, -6, -4, 1, 2,
    -- filter=223 channel=13
    6, -4, -7, -2, 3, -1, -6, -1, 0,
    -- filter=223 channel=14
    -6, 0, -4, -5, -2, -6, 1, -3, -4,
    -- filter=223 channel=15
    2, -6, -2, -5, -2, 0, -4, -4, 0,
    -- filter=223 channel=16
    -2, 5, 4, 3, -6, 6, -2, -3, 7,
    -- filter=223 channel=17
    -1, -4, 1, 5, 1, 2, -1, -3, 4,
    -- filter=223 channel=18
    1, -4, 1, 1, 6, 6, 5, -4, -3,
    -- filter=223 channel=19
    -6, -7, -5, -5, 0, -7, -5, 7, 4,
    -- filter=223 channel=20
    -5, 6, -3, 0, 2, 5, 5, 6, 3,
    -- filter=223 channel=21
    0, 3, 3, -3, 3, -1, 6, 5, -5,
    -- filter=223 channel=22
    -7, 0, -3, 4, -3, 4, 2, -6, 2,
    -- filter=223 channel=23
    3, 4, 4, -4, 4, 6, 0, 2, 6,
    -- filter=223 channel=24
    5, -5, 6, -3, 1, -2, 1, 0, -3,
    -- filter=223 channel=25
    -5, -3, -1, -2, 5, -2, 0, -4, 0,
    -- filter=223 channel=26
    -4, 0, -2, -1, -3, -2, -2, -5, 4,
    -- filter=223 channel=27
    2, -7, 4, -3, 5, -4, -5, 1, -1,
    -- filter=223 channel=28
    -3, 0, 5, -4, 6, 3, 1, -7, 2,
    -- filter=223 channel=29
    -2, -1, 5, -2, -1, 0, -5, 0, -5,
    -- filter=223 channel=30
    2, 0, 3, 5, 5, 6, -1, 6, 0,
    -- filter=223 channel=31
    -4, 1, -2, 6, -7, 6, -2, -4, 6,
    -- filter=223 channel=32
    -6, 5, -1, -2, -7, 2, -3, 0, 6,
    -- filter=223 channel=33
    5, 0, 0, 4, -3, 0, -3, -6, -7,
    -- filter=223 channel=34
    1, -5, -5, 0, 3, 1, -3, 3, 0,
    -- filter=223 channel=35
    2, 1, 2, 1, 5, -3, 3, -3, -6,
    -- filter=223 channel=36
    0, -3, 0, 6, 0, -1, -3, 3, 0,
    -- filter=223 channel=37
    -5, -8, 0, 0, -7, 4, 3, -6, 5,
    -- filter=223 channel=38
    6, 4, -5, 1, 1, 3, -7, 5, 0,
    -- filter=223 channel=39
    0, 0, 7, 7, 5, 1, 0, 7, -2,
    -- filter=223 channel=40
    -6, 2, -6, 3, -3, 1, 7, -6, 7,
    -- filter=223 channel=41
    -6, -7, 3, 0, 5, -6, 5, 1, -3,
    -- filter=223 channel=42
    1, -3, -7, -5, 3, 2, 3, -2, -2,
    -- filter=223 channel=43
    5, 7, -2, 1, 0, 7, 4, -3, -1,
    -- filter=223 channel=44
    -1, -5, 0, -3, 1, 5, 6, 0, -2,
    -- filter=223 channel=45
    -5, 2, 7, 3, -1, 0, 1, -5, 2,
    -- filter=223 channel=46
    6, 6, 5, -6, 5, 4, 1, 0, -5,
    -- filter=223 channel=47
    4, 0, -1, 3, -5, 6, -5, -5, -2,
    -- filter=223 channel=48
    -6, -4, 0, -7, -2, 6, -2, 3, 4,
    -- filter=223 channel=49
    5, 0, -2, -5, 1, 0, 2, 4, -6,
    -- filter=223 channel=50
    2, 0, 5, -1, 3, 5, -6, 6, -2,
    -- filter=223 channel=51
    2, -1, 5, -2, 2, -4, -5, -4, 3,
    -- filter=223 channel=52
    6, 0, 4, -6, -5, 4, -2, 0, -4,
    -- filter=223 channel=53
    -1, 1, -5, -4, -6, 2, -1, 5, 1,
    -- filter=223 channel=54
    2, 2, 5, -1, 6, 2, -1, 3, 5,
    -- filter=223 channel=55
    0, 6, -5, -3, 3, -2, -5, 6, -5,
    -- filter=223 channel=56
    -1, -2, 3, -1, -5, 1, -4, 2, 6,
    -- filter=223 channel=57
    -3, 2, -2, 0, -2, 4, 5, 5, 1,
    -- filter=223 channel=58
    -3, 3, 1, -1, 3, -3, -4, -6, 5,
    -- filter=223 channel=59
    -2, -2, 5, 2, -6, 1, 0, -2, -4,
    -- filter=223 channel=60
    -1, 0, 5, 1, 5, 2, 0, 2, -4,
    -- filter=223 channel=61
    1, 1, 0, 5, -6, 5, 1, -6, -3,
    -- filter=223 channel=62
    2, -6, 6, 0, 1, 7, 0, 7, 6,
    -- filter=223 channel=63
    -1, -5, 2, 5, -3, 3, 6, 3, 0,
    -- filter=223 channel=64
    -1, 5, -3, 5, 6, 4, 0, 6, 3,
    -- filter=223 channel=65
    2, -3, -1, 0, 5, 7, 4, 0, -7,
    -- filter=223 channel=66
    -6, -6, 1, -2, 4, 6, -4, -4, 0,
    -- filter=223 channel=67
    -4, 5, 4, 0, -4, -2, 1, 4, 2,
    -- filter=223 channel=68
    2, 3, 3, -5, -4, 7, -3, -6, -4,
    -- filter=223 channel=69
    -7, 1, -4, -6, -6, 6, -2, -4, -6,
    -- filter=223 channel=70
    -1, -2, -3, 6, -5, -1, -3, -8, 0,
    -- filter=223 channel=71
    0, 7, 1, -6, 4, -5, -4, -3, -1,
    -- filter=223 channel=72
    -3, -6, -2, -6, -7, 5, 4, -4, -3,
    -- filter=223 channel=73
    -4, 0, -3, 7, -2, 0, 2, -6, 2,
    -- filter=223 channel=74
    5, -5, 1, 5, 1, -5, -5, 0, -5,
    -- filter=223 channel=75
    0, 0, 0, -2, -2, 5, -3, -3, 0,
    -- filter=223 channel=76
    -6, 0, -1, 7, 0, 1, -2, 2, 0,
    -- filter=223 channel=77
    0, 4, -2, -3, 0, 5, 2, -4, 1,
    -- filter=223 channel=78
    -4, 6, 1, -6, -4, 3, -1, -3, 5,
    -- filter=223 channel=79
    -1, -6, 1, 2, 1, 4, -4, 0, 3,
    -- filter=223 channel=80
    3, -6, -4, 0, 1, -6, 0, -6, 2,
    -- filter=223 channel=81
    2, 6, 0, -3, -3, 5, 0, 1, -4,
    -- filter=223 channel=82
    0, 0, 0, -4, 4, -6, 4, -4, -4,
    -- filter=223 channel=83
    5, 5, -4, -7, -1, -3, 5, -2, -2,
    -- filter=223 channel=84
    -4, -2, 5, -2, 3, -3, 3, 2, 5,
    -- filter=223 channel=85
    3, 5, -3, -1, -4, 0, -6, 3, -7,
    -- filter=223 channel=86
    -1, 0, -1, -5, 1, -6, 0, -4, -7,
    -- filter=223 channel=87
    6, 1, 1, 6, 2, -3, -4, -7, -3,
    -- filter=223 channel=88
    -4, -2, 5, -1, 0, -3, 4, -5, -5,
    -- filter=223 channel=89
    -2, -6, 1, -6, -7, 1, -2, -4, -2,
    -- filter=223 channel=90
    -4, -6, 8, 5, 6, 0, 6, -5, -1,
    -- filter=223 channel=91
    0, -7, -2, -4, -3, 1, 3, 2, 5,
    -- filter=223 channel=92
    2, -3, 0, -4, -3, 0, 4, -2, -3,
    -- filter=223 channel=93
    -7, -1, -3, 5, 1, 0, -4, 5, 6,
    -- filter=223 channel=94
    -6, -1, 2, 3, 1, 7, -3, -4, -4,
    -- filter=223 channel=95
    -4, -5, 6, 5, 3, 2, -5, -5, 4,
    -- filter=223 channel=96
    3, 2, 6, 0, -2, -5, -5, 3, -6,
    -- filter=223 channel=97
    -3, -4, -4, 5, -2, -3, -6, 6, 6,
    -- filter=223 channel=98
    4, -7, -4, 4, 2, -6, -7, -1, 0,
    -- filter=223 channel=99
    6, 1, -5, 7, 2, 7, 5, -4, 3,
    -- filter=223 channel=100
    3, -4, 0, -6, -1, -6, -7, -3, -7,
    -- filter=223 channel=101
    -6, -6, 0, -4, -5, 1, -7, -2, -7,
    -- filter=223 channel=102
    -4, -3, 0, -2, 2, 6, -6, -2, 1,
    -- filter=223 channel=103
    -3, 6, -3, 0, 3, -1, -6, 0, -1,
    -- filter=223 channel=104
    -4, 6, 1, 7, 0, 7, -4, -4, 5,
    -- filter=223 channel=105
    1, 1, 0, -5, 5, -2, -2, 0, 4,
    -- filter=223 channel=106
    -6, 0, -1, 0, 4, 1, 7, -4, -3,
    -- filter=223 channel=107
    -1, 5, -4, 0, 6, 7, 3, -1, 2,
    -- filter=223 channel=108
    1, -5, 0, 0, 4, 4, -3, 4, 6,
    -- filter=223 channel=109
    -5, 5, 5, -1, -3, -6, 4, -2, -5,
    -- filter=223 channel=110
    -1, -2, -4, 1, 7, -3, 1, 2, -7,
    -- filter=223 channel=111
    6, 2, -5, -4, 0, 6, 0, 4, -7,
    -- filter=223 channel=112
    4, -1, -4, -1, 2, 6, -2, -5, 0,
    -- filter=223 channel=113
    1, -2, 0, -3, -7, 4, -7, -3, -1,
    -- filter=223 channel=114
    -1, -5, 5, 6, 4, -7, 4, 1, -4,
    -- filter=223 channel=115
    -1, 7, 6, 7, -2, -5, 5, -7, 2,
    -- filter=223 channel=116
    3, -7, -6, -4, 4, -7, -1, -4, -7,
    -- filter=223 channel=117
    6, 4, 4, 0, 6, -6, -2, 6, 2,
    -- filter=223 channel=118
    -5, 1, 0, 5, 6, 2, 0, 0, 4,
    -- filter=223 channel=119
    2, 6, -5, -5, -6, 3, -3, 0, 1,
    -- filter=223 channel=120
    1, 0, -3, -5, -6, 1, -7, -6, 1,
    -- filter=223 channel=121
    5, 0, 4, 3, -3, -5, 0, -6, 2,
    -- filter=223 channel=122
    -2, 5, 7, -2, 0, 0, -3, -1, 0,
    -- filter=223 channel=123
    -1, 2, -3, -6, 1, 4, 4, 4, -1,
    -- filter=223 channel=124
    -6, -1, 4, 4, 7, -5, -1, 0, -3,
    -- filter=223 channel=125
    -3, -6, 5, 6, -6, 3, 2, -2, 0,
    -- filter=223 channel=126
    -1, 3, -4, -3, -3, 2, -5, -4, -4,
    -- filter=223 channel=127
    -4, -4, -4, -4, -2, 0, -5, 0, -7,
    -- filter=224 channel=0
    -15, -18, 0, -11, -13, -6, -8, -9, 0,
    -- filter=224 channel=1
    -13, -8, -2, -4, -18, -5, -5, 1, 2,
    -- filter=224 channel=2
    0, 7, 4, 1, 6, 3, 4, -3, 7,
    -- filter=224 channel=3
    9, 0, 7, -6, -6, -4, 12, 6, 0,
    -- filter=224 channel=4
    0, -2, -4, 0, -6, 9, 0, 10, 6,
    -- filter=224 channel=5
    0, -7, -3, -5, -7, -11, -8, -7, -6,
    -- filter=224 channel=6
    0, 0, -7, -6, 2, -1, 0, -5, -8,
    -- filter=224 channel=7
    2, -1, 6, 0, 3, 6, 6, -2, 0,
    -- filter=224 channel=8
    0, -2, -1, 12, 8, 0, 6, 7, 0,
    -- filter=224 channel=9
    0, -3, 1, 4, -5, -8, -4, -4, -7,
    -- filter=224 channel=10
    12, 9, -6, 11, 5, -1, -5, 8, 2,
    -- filter=224 channel=11
    0, -1, -3, 8, 5, -10, -5, -7, -11,
    -- filter=224 channel=12
    10, 10, 8, 4, 2, 0, 1, 4, -5,
    -- filter=224 channel=13
    8, 0, 8, 7, 1, -2, 0, 11, -2,
    -- filter=224 channel=14
    -1, 0, -6, -6, 0, -6, -5, -6, 0,
    -- filter=224 channel=15
    -2, -13, -8, -2, -1, 2, 7, 3, 3,
    -- filter=224 channel=16
    -4, 4, 5, 9, 6, -3, -1, 5, 2,
    -- filter=224 channel=17
    0, -2, -5, 0, 3, 1, 6, -7, -3,
    -- filter=224 channel=18
    -7, -15, -13, -11, -21, -11, 0, -10, -8,
    -- filter=224 channel=19
    5, 2, 7, 0, -2, 0, 4, 6, 2,
    -- filter=224 channel=20
    10, 2, -10, 4, -4, -5, 5, 0, -13,
    -- filter=224 channel=21
    4, 6, -8, 11, 9, -8, -6, 3, -1,
    -- filter=224 channel=22
    -8, -11, 5, -7, -5, 0, -2, -2, -5,
    -- filter=224 channel=23
    5, -3, -7, 9, -2, -4, 4, -5, -4,
    -- filter=224 channel=24
    4, -2, -3, 5, 3, -4, -1, -6, 0,
    -- filter=224 channel=25
    5, 5, 0, 8, -1, 1, -2, 6, -5,
    -- filter=224 channel=26
    -5, 0, 5, 5, -2, -1, -1, 5, -6,
    -- filter=224 channel=27
    -11, -3, 0, -6, -15, -6, 1, 2, -1,
    -- filter=224 channel=28
    -4, -2, 1, 6, -3, -6, 0, 4, 6,
    -- filter=224 channel=29
    8, -4, -13, 9, -5, -7, -1, 5, -10,
    -- filter=224 channel=30
    -11, -1, -5, -1, -13, -12, -7, -4, -1,
    -- filter=224 channel=31
    5, 6, -5, 14, 9, -3, -3, 0, -17,
    -- filter=224 channel=32
    2, -4, 0, -2, -9, -7, -2, -1, -1,
    -- filter=224 channel=33
    2, -2, 1, -1, -5, 1, 2, -6, 6,
    -- filter=224 channel=34
    11, 0, 16, 9, 4, 8, 15, -1, 10,
    -- filter=224 channel=35
    2, -2, -6, 7, -2, -5, 3, 6, 4,
    -- filter=224 channel=36
    11, 3, 0, 16, 6, -3, 1, 4, 0,
    -- filter=224 channel=37
    -3, -15, -4, -15, -16, 3, -7, -4, 0,
    -- filter=224 channel=38
    -3, 6, 6, 3, 2, -2, 1, -6, 1,
    -- filter=224 channel=39
    5, -1, -6, 0, 3, 1, 5, -5, -1,
    -- filter=224 channel=40
    0, 5, -1, 0, -1, -7, 4, 2, -4,
    -- filter=224 channel=41
    10, 11, 5, 13, 4, 7, 1, 8, 18,
    -- filter=224 channel=42
    -3, -7, 0, -8, -2, -10, -10, -4, -5,
    -- filter=224 channel=43
    8, 3, 1, 0, 0, -4, 9, -4, -3,
    -- filter=224 channel=44
    -2, -5, 1, -10, 0, 4, -4, -4, 1,
    -- filter=224 channel=45
    -11, -7, 3, -10, 1, -6, -7, 0, -9,
    -- filter=224 channel=46
    -3, 0, 4, -5, 4, 6, -2, 0, 4,
    -- filter=224 channel=47
    -4, 9, -7, 1, 0, -4, 0, 0, -6,
    -- filter=224 channel=48
    -6, -6, -4, 5, -4, 1, 0, -4, 0,
    -- filter=224 channel=49
    0, -12, -1, 1, -4, -6, 0, -4, -7,
    -- filter=224 channel=50
    -1, -13, 2, 2, -13, -4, -8, 0, -6,
    -- filter=224 channel=51
    -5, 0, 1, -6, 0, -5, -6, -3, -4,
    -- filter=224 channel=52
    9, 6, 10, 10, 5, 5, 7, 0, -1,
    -- filter=224 channel=53
    0, 2, 3, 10, 6, -9, -1, -6, 3,
    -- filter=224 channel=54
    -6, 5, -4, 5, -3, 4, -3, -4, -4,
    -- filter=224 channel=55
    1, -2, 2, 9, 2, -11, 9, 4, 1,
    -- filter=224 channel=56
    -4, 0, 0, 10, 4, 3, 0, 5, 8,
    -- filter=224 channel=57
    -3, 3, 5, -2, 3, 0, 5, 4, 6,
    -- filter=224 channel=58
    1, -3, 0, 0, -3, -8, -7, -5, 5,
    -- filter=224 channel=59
    1, 9, 3, -4, 5, -1, -7, -1, -2,
    -- filter=224 channel=60
    0, 7, 2, -4, 0, 3, -1, -5, -1,
    -- filter=224 channel=61
    10, 10, 6, 14, 7, -5, 10, 0, 5,
    -- filter=224 channel=62
    -4, 5, -2, 6, 0, 1, 0, -3, 1,
    -- filter=224 channel=63
    -1, 5, -7, 1, 4, -10, 3, -2, 0,
    -- filter=224 channel=64
    5, 0, -4, 8, 3, 3, 8, 1, -2,
    -- filter=224 channel=65
    -2, -2, 1, 5, -2, 4, 6, 0, 3,
    -- filter=224 channel=66
    8, 8, 8, 14, -1, -6, 11, -2, 4,
    -- filter=224 channel=67
    2, 2, -2, 0, 4, 6, -4, 5, 3,
    -- filter=224 channel=68
    5, -4, -7, 5, -5, 0, -1, 0, -7,
    -- filter=224 channel=69
    2, -6, -2, -2, -4, -6, -6, -4, 3,
    -- filter=224 channel=70
    0, -7, 0, 1, -9, 2, 7, -2, -2,
    -- filter=224 channel=71
    2, 3, 9, 6, 0, -5, -5, 1, 4,
    -- filter=224 channel=72
    1, 6, -3, 2, 2, -1, -4, 2, -8,
    -- filter=224 channel=73
    -2, 1, -6, 0, -7, 0, 2, -4, -5,
    -- filter=224 channel=74
    3, -9, 4, 4, -3, 6, 8, -5, 1,
    -- filter=224 channel=75
    -8, -5, 7, -8, -8, -4, -9, -4, -2,
    -- filter=224 channel=76
    0, -8, -6, 5, -4, 0, -5, -3, 0,
    -- filter=224 channel=77
    0, 3, -7, -1, 4, -3, 5, 2, 0,
    -- filter=224 channel=78
    2, -4, -8, 1, -6, -5, -5, 0, -7,
    -- filter=224 channel=79
    -14, -6, 2, -10, -16, -1, 0, 0, -3,
    -- filter=224 channel=80
    9, 10, -4, -3, 8, -10, -6, 0, -4,
    -- filter=224 channel=81
    -1, -3, 0, 0, -2, 7, -6, 4, -4,
    -- filter=224 channel=82
    5, -2, 0, -6, 0, 5, -6, 4, 4,
    -- filter=224 channel=83
    4, 2, -1, 1, 1, -1, -4, -7, 4,
    -- filter=224 channel=84
    -3, 0, 3, 0, -1, 1, -2, 0, -4,
    -- filter=224 channel=85
    -3, 1, 6, 3, 0, 5, 5, -4, 0,
    -- filter=224 channel=86
    -1, 1, -4, 6, -5, 6, -3, 1, 5,
    -- filter=224 channel=87
    11, 8, 0, 10, -2, 8, 0, 4, 3,
    -- filter=224 channel=88
    7, 10, 3, 17, 7, -1, 9, 0, -5,
    -- filter=224 channel=89
    5, 10, -10, 3, -5, -5, -4, 5, 2,
    -- filter=224 channel=90
    15, 15, 6, 14, 9, -1, 10, 7, -4,
    -- filter=224 channel=91
    -8, -4, -7, 2, -2, -5, -3, -5, 5,
    -- filter=224 channel=92
    -1, 10, -2, 7, 7, 1, -3, 4, -4,
    -- filter=224 channel=93
    -4, -4, -1, -5, 1, -11, -6, -3, -1,
    -- filter=224 channel=94
    0, 2, -3, -4, 5, 2, 7, 3, -5,
    -- filter=224 channel=95
    2, 6, 6, 2, 3, -5, 7, 8, -3,
    -- filter=224 channel=96
    1, -2, -2, 5, -3, 0, 0, 0, 1,
    -- filter=224 channel=97
    6, 1, 10, 1, -3, 0, 2, -5, -6,
    -- filter=224 channel=98
    -4, -8, -11, -3, -6, -2, 3, 1, 1,
    -- filter=224 channel=99
    17, 7, 1, 19, 12, -6, 6, 1, 0,
    -- filter=224 channel=100
    6, 6, 4, 8, 1, -1, -5, 0, -3,
    -- filter=224 channel=101
    7, 0, -3, 9, 5, 0, -1, 8, -3,
    -- filter=224 channel=102
    -1, 2, -1, 6, -4, 7, -4, -1, 1,
    -- filter=224 channel=103
    -2, -3, 1, 0, -3, -9, -1, 0, -10,
    -- filter=224 channel=104
    10, 10, 3, 1, 0, -9, -7, 6, -9,
    -- filter=224 channel=105
    5, -2, -5, 1, -4, -8, 6, -2, 2,
    -- filter=224 channel=106
    5, -6, 1, 4, 2, -1, 0, 0, 3,
    -- filter=224 channel=107
    -6, -6, -11, -7, -5, 0, -6, -9, -2,
    -- filter=224 channel=108
    0, -1, -2, 0, 0, -7, 1, 0, 8,
    -- filter=224 channel=109
    -5, -1, 1, 6, -2, -8, 1, 8, -2,
    -- filter=224 channel=110
    11, 14, 1, 15, 12, 0, 4, 8, -10,
    -- filter=224 channel=111
    -2, 4, -2, -1, 8, 0, -1, -2, 1,
    -- filter=224 channel=112
    -2, 0, 1, 2, -5, -7, 5, 4, -5,
    -- filter=224 channel=113
    0, 0, 9, -5, 2, 6, 5, -2, 1,
    -- filter=224 channel=114
    -14, -16, -18, -15, -33, -5, -1, -8, -6,
    -- filter=224 channel=115
    1, -4, 2, -2, 6, 4, 3, -2, -4,
    -- filter=224 channel=116
    8, 6, -2, -1, -5, -3, -4, 4, 2,
    -- filter=224 channel=117
    1, 3, -2, 3, 0, 4, 0, 2, 0,
    -- filter=224 channel=118
    7, 0, -4, 2, 0, 4, -6, 4, 5,
    -- filter=224 channel=119
    5, 3, 14, 17, -2, 14, 1, -1, 0,
    -- filter=224 channel=120
    -8, -12, 0, 2, -5, 0, 8, 5, -9,
    -- filter=224 channel=121
    3, 9, 4, 2, 11, 1, 5, 5, 4,
    -- filter=224 channel=122
    7, 14, 8, 0, 12, -11, 1, -1, -8,
    -- filter=224 channel=123
    1, -2, -1, 13, 2, 0, 8, 0, 6,
    -- filter=224 channel=124
    0, 0, -1, 7, -1, 1, 3, -6, -5,
    -- filter=224 channel=125
    5, 11, 2, 11, 7, -12, 7, 7, -11,
    -- filter=224 channel=126
    1, 5, -6, 1, 0, -6, 0, 0, -3,
    -- filter=224 channel=127
    2, 6, 7, 0, 5, 1, -2, -5, 6,
    -- filter=225 channel=0
    8, -7, -4, -2, 1, 0, 16, 11, 3,
    -- filter=225 channel=1
    3, -5, -6, -3, 0, -8, 8, 0, 6,
    -- filter=225 channel=2
    -8, -2, 7, 2, 2, -2, -1, -2, 0,
    -- filter=225 channel=3
    -4, 3, 1, 1, 10, 10, 0, 6, -1,
    -- filter=225 channel=4
    -15, -11, -3, 5, -2, -1, -11, -6, 4,
    -- filter=225 channel=5
    -4, 2, 2, 1, -7, -2, 4, 5, 4,
    -- filter=225 channel=6
    2, -3, -12, 0, -3, -4, -1, 10, -3,
    -- filter=225 channel=7
    -5, 2, -6, -3, -1, 1, 2, 1, 0,
    -- filter=225 channel=8
    4, 0, -3, -8, -3, -6, 4, 1, 3,
    -- filter=225 channel=9
    5, 5, 7, 2, -4, 1, -4, 0, -6,
    -- filter=225 channel=10
    7, 8, 6, -7, 0, 0, -2, -7, 0,
    -- filter=225 channel=11
    -5, -7, -2, 4, 2, -3, 6, 6, 7,
    -- filter=225 channel=12
    0, 0, 0, -8, -6, -7, -3, 0, -4,
    -- filter=225 channel=13
    -7, -5, -8, -5, 8, -1, -2, -9, 0,
    -- filter=225 channel=14
    7, -2, -2, 3, -2, -4, 6, 0, 3,
    -- filter=225 channel=15
    5, 0, -14, -2, 4, 5, 8, 0, 7,
    -- filter=225 channel=16
    1, 7, 4, -8, -4, 0, -14, -6, -9,
    -- filter=225 channel=17
    -6, -7, 1, -7, 1, 6, 3, 0, 0,
    -- filter=225 channel=18
    -5, -4, -18, 8, 12, -4, 9, 8, 2,
    -- filter=225 channel=19
    -2, 2, 5, 3, -3, -7, -4, -5, 6,
    -- filter=225 channel=20
    0, -4, -11, 5, 10, 3, 0, 13, 0,
    -- filter=225 channel=21
    10, 14, 9, -4, 0, 8, -12, -16, -13,
    -- filter=225 channel=22
    4, -8, -10, 7, -5, 5, 5, 0, 3,
    -- filter=225 channel=23
    13, -7, -8, 7, 9, 9, 3, -7, -7,
    -- filter=225 channel=24
    0, 5, 0, 1, -6, -4, -2, 5, 0,
    -- filter=225 channel=25
    6, 6, 1, -1, 8, 7, -7, -8, -7,
    -- filter=225 channel=26
    2, 3, 2, -7, 1, -3, -10, 0, 0,
    -- filter=225 channel=27
    4, 2, 0, 13, 10, 4, 0, -2, -9,
    -- filter=225 channel=28
    -6, -7, -4, 0, 0, 5, -3, -6, 0,
    -- filter=225 channel=29
    1, -1, -2, -5, -2, -7, -3, -1, 8,
    -- filter=225 channel=30
    1, 0, 7, 8, 7, 0, -2, -7, 2,
    -- filter=225 channel=31
    9, 14, 26, -5, 1, 14, -16, -28, -6,
    -- filter=225 channel=32
    5, -4, -7, 8, 10, 4, 7, 8, -8,
    -- filter=225 channel=33
    0, 4, -6, 5, 4, 11, 6, -1, -9,
    -- filter=225 channel=34
    -2, -5, -1, -3, -9, -1, -9, -5, 0,
    -- filter=225 channel=35
    0, -2, 5, 1, 2, -3, 0, 0, -3,
    -- filter=225 channel=36
    4, -7, 8, -9, -9, 0, -12, -14, 4,
    -- filter=225 channel=37
    2, 0, -1, 6, -1, -5, -4, 6, 8,
    -- filter=225 channel=38
    2, 8, 5, 4, 6, 3, 0, 0, -6,
    -- filter=225 channel=39
    -5, 2, 3, 1, 0, -1, -2, 0, 0,
    -- filter=225 channel=40
    -5, 5, -4, 3, 2, 7, 0, 8, 6,
    -- filter=225 channel=41
    -1, -3, -8, -11, -22, -17, -9, -10, -5,
    -- filter=225 channel=42
    1, 2, 6, 3, -3, -2, -2, -3, -1,
    -- filter=225 channel=43
    -4, -6, -5, -4, -1, -5, 2, 10, -3,
    -- filter=225 channel=44
    6, 3, 2, 5, 3, 8, -4, -3, -9,
    -- filter=225 channel=45
    -3, 4, -7, 4, 4, -7, 8, -1, -4,
    -- filter=225 channel=46
    5, -3, -1, 3, 3, 1, 4, 2, 0,
    -- filter=225 channel=47
    -3, 6, 17, 0, -2, 8, -11, -18, -14,
    -- filter=225 channel=48
    6, 5, 16, -4, 3, 2, -3, -7, -9,
    -- filter=225 channel=49
    2, 0, -11, -2, 1, -8, -3, 4, 1,
    -- filter=225 channel=50
    11, 5, -3, 1, 0, 11, 2, -10, -3,
    -- filter=225 channel=51
    -1, -5, -6, -6, 3, 4, 3, -1, 0,
    -- filter=225 channel=52
    3, 0, -7, -2, 2, -5, -8, 4, 0,
    -- filter=225 channel=53
    4, 0, 5, 6, 6, 0, -7, -3, 4,
    -- filter=225 channel=54
    -4, -2, 1, -5, -5, 0, -2, -2, -3,
    -- filter=225 channel=55
    1, -5, -11, 0, 8, -1, -5, 0, 3,
    -- filter=225 channel=56
    1, 1, -5, -7, 1, -3, -2, -8, -6,
    -- filter=225 channel=57
    2, 1, -9, 0, 1, -1, -7, -10, 4,
    -- filter=225 channel=58
    3, -2, 0, -7, 0, -3, -2, 0, 6,
    -- filter=225 channel=59
    -4, 9, 1, 6, 1, 0, -5, -10, -2,
    -- filter=225 channel=60
    7, 3, 5, -2, -2, 1, -1, 0, 0,
    -- filter=225 channel=61
    0, 3, 1, -1, -6, 1, -4, -8, -2,
    -- filter=225 channel=62
    0, -5, 5, 0, 4, -6, 7, 0, 5,
    -- filter=225 channel=63
    3, -6, 6, 0, -1, -3, -6, -1, -9,
    -- filter=225 channel=64
    -3, 6, -3, -9, 5, 5, -4, 1, 2,
    -- filter=225 channel=65
    0, -4, 6, 2, 3, 0, 0, -6, 7,
    -- filter=225 channel=66
    -5, -7, -4, -7, -1, -6, 0, -9, -11,
    -- filter=225 channel=67
    -3, 0, -7, 0, -3, -3, -1, -3, -5,
    -- filter=225 channel=68
    4, 0, -7, -3, 4, -7, -1, -4, 7,
    -- filter=225 channel=69
    -7, 0, -8, -3, 3, 1, 0, -2, 2,
    -- filter=225 channel=70
    4, -8, -1, 0, 0, 5, -4, 5, 1,
    -- filter=225 channel=71
    -4, -5, 0, 0, -5, 3, -5, 0, 3,
    -- filter=225 channel=72
    3, 1, 12, -2, 5, 10, -16, -12, -4,
    -- filter=225 channel=73
    -7, 0, -10, 4, -3, -5, 2, 0, 0,
    -- filter=225 channel=74
    6, 5, -4, 2, -5, 0, 3, -2, -4,
    -- filter=225 channel=75
    2, 0, -4, -9, -6, 7, 9, 9, 1,
    -- filter=225 channel=76
    -4, -6, -12, 4, -4, 5, 3, 10, 1,
    -- filter=225 channel=77
    0, -8, -3, 0, 6, 3, -3, 2, 0,
    -- filter=225 channel=78
    -2, -3, 9, -8, -3, 3, 2, -9, -7,
    -- filter=225 channel=79
    -3, -3, -15, 5, 2, 3, 14, 5, -11,
    -- filter=225 channel=80
    2, 7, 24, 6, 4, 5, -17, -20, -7,
    -- filter=225 channel=81
    -4, 5, -6, -7, -6, 2, 1, 4, 2,
    -- filter=225 channel=82
    0, 0, 6, -1, 1, -4, -2, -3, -1,
    -- filter=225 channel=83
    0, 6, 8, 2, 1, -2, 2, -11, 0,
    -- filter=225 channel=84
    -9, 0, -12, -2, 7, -9, -2, 4, -5,
    -- filter=225 channel=85
    -3, -1, 5, -5, -5, 4, -5, -3, 0,
    -- filter=225 channel=86
    8, -12, -1, 0, -4, -10, -3, -2, -2,
    -- filter=225 channel=87
    -4, -13, -8, -6, 3, 0, 0, 4, -3,
    -- filter=225 channel=88
    7, 6, 14, -8, 4, 1, -5, -3, -8,
    -- filter=225 channel=89
    0, 8, 5, 1, 4, -1, 4, -12, -7,
    -- filter=225 channel=90
    -6, -2, 13, -11, -2, 6, -8, -14, 4,
    -- filter=225 channel=91
    -7, 3, -9, 13, 2, 4, 4, -1, -5,
    -- filter=225 channel=92
    2, -3, -8, 1, -7, 4, -3, 3, 0,
    -- filter=225 channel=93
    2, 8, 12, -6, 1, 4, -14, -8, 2,
    -- filter=225 channel=94
    2, -5, 1, -4, -4, 2, 4, 6, 3,
    -- filter=225 channel=95
    -1, -5, 5, -2, 2, 5, 2, -4, -2,
    -- filter=225 channel=96
    0, -4, -3, 7, -1, -5, 6, 2, 1,
    -- filter=225 channel=97
    -6, 0, -5, -3, 0, -3, 5, 9, 8,
    -- filter=225 channel=98
    10, 10, 9, 12, 0, 13, 1, -1, -16,
    -- filter=225 channel=99
    -2, -6, 11, 3, -1, 1, -22, -21, -1,
    -- filter=225 channel=100
    4, 1, -8, 0, -7, -6, -11, -6, -7,
    -- filter=225 channel=101
    -11, -4, -2, -2, -3, 6, 4, 1, 7,
    -- filter=225 channel=102
    -5, -3, 0, -7, -3, 5, -5, 5, 3,
    -- filter=225 channel=103
    5, 9, 8, -9, 0, 6, 0, -3, -4,
    -- filter=225 channel=104
    0, 15, 17, 3, -2, 0, -6, -22, -4,
    -- filter=225 channel=105
    3, -1, -6, -2, -5, -6, 6, 10, -4,
    -- filter=225 channel=106
    -7, 2, -6, 6, 4, 6, 1, -6, 4,
    -- filter=225 channel=107
    3, -8, -13, -2, -1, 1, 12, 3, 7,
    -- filter=225 channel=108
    -4, -1, 2, 0, 3, -1, 6, 0, 2,
    -- filter=225 channel=109
    -4, -2, 4, 13, 8, 4, -8, -6, -2,
    -- filter=225 channel=110
    -7, 2, 1, 1, 0, 9, -1, -8, -4,
    -- filter=225 channel=111
    -4, 0, -6, 2, 0, -8, -7, 1, 0,
    -- filter=225 channel=112
    3, -2, -3, 9, 1, 2, -2, -6, 3,
    -- filter=225 channel=113
    8, 2, 4, 7, -1, 5, 2, -5, 0,
    -- filter=225 channel=114
    -8, -7, -20, 8, 10, -4, 7, 6, -9,
    -- filter=225 channel=115
    -1, 1, -4, 2, -6, 3, 6, -1, -1,
    -- filter=225 channel=116
    -2, 4, -2, 8, 5, 5, -15, -15, -5,
    -- filter=225 channel=117
    4, 5, 0, 5, 0, -3, -4, 0, -1,
    -- filter=225 channel=118
    2, 0, -5, 0, 4, 2, 6, 2, 2,
    -- filter=225 channel=119
    -6, -11, -6, -12, 1, 0, -2, -16, 1,
    -- filter=225 channel=120
    12, -11, 0, 5, 9, 3, -2, -2, -2,
    -- filter=225 channel=121
    5, -3, 1, -7, -6, 8, -1, -12, -10,
    -- filter=225 channel=122
    6, 16, 33, -5, -7, 6, -12, -15, -7,
    -- filter=225 channel=123
    4, 4, 3, 2, 0, 3, -2, -6, 1,
    -- filter=225 channel=124
    -6, -4, -8, -3, 1, -3, 0, -1, 6,
    -- filter=225 channel=125
    -3, 3, 15, 5, -2, 6, -17, -20, -4,
    -- filter=225 channel=126
    0, 4, -9, 1, 2, 0, 8, 0, 4,
    -- filter=225 channel=127
    -1, -1, 4, -8, -1, 0, 5, 5, -9,
    -- filter=226 channel=0
    4, -6, -10, -5, -25, -17, -5, -32, -10,
    -- filter=226 channel=1
    7, 2, -5, 5, -21, -16, 0, -17, -1,
    -- filter=226 channel=2
    4, 4, 8, 0, -4, 4, -4, 4, 1,
    -- filter=226 channel=3
    3, 6, 1, -9, -12, -5, 2, -9, -5,
    -- filter=226 channel=4
    0, 6, 9, -6, -10, -2, 0, -2, 10,
    -- filter=226 channel=5
    -6, -11, -9, 3, -10, -8, 2, -8, -5,
    -- filter=226 channel=6
    -1, 2, 4, -5, -10, -1, -4, -6, -10,
    -- filter=226 channel=7
    6, -4, -7, 3, 1, 5, -2, -1, 0,
    -- filter=226 channel=8
    3, 0, 8, 5, -4, -1, -5, 5, 5,
    -- filter=226 channel=9
    -7, -3, -3, 5, -2, 0, -4, 5, -3,
    -- filter=226 channel=10
    -8, -8, -3, -4, 9, 11, 2, 16, 7,
    -- filter=226 channel=11
    9, 3, 7, 3, 0, 4, -4, 8, 3,
    -- filter=226 channel=12
    1, -3, 9, -6, 1, -4, -2, -8, 7,
    -- filter=226 channel=13
    -5, 1, 4, 2, 0, 2, 2, 4, 0,
    -- filter=226 channel=14
    0, 5, 3, -1, 4, -2, -3, 0, -7,
    -- filter=226 channel=15
    1, 10, 9, -2, -8, -7, 2, -10, 2,
    -- filter=226 channel=16
    -15, -15, -5, -7, 6, -1, -1, 8, 5,
    -- filter=226 channel=17
    3, -1, 4, -4, 3, 0, 0, -1, 1,
    -- filter=226 channel=18
    15, 5, 5, -2, -20, -7, -2, -16, -12,
    -- filter=226 channel=19
    2, -4, 0, -6, 1, 7, 5, -5, 3,
    -- filter=226 channel=20
    -2, 18, 4, 6, -1, 4, -6, 0, 4,
    -- filter=226 channel=21
    -10, -12, -5, 8, 15, 11, 0, 23, 6,
    -- filter=226 channel=22
    0, -3, 1, -9, -16, -12, -6, -6, -11,
    -- filter=226 channel=23
    8, 15, -2, 3, -3, 1, -3, 0, 2,
    -- filter=226 channel=24
    6, 3, 3, 7, -1, 2, 4, -1, -5,
    -- filter=226 channel=25
    3, -6, 7, 1, 3, -1, 0, 1, -2,
    -- filter=226 channel=26
    -15, -10, -8, -4, -1, -4, -6, 0, 8,
    -- filter=226 channel=27
    10, 1, 3, 1, -13, -8, 0, -11, -6,
    -- filter=226 channel=28
    -7, -2, 1, 1, -6, 7, -2, -5, -6,
    -- filter=226 channel=29
    1, 9, 0, -1, -3, -2, -2, -3, 0,
    -- filter=226 channel=30
    -4, -9, -2, 7, 0, -5, -2, 0, -2,
    -- filter=226 channel=31
    -15, 0, -10, 8, 32, 5, 11, 26, 10,
    -- filter=226 channel=32
    11, 9, 12, 4, -14, -6, 2, -13, -9,
    -- filter=226 channel=33
    -1, -2, 6, -3, -8, 0, -4, 2, -6,
    -- filter=226 channel=34
    -9, -1, 4, -2, -5, -5, 0, 0, 6,
    -- filter=226 channel=35
    6, -1, -6, 5, -1, -6, -1, 3, -6,
    -- filter=226 channel=36
    -9, 1, -4, 3, 20, 9, -1, 6, 7,
    -- filter=226 channel=37
    -4, -6, -5, 4, -11, -3, -6, -7, 1,
    -- filter=226 channel=38
    -2, -2, 8, -1, 6, -2, 0, 8, -1,
    -- filter=226 channel=39
    0, 4, 3, 2, -1, -3, 3, -4, 7,
    -- filter=226 channel=40
    2, 6, 1, -3, -8, 6, 0, 4, 0,
    -- filter=226 channel=41
    -5, 7, 8, 1, 1, -2, -8, -10, 2,
    -- filter=226 channel=42
    5, -1, -8, 6, -7, -9, 0, 3, 0,
    -- filter=226 channel=43
    -1, 0, -2, -14, -6, -3, -9, -14, 0,
    -- filter=226 channel=44
    -7, -9, -9, -8, -8, -3, -4, 0, -2,
    -- filter=226 channel=45
    4, 6, -2, 5, -4, 0, -1, -4, 1,
    -- filter=226 channel=46
    0, 1, -7, 5, -2, 4, -8, -2, 0,
    -- filter=226 channel=47
    -8, -12, -16, -3, 0, 2, -2, 18, 0,
    -- filter=226 channel=48
    0, -9, -6, -1, 10, -3, 3, 4, -2,
    -- filter=226 channel=49
    13, 0, 0, 0, -5, 3, 0, -11, 0,
    -- filter=226 channel=50
    9, -7, -10, 4, 1, -6, 8, 3, -8,
    -- filter=226 channel=51
    0, 2, -6, 1, 4, 4, -7, 4, 5,
    -- filter=226 channel=52
    0, 0, 9, 2, -7, 5, -5, 1, 0,
    -- filter=226 channel=53
    -2, 12, 0, -1, 5, -1, -3, -3, 1,
    -- filter=226 channel=54
    -4, 3, 0, 7, 2, 1, 4, -1, 3,
    -- filter=226 channel=55
    13, 11, 4, -5, 0, 0, 1, 0, -3,
    -- filter=226 channel=56
    -3, 3, 7, -2, -3, 3, -3, 6, 2,
    -- filter=226 channel=57
    0, 4, -1, -7, -5, -2, -7, 3, -1,
    -- filter=226 channel=58
    -3, -1, -10, 0, -9, -1, -5, -8, 0,
    -- filter=226 channel=59
    -4, 2, -2, -1, 8, -4, 0, 14, 7,
    -- filter=226 channel=60
    -3, -1, 6, 5, 2, -6, -2, 1, -3,
    -- filter=226 channel=61
    -4, 0, 2, -5, 3, 9, 6, 9, 12,
    -- filter=226 channel=62
    -5, -1, 2, -1, 2, 1, -4, 6, 3,
    -- filter=226 channel=63
    -1, 1, -7, -4, 1, -2, 3, -2, 1,
    -- filter=226 channel=64
    -6, -1, 4, 3, 6, -3, -1, 3, 9,
    -- filter=226 channel=65
    4, -2, 5, 2, -3, 1, 0, -5, -6,
    -- filter=226 channel=66
    -8, 1, 13, -2, -2, -3, 0, -6, 2,
    -- filter=226 channel=67
    -1, 3, 0, 5, -6, -5, -2, 0, -7,
    -- filter=226 channel=68
    5, -3, 6, 7, 6, -1, 6, 3, 0,
    -- filter=226 channel=69
    0, -5, 1, 8, 4, 0, -1, -3, -5,
    -- filter=226 channel=70
    7, 3, 6, -6, -4, -7, 0, -3, -8,
    -- filter=226 channel=71
    -2, -2, 5, -3, -2, 4, -3, 2, -5,
    -- filter=226 channel=72
    -14, 4, -14, 9, 16, 4, 13, 16, 3,
    -- filter=226 channel=73
    6, 7, 1, -3, -6, 6, 2, 3, 10,
    -- filter=226 channel=74
    -4, -3, -5, 5, -2, 5, -5, 9, 10,
    -- filter=226 channel=75
    12, 5, 1, 1, -7, -11, -3, -19, -1,
    -- filter=226 channel=76
    7, 11, 5, -1, -1, 3, 6, 3, 0,
    -- filter=226 channel=77
    2, -7, -6, 6, 2, -2, 7, 3, 7,
    -- filter=226 channel=78
    -4, -2, 2, 3, -2, 3, 4, 5, 0,
    -- filter=226 channel=79
    9, -4, 0, -10, -18, -10, -12, -26, -1,
    -- filter=226 channel=80
    -7, -5, -14, 14, 18, 8, 5, 29, 9,
    -- filter=226 channel=81
    -3, 5, 2, -3, 0, -2, 7, 0, -1,
    -- filter=226 channel=82
    3, 4, -4, -4, 0, -6, 0, -1, -4,
    -- filter=226 channel=83
    -5, 1, -1, -1, -1, 0, 8, 5, 13,
    -- filter=226 channel=84
    7, 6, 3, -4, -5, -8, 0, -15, 4,
    -- filter=226 channel=85
    -6, 3, -3, -6, -3, 0, 6, 4, 0,
    -- filter=226 channel=86
    -10, -6, 6, -6, 0, -5, -4, -2, 3,
    -- filter=226 channel=87
    6, 3, 6, 3, -5, 11, -4, 0, 10,
    -- filter=226 channel=88
    -10, 0, 2, 0, 19, 11, 0, 18, 1,
    -- filter=226 channel=89
    8, 3, 4, 8, 12, -3, 8, 9, 4,
    -- filter=226 channel=90
    -9, 1, 1, -4, 8, 9, 3, 14, 13,
    -- filter=226 channel=91
    4, 1, 1, -3, -3, -3, -4, -6, 8,
    -- filter=226 channel=92
    6, 1, 0, 3, 0, -3, -2, -10, -5,
    -- filter=226 channel=93
    -7, -15, -11, -4, 0, -1, 0, 0, 8,
    -- filter=226 channel=94
    -6, -3, -4, -1, -6, -1, -3, 6, 1,
    -- filter=226 channel=95
    -7, -5, -1, -4, -1, 0, -7, 0, -1,
    -- filter=226 channel=96
    -5, -3, 5, 5, 5, -4, 6, 2, -6,
    -- filter=226 channel=97
    1, 5, -2, 4, -6, 8, -7, -3, -7,
    -- filter=226 channel=98
    -6, -4, 1, -5, 8, 6, 2, 0, -5,
    -- filter=226 channel=99
    -9, -1, -5, 7, 23, 5, 2, 19, 18,
    -- filter=226 channel=100
    -6, -1, 3, 7, 4, 2, -6, -6, 3,
    -- filter=226 channel=101
    1, 4, 1, -2, -8, 4, -2, 5, 15,
    -- filter=226 channel=102
    3, 0, -7, 7, 2, -3, 6, -3, -5,
    -- filter=226 channel=103
    -12, -3, -5, 6, 10, 0, 0, 14, 8,
    -- filter=226 channel=104
    -19, -1, -16, -1, 26, 0, 9, 15, 13,
    -- filter=226 channel=105
    0, 8, 9, 0, -9, 5, 8, 0, -1,
    -- filter=226 channel=106
    2, -2, -4, -4, 3, -5, -1, 4, -4,
    -- filter=226 channel=107
    7, 7, -1, -13, -19, -13, -9, -15, -7,
    -- filter=226 channel=108
    1, 3, 0, -4, -5, -5, -10, 3, 5,
    -- filter=226 channel=109
    -1, -3, 9, 4, 2, 0, -4, 2, 1,
    -- filter=226 channel=110
    -11, 3, 0, -7, 18, 0, 1, 15, 0,
    -- filter=226 channel=111
    -4, -1, 10, 4, -4, 8, 4, 2, 9,
    -- filter=226 channel=112
    -4, -1, -1, 3, -7, -5, -6, -5, 1,
    -- filter=226 channel=113
    5, 6, 3, -6, 6, 2, -2, 0, 6,
    -- filter=226 channel=114
    13, -2, -3, -6, -45, -16, -9, -37, -16,
    -- filter=226 channel=115
    -7, 3, -6, 0, 6, 6, 5, -4, -7,
    -- filter=226 channel=116
    -5, -3, -2, 13, 12, 0, 13, 1, 12,
    -- filter=226 channel=117
    3, -1, -8, -3, 8, 4, 0, 9, 0,
    -- filter=226 channel=118
    -2, 6, 6, 2, 0, 3, -1, 0, -4,
    -- filter=226 channel=119
    -8, -6, -1, -5, -1, -4, 0, 3, 6,
    -- filter=226 channel=120
    -7, 4, 13, -3, -4, 4, -10, -1, 3,
    -- filter=226 channel=121
    -2, -6, 0, 4, 8, 2, 7, 9, 9,
    -- filter=226 channel=122
    -34, -29, -30, -1, 10, 13, 0, 18, 12,
    -- filter=226 channel=123
    -5, -5, 4, -6, 0, -3, -4, 4, -5,
    -- filter=226 channel=124
    0, 6, 6, -2, -1, -5, -3, -1, -3,
    -- filter=226 channel=125
    -7, -5, 0, 0, 23, 0, 10, 20, 15,
    -- filter=226 channel=126
    8, 0, 1, 7, 3, -2, 7, -2, -7,
    -- filter=226 channel=127
    -3, 0, -3, -6, -4, 7, -1, 0, 6,
    -- filter=227 channel=0
    -7, -10, 1, -23, 0, 1, -18, 2, 0,
    -- filter=227 channel=1
    -5, -16, -8, -20, -9, 2, -13, -6, 8,
    -- filter=227 channel=2
    -1, 4, -8, 5, 0, -5, 1, 2, 3,
    -- filter=227 channel=3
    -2, -10, 0, 5, -11, -8, -3, 0, -6,
    -- filter=227 channel=4
    -1, -4, -14, -1, -6, -6, 1, -20, 0,
    -- filter=227 channel=5
    -12, -14, 0, -11, -12, -3, -7, 0, 9,
    -- filter=227 channel=6
    -2, 6, 8, -7, 1, 4, 3, -7, -1,
    -- filter=227 channel=7
    -2, 7, 0, 5, 3, 7, 2, 6, 1,
    -- filter=227 channel=8
    3, -5, -4, 4, -3, -1, -5, -4, -8,
    -- filter=227 channel=9
    2, -3, 9, 0, 1, 8, 0, 1, 5,
    -- filter=227 channel=10
    0, 0, 0, 3, 8, 0, 3, 0, 7,
    -- filter=227 channel=11
    6, 5, 6, 6, 1, 0, -7, -8, 11,
    -- filter=227 channel=12
    -10, -10, -10, -3, 0, 0, -2, -6, -2,
    -- filter=227 channel=13
    -4, 1, -8, -16, -3, -6, -4, -11, 4,
    -- filter=227 channel=14
    -4, 2, -2, 1, -5, 4, 0, -2, 0,
    -- filter=227 channel=15
    -6, 6, 11, -8, -1, 3, -14, -6, 12,
    -- filter=227 channel=16
    -8, -13, -13, 0, -5, -5, -4, 8, -2,
    -- filter=227 channel=17
    0, 5, -3, 1, -1, 5, 1, 7, -7,
    -- filter=227 channel=18
    -1, 13, 15, -24, 7, 18, -25, -14, 8,
    -- filter=227 channel=19
    3, -1, 6, 3, -6, 6, 0, -1, 0,
    -- filter=227 channel=20
    4, 4, 5, 4, -7, 3, 1, -11, 9,
    -- filter=227 channel=21
    -5, -11, -3, 4, 8, -5, 2, 7, 0,
    -- filter=227 channel=22
    -8, -1, -6, -1, -2, 1, 4, -2, 6,
    -- filter=227 channel=23
    6, 5, 0, 4, 19, -1, 2, 5, -3,
    -- filter=227 channel=24
    -3, -1, -5, -6, 1, 6, 0, 7, 1,
    -- filter=227 channel=25
    -8, 0, 4, -15, 4, 8, -5, 0, 17,
    -- filter=227 channel=26
    -8, -1, -8, -1, -8, -4, -7, 1, 1,
    -- filter=227 channel=27
    -12, 8, 6, -14, 17, 18, -11, 6, 21,
    -- filter=227 channel=28
    3, 2, 3, -3, 3, 6, -3, -5, 0,
    -- filter=227 channel=29
    -1, -3, 10, -3, -6, -2, -3, -8, 6,
    -- filter=227 channel=30
    -11, 1, 1, -10, 0, 9, -4, 3, 9,
    -- filter=227 channel=31
    9, 3, -5, 8, 22, -8, 0, 27, 14,
    -- filter=227 channel=32
    -8, -2, 12, -12, 11, 7, -20, 0, 3,
    -- filter=227 channel=33
    -2, -2, 3, -2, 13, 13, -15, 3, 14,
    -- filter=227 channel=34
    -9, -11, 4, -4, -7, -8, 0, -2, -8,
    -- filter=227 channel=35
    1, 0, -7, -7, -2, 3, -1, -4, -3,
    -- filter=227 channel=36
    -1, -5, -10, -1, -5, -6, 0, -6, -1,
    -- filter=227 channel=37
    -18, -8, -5, -10, -3, -5, -11, -6, 2,
    -- filter=227 channel=38
    8, -3, 7, 6, 1, 8, -3, 6, 12,
    -- filter=227 channel=39
    -2, -4, -4, -5, 5, 1, -2, -4, 2,
    -- filter=227 channel=40
    -1, -1, 0, 2, 2, -10, 5, 3, -2,
    -- filter=227 channel=41
    -19, -13, -17, -25, -22, -15, -27, -34, -13,
    -- filter=227 channel=42
    -6, -1, -5, -6, -2, 9, -9, 6, 4,
    -- filter=227 channel=43
    0, -14, -8, 0, 0, -2, 0, -9, -1,
    -- filter=227 channel=44
    -10, -13, -12, -4, 1, -1, 0, 0, 1,
    -- filter=227 channel=45
    -4, -4, 3, 5, 0, 4, 2, -4, 9,
    -- filter=227 channel=46
    0, -6, -8, 2, -4, 3, -8, 0, -6,
    -- filter=227 channel=47
    -12, -18, -7, 0, 2, -3, -3, 6, 4,
    -- filter=227 channel=48
    -5, -2, -1, 2, 7, 10, -2, 0, 11,
    -- filter=227 channel=49
    2, 14, 5, -10, 5, 11, -9, -10, 6,
    -- filter=227 channel=50
    -1, 9, 3, -1, 10, 8, -3, 17, 12,
    -- filter=227 channel=51
    5, 6, -1, -1, -3, -4, -6, 4, -6,
    -- filter=227 channel=52
    -7, 0, 0, 3, 0, -10, 0, -10, -10,
    -- filter=227 channel=53
    1, 0, 8, 4, -6, -4, 3, 0, 8,
    -- filter=227 channel=54
    -1, -3, 6, 0, -4, -3, 3, 2, 3,
    -- filter=227 channel=55
    0, 3, 10, 0, 8, 3, -3, -3, 11,
    -- filter=227 channel=56
    3, 1, -3, -7, -3, -12, -8, -7, -2,
    -- filter=227 channel=57
    -9, -2, 0, 0, -3, -4, 5, -9, -9,
    -- filter=227 channel=58
    -9, 0, -4, -8, -12, 4, 0, 0, -3,
    -- filter=227 channel=59
    -9, -4, 0, -10, 3, 0, -1, 0, 4,
    -- filter=227 channel=60
    -3, 0, 0, 5, 0, -1, -7, 5, 3,
    -- filter=227 channel=61
    -2, 3, -2, -4, -4, -2, -2, -6, -5,
    -- filter=227 channel=62
    -7, -4, 1, -3, -7, 0, 0, -7, -6,
    -- filter=227 channel=63
    3, -7, -3, -5, -3, -8, 0, 7, -4,
    -- filter=227 channel=64
    -3, -4, 1, -4, -6, -5, 3, -5, -3,
    -- filter=227 channel=65
    1, 4, -4, -4, 4, 4, -6, 0, -6,
    -- filter=227 channel=66
    -7, 1, -1, -6, -8, -6, -1, -17, -11,
    -- filter=227 channel=67
    1, -6, -4, 5, 4, 5, -4, -9, -4,
    -- filter=227 channel=68
    1, 1, 3, 3, 3, 0, 5, 2, 2,
    -- filter=227 channel=69
    4, -6, -5, 1, 2, 4, -6, 4, -6,
    -- filter=227 channel=70
    -4, 7, 0, -2, 11, -4, -12, 2, 7,
    -- filter=227 channel=71
    5, -9, 0, 8, -1, -7, -2, 6, 0,
    -- filter=227 channel=72
    -2, 6, 1, 4, 20, 8, -2, 6, 13,
    -- filter=227 channel=73
    -3, 9, 5, -3, 9, 0, -4, -4, 9,
    -- filter=227 channel=74
    -8, -4, -3, 3, 7, -5, -3, 4, 0,
    -- filter=227 channel=75
    -6, -5, -3, -21, -10, -5, -12, 3, 7,
    -- filter=227 channel=76
    -9, 0, 4, -10, -12, 2, -9, -13, -2,
    -- filter=227 channel=77
    2, 0, 2, -1, 5, -2, -4, 4, -2,
    -- filter=227 channel=78
    0, -3, 5, -1, -4, 6, 3, -3, 2,
    -- filter=227 channel=79
    -6, 11, 7, -18, 13, 14, -25, -14, 14,
    -- filter=227 channel=80
    0, 3, -1, 10, 20, 3, 7, 18, 15,
    -- filter=227 channel=81
    -5, -1, 3, -5, -3, -6, -4, 5, 5,
    -- filter=227 channel=82
    1, -3, 3, -2, -8, 0, 4, -6, 1,
    -- filter=227 channel=83
    9, 0, 5, 5, 3, 5, 2, -6, 4,
    -- filter=227 channel=84
    -3, 9, 8, -17, 0, 6, -14, -2, 0,
    -- filter=227 channel=85
    -3, 1, -3, -3, 2, -2, 1, 4, -7,
    -- filter=227 channel=86
    -6, -4, 0, -3, -8, -6, -7, -6, -11,
    -- filter=227 channel=87
    -6, -7, -7, -10, 1, -5, 0, -7, 0,
    -- filter=227 channel=88
    3, -4, -6, 9, -6, -8, 9, -6, -12,
    -- filter=227 channel=89
    2, 8, -1, -11, 0, 13, 0, 0, 15,
    -- filter=227 channel=90
    6, -5, -11, 9, 1, -14, -2, 7, -6,
    -- filter=227 channel=91
    3, 16, 3, -15, 6, 6, -5, -5, 8,
    -- filter=227 channel=92
    2, -9, 0, 3, 1, 0, 5, -5, -5,
    -- filter=227 channel=93
    -12, -14, -9, -5, 0, -5, -9, 0, 0,
    -- filter=227 channel=94
    5, -6, 4, 3, 7, 0, -3, 7, 2,
    -- filter=227 channel=95
    5, -2, 3, -2, -2, -4, 2, -5, 5,
    -- filter=227 channel=96
    -2, -1, 5, 3, 1, 1, -9, 1, 0,
    -- filter=227 channel=97
    -2, -9, -5, 3, -3, -4, 2, 2, -4,
    -- filter=227 channel=98
    1, -1, 8, 3, 22, 14, 0, 10, 17,
    -- filter=227 channel=99
    1, 9, 0, 12, 19, 5, 6, 5, 0,
    -- filter=227 channel=100
    2, 3, -5, -1, 1, 0, -2, -12, -12,
    -- filter=227 channel=101
    4, -4, -8, 0, -6, -10, -6, -4, -5,
    -- filter=227 channel=102
    0, 2, 4, 0, 0, 6, 0, 3, -2,
    -- filter=227 channel=103
    -4, 0, 7, -5, -4, -10, 5, 13, 2,
    -- filter=227 channel=104
    3, 0, -10, 4, 5, -3, 0, 13, 11,
    -- filter=227 channel=105
    -4, 0, -2, -2, -3, -3, -2, -7, -5,
    -- filter=227 channel=106
    -9, -6, 3, -9, -1, -8, 2, -9, -2,
    -- filter=227 channel=107
    4, 6, 8, 0, 0, -1, -3, -4, 11,
    -- filter=227 channel=108
    -12, -2, 0, -8, -11, -8, 0, -11, 0,
    -- filter=227 channel=109
    -12, 7, 9, -4, 11, 11, -20, 5, 11,
    -- filter=227 channel=110
    7, 2, -6, 4, 9, -11, -4, 6, -3,
    -- filter=227 channel=111
    -5, -1, -2, -1, 0, -3, -6, -4, 1,
    -- filter=227 channel=112
    -3, 0, 8, 2, 9, 3, 1, 13, 8,
    -- filter=227 channel=113
    6, -3, 8, 9, 13, -4, 0, 14, -3,
    -- filter=227 channel=114
    -8, 17, 12, -26, 6, 11, -28, -10, 11,
    -- filter=227 channel=115
    0, 0, 4, 3, -3, -4, 6, 5, 1,
    -- filter=227 channel=116
    4, 2, 0, -7, 17, 11, -8, 2, 14,
    -- filter=227 channel=117
    -3, 0, -10, 3, -1, 6, 6, -3, 4,
    -- filter=227 channel=118
    0, 6, 2, 0, 6, 4, 0, -5, 0,
    -- filter=227 channel=119
    -4, -10, -4, -11, -8, -6, -5, 0, 0,
    -- filter=227 channel=120
    3, 5, 7, 1, 15, 15, -6, 14, 11,
    -- filter=227 channel=121
    -10, 0, -6, -3, -10, -2, -8, -2, -5,
    -- filter=227 channel=122
    -2, -19, -18, 0, -5, -11, 8, 15, 4,
    -- filter=227 channel=123
    -9, -4, -2, -4, -8, -7, -6, -7, -5,
    -- filter=227 channel=124
    4, 0, -3, -1, -6, -6, 2, -10, 2,
    -- filter=227 channel=125
    3, 5, 4, -6, 22, -1, -4, 4, 11,
    -- filter=227 channel=126
    -12, -11, -5, -15, -8, 9, -5, -6, -2,
    -- filter=227 channel=127
    -1, -5, -5, -6, -5, -10, -5, 3, -1,
    -- filter=228 channel=0
    2, 3, -6, -8, -17, -18, -6, -23, -12,
    -- filter=228 channel=1
    8, 3, -12, 1, -16, -21, -4, -20, -23,
    -- filter=228 channel=2
    -7, -4, 6, -2, 5, -9, 0, -4, -1,
    -- filter=228 channel=3
    -4, 2, 5, -3, 8, 2, -3, 0, 0,
    -- filter=228 channel=4
    -2, 0, 5, 0, 2, -1, -15, -7, 6,
    -- filter=228 channel=5
    8, 10, -4, 0, -10, -2, -3, -3, -11,
    -- filter=228 channel=6
    0, -8, -1, 4, -7, -4, -4, 7, 8,
    -- filter=228 channel=7
    -3, -4, -5, 4, 0, 3, -5, -2, -4,
    -- filter=228 channel=8
    5, -6, -2, 4, -4, -9, 0, -9, 3,
    -- filter=228 channel=9
    3, 2, 7, -1, -1, 0, 7, 2, -7,
    -- filter=228 channel=10
    2, 15, 4, 8, 11, 2, 11, 3, 2,
    -- filter=228 channel=11
    -2, -13, -5, 5, 3, 2, 0, 9, 9,
    -- filter=228 channel=12
    -7, -6, 2, 5, -4, -11, 0, -7, -9,
    -- filter=228 channel=13
    -1, -3, 1, 1, 0, -5, 6, -6, -1,
    -- filter=228 channel=14
    1, 3, 0, -7, -2, -5, -1, 2, -6,
    -- filter=228 channel=15
    0, -5, 9, -4, -8, 2, 4, 4, -2,
    -- filter=228 channel=16
    5, 0, -4, 6, -4, -6, -3, -7, -8,
    -- filter=228 channel=17
    -7, 0, 1, -1, 1, 6, -2, 1, 5,
    -- filter=228 channel=18
    -2, 8, 7, 8, -9, 0, 12, -9, -7,
    -- filter=228 channel=19
    -4, 2, -1, -2, 5, 0, 5, 6, -6,
    -- filter=228 channel=20
    -15, -14, 4, -8, -7, 16, 6, 11, 5,
    -- filter=228 channel=21
    1, 4, 1, -2, 5, 0, -1, 5, -10,
    -- filter=228 channel=22
    0, -3, 2, 0, -3, 0, -1, -9, -4,
    -- filter=228 channel=23
    9, 7, 17, -3, 0, 3, 1, -5, -5,
    -- filter=228 channel=24
    -2, -6, -2, 2, -1, -4, -3, 3, 5,
    -- filter=228 channel=25
    3, 10, -1, 0, 0, -6, 0, -9, -7,
    -- filter=228 channel=26
    -5, -1, 0, 0, 6, 4, 6, -4, 5,
    -- filter=228 channel=27
    5, 18, 12, 6, 0, -12, 0, -12, -9,
    -- filter=228 channel=28
    2, -3, -1, -2, 0, -5, 0, -3, 4,
    -- filter=228 channel=29
    0, -1, -2, 4, 1, 5, 4, 3, 13,
    -- filter=228 channel=30
    4, 8, -4, 5, -4, -7, -6, -8, -12,
    -- filter=228 channel=31
    -4, 8, 7, 0, 0, 0, -4, 1, -10,
    -- filter=228 channel=32
    2, 10, 4, -1, -8, -5, 7, -4, -5,
    -- filter=228 channel=33
    3, 7, 11, 1, 7, 4, 0, -8, -6,
    -- filter=228 channel=34
    11, 0, -8, -3, -14, -5, -5, -5, -3,
    -- filter=228 channel=35
    2, 0, 0, 2, 4, 5, 0, 0, -3,
    -- filter=228 channel=36
    -1, -6, -9, 3, -6, -3, -2, -6, -1,
    -- filter=228 channel=37
    10, -6, -9, 6, -7, -9, -8, -23, -16,
    -- filter=228 channel=38
    0, 6, 9, -5, 4, -1, -1, -5, -7,
    -- filter=228 channel=39
    -9, 0, -6, -4, 3, 9, -2, 0, 8,
    -- filter=228 channel=40
    -10, -6, -7, -7, -1, -2, 2, 3, 4,
    -- filter=228 channel=41
    -4, -15, -21, -2, -4, -15, 0, 6, -15,
    -- filter=228 channel=42
    -4, 1, -1, -4, 2, -3, 0, -4, -1,
    -- filter=228 channel=43
    9, 0, 9, -1, -7, 5, 0, 2, 4,
    -- filter=228 channel=44
    -2, 11, 3, -4, -6, -7, 1, -6, -4,
    -- filter=228 channel=45
    0, -4, 0, -2, -10, 4, -9, -9, 5,
    -- filter=228 channel=46
    -3, 2, -5, 4, -8, 4, -4, 0, -5,
    -- filter=228 channel=47
    -3, 10, 11, 2, -1, -3, 3, -2, -9,
    -- filter=228 channel=48
    0, 2, -1, 6, -4, -11, 3, -11, -11,
    -- filter=228 channel=49
    -1, -1, 8, -5, -10, -7, 0, 0, -4,
    -- filter=228 channel=50
    -2, 8, 4, 6, 1, -8, -1, -3, -10,
    -- filter=228 channel=51
    3, -1, -5, 0, -3, -3, -6, 6, 4,
    -- filter=228 channel=52
    2, -2, 3, -8, -8, -5, 4, 2, -4,
    -- filter=228 channel=53
    -4, -1, -2, -1, 1, 9, 8, -2, 9,
    -- filter=228 channel=54
    0, 0, -5, 6, 3, 2, 0, 4, 1,
    -- filter=228 channel=55
    -1, -4, -1, 5, -2, 0, 6, 6, 5,
    -- filter=228 channel=56
    0, -2, -6, 6, 0, -8, 2, -9, -7,
    -- filter=228 channel=57
    -4, 4, 0, -4, -4, -1, -4, -9, -1,
    -- filter=228 channel=58
    8, 4, -2, -6, -3, -7, 4, 0, 0,
    -- filter=228 channel=59
    0, 14, 8, 0, 2, -12, 0, 2, -4,
    -- filter=228 channel=60
    -6, -3, 4, -3, 0, -6, 7, 0, 2,
    -- filter=228 channel=61
    -2, -10, -9, -1, -3, 4, 5, 5, -6,
    -- filter=228 channel=62
    4, 1, 1, 6, 2, -4, -3, -2, 6,
    -- filter=228 channel=63
    -3, -4, -4, 0, 0, -5, -6, 6, 0,
    -- filter=228 channel=64
    -8, -5, -10, -5, 2, 2, -3, -1, -4,
    -- filter=228 channel=65
    -6, -1, -5, 6, 0, 7, 1, 4, -5,
    -- filter=228 channel=66
    6, -3, -6, 2, -4, -9, 7, 0, -11,
    -- filter=228 channel=67
    1, -4, 5, 2, 4, 6, -4, -6, 4,
    -- filter=228 channel=68
    1, -7, 2, 5, -1, -3, -8, -3, 1,
    -- filter=228 channel=69
    0, 0, -6, -7, 1, -5, -6, 0, -2,
    -- filter=228 channel=70
    4, 3, 7, -8, -10, -6, -10, -3, -7,
    -- filter=228 channel=71
    7, 3, 11, -6, 6, 9, -2, 1, 0,
    -- filter=228 channel=72
    -4, 4, 7, 3, 9, 1, 5, 8, -3,
    -- filter=228 channel=73
    5, 2, 8, -1, -6, -8, 6, 3, 3,
    -- filter=228 channel=74
    7, 7, 2, -4, -2, -6, -9, -1, -4,
    -- filter=228 channel=75
    -2, 0, 7, -9, -3, -13, -2, -22, -14,
    -- filter=228 channel=76
    -4, -3, -9, 0, 0, 7, 1, 3, 0,
    -- filter=228 channel=77
    -2, -7, -3, 6, 3, -3, -1, 4, -2,
    -- filter=228 channel=78
    -3, 4, 5, 9, 6, -6, 3, 0, 4,
    -- filter=228 channel=79
    -1, 13, 13, -4, -5, -4, 0, -9, -8,
    -- filter=228 channel=80
    6, 18, 14, 5, 10, -10, -2, 5, -9,
    -- filter=228 channel=81
    -2, -1, 6, 3, -6, 4, -5, -6, 4,
    -- filter=228 channel=82
    1, 5, 0, -1, 4, 4, -6, 5, -3,
    -- filter=228 channel=83
    0, 2, 8, 0, 4, -2, 0, -7, 4,
    -- filter=228 channel=84
    0, 3, -6, 3, -8, 0, 1, -3, -5,
    -- filter=228 channel=85
    5, 0, 3, 4, 4, -3, 2, -1, -6,
    -- filter=228 channel=86
    0, -7, 0, -1, -5, -6, -1, 0, -11,
    -- filter=228 channel=87
    -1, -7, -9, -5, -4, 2, -1, 1, 0,
    -- filter=228 channel=88
    -5, 0, -10, -7, -10, -9, -10, 5, -4,
    -- filter=228 channel=89
    1, 9, 10, 0, 7, 4, 3, 0, -1,
    -- filter=228 channel=90
    -8, -3, -7, -11, 0, -6, -7, -1, -5,
    -- filter=228 channel=91
    4, 7, 8, -2, -6, -9, -8, -10, 0,
    -- filter=228 channel=92
    8, -3, -5, -2, 2, -8, -4, 0, -4,
    -- filter=228 channel=93
    2, 12, 7, 2, 3, -14, -2, 0, -6,
    -- filter=228 channel=94
    -4, 2, 2, -7, 6, 6, 6, -6, 0,
    -- filter=228 channel=95
    6, 9, 1, -2, -3, 5, -6, 0, 0,
    -- filter=228 channel=96
    -2, 0, 1, 5, -6, 7, 0, -1, -5,
    -- filter=228 channel=97
    -3, 4, 3, 0, 6, -3, 4, 3, 2,
    -- filter=228 channel=98
    1, 20, 18, 8, 12, -8, 4, 1, -8,
    -- filter=228 channel=99
    -2, 4, 10, 4, -2, -7, 6, 5, 5,
    -- filter=228 channel=100
    3, 0, 1, 0, 1, -7, 0, 2, 3,
    -- filter=228 channel=101
    0, -1, 7, 3, 0, 1, -8, -7, -5,
    -- filter=228 channel=102
    -2, -1, 0, 0, 5, -2, 4, 3, 4,
    -- filter=228 channel=103
    10, 15, 4, 1, -1, -9, -7, -3, -14,
    -- filter=228 channel=104
    8, 7, 12, 1, 10, -2, 4, -4, -6,
    -- filter=228 channel=105
    -5, -11, 1, 4, -4, 13, 0, 3, 14,
    -- filter=228 channel=106
    -10, 0, 2, -4, -6, -5, -3, 7, 6,
    -- filter=228 channel=107
    -10, 1, 6, 0, -4, -1, -3, -1, 8,
    -- filter=228 channel=108
    6, 1, -8, 2, -6, -3, 2, 2, -2,
    -- filter=228 channel=109
    8, 16, 1, 8, 3, 0, -1, -3, -2,
    -- filter=228 channel=110
    6, 13, 6, -1, 0, 9, 1, -2, 2,
    -- filter=228 channel=111
    -5, 3, -4, -1, -3, 4, 2, 0, -7,
    -- filter=228 channel=112
    6, 1, -3, 2, 2, -6, 4, -10, -5,
    -- filter=228 channel=113
    12, 11, 11, 5, 8, -5, -3, -3, 0,
    -- filter=228 channel=114
    1, 5, 11, -4, -11, -4, -2, -10, -17,
    -- filter=228 channel=115
    -1, 6, 6, -6, 4, 0, -2, 5, 1,
    -- filter=228 channel=116
    6, 10, 4, 7, -5, -10, 2, 2, 2,
    -- filter=228 channel=117
    -6, -4, -4, -3, 2, -1, -4, -7, -6,
    -- filter=228 channel=118
    -7, -6, 6, 4, 2, 5, 5, 0, -2,
    -- filter=228 channel=119
    4, 0, 0, 2, -7, -4, -6, -5, -10,
    -- filter=228 channel=120
    11, 10, 6, -2, 0, -3, -4, -1, 2,
    -- filter=228 channel=121
    3, 1, 1, 5, 4, 2, 8, -6, -9,
    -- filter=228 channel=122
    -2, 5, -2, -4, 2, -7, -14, 1, -12,
    -- filter=228 channel=123
    6, -2, -3, 0, -6, -2, -9, 0, -3,
    -- filter=228 channel=124
    6, -2, -5, 0, 3, 12, 8, 5, 6,
    -- filter=228 channel=125
    5, 3, -2, 0, 0, -9, -6, -5, 2,
    -- filter=228 channel=126
    -1, 8, 2, 2, -1, 4, 7, 4, -1,
    -- filter=228 channel=127
    -1, 1, -1, 0, 2, 0, -1, 6, -1,
    -- filter=229 channel=0
    -23, 1, 2, 2, -1, -12, 0, 8, 0,
    -- filter=229 channel=1
    -10, 2, 1, 7, 18, -10, 5, -4, -4,
    -- filter=229 channel=2
    -5, -3, 3, 0, 4, 1, -4, 13, 6,
    -- filter=229 channel=3
    -2, 9, 10, 0, -2, 0, 11, 5, 16,
    -- filter=229 channel=4
    -6, -1, 11, -15, 24, 20, 18, 21, 22,
    -- filter=229 channel=5
    -10, 8, 6, -2, 1, 8, 1, -6, -10,
    -- filter=229 channel=6
    4, 1, -3, -8, -6, -1, -1, 8, 2,
    -- filter=229 channel=7
    -5, -3, -7, -5, -5, -5, 3, -3, -7,
    -- filter=229 channel=8
    0, -10, 11, 0, 1, 7, -4, 11, 1,
    -- filter=229 channel=9
    1, 9, -6, 1, -6, -2, -2, 5, 0,
    -- filter=229 channel=10
    1, 11, -5, 6, -3, -8, -2, 3, 8,
    -- filter=229 channel=11
    4, -7, -2, -13, -10, -1, -6, 7, 27,
    -- filter=229 channel=12
    0, -3, -2, 10, -4, 1, -2, 7, -7,
    -- filter=229 channel=13
    5, 2, -18, 8, -4, -13, -10, 5, 19,
    -- filter=229 channel=14
    -2, -7, 7, 1, -2, 6, -1, -2, -6,
    -- filter=229 channel=15
    5, -7, -14, -7, -25, -8, 1, 16, 21,
    -- filter=229 channel=16
    -4, 16, 5, 4, 9, -4, -11, -18, -18,
    -- filter=229 channel=17
    -6, 5, 0, 6, 4, -3, 6, -4, 0,
    -- filter=229 channel=18
    3, -7, -34, 0, -15, -10, -8, 16, 37,
    -- filter=229 channel=19
    -3, -2, 3, -4, -3, 3, -2, -3, -2,
    -- filter=229 channel=20
    12, -24, -11, -19, -21, 7, 0, 22, 29,
    -- filter=229 channel=21
    13, 28, 17, 3, 4, -5, -9, -20, -11,
    -- filter=229 channel=22
    1, 1, -6, 5, -1, -8, 1, 11, 3,
    -- filter=229 channel=23
    10, -28, -18, -10, -37, -15, -11, 35, 23,
    -- filter=229 channel=24
    0, 1, -3, 6, 0, 0, -3, 3, 4,
    -- filter=229 channel=25
    4, 0, -12, 10, -6, -11, -13, 3, 5,
    -- filter=229 channel=26
    -1, 8, 16, 5, 21, 14, -1, -4, -7,
    -- filter=229 channel=27
    18, -15, -26, -9, -13, -4, -11, 33, 23,
    -- filter=229 channel=28
    5, 3, -1, -1, -5, -1, 5, 1, -2,
    -- filter=229 channel=29
    15, -22, -13, -12, -19, 13, -5, 13, 23,
    -- filter=229 channel=30
    -8, -8, -5, 3, 7, 8, -2, 8, -2,
    -- filter=229 channel=31
    14, -4, -1, 0, -7, -10, -21, 5, 2,
    -- filter=229 channel=32
    3, -9, -19, 0, -18, 0, -9, 13, 34,
    -- filter=229 channel=33
    -7, -8, -21, 7, -13, -22, -4, 12, 14,
    -- filter=229 channel=34
    3, -4, -2, 3, 2, -8, 2, 24, -5,
    -- filter=229 channel=35
    2, 2, 1, -3, -4, -5, 1, 4, -2,
    -- filter=229 channel=36
    3, -1, 5, 0, -2, 7, 1, 5, -9,
    -- filter=229 channel=37
    -14, -1, 2, -1, 13, 1, 2, 4, -18,
    -- filter=229 channel=38
    9, 6, -11, 3, -3, -16, 0, 8, 1,
    -- filter=229 channel=39
    0, -5, 2, -9, -8, 3, 0, 1, 20,
    -- filter=229 channel=40
    6, 1, 0, -8, -15, -3, -5, 5, 12,
    -- filter=229 channel=41
    -13, 24, -17, 2, 21, -18, 3, -4, 12,
    -- filter=229 channel=42
    -3, -6, 5, -10, 0, 12, -10, -7, -7,
    -- filter=229 channel=43
    -9, 3, -4, -4, -6, -6, 6, 7, 15,
    -- filter=229 channel=44
    0, 5, 7, 0, 8, 2, -10, 0, -6,
    -- filter=229 channel=45
    5, 3, 0, -8, 1, 5, -6, -1, 4,
    -- filter=229 channel=46
    -7, 4, -2, 6, 3, 5, 0, 5, 0,
    -- filter=229 channel=47
    3, 25, 11, 14, 9, 0, -16, -23, -9,
    -- filter=229 channel=48
    2, -5, -8, -6, 0, 10, -7, 5, 5,
    -- filter=229 channel=49
    2, -12, -1, -17, 8, 15, 0, 7, 21,
    -- filter=229 channel=50
    3, -16, -4, 0, 0, 1, -8, 5, 9,
    -- filter=229 channel=51
    -2, -2, -7, -3, -6, -4, -3, -4, -1,
    -- filter=229 channel=52
    5, -15, 3, -6, -1, 4, 7, 17, 0,
    -- filter=229 channel=53
    4, -13, -10, -1, -1, 5, -1, 10, 16,
    -- filter=229 channel=54
    0, 5, 5, -3, -7, -6, -5, 0, 1,
    -- filter=229 channel=55
    7, -12, -22, -12, -22, -3, -15, 19, 38,
    -- filter=229 channel=56
    6, 3, -3, -5, 4, 1, 5, 11, 3,
    -- filter=229 channel=57
    0, 0, -1, -10, -1, 0, 7, 0, -1,
    -- filter=229 channel=58
    -4, 2, 3, 6, 12, 6, 2, -1, -6,
    -- filter=229 channel=59
    0, 1, -8, 4, 3, 0, -5, -4, 5,
    -- filter=229 channel=60
    -4, -5, 2, 0, -1, 1, -6, 3, -4,
    -- filter=229 channel=61
    -2, 4, -4, -5, 9, -2, 7, -2, -1,
    -- filter=229 channel=62
    -6, 0, 5, -5, -3, 1, 5, 8, -3,
    -- filter=229 channel=63
    -7, 13, 16, 7, 2, 4, 1, -4, -14,
    -- filter=229 channel=64
    -5, 2, -4, -7, 3, -3, -1, 0, 1,
    -- filter=229 channel=65
    3, 0, 5, -5, -7, -5, 0, -7, 6,
    -- filter=229 channel=66
    -1, 18, 0, 7, -2, -9, -1, -2, -4,
    -- filter=229 channel=67
    2, 2, -3, -3, 3, -4, -2, -5, -6,
    -- filter=229 channel=68
    6, -7, -4, -7, -1, 9, 0, 7, 8,
    -- filter=229 channel=69
    -2, -1, 0, 10, 8, 1, -4, -9, -5,
    -- filter=229 channel=70
    0, -22, -7, -12, -10, -11, -9, 10, 6,
    -- filter=229 channel=71
    -3, 7, -1, -2, -5, -13, 3, -9, -3,
    -- filter=229 channel=72
    16, 6, -16, 4, -14, -6, -10, -5, 13,
    -- filter=229 channel=73
    14, -12, -15, -10, -7, 7, -8, 21, 23,
    -- filter=229 channel=74
    -1, -19, -11, -5, 11, 8, 2, 24, 2,
    -- filter=229 channel=75
    -16, 10, -3, 11, 2, -23, 0, -18, -6,
    -- filter=229 channel=76
    14, -5, -9, -8, -25, 1, -11, 12, 31,
    -- filter=229 channel=77
    6, 2, 5, 5, 3, -5, -3, -3, -4,
    -- filter=229 channel=78
    5, 10, 11, -5, -2, 11, -2, 6, -3,
    -- filter=229 channel=79
    -3, -9, -28, -10, -25, -6, -13, 21, 40,
    -- filter=229 channel=80
    10, 12, -8, 13, 4, -12, -17, -8, -2,
    -- filter=229 channel=81
    -4, -2, 1, 0, -6, -5, 7, 3, -2,
    -- filter=229 channel=82
    0, 4, -1, 4, -1, -10, 0, 1, 1,
    -- filter=229 channel=83
    7, -10, -4, -8, 2, 2, -2, 4, 9,
    -- filter=229 channel=84
    9, -12, -10, -8, -2, 5, 5, 20, 19,
    -- filter=229 channel=85
    5, -5, 2, -3, -6, -4, 1, -3, 0,
    -- filter=229 channel=86
    -2, 0, 5, -7, 6, -7, 0, 0, -6,
    -- filter=229 channel=87
    4, -8, 3, -11, -7, 0, -5, 5, 17,
    -- filter=229 channel=88
    1, -6, 7, 1, 1, 10, 0, 0, -13,
    -- filter=229 channel=89
    3, -1, -21, 1, -30, -17, -17, 9, 29,
    -- filter=229 channel=90
    3, -2, 15, 0, -5, 0, 0, -2, -13,
    -- filter=229 channel=91
    14, -26, -7, -9, 0, 2, -2, 18, 28,
    -- filter=229 channel=92
    -4, 0, 2, -11, -2, 0, -5, -3, 0,
    -- filter=229 channel=93
    -10, 10, 10, -4, 20, 13, -11, 2, -9,
    -- filter=229 channel=94
    -5, 0, 6, 2, -5, -2, -1, 4, 1,
    -- filter=229 channel=95
    3, 7, -2, 1, -1, 4, -2, 0, 6,
    -- filter=229 channel=96
    0, -2, 1, -5, -3, -2, 1, -8, 3,
    -- filter=229 channel=97
    -3, 3, 8, -4, 0, -12, 2, 0, -3,
    -- filter=229 channel=98
    10, 0, -17, 9, -14, -4, -16, 8, 6,
    -- filter=229 channel=99
    17, -18, -8, -4, -12, -4, -11, 29, 9,
    -- filter=229 channel=100
    -3, 0, -5, -1, 4, 4, -2, -2, 1,
    -- filter=229 channel=101
    5, -4, 6, -8, 17, 13, 10, 18, 7,
    -- filter=229 channel=102
    -5, -5, 6, -6, -5, 5, -5, -1, -7,
    -- filter=229 channel=103
    -3, 12, -1, 7, 5, -7, -15, -22, -15,
    -- filter=229 channel=104
    14, 6, 0, 11, 10, 6, -17, -6, -4,
    -- filter=229 channel=105
    9, -6, 0, -14, -14, 1, -9, 14, 14,
    -- filter=229 channel=106
    -3, -2, -8, 2, -8, -1, -2, 2, 5,
    -- filter=229 channel=107
    2, -23, -9, -16, -20, 7, 2, 17, 22,
    -- filter=229 channel=108
    -10, 7, -5, 10, 12, 1, 3, -8, 8,
    -- filter=229 channel=109
    21, -16, -25, -7, -1, 8, -3, 17, 20,
    -- filter=229 channel=110
    10, -5, 5, -6, -2, -2, -4, -2, 0,
    -- filter=229 channel=111
    1, 2, 4, -1, 0, 1, 7, 6, 2,
    -- filter=229 channel=112
    6, -14, -6, -1, 3, 1, 5, 6, 5,
    -- filter=229 channel=113
    -5, 5, -7, 0, -15, -21, -7, 7, 0,
    -- filter=229 channel=114
    6, -21, -27, -16, -14, 8, 3, 29, 34,
    -- filter=229 channel=115
    -5, -4, -1, 0, 1, 3, 1, -5, 5,
    -- filter=229 channel=116
    2, -11, -16, -2, 4, 5, -10, 6, 26,
    -- filter=229 channel=117
    9, 2, -2, -5, -1, -4, 2, -7, 7,
    -- filter=229 channel=118
    -3, -7, -2, -1, -5, 8, 5, -5, 1,
    -- filter=229 channel=119
    1, -1, 6, -3, 9, -9, 7, 9, -11,
    -- filter=229 channel=120
    23, -27, -18, -7, -7, 18, -6, 43, 28,
    -- filter=229 channel=121
    4, 11, -5, 2, -2, -11, 0, -9, 1,
    -- filter=229 channel=122
    4, 37, 20, 11, 21, 2, -19, -28, -38,
    -- filter=229 channel=123
    -4, -6, 0, 1, -1, -8, 1, 6, -1,
    -- filter=229 channel=124
    3, -3, -3, 0, -6, 1, -1, 12, 13,
    -- filter=229 channel=125
    9, 1, -15, 4, -2, 8, -8, 9, 13,
    -- filter=229 channel=126
    0, 16, -5, 6, -6, -19, -3, -1, 13,
    -- filter=229 channel=127
    -6, 9, -5, 6, 5, 0, 0, 4, 0,
    -- filter=230 channel=0
    -4, 9, -6, -20, 13, -1, -9, 13, 12,
    -- filter=230 channel=1
    -7, 14, -9, -10, 20, 14, -6, 5, 3,
    -- filter=230 channel=2
    -9, 6, 5, 7, 4, 5, 2, -7, -3,
    -- filter=230 channel=3
    -1, -11, 4, -1, 2, -5, 0, 3, 0,
    -- filter=230 channel=4
    -6, 2, 0, -8, 1, 8, 6, 2, 13,
    -- filter=230 channel=5
    -6, 14, -9, -1, 24, -1, -2, 4, -2,
    -- filter=230 channel=6
    3, -3, 3, 0, 7, 7, -4, 7, 4,
    -- filter=230 channel=7
    -3, -5, 3, 5, 6, -4, -6, 7, -7,
    -- filter=230 channel=8
    -1, -10, -6, 5, 4, -7, -5, 0, -5,
    -- filter=230 channel=9
    -2, 6, -4, 3, 3, -6, -3, 7, -7,
    -- filter=230 channel=10
    7, -8, 0, 1, 4, 0, -2, 1, 3,
    -- filter=230 channel=11
    1, 3, 10, 4, -3, 5, 4, 1, 4,
    -- filter=230 channel=12
    -1, 0, 2, 1, 1, -2, 8, 4, 0,
    -- filter=230 channel=13
    0, -2, 0, -8, 8, 2, 2, 1, 4,
    -- filter=230 channel=14
    -2, 0, 2, 6, -3, -6, 5, 0, -5,
    -- filter=230 channel=15
    1, 2, -6, -1, 10, -13, 6, 2, 3,
    -- filter=230 channel=16
    0, 0, -6, 3, 10, -9, -5, 9, 2,
    -- filter=230 channel=17
    -2, -7, 7, 4, 0, 6, -5, -6, 0,
    -- filter=230 channel=18
    6, 4, -11, 0, 9, 2, -8, 5, -1,
    -- filter=230 channel=19
    -1, -3, -5, 3, -6, -5, -5, 6, 0,
    -- filter=230 channel=20
    11, 9, 11, 8, 7, -5, 12, 0, 1,
    -- filter=230 channel=21
    -2, -2, -8, -8, 12, -9, 3, -4, -6,
    -- filter=230 channel=22
    3, -4, 0, 4, 3, -12, 4, 11, 3,
    -- filter=230 channel=23
    14, -12, -10, 1, 12, -25, -2, 6, -2,
    -- filter=230 channel=24
    5, 4, -3, 7, 0, 0, -3, -1, 5,
    -- filter=230 channel=25
    -2, 1, -18, -14, 10, -6, 0, 5, -6,
    -- filter=230 channel=26
    -2, 3, 3, -4, 11, 1, 2, 1, -5,
    -- filter=230 channel=27
    0, -8, -21, -1, 17, -21, 0, 2, -5,
    -- filter=230 channel=28
    -5, -3, 5, 1, -4, -5, -2, -7, -4,
    -- filter=230 channel=29
    8, -2, 6, -1, 0, -2, 8, 2, 4,
    -- filter=230 channel=30
    5, 5, 0, -8, 11, 2, -10, 0, 5,
    -- filter=230 channel=31
    6, 0, -15, -5, 3, -20, -7, 2, -8,
    -- filter=230 channel=32
    9, 5, -10, -12, 7, -1, 0, 4, 2,
    -- filter=230 channel=33
    -2, -5, -14, -4, 0, -8, 1, 3, -4,
    -- filter=230 channel=34
    12, -5, 13, 2, 16, -3, 3, 8, 0,
    -- filter=230 channel=35
    2, 1, -5, -7, -3, 3, -6, -1, 1,
    -- filter=230 channel=36
    7, 5, -1, 0, -3, -1, 7, 0, 5,
    -- filter=230 channel=37
    -14, 14, 0, -13, 13, 9, -13, 12, 3,
    -- filter=230 channel=38
    11, 4, -13, -3, 6, -2, -1, 6, 3,
    -- filter=230 channel=39
    5, 2, 0, 0, -1, -6, 7, -8, -2,
    -- filter=230 channel=40
    10, 6, -1, 3, 2, -3, 5, 2, -6,
    -- filter=230 channel=41
    -9, 10, 1, -9, 2, 32, 0, -8, 15,
    -- filter=230 channel=42
    0, 0, 4, 1, 8, 12, -8, -7, 7,
    -- filter=230 channel=43
    7, -9, 3, -6, -3, -4, -7, 3, 4,
    -- filter=230 channel=44
    -2, 0, -1, -11, 13, -11, -10, 2, 2,
    -- filter=230 channel=45
    2, 0, -3, -5, -3, -1, -6, 7, -1,
    -- filter=230 channel=46
    1, -4, 6, 2, 0, -1, 5, 7, 5,
    -- filter=230 channel=47
    5, 11, -6, -5, 9, -9, -6, 1, -6,
    -- filter=230 channel=48
    0, 8, -5, -4, 4, 1, -10, 9, -1,
    -- filter=230 channel=49
    -1, 3, -4, 2, 0, -6, 0, 2, 7,
    -- filter=230 channel=50
    0, -8, -10, -1, -1, -13, -3, -4, -7,
    -- filter=230 channel=51
    -5, 3, 0, -4, 5, -5, 0, -2, 0,
    -- filter=230 channel=52
    10, 4, -3, 3, 2, -3, 6, 2, -4,
    -- filter=230 channel=53
    -2, -1, 3, 2, 7, -7, -4, 3, 2,
    -- filter=230 channel=54
    -5, 0, -7, -4, 1, 6, 4, -2, 0,
    -- filter=230 channel=55
    6, 3, 0, 2, -1, -8, 0, -2, -5,
    -- filter=230 channel=56
    -1, 3, -6, 0, 9, -6, 1, 0, -5,
    -- filter=230 channel=57
    -8, 5, 4, 1, 5, 11, 6, -4, 7,
    -- filter=230 channel=58
    0, 13, 5, -10, 13, 0, -4, -3, 0,
    -- filter=230 channel=59
    5, -1, -10, 2, -1, -9, -7, -2, 3,
    -- filter=230 channel=60
    5, 6, -5, -1, 0, 0, -4, 3, 0,
    -- filter=230 channel=61
    3, 8, 0, -2, 7, 4, 3, 1, 2,
    -- filter=230 channel=62
    -2, 3, -3, 6, 5, -4, 0, -4, 4,
    -- filter=230 channel=63
    -3, 13, 2, -5, 1, 9, 1, 0, 2,
    -- filter=230 channel=64
    6, -5, 1, 0, -2, -3, -5, -5, 7,
    -- filter=230 channel=65
    -1, -6, 4, -2, 0, -1, 6, -3, 4,
    -- filter=230 channel=66
    -3, 9, -5, 7, 6, 5, 6, 2, -1,
    -- filter=230 channel=67
    0, 5, 0, 7, 0, -7, -4, 6, 0,
    -- filter=230 channel=68
    -4, -2, 1, 3, -9, 3, 5, -3, 7,
    -- filter=230 channel=69
    -6, -2, -5, -3, 0, 5, -1, 0, -4,
    -- filter=230 channel=70
    -2, -3, -12, -7, 7, -15, -8, 1, -4,
    -- filter=230 channel=71
    2, -9, -6, 7, -1, -5, -6, -5, 6,
    -- filter=230 channel=72
    5, 0, -3, 1, -5, -15, -1, 6, -8,
    -- filter=230 channel=73
    0, -5, -8, -6, -7, 0, -9, -5, 0,
    -- filter=230 channel=74
    7, -12, -8, -4, 2, -11, -6, 3, 0,
    -- filter=230 channel=75
    -6, 7, -7, -19, 27, 6, -5, 15, 15,
    -- filter=230 channel=76
    3, 12, 11, 12, -5, -3, 10, -7, 0,
    -- filter=230 channel=77
    -6, 6, -2, 0, -4, -3, 0, -6, -6,
    -- filter=230 channel=78
    3, 6, -3, 1, -1, 5, 4, 6, 7,
    -- filter=230 channel=79
    -2, 9, -21, -8, 8, -14, -8, 2, 10,
    -- filter=230 channel=80
    -1, -1, -17, -2, 4, -10, -2, 5, 7,
    -- filter=230 channel=81
    4, 4, -1, -1, 2, 0, 2, 5, 5,
    -- filter=230 channel=82
    2, -7, 0, 1, 3, -6, 6, 0, -2,
    -- filter=230 channel=83
    -5, 6, -10, 0, 0, -2, -3, -3, 0,
    -- filter=230 channel=84
    -2, 5, -4, -6, 2, 4, 0, 7, -2,
    -- filter=230 channel=85
    0, -5, 6, 0, -4, -4, 0, -7, -4,
    -- filter=230 channel=86
    -1, 0, -7, 4, 8, 4, -2, 8, -4,
    -- filter=230 channel=87
    9, 4, 3, 5, 5, -8, -3, -2, 3,
    -- filter=230 channel=88
    8, -9, 0, -1, 4, 2, 0, 0, -6,
    -- filter=230 channel=89
    4, -1, -11, -11, -9, 0, 2, -12, -7,
    -- filter=230 channel=90
    3, -8, -3, 2, 0, 2, 2, -1, 0,
    -- filter=230 channel=91
    0, 3, -17, -5, -2, -12, -9, 8, 0,
    -- filter=230 channel=92
    6, -2, 5, 0, 0, 0, -6, 8, 3,
    -- filter=230 channel=93
    -11, 11, -9, -12, 3, -3, -7, 1, -1,
    -- filter=230 channel=94
    -4, 0, 4, 5, -6, 0, -5, 1, -2,
    -- filter=230 channel=95
    5, 0, -3, 3, 1, 6, 6, 0, -3,
    -- filter=230 channel=96
    -2, 0, -3, 1, -1, 0, -4, -8, 2,
    -- filter=230 channel=97
    -5, -5, 6, -3, -6, 1, 4, -5, -1,
    -- filter=230 channel=98
    -2, 0, -14, -3, 14, -3, -4, -5, 5,
    -- filter=230 channel=99
    14, -1, 0, -1, 15, -16, -2, 3, 0,
    -- filter=230 channel=100
    1, -4, 10, 1, -2, -2, 3, 8, -1,
    -- filter=230 channel=101
    -11, -5, -5, 1, 0, 8, 1, -7, -2,
    -- filter=230 channel=102
    -2, 0, -7, 4, 4, 2, -3, -4, 1,
    -- filter=230 channel=103
    6, 4, -13, -7, 10, -2, -11, 5, -6,
    -- filter=230 channel=104
    5, -5, -8, -8, 4, -14, 2, -1, -3,
    -- filter=230 channel=105
    1, 0, 3, 2, 2, 4, 1, 4, -3,
    -- filter=230 channel=106
    -2, -3, -2, 4, 1, 4, -2, -4, -4,
    -- filter=230 channel=107
    10, 0, 0, -1, 1, 0, -1, -4, -7,
    -- filter=230 channel=108
    2, 11, 1, -6, 10, 9, 5, -4, 3,
    -- filter=230 channel=109
    0, -6, -18, -2, 15, -22, 3, 5, -6,
    -- filter=230 channel=110
    8, 2, -2, 0, 5, -7, 0, 3, -4,
    -- filter=230 channel=111
    -6, -2, -7, -6, 4, -3, 0, -1, 0,
    -- filter=230 channel=112
    -1, 2, -9, -4, 10, -15, -4, 2, 0,
    -- filter=230 channel=113
    8, -10, -13, -2, 3, -14, -6, 10, 0,
    -- filter=230 channel=114
    -2, 18, -20, -14, 19, -5, -5, 2, -5,
    -- filter=230 channel=115
    1, -3, -1, -1, -5, -3, -4, 7, -3,
    -- filter=230 channel=116
    0, -4, -15, 0, 5, 4, -4, -6, 0,
    -- filter=230 channel=117
    1, 3, -4, 5, -4, -2, 4, -5, -1,
    -- filter=230 channel=118
    -5, 0, -4, -6, -4, 6, -4, -7, -5,
    -- filter=230 channel=119
    4, 5, 7, 7, 7, 1, 4, 9, -5,
    -- filter=230 channel=120
    7, -10, -18, -5, 7, -26, -9, 10, -9,
    -- filter=230 channel=121
    8, -2, 1, -3, -6, 0, -1, -6, 0,
    -- filter=230 channel=122
    -6, 1, -4, -10, 15, -11, -10, 11, -4,
    -- filter=230 channel=123
    8, -2, -3, 7, 10, -4, -8, 5, -3,
    -- filter=230 channel=124
    7, 5, 2, 4, -3, 0, 2, 4, 4,
    -- filter=230 channel=125
    9, -4, -18, 0, 1, -4, -5, 11, -1,
    -- filter=230 channel=126
    -2, 11, -6, -1, -5, 4, 4, 2, -4,
    -- filter=230 channel=127
    2, 4, 4, 0, 0, 3, -4, -6, 0,
    -- filter=231 channel=0
    -11, -11, -4, -2, 0, -8, 4, 9, -2,
    -- filter=231 channel=1
    -8, -7, -13, 3, 0, -7, -1, 7, -5,
    -- filter=231 channel=2
    -2, 3, -2, 4, 0, -3, 4, -2, -7,
    -- filter=231 channel=3
    -11, -1, -7, 2, -3, 6, 8, 1, 3,
    -- filter=231 channel=4
    -2, -4, 3, -1, 6, 6, -4, 0, 0,
    -- filter=231 channel=5
    1, -4, -1, 0, -2, -9, 9, 10, -4,
    -- filter=231 channel=6
    0, 0, -6, -1, 1, -3, 0, -4, 4,
    -- filter=231 channel=7
    0, 0, 3, -3, -4, 4, 6, -4, 3,
    -- filter=231 channel=8
    4, -3, 2, 0, 3, -3, -2, -4, -2,
    -- filter=231 channel=9
    -6, -5, 3, 0, 9, 6, 1, 8, 2,
    -- filter=231 channel=10
    -4, 0, 5, 0, 9, 9, 9, 8, 5,
    -- filter=231 channel=11
    0, 2, 9, -3, 11, 1, -3, -5, 5,
    -- filter=231 channel=12
    0, -5, 0, 5, -7, 3, 1, 6, -6,
    -- filter=231 channel=13
    -7, -3, -4, 5, -2, 11, 3, 0, -3,
    -- filter=231 channel=14
    -4, -2, 3, 0, 2, 4, 4, 5, -7,
    -- filter=231 channel=15
    -12, -3, -8, 9, 9, 6, 4, 4, 5,
    -- filter=231 channel=16
    0, 7, -4, 3, 8, -4, -1, 0, -6,
    -- filter=231 channel=17
    -1, 7, -6, -1, 0, -2, 1, 3, -2,
    -- filter=231 channel=18
    -12, -11, -9, 15, 10, 2, 7, 3, 0,
    -- filter=231 channel=19
    3, 1, -4, -5, -6, -4, 1, 4, -4,
    -- filter=231 channel=20
    -3, 11, 9, -2, 10, 0, -8, -8, -4,
    -- filter=231 channel=21
    -3, 7, 1, -7, 15, 8, 0, 6, 0,
    -- filter=231 channel=22
    -8, -6, -11, 4, -9, -5, -1, 0, -7,
    -- filter=231 channel=23
    -13, -11, 1, 6, 5, -7, 10, -2, -11,
    -- filter=231 channel=24
    -5, -1, 6, -5, 1, 5, 0, 2, -5,
    -- filter=231 channel=25
    -8, -3, -10, 12, 17, -1, 11, 3, -3,
    -- filter=231 channel=26
    5, 6, -3, 2, -3, 0, 0, -1, 0,
    -- filter=231 channel=27
    0, -11, -5, 16, 10, -2, 11, -16, -20,
    -- filter=231 channel=28
    0, 4, -1, 1, -1, 6, -3, 7, -2,
    -- filter=231 channel=29
    -6, 8, 5, 7, 1, -1, -7, 1, 4,
    -- filter=231 channel=30
    -9, -7, 0, 2, 5, -6, -2, 1, -10,
    -- filter=231 channel=31
    -9, 6, -2, 8, 11, -10, -5, -9, -19,
    -- filter=231 channel=32
    -2, -15, -9, 16, 3, 5, 7, 0, -11,
    -- filter=231 channel=33
    -14, -10, -7, 1, 7, 1, 12, -1, -4,
    -- filter=231 channel=34
    2, -14, -8, -8, -14, -1, -2, -3, 4,
    -- filter=231 channel=35
    0, 1, 5, -6, -4, 0, -3, 1, 0,
    -- filter=231 channel=36
    -2, 5, 0, -3, 3, 6, -13, -14, -2,
    -- filter=231 channel=37
    -1, 0, -15, -5, 2, -11, -8, -2, -8,
    -- filter=231 channel=38
    -1, -9, 0, 3, -3, 4, 7, 6, -8,
    -- filter=231 channel=39
    3, 0, -3, 5, 0, -1, 2, 1, -6,
    -- filter=231 channel=40
    -8, 3, 7, 0, -1, 0, 2, -4, -2,
    -- filter=231 channel=41
    6, -5, -7, 1, 1, -7, 13, 3, 10,
    -- filter=231 channel=42
    0, -4, 0, 5, 4, 6, 6, 2, 2,
    -- filter=231 channel=43
    -3, -3, 1, -4, -7, 0, 4, 9, 1,
    -- filter=231 channel=44
    4, 3, 3, -3, 4, -10, -3, 0, -7,
    -- filter=231 channel=45
    -7, -3, 0, -5, 0, -5, -4, 1, -3,
    -- filter=231 channel=46
    3, -2, 4, 0, 1, 4, 7, -6, 2,
    -- filter=231 channel=47
    1, 8, -4, -4, 9, -2, 12, 16, -3,
    -- filter=231 channel=48
    -7, 6, 3, 6, 19, 9, 2, -4, -16,
    -- filter=231 channel=49
    0, -8, -5, 6, 3, -3, -7, -9, -1,
    -- filter=231 channel=50
    -6, -6, -5, 0, 4, -4, 5, -5, -10,
    -- filter=231 channel=51
    -6, -1, 1, -1, 5, 6, 2, 2, 4,
    -- filter=231 channel=52
    -6, -8, 3, -6, 0, -5, 3, 0, -10,
    -- filter=231 channel=53
    5, 4, 9, -1, 5, -1, 0, -2, -7,
    -- filter=231 channel=54
    -1, -3, -6, -6, 2, 0, 5, 1, -3,
    -- filter=231 channel=55
    2, 4, -1, 1, 11, 3, 14, 4, -4,
    -- filter=231 channel=56
    0, -1, -2, 7, 1, -9, -1, 0, -6,
    -- filter=231 channel=57
    -3, 6, -5, 1, 1, -2, 5, 4, 6,
    -- filter=231 channel=58
    1, 4, -1, -4, -2, 6, -5, 12, -3,
    -- filter=231 channel=59
    -9, 0, 0, 15, 15, 1, 13, 5, -8,
    -- filter=231 channel=60
    -2, -7, 6, -1, -3, -6, -5, 6, -2,
    -- filter=231 channel=61
    1, 5, 4, 4, 5, 2, 0, -2, -2,
    -- filter=231 channel=62
    3, 1, -2, -4, -5, 6, 7, -1, 5,
    -- filter=231 channel=63
    2, 0, -5, -1, 0, -6, -2, 9, 3,
    -- filter=231 channel=64
    5, 0, 7, -9, 6, -1, 0, 0, -2,
    -- filter=231 channel=65
    -2, -1, -4, 6, -5, -4, 3, -5, 3,
    -- filter=231 channel=66
    0, -10, -5, 2, -8, 0, 3, -2, 0,
    -- filter=231 channel=67
    4, -5, -8, 1, 0, 5, -3, 5, -5,
    -- filter=231 channel=68
    4, 4, 3, 0, 5, -6, 4, 1, -8,
    -- filter=231 channel=69
    2, 1, 3, 2, 3, -2, 1, 3, 1,
    -- filter=231 channel=70
    -9, -11, -11, 4, 4, -11, 1, -10, -10,
    -- filter=231 channel=71
    -12, -2, 2, -11, 1, 0, 4, 0, 7,
    -- filter=231 channel=72
    3, 5, 5, 13, 16, 8, -2, -8, -5,
    -- filter=231 channel=73
    2, -5, -8, 14, 6, 8, 5, -12, -15,
    -- filter=231 channel=74
    0, 0, -10, 11, -7, -1, 2, -13, -14,
    -- filter=231 channel=75
    -14, -16, -6, 4, -4, 1, 7, 21, 7,
    -- filter=231 channel=76
    2, 0, 3, 5, 0, 9, 6, -3, -2,
    -- filter=231 channel=77
    1, -1, -1, -4, 3, -1, -1, 0, -5,
    -- filter=231 channel=78
    -7, 7, -6, 8, 0, 0, -5, 10, -2,
    -- filter=231 channel=79
    -10, -16, -4, 15, 0, -6, 11, -7, -4,
    -- filter=231 channel=80
    0, 0, -3, 9, 15, 10, 15, 1, -10,
    -- filter=231 channel=81
    -3, -6, 6, 7, 4, 4, -4, -3, -2,
    -- filter=231 channel=82
    -10, -7, -8, 0, -7, 0, 4, 4, 4,
    -- filter=231 channel=83
    -4, 0, 2, 0, 11, -2, 2, -9, -12,
    -- filter=231 channel=84
    6, 3, -4, 13, 12, 5, -8, -1, -14,
    -- filter=231 channel=85
    -5, 6, -5, -6, -3, -1, -5, 2, -3,
    -- filter=231 channel=86
    0, -9, -2, -4, -6, -5, -3, 4, 2,
    -- filter=231 channel=87
    4, -6, 1, -3, 2, -6, 3, 6, 0,
    -- filter=231 channel=88
    -3, 5, 0, -3, 5, -2, -12, -6, -2,
    -- filter=231 channel=89
    -5, -9, -1, 4, 8, 12, 8, 3, -10,
    -- filter=231 channel=90
    -1, 0, 0, -6, -1, -10, -11, 0, -7,
    -- filter=231 channel=91
    -3, -9, -4, 12, 5, 0, -2, -7, -19,
    -- filter=231 channel=92
    3, 0, -5, 3, -4, -3, 2, -7, 5,
    -- filter=231 channel=93
    -7, -3, 0, 11, 3, 3, -4, 7, -2,
    -- filter=231 channel=94
    1, -7, -7, -1, 4, 5, 2, -3, 3,
    -- filter=231 channel=95
    -4, 4, -5, 0, -6, 0, 5, 0, 0,
    -- filter=231 channel=96
    6, -5, 0, -7, -4, 3, 6, 5, -5,
    -- filter=231 channel=97
    -12, -12, -7, 2, -9, 1, 3, 0, 6,
    -- filter=231 channel=98
    -4, -4, -1, 15, 19, 0, 12, 0, -12,
    -- filter=231 channel=99
    -1, -1, 6, 12, 15, 1, 7, -10, -21,
    -- filter=231 channel=100
    2, 4, 2, -2, -6, -3, 4, -3, -1,
    -- filter=231 channel=101
    2, -5, 5, -3, 6, -4, -3, 0, -5,
    -- filter=231 channel=102
    -6, 7, -6, 0, -4, -2, 2, 1, -6,
    -- filter=231 channel=103
    -8, -8, -9, -9, 10, 2, 2, 15, -6,
    -- filter=231 channel=104
    1, 3, 6, 3, 12, -3, -6, 3, -17,
    -- filter=231 channel=105
    4, 7, 9, -2, 0, 9, 2, 2, 7,
    -- filter=231 channel=106
    -2, -5, 0, -6, -2, 4, 1, -5, 7,
    -- filter=231 channel=107
    -1, 1, -4, -3, -3, -2, 1, -1, 2,
    -- filter=231 channel=108
    -6, 2, -1, -4, 3, 1, 5, 0, 0,
    -- filter=231 channel=109
    -3, -5, -5, 19, 18, 9, 14, -11, -11,
    -- filter=231 channel=110
    -7, 0, 2, 0, -2, 0, 2, -3, 1,
    -- filter=231 channel=111
    -3, 1, -5, -2, -8, -3, -5, 3, -3,
    -- filter=231 channel=112
    0, -8, -7, 0, -1, -11, 0, 1, -4,
    -- filter=231 channel=113
    -13, -11, -3, 2, -2, 5, 11, 12, 1,
    -- filter=231 channel=114
    -7, -12, -15, 13, 0, -5, 2, -5, -19,
    -- filter=231 channel=115
    2, 1, 6, 4, 5, 3, -2, 4, 1,
    -- filter=231 channel=116
    -5, -2, 6, 12, 19, 12, -2, -3, -8,
    -- filter=231 channel=117
    4, 1, 2, 4, -3, -1, 0, -2, 0,
    -- filter=231 channel=118
    -3, -6, 6, 0, 5, 1, -6, -2, 0,
    -- filter=231 channel=119
    0, 0, -9, 7, -3, -13, -1, 2, -11,
    -- filter=231 channel=120
    -1, -2, -2, 17, 14, -5, -1, -6, -19,
    -- filter=231 channel=121
    -2, -11, 2, 6, -2, -4, 1, 1, -2,
    -- filter=231 channel=122
    -3, 0, 3, -3, 15, 0, 0, 6, -9,
    -- filter=231 channel=123
    0, 0, 3, 1, 2, -8, 4, 0, 6,
    -- filter=231 channel=124
    0, 5, 2, 3, 3, 0, -2, 0, 8,
    -- filter=231 channel=125
    -2, 0, -5, 20, 19, 5, -1, -11, -19,
    -- filter=231 channel=126
    -10, -11, -6, 6, 1, 3, 20, 17, 13,
    -- filter=231 channel=127
    -2, -6, 4, 3, -6, -5, -3, -6, 0,
    -- filter=232 channel=0
    4, 1, 0, 6, 4, 6, 1, 0, -1,
    -- filter=232 channel=1
    -1, -6, 7, 0, -1, -2, 5, -3, 2,
    -- filter=232 channel=2
    -6, -6, -6, 0, -5, -6, -2, 6, 6,
    -- filter=232 channel=3
    -1, 4, 0, 1, 5, 7, -2, -3, 0,
    -- filter=232 channel=4
    4, 5, 8, -3, -6, 5, -6, 3, 7,
    -- filter=232 channel=5
    2, 7, -3, 5, 1, 5, 0, -5, 5,
    -- filter=232 channel=6
    7, 1, -6, 2, -2, 3, -2, 0, 6,
    -- filter=232 channel=7
    4, 0, -6, 6, 1, -6, 4, 5, -4,
    -- filter=232 channel=8
    0, -3, 2, -4, 2, 3, -3, 5, -2,
    -- filter=232 channel=9
    0, 3, 0, 5, 5, -4, -2, 5, 0,
    -- filter=232 channel=10
    5, -3, 2, 0, -8, -5, 0, -8, 0,
    -- filter=232 channel=11
    8, -2, 4, 3, 1, 0, 3, -3, 6,
    -- filter=232 channel=12
    0, -4, 5, -3, 1, 4, 0, -3, -4,
    -- filter=232 channel=13
    0, -3, -9, 5, -4, 3, -9, 2, -1,
    -- filter=232 channel=14
    -6, -7, -6, 0, -5, 4, -1, -4, 5,
    -- filter=232 channel=15
    3, -1, -1, 1, -7, 2, -3, 2, 5,
    -- filter=232 channel=16
    4, 6, 3, -3, -4, 6, 1, 7, -4,
    -- filter=232 channel=17
    4, 3, 7, -6, -3, -4, 6, 6, -7,
    -- filter=232 channel=18
    -5, 0, -9, 4, -5, -4, -4, 0, 3,
    -- filter=232 channel=19
    -4, -3, 0, -5, 2, -5, 7, -2, 1,
    -- filter=232 channel=20
    0, -2, 5, 11, 5, 6, 6, 1, -3,
    -- filter=232 channel=21
    2, -3, 5, 4, 0, -5, -4, 2, 0,
    -- filter=232 channel=22
    -5, -1, -3, 4, 0, 6, 2, 1, 9,
    -- filter=232 channel=23
    0, -4, 5, -1, 0, 0, 4, -4, 3,
    -- filter=232 channel=24
    -7, -1, -4, 4, -4, -7, 4, 0, 1,
    -- filter=232 channel=25
    -3, 3, 4, -1, -7, -4, -1, -5, -2,
    -- filter=232 channel=26
    -5, 0, -3, 3, 7, 1, -5, 3, 2,
    -- filter=232 channel=27
    -5, -3, -2, -15, -10, 6, -14, -5, -5,
    -- filter=232 channel=28
    -1, 7, 6, 0, -6, 2, -6, -1, -3,
    -- filter=232 channel=29
    1, 0, 0, 9, 7, 1, -3, 0, -5,
    -- filter=232 channel=30
    2, -6, 8, -7, -7, 8, -9, 5, -5,
    -- filter=232 channel=31
    3, -6, 3, -9, -4, 3, -8, -7, 0,
    -- filter=232 channel=32
    3, -8, 5, -6, -9, 2, 3, 0, 0,
    -- filter=232 channel=33
    1, 1, -4, -6, 0, -1, -9, -9, 0,
    -- filter=232 channel=34
    -6, -1, 4, -8, 7, 5, 4, 2, 1,
    -- filter=232 channel=35
    -3, 5, 3, 4, 2, 1, 4, 1, -5,
    -- filter=232 channel=36
    5, 5, -1, 1, -4, -4, 6, 6, -6,
    -- filter=232 channel=37
    5, -7, 10, 7, 0, 2, 4, 3, 5,
    -- filter=232 channel=38
    -4, -3, -5, -3, 5, 0, 4, -8, -1,
    -- filter=232 channel=39
    2, 6, -4, 0, 4, 5, 0, 7, 7,
    -- filter=232 channel=40
    -2, 1, 3, 7, 2, -4, -2, 7, -4,
    -- filter=232 channel=41
    -2, -9, -6, 4, 1, 4, 2, -10, -3,
    -- filter=232 channel=42
    -7, 6, 3, 6, -2, -7, 0, -7, -6,
    -- filter=232 channel=43
    -1, -1, 5, 8, -2, -2, 4, 6, -3,
    -- filter=232 channel=44
    -4, -5, -2, -9, -5, 0, -4, -2, 4,
    -- filter=232 channel=45
    5, 8, 4, -2, 8, 6, 8, 5, 5,
    -- filter=232 channel=46
    2, 0, 3, -1, -3, 4, 4, 4, -2,
    -- filter=232 channel=47
    -1, 0, -1, 2, 4, -1, 1, -4, 6,
    -- filter=232 channel=48
    -2, 2, -5, -2, -9, -4, -6, -2, -6,
    -- filter=232 channel=49
    5, -1, 5, -5, 6, 1, -6, 0, 5,
    -- filter=232 channel=50
    -1, 6, 8, -8, -5, -4, 3, -7, -1,
    -- filter=232 channel=51
    -2, 3, -3, 5, -6, 2, 5, -1, -4,
    -- filter=232 channel=52
    6, -7, 0, -3, 4, 8, -1, -1, 0,
    -- filter=232 channel=53
    -6, -5, 5, 0, 0, -3, 5, 4, -6,
    -- filter=232 channel=54
    -5, -4, 0, -7, 6, 5, 3, -6, 1,
    -- filter=232 channel=55
    -2, -2, 0, 6, -8, -7, 1, 3, -1,
    -- filter=232 channel=56
    3, -5, -4, -6, -5, 5, -8, 4, 0,
    -- filter=232 channel=57
    2, 5, 4, -2, -6, 3, 0, 1, -3,
    -- filter=232 channel=58
    -3, -3, 2, -3, -1, -3, -1, 1, -5,
    -- filter=232 channel=59
    -4, -7, -1, -4, 0, 0, -7, -10, 3,
    -- filter=232 channel=60
    5, 4, -3, -4, -4, 1, 4, 0, -4,
    -- filter=232 channel=61
    0, 2, -3, 3, 3, -4, -5, -2, -1,
    -- filter=232 channel=62
    6, 3, -5, 4, -5, -2, -1, -4, -5,
    -- filter=232 channel=63
    2, 0, -4, 4, 0, -4, -5, 0, 6,
    -- filter=232 channel=64
    4, 5, 4, 7, 6, -2, 0, 5, 5,
    -- filter=232 channel=65
    5, -5, 1, 5, 1, 5, 0, 2, 0,
    -- filter=232 channel=66
    -5, -9, 6, 7, 0, -5, -8, 0, -5,
    -- filter=232 channel=67
    4, 0, 0, 1, -6, -1, 1, 2, 3,
    -- filter=232 channel=68
    0, 7, -1, 1, 3, 2, 4, -5, -5,
    -- filter=232 channel=69
    0, -6, -3, -5, -7, 3, -2, 6, -1,
    -- filter=232 channel=70
    -4, -8, 5, -10, -7, 4, -5, 5, 4,
    -- filter=232 channel=71
    -4, -4, 5, -1, -2, 7, 7, 0, 0,
    -- filter=232 channel=72
    0, -2, -6, -1, -7, -6, -7, 0, -8,
    -- filter=232 channel=73
    -3, -8, -6, 1, 1, 0, 0, -6, -3,
    -- filter=232 channel=74
    0, 4, 0, -10, -6, 0, 1, 2, 2,
    -- filter=232 channel=75
    -1, 3, 7, 5, 0, -1, -6, 3, 7,
    -- filter=232 channel=76
    1, 5, -1, 12, 6, -4, 11, 3, -2,
    -- filter=232 channel=77
    4, -1, 0, 6, -5, -3, -3, -5, 6,
    -- filter=232 channel=78
    5, -1, 6, 0, -5, -5, -3, 6, 5,
    -- filter=232 channel=79
    -8, -10, -6, -4, -9, 1, -10, 0, 0,
    -- filter=232 channel=80
    -2, -4, -1, 3, -6, 2, 0, 2, 2,
    -- filter=232 channel=81
    0, 1, 0, 1, -7, 0, 6, -7, 6,
    -- filter=232 channel=82
    0, 0, 1, 2, 3, 8, 2, 1, 6,
    -- filter=232 channel=83
    1, 0, 2, 6, 5, 6, 0, -6, 0,
    -- filter=232 channel=84
    1, 0, -3, 0, -8, 3, 1, 6, 0,
    -- filter=232 channel=85
    -6, 1, -1, -7, 6, -5, 1, -4, -4,
    -- filter=232 channel=86
    3, -1, 1, -7, 3, 5, 5, 5, 2,
    -- filter=232 channel=87
    -3, -1, 7, -2, -1, 7, 3, 5, 6,
    -- filter=232 channel=88
    -1, 7, 1, 7, 2, 1, 0, -3, -3,
    -- filter=232 channel=89
    -5, 1, -3, -8, -9, 2, -7, -11, 0,
    -- filter=232 channel=90
    6, 4, 2, -2, 1, 0, 0, 4, 2,
    -- filter=232 channel=91
    0, 0, 8, -4, 0, 4, -7, -9, 0,
    -- filter=232 channel=92
    -1, 0, -5, 0, 2, 3, -7, 3, 0,
    -- filter=232 channel=93
    -7, 2, -4, 1, 4, 4, -4, -1, 3,
    -- filter=232 channel=94
    -5, -5, -2, 6, -3, 6, -3, -6, -6,
    -- filter=232 channel=95
    -4, 1, 6, 0, -4, -7, -6, 4, 5,
    -- filter=232 channel=96
    3, 0, 0, -5, -5, 6, -4, -1, -3,
    -- filter=232 channel=97
    -6, 0, -3, -4, 3, -6, -2, 0, -4,
    -- filter=232 channel=98
    3, 3, 2, -6, -3, 3, -7, -2, -2,
    -- filter=232 channel=99
    -2, -4, 0, 2, -8, 7, -5, -3, 2,
    -- filter=232 channel=100
    -8, -8, -3, -4, -6, -6, 3, 1, -7,
    -- filter=232 channel=101
    -3, 5, 6, -4, 0, -6, 5, 1, -3,
    -- filter=232 channel=102
    5, -1, -5, 2, 3, 7, -5, 4, 2,
    -- filter=232 channel=103
    -1, 2, 0, -2, -7, 2, -4, -4, 3,
    -- filter=232 channel=104
    -7, -8, -6, 5, -9, 4, -1, 1, -9,
    -- filter=232 channel=105
    7, -1, 6, 5, -1, -7, -1, 0, 0,
    -- filter=232 channel=106
    -1, 1, 1, 5, 8, -7, -1, -5, 6,
    -- filter=232 channel=107
    7, 1, 4, 10, 11, 8, 10, 7, 0,
    -- filter=232 channel=108
    7, 7, -6, 0, -1, 7, 6, -7, 3,
    -- filter=232 channel=109
    -1, -1, 1, -2, -1, -5, 0, -4, -5,
    -- filter=232 channel=110
    -5, 0, -1, 0, 0, -7, -1, 4, 4,
    -- filter=232 channel=111
    6, 2, 5, -5, 7, -4, 5, -2, -1,
    -- filter=232 channel=112
    -8, 2, 1, 1, 3, 2, -2, -5, -3,
    -- filter=232 channel=113
    3, 0, -5, -1, -7, 0, -4, -3, -5,
    -- filter=232 channel=114
    -3, -6, -5, -6, 1, 5, -7, 2, 8,
    -- filter=232 channel=115
    0, -3, -3, 2, 4, 3, -3, 0, 7,
    -- filter=232 channel=116
    0, -3, -6, 3, -7, 2, -10, 0, -5,
    -- filter=232 channel=117
    3, -7, 6, 3, 3, 0, -1, -4, 5,
    -- filter=232 channel=118
    1, -2, 0, -1, -5, -4, -4, 2, 0,
    -- filter=232 channel=119
    -8, -3, -2, 1, 3, 1, -1, -1, 3,
    -- filter=232 channel=120
    -3, 3, 2, 0, 0, 6, -4, 3, 4,
    -- filter=232 channel=121
    3, 4, 4, 1, -1, 0, 1, -4, -2,
    -- filter=232 channel=122
    8, 4, 4, -7, 3, 4, 3, -6, -5,
    -- filter=232 channel=123
    0, 6, -5, 0, 0, 9, 3, -1, 8,
    -- filter=232 channel=124
    0, 3, 6, -3, -4, 7, 3, 2, 7,
    -- filter=232 channel=125
    -5, -2, -1, -5, -6, -7, -5, -8, 2,
    -- filter=232 channel=126
    -5, -1, 1, 1, -4, -4, 2, 2, 0,
    -- filter=232 channel=127
    -1, -5, 0, 2, 0, 3, 5, -1, -1,
    -- filter=233 channel=0
    -10, -10, 0, -5, -25, -18, -10, -21, -13,
    -- filter=233 channel=1
    -8, -22, -4, -19, -24, -6, -9, -20, -7,
    -- filter=233 channel=2
    -1, 2, -3, 6, 3, -5, 7, 1, 5,
    -- filter=233 channel=3
    4, 3, 6, -4, 3, 0, 3, 7, 3,
    -- filter=233 channel=4
    -6, -4, 10, -5, -3, 0, 5, -1, -2,
    -- filter=233 channel=5
    -3, 0, 7, -13, -9, 2, 0, -9, -1,
    -- filter=233 channel=6
    3, 0, 0, 8, -6, -6, 1, 4, -10,
    -- filter=233 channel=7
    -4, 0, 0, 3, -4, 5, -2, -6, 0,
    -- filter=233 channel=8
    2, 1, 0, -3, 3, -2, -7, 0, -3,
    -- filter=233 channel=9
    -8, 5, 10, -4, 9, 11, 0, 7, 0,
    -- filter=233 channel=10
    2, 3, 12, 0, -4, 12, -2, 3, 0,
    -- filter=233 channel=11
    2, 7, -1, -6, 5, 8, -1, 4, -3,
    -- filter=233 channel=12
    8, -8, 0, 8, -5, -4, 6, -1, -7,
    -- filter=233 channel=13
    0, 2, -3, 4, -6, -5, 0, 0, -9,
    -- filter=233 channel=14
    6, -4, 3, 3, -6, 2, 5, -5, 4,
    -- filter=233 channel=15
    10, 6, 1, 6, 6, -13, 6, -4, -11,
    -- filter=233 channel=16
    -1, -14, -4, -16, -14, 4, 0, -6, 8,
    -- filter=233 channel=17
    4, -3, -3, 0, 4, -4, -5, 3, 0,
    -- filter=233 channel=18
    11, 5, -6, 12, 6, -6, 13, 4, -8,
    -- filter=233 channel=19
    1, -6, 1, 3, 2, 0, 4, 5, -7,
    -- filter=233 channel=20
    4, 8, 1, -6, 4, 0, 4, 7, -4,
    -- filter=233 channel=21
    -11, -7, 5, -5, -8, 8, -7, -3, 11,
    -- filter=233 channel=22
    -4, 0, -1, 0, -1, -7, 0, 4, -9,
    -- filter=233 channel=23
    7, 13, -9, 3, 9, -7, -3, 7, -11,
    -- filter=233 channel=24
    -5, 4, -3, 6, -6, 7, 1, 5, -1,
    -- filter=233 channel=25
    0, -10, 3, -5, -1, 7, 11, 0, 1,
    -- filter=233 channel=26
    -1, -1, 6, -1, -4, 3, -4, 2, -2,
    -- filter=233 channel=27
    -6, 13, 0, 2, 3, 3, -1, 0, -10,
    -- filter=233 channel=28
    -6, 0, 3, -4, -4, -1, 7, 4, -6,
    -- filter=233 channel=29
    6, 14, -3, 8, 10, -4, 4, 7, -6,
    -- filter=233 channel=30
    -12, -1, -6, -11, 0, 6, 4, -1, -2,
    -- filter=233 channel=31
    -3, 7, -1, -12, 17, 18, -7, 7, 14,
    -- filter=233 channel=32
    0, 5, 2, -8, 7, -10, 11, -8, -6,
    -- filter=233 channel=33
    2, 8, 4, -4, 0, -8, 6, 6, -2,
    -- filter=233 channel=34
    5, 4, -3, -2, -6, -25, 2, -13, -17,
    -- filter=233 channel=35
    5, -3, -3, -2, -3, -5, 0, 2, 1,
    -- filter=233 channel=36
    1, -5, -3, -2, 5, -3, -2, -4, 1,
    -- filter=233 channel=37
    -20, -21, -9, -20, -20, -10, -14, -21, -6,
    -- filter=233 channel=38
    4, 6, 8, -3, 10, 10, 0, 9, 11,
    -- filter=233 channel=39
    -4, 5, 2, 7, 0, 1, -1, 3, -2,
    -- filter=233 channel=40
    0, -7, -3, -3, -1, 3, -6, 0, -11,
    -- filter=233 channel=41
    -4, -11, -2, 7, -13, -22, 3, -11, -10,
    -- filter=233 channel=42
    -11, 2, 0, 2, 0, 0, 3, 2, -6,
    -- filter=233 channel=43
    3, 10, -8, -3, 0, -6, -6, -3, -4,
    -- filter=233 channel=44
    -15, -6, -8, -16, -17, 0, -7, -7, 0,
    -- filter=233 channel=45
    0, 3, -1, 0, 1, 5, -1, -7, -4,
    -- filter=233 channel=46
    0, 0, -6, 0, 0, -5, 1, -6, -6,
    -- filter=233 channel=47
    -8, -21, 5, -20, -17, 12, -13, -10, 9,
    -- filter=233 channel=48
    -8, -2, 6, -5, -5, 7, 4, 5, 4,
    -- filter=233 channel=49
    4, 9, 2, 2, 15, -8, 13, 2, -1,
    -- filter=233 channel=50
    -3, 12, -5, 3, 6, 5, 1, 3, -4,
    -- filter=233 channel=51
    0, -3, -3, 1, -4, -3, -1, -6, 3,
    -- filter=233 channel=52
    -4, 1, -6, -7, -5, -13, -1, -3, -12,
    -- filter=233 channel=53
    -7, 9, -5, -3, 11, -2, 1, 7, 4,
    -- filter=233 channel=54
    1, 6, 7, -4, 2, -7, 3, -3, 1,
    -- filter=233 channel=55
    12, 13, 5, 6, 12, -4, 6, 8, -10,
    -- filter=233 channel=56
    -6, -4, -10, -5, -4, -3, -1, 2, -10,
    -- filter=233 channel=57
    -3, 0, 2, 2, -8, 0, 3, 3, -5,
    -- filter=233 channel=58
    4, 2, 1, -7, -10, -6, -9, -9, -8,
    -- filter=233 channel=59
    0, -2, 1, -5, -7, 17, 7, 5, 6,
    -- filter=233 channel=60
    5, -5, -7, 5, -5, 7, -5, -3, -2,
    -- filter=233 channel=61
    -8, -8, 0, 2, -7, 5, -4, -8, -7,
    -- filter=233 channel=62
    1, 7, -2, 0, 8, -1, 3, 0, -4,
    -- filter=233 channel=63
    1, -8, 4, 3, 2, -1, -4, 0, 4,
    -- filter=233 channel=64
    -1, 0, -7, -1, -7, 0, -3, 0, -6,
    -- filter=233 channel=65
    -4, 6, 6, -1, 1, -2, 4, 0, -7,
    -- filter=233 channel=66
    0, -11, 0, 11, -12, 0, 0, -14, 3,
    -- filter=233 channel=67
    4, 4, 3, 3, 0, 3, 6, -5, 3,
    -- filter=233 channel=68
    -4, 4, 1, 4, -5, 3, -4, 2, 0,
    -- filter=233 channel=69
    5, -3, 2, 0, -10, -4, 3, -3, 1,
    -- filter=233 channel=70
    0, 7, -12, 1, 2, -11, 0, 3, -8,
    -- filter=233 channel=71
    -4, -2, 5, 4, -5, 0, -4, -3, 7,
    -- filter=233 channel=72
    2, 4, 0, 3, 6, 6, 6, 1, 12,
    -- filter=233 channel=73
    5, 1, 3, 7, 6, 0, 7, 2, -9,
    -- filter=233 channel=74
    0, 4, -14, -9, 8, -4, 0, 7, -2,
    -- filter=233 channel=75
    -8, -15, 6, -24, -24, -4, -4, -17, 3,
    -- filter=233 channel=76
    -7, 7, -2, 5, -1, -6, 1, 3, -4,
    -- filter=233 channel=77
    4, -4, 0, 3, 5, -5, 6, 2, 6,
    -- filter=233 channel=78
    0, 0, 3, 0, -5, -1, 6, 0, 6,
    -- filter=233 channel=79
    0, 9, -3, 3, 4, -8, 14, -2, -19,
    -- filter=233 channel=80
    -7, 2, 4, -8, -5, 26, 8, 5, 21,
    -- filter=233 channel=81
    2, 4, -5, 3, -6, -6, 0, 1, -4,
    -- filter=233 channel=82
    2, -4, 6, -5, 3, 4, 0, 6, 5,
    -- filter=233 channel=83
    0, 8, -2, 5, 4, 1, 1, -1, 9,
    -- filter=233 channel=84
    2, -2, 0, 3, -4, 0, -3, -3, -17,
    -- filter=233 channel=85
    5, 7, 2, -2, -3, -1, 5, -7, 7,
    -- filter=233 channel=86
    -6, -5, -1, 1, -9, -10, 1, -14, -11,
    -- filter=233 channel=87
    -3, 2, -2, -4, -8, -12, -1, 0, -11,
    -- filter=233 channel=88
    -6, -8, 0, -8, -2, -2, -6, -6, 3,
    -- filter=233 channel=89
    14, 0, 8, 8, 13, 1, 10, 11, 1,
    -- filter=233 channel=90
    -7, -5, -7, -7, -2, -5, -4, -7, -7,
    -- filter=233 channel=91
    -2, 2, -5, 9, 10, -7, 1, 9, -10,
    -- filter=233 channel=92
    -1, 5, -6, 1, 0, -5, 2, 1, 2,
    -- filter=233 channel=93
    -20, -21, -3, -5, -19, -1, -12, -4, 6,
    -- filter=233 channel=94
    0, -2, -6, -6, -5, -3, 0, 1, 5,
    -- filter=233 channel=95
    5, 6, -4, -4, -7, 2, -7, 0, 4,
    -- filter=233 channel=96
    2, -3, 0, 6, 2, 7, 8, 6, 4,
    -- filter=233 channel=97
    -6, -4, -3, 1, -2, -5, -10, -2, 11,
    -- filter=233 channel=98
    3, 9, 3, -7, 15, 15, 3, 9, 4,
    -- filter=233 channel=99
    3, 15, 5, -4, 20, 1, -1, 10, -1,
    -- filter=233 channel=100
    0, 7, -4, 4, -7, 0, 9, 5, -2,
    -- filter=233 channel=101
    -3, 2, -1, -8, -1, 4, -1, 5, 0,
    -- filter=233 channel=102
    -5, 0, 0, 0, 3, 1, -5, -1, 4,
    -- filter=233 channel=103
    -6, -11, 13, -15, -12, 1, -18, -5, 19,
    -- filter=233 channel=104
    -14, -7, 12, -7, 0, 20, -4, 2, 19,
    -- filter=233 channel=105
    3, -1, -4, 0, -2, -12, 2, -3, -11,
    -- filter=233 channel=106
    -5, -7, 0, -1, 0, -7, -5, 7, -1,
    -- filter=233 channel=107
    -4, 5, -9, 1, 4, -8, 4, -1, -9,
    -- filter=233 channel=108
    -7, 3, -1, 5, -7, -6, 3, -1, 3,
    -- filter=233 channel=109
    0, 0, 0, -3, 7, 0, 8, -4, -10,
    -- filter=233 channel=110
    5, 1, 7, -10, 6, -2, -8, -1, 12,
    -- filter=233 channel=111
    0, -4, 0, 5, -1, -8, 0, -1, 1,
    -- filter=233 channel=112
    -3, 11, -9, -1, 5, 1, 6, 10, -5,
    -- filter=233 channel=113
    0, 0, 3, -8, 2, -4, -3, 0, 6,
    -- filter=233 channel=114
    5, 5, 0, -3, -8, -19, 16, -2, -22,
    -- filter=233 channel=115
    7, -3, -2, 0, 0, 0, -2, -3, -4,
    -- filter=233 channel=116
    0, -3, -1, 4, 11, 14, 7, 8, 0,
    -- filter=233 channel=117
    -7, 3, 6, -4, -2, 7, 6, 3, -1,
    -- filter=233 channel=118
    3, 3, -2, 5, 1, -2, -1, 0, 6,
    -- filter=233 channel=119
    2, -6, -9, -1, 0, -20, 1, -7, -6,
    -- filter=233 channel=120
    -3, 16, -6, -5, 17, -10, 2, 15, -9,
    -- filter=233 channel=121
    4, 0, 1, 0, -4, 0, 0, 2, 1,
    -- filter=233 channel=122
    -20, -26, 0, -25, -24, 14, -19, -17, 13,
    -- filter=233 channel=123
    2, 1, 1, 4, -4, -1, 3, 0, 0,
    -- filter=233 channel=124
    4, 0, -2, -2, -6, -10, -5, 5, -10,
    -- filter=233 channel=125
    2, 0, 1, -10, 13, 8, 2, -2, 0,
    -- filter=233 channel=126
    9, 0, 8, 9, -3, 6, 11, 7, 11,
    -- filter=233 channel=127
    2, 5, -4, -5, -5, 2, -3, 0, 0,
    -- filter=234 channel=0
    -2, -4, 0, 5, -5, -1, -6, -6, -7,
    -- filter=234 channel=1
    -5, 1, -1, 3, 0, -7, -5, 3, -2,
    -- filter=234 channel=2
    0, 4, -5, -6, -7, 3, 0, 2, 6,
    -- filter=234 channel=3
    -6, 0, 4, 2, 2, 2, -3, 2, 1,
    -- filter=234 channel=4
    3, -2, -4, 2, 5, -1, 2, 0, 4,
    -- filter=234 channel=5
    7, 5, 0, 7, -5, -3, -3, -1, 1,
    -- filter=234 channel=6
    4, -5, 1, -6, 5, -5, 0, -7, 3,
    -- filter=234 channel=7
    -5, -4, -1, -5, 7, -1, -6, -2, 0,
    -- filter=234 channel=8
    -2, 0, 3, -2, 7, 1, 0, -7, 4,
    -- filter=234 channel=9
    2, 2, -2, -1, -3, -5, 7, 4, -6,
    -- filter=234 channel=10
    -3, 0, -6, -4, -1, 0, 3, -3, -2,
    -- filter=234 channel=11
    2, -4, 1, 7, -4, 5, 0, -7, 2,
    -- filter=234 channel=12
    -5, -3, -6, 0, 0, 3, 0, 1, -2,
    -- filter=234 channel=13
    -4, 5, -1, -4, -3, 6, -2, 3, 3,
    -- filter=234 channel=14
    -4, -2, -3, -4, 1, -3, 1, -5, 3,
    -- filter=234 channel=15
    4, 0, 0, 5, -6, -3, 0, -5, -5,
    -- filter=234 channel=16
    -1, 5, 1, 3, 0, 2, 2, -6, -1,
    -- filter=234 channel=17
    1, -2, 1, -3, -6, 0, 5, 1, 7,
    -- filter=234 channel=18
    -2, -1, 3, 0, -1, 1, 3, 1, 2,
    -- filter=234 channel=19
    -6, -3, -4, 2, 6, -2, -3, -4, 6,
    -- filter=234 channel=20
    5, 1, 2, 3, 2, -6, -7, 5, 5,
    -- filter=234 channel=21
    -7, 0, 4, -1, 1, 5, 0, -7, 4,
    -- filter=234 channel=22
    0, 5, 1, 7, 1, 1, 5, 0, 2,
    -- filter=234 channel=23
    -1, -5, 6, -1, -3, -3, -5, -3, 2,
    -- filter=234 channel=24
    -5, -4, -3, -3, -5, 5, 4, -4, 0,
    -- filter=234 channel=25
    0, -4, 3, -4, -5, 4, 4, -6, -3,
    -- filter=234 channel=26
    5, 7, 4, -4, 1, -3, -4, -3, -6,
    -- filter=234 channel=27
    -3, -4, 0, -2, -3, -1, 1, -2, -2,
    -- filter=234 channel=28
    3, -5, 1, 4, 4, 6, 6, 2, 6,
    -- filter=234 channel=29
    3, -5, 0, -5, -3, 4, 1, 0, 0,
    -- filter=234 channel=30
    5, 3, 0, 1, -2, 2, 0, 4, 0,
    -- filter=234 channel=31
    -2, -6, 0, 0, 2, 0, -1, 0, -6,
    -- filter=234 channel=32
    6, -7, 0, 4, -2, 5, -5, -7, -2,
    -- filter=234 channel=33
    2, -5, -7, -4, 5, -6, -5, 5, 0,
    -- filter=234 channel=34
    -4, 4, -4, -6, 1, -1, 3, 0, -3,
    -- filter=234 channel=35
    -1, 4, 4, 1, 5, 2, 3, -5, -4,
    -- filter=234 channel=36
    3, -2, -7, 3, -3, 0, 5, 1, 4,
    -- filter=234 channel=37
    -4, 0, 6, 0, -7, 1, -1, 0, 6,
    -- filter=234 channel=38
    5, 3, -5, 4, 0, -7, -1, 0, -1,
    -- filter=234 channel=39
    -5, 4, -1, 0, 2, 6, -7, -4, 3,
    -- filter=234 channel=40
    7, -6, -1, 0, -5, 0, -5, 0, 6,
    -- filter=234 channel=41
    3, -6, 5, -7, -4, 0, -4, -4, -2,
    -- filter=234 channel=42
    3, 4, -1, 3, -6, 0, 2, 2, 2,
    -- filter=234 channel=43
    -1, 0, -4, -6, -1, -5, 6, -1, 5,
    -- filter=234 channel=44
    -3, 2, 0, 0, -2, 6, 7, -2, -7,
    -- filter=234 channel=45
    1, 2, 0, -5, -2, 2, 1, -4, 1,
    -- filter=234 channel=46
    6, 5, 4, 1, 2, -3, -4, -6, -7,
    -- filter=234 channel=47
    -6, -2, 1, 5, 5, 0, 3, -4, 0,
    -- filter=234 channel=48
    1, 2, 6, -3, 1, 0, 0, -2, -5,
    -- filter=234 channel=49
    1, -6, 1, -5, -5, 5, 7, -6, 1,
    -- filter=234 channel=50
    -4, 0, 0, -4, -7, -5, 6, 4, -5,
    -- filter=234 channel=51
    -2, 2, 7, 0, -2, -3, 3, -1, -5,
    -- filter=234 channel=52
    -2, 4, -3, 0, -2, 3, -3, 7, -7,
    -- filter=234 channel=53
    -5, 6, 0, -2, -3, -4, 3, -4, -4,
    -- filter=234 channel=54
    -4, 6, -4, -5, -1, 4, 2, 5, -2,
    -- filter=234 channel=55
    0, 0, 0, 0, 5, 3, 5, 5, 7,
    -- filter=234 channel=56
    -3, 6, 2, 5, 2, -2, 5, 2, -1,
    -- filter=234 channel=57
    -7, 3, -5, -7, -6, 4, 5, 0, -6,
    -- filter=234 channel=58
    3, 3, -2, 4, -4, -3, 5, 5, 0,
    -- filter=234 channel=59
    0, -3, -7, 7, -6, 3, -1, 2, 5,
    -- filter=234 channel=60
    -2, -4, -2, -3, 0, 0, -1, -5, 6,
    -- filter=234 channel=61
    2, -3, -3, 4, 4, -6, 0, -1, 4,
    -- filter=234 channel=62
    6, 0, 7, 1, -3, -5, 0, -5, 4,
    -- filter=234 channel=63
    -4, -6, -6, 3, -5, 2, 2, -4, -5,
    -- filter=234 channel=64
    -5, -6, -2, 3, 3, -3, 5, -2, 3,
    -- filter=234 channel=65
    -5, 0, 6, 2, 3, -5, -4, -6, 4,
    -- filter=234 channel=66
    1, -1, -1, -2, 5, -3, -2, 7, -1,
    -- filter=234 channel=67
    -3, -1, -5, -6, 7, -2, 0, 2, 1,
    -- filter=234 channel=68
    0, -2, -2, 2, -4, -6, 3, 0, -4,
    -- filter=234 channel=69
    0, -5, -4, 0, 3, 0, 1, -1, 4,
    -- filter=234 channel=70
    6, -3, -3, -6, -5, 6, 0, 3, 3,
    -- filter=234 channel=71
    -5, -2, 2, -5, -6, -3, 0, 0, 5,
    -- filter=234 channel=72
    -4, 0, -1, -5, -4, -6, -7, -2, -1,
    -- filter=234 channel=73
    -2, -4, -1, 5, -2, -2, 3, 0, 6,
    -- filter=234 channel=74
    0, 2, 2, -7, -6, -6, 6, -2, -2,
    -- filter=234 channel=75
    -4, -2, 7, 6, 4, 2, -1, 3, -5,
    -- filter=234 channel=76
    -5, 6, -2, -1, -3, -4, -4, 4, -1,
    -- filter=234 channel=77
    3, -3, -4, -5, 1, 5, 0, 0, 5,
    -- filter=234 channel=78
    -4, -3, 3, -7, -4, 3, 0, -3, -6,
    -- filter=234 channel=79
    0, -4, 5, 0, -1, 3, 0, -5, 3,
    -- filter=234 channel=80
    5, 3, 7, 0, -2, 1, -7, 1, 0,
    -- filter=234 channel=81
    1, 0, -1, 1, 6, 0, 4, -5, 4,
    -- filter=234 channel=82
    1, 4, -7, -3, 1, 3, -5, -5, 0,
    -- filter=234 channel=83
    6, 0, 5, 0, -6, -3, -6, 6, 6,
    -- filter=234 channel=84
    -7, -7, -3, 6, -7, 0, -4, -3, 3,
    -- filter=234 channel=85
    1, -4, 2, -2, 5, -5, -5, -2, -4,
    -- filter=234 channel=86
    -3, -2, -1, 0, -1, 5, -7, 5, 0,
    -- filter=234 channel=87
    -2, 0, -7, 4, -6, 4, 4, 0, 4,
    -- filter=234 channel=88
    -2, -3, 1, 0, 7, -5, 3, 5, 7,
    -- filter=234 channel=89
    -4, -3, -7, 1, 6, -2, 1, 2, -4,
    -- filter=234 channel=90
    -6, -5, -4, 1, -2, 4, -4, -6, 4,
    -- filter=234 channel=91
    -1, -6, 5, -2, 7, 0, -2, 1, -5,
    -- filter=234 channel=92
    2, 2, 6, -1, 1, -1, -3, 1, 4,
    -- filter=234 channel=93
    5, 5, 3, 1, 5, -5, 0, 3, 2,
    -- filter=234 channel=94
    -5, 3, 1, 0, 6, 0, -6, -5, 0,
    -- filter=234 channel=95
    3, 6, -7, 3, 0, -1, 0, -5, 6,
    -- filter=234 channel=96
    5, 6, -6, 7, 0, -1, -5, 3, 6,
    -- filter=234 channel=97
    -4, -2, 2, 5, 7, -6, -6, -6, 5,
    -- filter=234 channel=98
    -6, 4, -3, -4, -6, -2, 1, 5, 4,
    -- filter=234 channel=99
    1, 5, -6, 2, -6, 3, 0, -3, 6,
    -- filter=234 channel=100
    -1, 2, 0, 6, 2, 0, -2, 1, -6,
    -- filter=234 channel=101
    2, 0, 5, -2, 0, 2, -7, 4, -3,
    -- filter=234 channel=102
    2, -2, 4, 3, 4, 0, 5, -4, 5,
    -- filter=234 channel=103
    4, -3, 0, -1, -5, -6, 3, 6, -2,
    -- filter=234 channel=104
    3, -1, -6, 4, 3, -2, -6, -2, -1,
    -- filter=234 channel=105
    -6, -1, -7, -4, -3, 2, -1, -7, 5,
    -- filter=234 channel=106
    1, 6, -5, 2, 0, 1, 2, -3, 6,
    -- filter=234 channel=107
    -3, -2, 0, 3, 6, -1, 1, 6, 5,
    -- filter=234 channel=108
    -1, -3, -6, -4, -4, 0, 0, 0, 4,
    -- filter=234 channel=109
    3, 6, 5, 3, 0, 4, 3, 1, -8,
    -- filter=234 channel=110
    -5, 4, 5, -2, -1, 4, 0, 5, 1,
    -- filter=234 channel=111
    -2, 2, 6, -7, 7, 3, 2, 4, 6,
    -- filter=234 channel=112
    2, -1, -4, 3, 4, -5, 1, -5, 5,
    -- filter=234 channel=113
    7, -1, 6, 5, 0, 2, -2, -1, 7,
    -- filter=234 channel=114
    -5, 4, -6, 6, 2, -7, 5, 5, -2,
    -- filter=234 channel=115
    -1, 5, -5, 0, -2, -2, 6, 0, 1,
    -- filter=234 channel=116
    -6, 3, -2, 3, 0, 3, 0, -1, -5,
    -- filter=234 channel=117
    0, 0, 0, 3, 0, -4, 3, 3, -6,
    -- filter=234 channel=118
    6, -1, -4, 6, 3, -1, 5, -4, 5,
    -- filter=234 channel=119
    5, 0, -1, 0, -4, 5, -6, -3, -4,
    -- filter=234 channel=120
    7, -5, 3, -2, -2, -3, 0, 0, -4,
    -- filter=234 channel=121
    -4, 6, 2, -3, -4, -6, -7, -7, -7,
    -- filter=234 channel=122
    0, 3, 0, 5, 4, -3, -5, -6, -4,
    -- filter=234 channel=123
    6, -7, 2, 0, -1, 1, -4, 0, 4,
    -- filter=234 channel=124
    3, 0, 4, 3, 6, 1, -2, 0, -5,
    -- filter=234 channel=125
    -3, -3, -1, 2, -5, -3, 0, -2, 5,
    -- filter=234 channel=126
    -6, 6, 0, 5, 3, -5, -4, 0, -3,
    -- filter=234 channel=127
    -3, 1, 1, 2, -1, 3, 1, 0, -3,
    -- filter=235 channel=0
    16, 4, 3, 11, 6, -7, -3, -17, -20,
    -- filter=235 channel=1
    4, 16, 14, 3, 6, 6, -10, -9, -3,
    -- filter=235 channel=2
    2, 2, -1, 0, -11, -10, 3, 0, -2,
    -- filter=235 channel=3
    -4, -3, -2, -12, -2, -8, -4, 0, -2,
    -- filter=235 channel=4
    -1, 0, 4, -3, -8, -3, -13, -14, -1,
    -- filter=235 channel=5
    -3, -1, 6, 3, -1, 6, -13, -4, -13,
    -- filter=235 channel=6
    0, -4, -11, -5, -12, -9, -8, -11, 1,
    -- filter=235 channel=7
    2, 0, 5, 0, 4, 0, -5, -7, 4,
    -- filter=235 channel=8
    -5, 0, -3, 0, 2, -8, 0, -5, -6,
    -- filter=235 channel=9
    -3, 4, 4, 7, 1, 0, 2, 2, -6,
    -- filter=235 channel=10
    3, -7, -7, -7, 6, -6, 8, 1, 4,
    -- filter=235 channel=11
    -5, -8, -7, 2, -3, -3, 10, -3, -4,
    -- filter=235 channel=12
    1, 2, 3, -5, 1, 6, 3, -7, 7,
    -- filter=235 channel=13
    7, -5, 3, -6, 1, 4, 9, -5, 6,
    -- filter=235 channel=14
    -2, -5, 4, 7, 3, 5, 2, 0, 0,
    -- filter=235 channel=15
    17, 4, -4, 6, -8, -14, 8, -10, -14,
    -- filter=235 channel=16
    -17, 2, -2, -9, -1, 13, 0, 11, 12,
    -- filter=235 channel=17
    -5, 6, -7, -5, 6, 0, -4, 5, -5,
    -- filter=235 channel=18
    9, 9, -4, 0, -10, -22, 3, -17, -22,
    -- filter=235 channel=19
    -5, -5, 2, 3, -7, -3, -1, 6, 1,
    -- filter=235 channel=20
    1, -9, -16, 0, -4, -15, 7, -1, 0,
    -- filter=235 channel=21
    -20, -6, 8, 3, 4, 5, -4, 10, 18,
    -- filter=235 channel=22
    8, -1, -4, 2, -2, 0, -1, -6, 1,
    -- filter=235 channel=23
    5, -1, -11, -6, -3, -17, 4, -13, 0,
    -- filter=235 channel=24
    -7, 3, 6, -7, -1, -6, 5, -8, 4,
    -- filter=235 channel=25
    -2, 13, 3, -4, 0, -7, -2, 4, 4,
    -- filter=235 channel=26
    -13, -3, -7, -9, -3, 4, -3, -10, -6,
    -- filter=235 channel=27
    8, 21, 0, 9, 4, -16, 2, -1, -18,
    -- filter=235 channel=28
    1, 7, 0, -2, 6, 4, 0, -7, 1,
    -- filter=235 channel=29
    2, -10, -4, 0, -9, -13, 9, 1, 1,
    -- filter=235 channel=30
    4, 9, 0, -2, 4, -1, 0, -9, -8,
    -- filter=235 channel=31
    -24, -9, -7, 3, 6, -6, 3, 11, 11,
    -- filter=235 channel=32
    2, 5, -9, 8, -4, -15, 4, -11, -19,
    -- filter=235 channel=33
    4, 14, 1, -3, 2, -8, -2, -1, -12,
    -- filter=235 channel=34
    -9, -5, -2, -3, -12, 2, -1, -14, 1,
    -- filter=235 channel=35
    1, -1, 0, -6, 3, 6, 1, -1, -5,
    -- filter=235 channel=36
    -2, -15, -6, 0, -10, -5, 4, 0, 0,
    -- filter=235 channel=37
    5, 6, 9, 0, 12, 6, -7, -13, -9,
    -- filter=235 channel=38
    -2, 6, 0, 4, -4, -7, 6, -1, -6,
    -- filter=235 channel=39
    5, 3, -5, 3, -3, 1, 1, -4, -4,
    -- filter=235 channel=40
    6, -3, -10, -5, 5, -6, 4, 8, 0,
    -- filter=235 channel=41
    3, -7, 9, -6, -4, 17, 0, -10, 15,
    -- filter=235 channel=42
    9, 1, 8, 2, 6, -3, 4, 1, -3,
    -- filter=235 channel=43
    -1, 2, 1, -5, -13, -6, 4, -11, 0,
    -- filter=235 channel=44
    -12, 7, 6, 0, 13, 4, -2, 1, 0,
    -- filter=235 channel=45
    0, 0, 4, 4, 0, 1, 2, -3, 1,
    -- filter=235 channel=46
    2, 4, 0, 1, -4, 3, 0, -4, -6,
    -- filter=235 channel=47
    -17, 0, 3, -4, 19, 9, -2, 4, 10,
    -- filter=235 channel=48
    -8, 11, 9, 0, 1, 2, 0, 0, -7,
    -- filter=235 channel=49
    2, 5, -3, 0, -12, -17, -3, -6, -12,
    -- filter=235 channel=50
    0, 6, 4, 5, 7, 6, 0, 2, -9,
    -- filter=235 channel=51
    0, 5, 6, -5, 7, -4, -5, -3, -6,
    -- filter=235 channel=52
    3, -1, -7, -9, -9, -1, -3, -4, 1,
    -- filter=235 channel=53
    3, -3, -3, -3, -1, -5, 0, 1, -5,
    -- filter=235 channel=54
    7, 2, 0, -5, 1, -3, -6, 4, -2,
    -- filter=235 channel=55
    -1, -12, -12, -4, -4, -19, 2, 0, -10,
    -- filter=235 channel=56
    -1, -1, -1, 4, -11, 0, 3, -9, -4,
    -- filter=235 channel=57
    1, -10, 0, -1, 1, -4, -3, -5, 7,
    -- filter=235 channel=58
    -1, -1, -3, -8, 2, 0, -6, -2, -8,
    -- filter=235 channel=59
    0, 7, 8, -2, 12, 0, 7, -3, 5,
    -- filter=235 channel=60
    4, 3, 0, -6, -1, 0, 0, -7, 5,
    -- filter=235 channel=61
    -11, 1, -2, -10, -2, -6, -7, 0, -2,
    -- filter=235 channel=62
    -5, 0, 6, -5, -1, 1, 0, -6, 5,
    -- filter=235 channel=63
    -2, -10, -2, -6, 0, 6, 0, 1, -4,
    -- filter=235 channel=64
    0, -2, 0, -9, -11, 0, -3, 7, 6,
    -- filter=235 channel=65
    6, -3, 0, -5, 6, -5, -7, 3, -6,
    -- filter=235 channel=66
    -7, 3, 0, -2, -2, 4, -2, -9, 13,
    -- filter=235 channel=67
    -5, 6, 3, -6, -3, 4, 2, -4, 0,
    -- filter=235 channel=68
    0, -4, -3, 8, -6, -8, -1, 0, 7,
    -- filter=235 channel=69
    -2, -7, -1, 4, 2, 0, 2, -5, 5,
    -- filter=235 channel=70
    14, 13, 5, 7, -4, -3, 0, -4, 0,
    -- filter=235 channel=71
    0, 1, 8, 4, -1, 2, 3, 7, -4,
    -- filter=235 channel=72
    -2, 2, -6, -6, 0, 0, 9, 10, 0,
    -- filter=235 channel=73
    0, -7, -9, 4, 2, -5, -3, 1, -4,
    -- filter=235 channel=74
    3, -1, -7, 2, 0, -4, -4, 1, -2,
    -- filter=235 channel=75
    -1, 9, 8, 6, 16, 7, -11, 1, -4,
    -- filter=235 channel=76
    0, 1, -6, 1, -3, -16, 4, -3, -1,
    -- filter=235 channel=77
    -3, 0, 0, -7, 5, -1, 0, -2, 6,
    -- filter=235 channel=78
    1, -8, 2, -3, -7, 3, 0, -4, 0,
    -- filter=235 channel=79
    16, 14, -6, 14, 0, -13, 0, -3, -11,
    -- filter=235 channel=80
    -15, 5, 8, 6, 8, 12, 0, 16, 6,
    -- filter=235 channel=81
    3, 3, 0, -4, -4, 4, -3, 6, -1,
    -- filter=235 channel=82
    4, 0, 1, 5, 0, -1, 5, 0, 5,
    -- filter=235 channel=83
    0, -7, 7, 4, 0, -6, 4, 1, 0,
    -- filter=235 channel=84
    0, -1, 0, 5, -6, -14, -8, -11, -4,
    -- filter=235 channel=85
    -1, 3, 2, 0, -2, 5, -2, -5, 0,
    -- filter=235 channel=86
    -8, -6, 0, 3, -4, -8, -4, 0, -3,
    -- filter=235 channel=87
    -7, -9, 0, -2, 0, -3, -4, -6, 3,
    -- filter=235 channel=88
    -16, -10, -9, 2, 3, 0, -2, 4, 1,
    -- filter=235 channel=89
    0, 0, 1, 9, 8, -6, 5, -3, -2,
    -- filter=235 channel=90
    -10, -15, -8, -10, -3, -4, 5, 5, 6,
    -- filter=235 channel=91
    0, 12, -5, 4, 4, -12, -3, -5, -9,
    -- filter=235 channel=92
    -5, 0, -5, -3, -5, -2, -2, -7, -1,
    -- filter=235 channel=93
    -10, 5, 8, 2, 1, 9, 1, 0, 5,
    -- filter=235 channel=94
    3, 1, 3, -1, -2, 3, 7, -6, 2,
    -- filter=235 channel=95
    -4, 4, 6, 2, -6, -2, 5, -5, 4,
    -- filter=235 channel=96
    1, 0, 1, 1, 4, -4, 1, 5, -5,
    -- filter=235 channel=97
    -3, 7, 6, 0, -5, 10, 4, -3, 0,
    -- filter=235 channel=98
    -4, 5, 7, 0, 1, 2, -3, -7, -1,
    -- filter=235 channel=99
    -8, -17, -6, 1, -15, -13, 3, -7, -2,
    -- filter=235 channel=100
    -1, -7, 5, 1, -5, 4, -9, -4, 1,
    -- filter=235 channel=101
    -6, -2, -3, 1, -6, -9, -2, -5, 0,
    -- filter=235 channel=102
    5, 0, 1, 0, -4, -2, -2, 0, 6,
    -- filter=235 channel=103
    -12, -3, 8, 6, 12, 7, 1, 14, -1,
    -- filter=235 channel=104
    -14, -5, 7, 3, 11, 9, -1, 12, 8,
    -- filter=235 channel=105
    -2, -6, -9, 1, -6, 0, 2, -1, -7,
    -- filter=235 channel=106
    -3, 3, -7, 0, 1, -4, 8, 2, -5,
    -- filter=235 channel=107
    8, 6, -4, 8, -10, -13, -5, -4, -4,
    -- filter=235 channel=108
    -7, 0, 2, -7, -10, -2, -2, -6, 4,
    -- filter=235 channel=109
    11, 0, -1, 12, 8, -15, 2, -1, -6,
    -- filter=235 channel=110
    -13, -1, 1, 0, -11, -3, -6, 4, 2,
    -- filter=235 channel=111
    2, 0, 2, -4, -1, 0, 6, 2, 7,
    -- filter=235 channel=112
    0, 8, 0, 0, 5, -5, -5, -6, -6,
    -- filter=235 channel=113
    -3, 0, 3, 5, 11, 6, -2, -3, 4,
    -- filter=235 channel=114
    20, 13, -9, 9, -2, -21, -11, -26, -19,
    -- filter=235 channel=115
    2, 0, 4, -5, -6, 0, -1, 3, -2,
    -- filter=235 channel=116
    0, -11, 2, 0, -3, -7, 2, 2, -7,
    -- filter=235 channel=117
    -6, -3, 6, -1, -4, 6, 8, 5, 3,
    -- filter=235 channel=118
    2, 1, 7, 2, -7, 6, 3, 0, 0,
    -- filter=235 channel=119
    -7, -10, -3, -3, 0, 0, 0, 0, -2,
    -- filter=235 channel=120
    8, 8, -1, 3, -2, -10, -2, -6, -12,
    -- filter=235 channel=121
    -7, -9, 3, -4, -1, 0, -5, 5, -1,
    -- filter=235 channel=122
    -23, -8, 13, -4, 23, 27, -6, 20, 21,
    -- filter=235 channel=123
    -8, -2, -1, 0, 1, -5, -7, 3, -2,
    -- filter=235 channel=124
    7, 3, -11, -4, 3, 0, 4, -3, -1,
    -- filter=235 channel=125
    -10, -6, 1, -1, 4, -8, 5, -4, 5,
    -- filter=235 channel=126
    2, 4, 6, -5, 4, 7, 3, 6, -1,
    -- filter=235 channel=127
    -2, 5, 5, -6, 1, 5, -3, 1, 2,
    -- filter=236 channel=0
    6, 2, 14, 3, 1, -3, -12, 2, 3,
    -- filter=236 channel=1
    -4, -8, 3, 7, 2, -8, -11, -7, 0,
    -- filter=236 channel=2
    5, -8, -7, -5, 2, 4, -5, -1, -2,
    -- filter=236 channel=3
    -5, 22, 16, -2, -1, 6, -1, 1, -3,
    -- filter=236 channel=4
    8, -3, -4, 4, 25, 10, -3, 0, 7,
    -- filter=236 channel=5
    -4, 2, -1, 2, -6, 10, -1, -2, 0,
    -- filter=236 channel=6
    -5, 0, 6, -6, 0, -4, 0, 0, 4,
    -- filter=236 channel=7
    -1, 7, 4, 4, 2, 3, -5, 2, 4,
    -- filter=236 channel=8
    1, 0, -4, -7, 0, 5, 5, -5, -7,
    -- filter=236 channel=9
    -6, -6, 3, 9, 3, 2, 2, 8, -2,
    -- filter=236 channel=10
    -5, -4, -2, 6, 1, 1, 4, 7, -2,
    -- filter=236 channel=11
    -3, 7, 6, 0, 0, 1, -2, -4, -7,
    -- filter=236 channel=12
    2, -5, 0, -1, -6, -4, -5, 4, -2,
    -- filter=236 channel=13
    -9, -15, 13, 3, -3, -14, 0, 4, -4,
    -- filter=236 channel=14
    5, 5, -2, 1, -2, 2, -1, 5, -1,
    -- filter=236 channel=15
    -1, 7, 11, 5, -15, -8, 0, 8, -3,
    -- filter=236 channel=16
    -4, 7, 1, 1, 0, 1, 2, 14, -1,
    -- filter=236 channel=17
    -1, -3, 6, -7, 6, -3, -1, -6, -3,
    -- filter=236 channel=18
    -9, -6, 11, 8, -4, -3, -4, -6, -3,
    -- filter=236 channel=19
    -1, 0, -5, 5, -3, -4, -5, -6, -2,
    -- filter=236 channel=20
    -5, 9, 10, 10, -9, -3, 9, -4, -5,
    -- filter=236 channel=21
    2, 1, -4, -4, 0, 0, -2, 8, 4,
    -- filter=236 channel=22
    2, 3, 13, 0, -4, 7, 8, -3, -4,
    -- filter=236 channel=23
    -12, 11, 16, 16, -29, 7, 13, 13, -19,
    -- filter=236 channel=24
    3, -1, 1, -2, -1, -6, 5, 3, -1,
    -- filter=236 channel=25
    0, -12, -1, 16, 0, -14, -16, 3, 6,
    -- filter=236 channel=26
    6, 0, -7, -2, 5, -2, -5, -3, -3,
    -- filter=236 channel=27
    -13, -3, 16, 24, -6, -6, -2, 13, -6,
    -- filter=236 channel=28
    -3, 1, -6, 6, 0, -5, -4, -4, 3,
    -- filter=236 channel=29
    5, 3, 8, 4, -5, -2, 5, -7, 0,
    -- filter=236 channel=30
    -8, -9, 10, 2, 1, -6, 0, 0, -6,
    -- filter=236 channel=31
    -15, -1, -8, 18, -6, -3, 0, 20, -3,
    -- filter=236 channel=32
    1, 0, 15, 17, -5, 1, -11, -3, -6,
    -- filter=236 channel=33
    -11, 0, 19, 2, -15, -6, -9, 14, 0,
    -- filter=236 channel=34
    -2, 18, 7, 6, -17, 12, 15, 6, -9,
    -- filter=236 channel=35
    4, 5, -3, 7, 1, -7, -6, 0, 2,
    -- filter=236 channel=36
    -1, -7, -7, -1, 11, -1, -7, 5, -3,
    -- filter=236 channel=37
    -8, 4, -5, -8, 0, -4, -13, 4, -4,
    -- filter=236 channel=38
    3, 8, 0, 1, -11, 2, 0, 8, 0,
    -- filter=236 channel=39
    4, -7, 7, 9, -3, -8, -3, -6, -5,
    -- filter=236 channel=40
    2, 0, -1, -6, -10, -1, -1, -3, -8,
    -- filter=236 channel=41
    1, -16, -2, -1, 24, -13, -2, 0, 6,
    -- filter=236 channel=42
    -2, 3, 3, -5, -1, -7, 0, -1, -1,
    -- filter=236 channel=43
    -9, 11, 14, -6, -10, 1, 6, 8, -6,
    -- filter=236 channel=44
    0, 0, -8, 0, 5, 0, -11, -1, -2,
    -- filter=236 channel=45
    0, 3, 5, 5, -3, 2, -3, -3, 3,
    -- filter=236 channel=46
    1, -1, 1, -7, -1, -5, 2, -6, -5,
    -- filter=236 channel=47
    -7, 8, -1, 7, 10, -7, -13, 10, 9,
    -- filter=236 channel=48
    8, -15, -5, 10, 11, 0, -13, 3, 0,
    -- filter=236 channel=49
    -1, -10, 8, 3, 5, -6, -12, -1, 3,
    -- filter=236 channel=50
    -9, -2, 3, 15, -10, -10, -2, 0, -10,
    -- filter=236 channel=51
    5, 6, -1, -5, -6, 3, -1, -6, -2,
    -- filter=236 channel=52
    0, 8, -1, 8, -2, 7, -2, -2, 2,
    -- filter=236 channel=53
    -6, -5, 0, -1, 0, -3, 8, -6, 0,
    -- filter=236 channel=54
    2, -1, 0, -4, -5, 0, -2, -4, 3,
    -- filter=236 channel=55
    -5, 3, 1, 2, -7, -12, 1, -1, 3,
    -- filter=236 channel=56
    1, 0, 1, 5, -9, -5, 0, -3, 5,
    -- filter=236 channel=57
    6, 3, 4, -5, 10, 1, -1, 0, 9,
    -- filter=236 channel=58
    6, 6, 2, -6, 6, 5, -11, 6, 6,
    -- filter=236 channel=59
    7, -9, -6, 9, 7, -4, -14, 7, 9,
    -- filter=236 channel=60
    0, -5, 4, -7, 3, -4, 2, -4, 0,
    -- filter=236 channel=61
    0, -2, 3, 4, -4, 0, 5, -1, 0,
    -- filter=236 channel=62
    6, -1, 6, -6, 0, 3, -4, -6, 2,
    -- filter=236 channel=63
    2, 8, -4, 2, 2, 3, -7, 4, -1,
    -- filter=236 channel=64
    5, 0, -2, -7, -3, 2, -4, -3, 1,
    -- filter=236 channel=65
    -6, 1, -4, 3, 5, -5, -4, -2, 5,
    -- filter=236 channel=66
    4, -4, 0, 3, -2, -5, -1, 0, 8,
    -- filter=236 channel=67
    4, -2, -6, -6, -5, -6, -4, -2, 1,
    -- filter=236 channel=68
    -1, -5, 0, -5, 1, -8, -6, -3, 7,
    -- filter=236 channel=69
    -1, 3, 0, 2, -6, 0, -5, -2, 7,
    -- filter=236 channel=70
    -10, 4, 15, 8, -16, -4, -6, -2, -11,
    -- filter=236 channel=71
    -9, 0, 4, 2, -10, 0, 5, 3, 0,
    -- filter=236 channel=72
    -1, -12, -3, 12, 4, -16, -3, 13, 0,
    -- filter=236 channel=73
    5, 1, 4, 8, -3, 1, -7, 4, 2,
    -- filter=236 channel=74
    0, -8, -4, -3, -7, 7, 2, 7, 0,
    -- filter=236 channel=75
    1, 7, 9, 2, -10, 0, -3, 13, -7,
    -- filter=236 channel=76
    -6, 0, 6, -1, -10, 1, 1, -10, 1,
    -- filter=236 channel=77
    2, -1, -4, 5, 0, -1, -3, 2, 4,
    -- filter=236 channel=78
    -6, 0, -3, -3, 8, -1, 0, 5, -4,
    -- filter=236 channel=79
    -10, -13, 18, 12, -13, -1, -12, 3, -10,
    -- filter=236 channel=80
    1, -12, -10, 17, 0, -14, -11, 12, 7,
    -- filter=236 channel=81
    -4, 0, -4, 0, -4, -3, 3, 2, -7,
    -- filter=236 channel=82
    2, 3, 8, -3, 1, -5, 3, -3, 1,
    -- filter=236 channel=83
    3, -8, -1, 4, 2, -2, -11, 2, 6,
    -- filter=236 channel=84
    -2, -5, 10, 6, 0, -7, -6, 0, 1,
    -- filter=236 channel=85
    2, -1, 3, 7, -2, 3, -2, 6, 3,
    -- filter=236 channel=86
    -8, 3, 11, 6, -8, 0, 1, 7, 4,
    -- filter=236 channel=87
    -5, -1, 8, 1, -10, 6, 11, 0, 0,
    -- filter=236 channel=88
    -7, 3, -13, -3, 2, -1, 8, 3, 0,
    -- filter=236 channel=89
    2, -10, 6, 10, -7, -15, -2, 0, -6,
    -- filter=236 channel=90
    -4, 7, -7, -4, -3, 8, 1, 6, -2,
    -- filter=236 channel=91
    -1, -17, 3, 11, -4, -9, -4, -1, -2,
    -- filter=236 channel=92
    -2, 12, 5, -4, -4, 4, 13, 4, -6,
    -- filter=236 channel=93
    6, 0, -12, 3, 4, -1, -18, 4, 8,
    -- filter=236 channel=94
    -3, 1, 0, -1, 0, -6, -5, -3, 7,
    -- filter=236 channel=95
    0, 1, 7, 2, 4, 0, -2, 0, -6,
    -- filter=236 channel=96
    6, -6, -5, 2, -2, 3, 0, 1, -5,
    -- filter=236 channel=97
    0, 8, 6, -7, 0, 4, 7, 11, -4,
    -- filter=236 channel=98
    -7, -7, 7, 20, -7, 0, -7, 10, -1,
    -- filter=236 channel=99
    -9, 5, 6, 10, -16, 0, 14, 14, 2,
    -- filter=236 channel=100
    4, 5, 3, -8, 7, -3, 1, 0, 7,
    -- filter=236 channel=101
    0, 0, -6, 0, 18, 2, 3, 5, 8,
    -- filter=236 channel=102
    6, 0, 2, -4, -2, 2, -1, 2, 0,
    -- filter=236 channel=103
    6, 11, 3, -2, 1, 0, -3, 18, -5,
    -- filter=236 channel=104
    4, -1, -9, 5, 10, -6, 0, 7, -5,
    -- filter=236 channel=105
    1, -4, 8, -4, 1, 0, 8, -6, -3,
    -- filter=236 channel=106
    7, 4, 4, 3, -7, 3, -5, -2, -3,
    -- filter=236 channel=107
    -10, 5, 13, 5, -15, 1, 11, -3, -1,
    -- filter=236 channel=108
    -2, -3, 7, -4, 4, -7, -3, 6, -3,
    -- filter=236 channel=109
    -7, -4, -1, 20, -9, -11, -9, 4, -3,
    -- filter=236 channel=110
    -7, 5, 0, 9, 2, -6, -2, 12, -7,
    -- filter=236 channel=111
    6, 2, 0, 7, 6, -5, 3, -4, 5,
    -- filter=236 channel=112
    -5, -4, 9, 1, -2, 0, 3, 14, -9,
    -- filter=236 channel=113
    0, -1, 11, -3, -14, 0, 9, 7, -9,
    -- filter=236 channel=114
    -7, -13, 12, 8, -1, -1, -3, -7, 5,
    -- filter=236 channel=115
    0, 0, 6, 6, 3, -5, -5, 7, 5,
    -- filter=236 channel=116
    0, -16, 4, 8, 13, -17, -9, 3, 6,
    -- filter=236 channel=117
    -1, 0, -2, -1, 2, -8, -6, -6, 6,
    -- filter=236 channel=118
    -5, -4, 6, 0, -1, -1, 6, -1, 2,
    -- filter=236 channel=119
    -9, 9, 1, -3, 0, 5, 13, 0, -9,
    -- filter=236 channel=120
    0, -9, 11, 7, -19, -5, 1, 8, -6,
    -- filter=236 channel=121
    5, 0, 5, -2, 6, 2, 6, 7, 7,
    -- filter=236 channel=122
    -7, 0, -6, 9, 1, -4, -15, 13, 0,
    -- filter=236 channel=123
    -6, 12, 0, 0, -8, 0, 10, 5, 2,
    -- filter=236 channel=124
    -4, 7, 7, 5, -8, 3, 0, 6, -2,
    -- filter=236 channel=125
    -1, -4, 2, 15, 2, -5, -9, 6, -4,
    -- filter=236 channel=126
    -2, -1, -1, 1, 0, -8, -5, -1, -2,
    -- filter=236 channel=127
    -4, -4, 0, -4, 4, -6, -4, 2, 2,
    -- filter=237 channel=0
    -17, 12, -15, 8, 45, -6, 0, 16, -18,
    -- filter=237 channel=1
    -6, 5, -13, 6, 30, 0, 0, 10, -25,
    -- filter=237 channel=2
    5, 0, 2, 3, -8, -5, -1, 6, 0,
    -- filter=237 channel=3
    0, 0, 9, -1, 3, 4, -6, 6, -6,
    -- filter=237 channel=4
    -2, 8, 8, -2, 2, 9, 3, 2, -2,
    -- filter=237 channel=5
    -8, 6, -11, 14, 42, -10, -4, 12, -9,
    -- filter=237 channel=6
    -5, 5, 0, -7, 0, -5, 2, -4, -2,
    -- filter=237 channel=7
    2, 5, 3, -6, 0, -2, -7, -3, -3,
    -- filter=237 channel=8
    0, 4, 7, -3, 3, 6, 2, 1, -1,
    -- filter=237 channel=9
    -3, 2, -3, 8, 4, 0, -2, -3, -7,
    -- filter=237 channel=10
    8, -8, 4, -3, -6, 0, -2, -2, 12,
    -- filter=237 channel=11
    1, -6, 8, -12, -7, -5, 0, 7, 5,
    -- filter=237 channel=12
    0, -8, 5, 4, -9, 2, 0, 3, 3,
    -- filter=237 channel=13
    0, -9, -3, -1, -15, 4, 5, 0, 5,
    -- filter=237 channel=14
    5, -4, 3, -1, 1, 0, -3, -2, -3,
    -- filter=237 channel=15
    4, -6, -1, -9, -9, -9, 8, -2, 5,
    -- filter=237 channel=16
    0, -3, 0, 0, 14, -3, -11, 1, -8,
    -- filter=237 channel=17
    -4, -6, 7, -2, 0, 3, 3, 3, 6,
    -- filter=237 channel=18
    2, 0, -1, -4, -9, -7, 2, -3, -5,
    -- filter=237 channel=19
    7, 0, -2, 1, 4, 1, 2, -3, 6,
    -- filter=237 channel=20
    14, -2, 3, -6, -15, 2, 15, 0, 10,
    -- filter=237 channel=21
    -2, -6, -5, 3, 7, 9, -8, -6, 1,
    -- filter=237 channel=22
    7, 3, -6, 10, 4, -6, 9, 5, 1,
    -- filter=237 channel=23
    3, 7, 10, -11, -22, 2, 5, 1, 9,
    -- filter=237 channel=24
    -3, 4, -3, -1, 6, -6, -5, 1, 6,
    -- filter=237 channel=25
    0, 2, -2, 8, 4, -7, -1, -9, -4,
    -- filter=237 channel=26
    -6, 8, -3, 7, 8, 0, -6, -4, -9,
    -- filter=237 channel=27
    -9, -5, 1, -1, 0, -2, 6, 7, -6,
    -- filter=237 channel=28
    4, 1, 5, 5, -4, -6, -5, -6, 4,
    -- filter=237 channel=29
    8, 0, 5, -10, -18, -4, 10, 9, 17,
    -- filter=237 channel=30
    -12, 4, -5, 4, 12, 2, -6, 3, 2,
    -- filter=237 channel=31
    -5, -9, 4, -13, -3, 14, -11, -5, 3,
    -- filter=237 channel=32
    0, -3, -2, 2, -4, 0, -1, 4, -4,
    -- filter=237 channel=33
    5, -3, -7, -5, 1, 1, -8, -6, -2,
    -- filter=237 channel=34
    3, 4, -4, 10, 8, -12, 8, 4, 5,
    -- filter=237 channel=35
    -6, -6, -2, -6, 6, 6, 3, 2, -7,
    -- filter=237 channel=36
    -7, -10, 8, 0, -19, 10, 4, -6, 8,
    -- filter=237 channel=37
    -11, 9, -6, 10, 39, -4, -6, 11, -16,
    -- filter=237 channel=38
    -1, 6, -1, 3, 3, -8, 3, -2, -1,
    -- filter=237 channel=39
    5, -6, 2, -11, -12, -1, 7, 8, 14,
    -- filter=237 channel=40
    8, -5, 4, 1, -11, 1, 9, 0, 0,
    -- filter=237 channel=41
    0, 3, -9, -6, -5, -18, 0, -12, -20,
    -- filter=237 channel=42
    -14, -3, -3, -7, 8, 5, 0, -2, 5,
    -- filter=237 channel=43
    -3, 1, 5, -4, -1, 5, -3, -4, -6,
    -- filter=237 channel=44
    -15, -1, -7, 11, 26, 2, -13, 4, -3,
    -- filter=237 channel=45
    -5, -2, 3, -2, 10, 1, 5, 0, -3,
    -- filter=237 channel=46
    3, -6, -4, 5, -2, -1, 6, 3, -3,
    -- filter=237 channel=47
    1, -4, 1, 3, 13, 5, -8, 5, 0,
    -- filter=237 channel=48
    2, 6, -2, 9, 14, -4, 1, 4, -3,
    -- filter=237 channel=49
    -5, 1, 2, -7, 1, 2, -1, 7, -1,
    -- filter=237 channel=50
    4, 2, -3, 1, 1, 5, -3, -5, 0,
    -- filter=237 channel=51
    0, 1, 0, -4, -5, 7, 7, -1, 0,
    -- filter=237 channel=52
    0, -5, -1, 5, -4, 0, -2, 0, 3,
    -- filter=237 channel=53
    2, 6, 10, -4, -10, -6, -4, -4, 1,
    -- filter=237 channel=54
    2, 2, -3, -5, 1, 3, -6, -6, 4,
    -- filter=237 channel=55
    4, -8, 17, -12, -32, -3, 3, -1, 19,
    -- filter=237 channel=56
    2, 0, 3, -4, 1, 0, 3, 1, -5,
    -- filter=237 channel=57
    -8, 5, 4, -8, 2, -3, 0, -4, -2,
    -- filter=237 channel=58
    -12, 4, -5, -4, 19, 0, -10, 8, 1,
    -- filter=237 channel=59
    4, 4, 1, 6, 5, 3, 3, -7, -4,
    -- filter=237 channel=60
    -1, 4, 6, 0, 7, 2, 0, 0, -1,
    -- filter=237 channel=61
    5, -1, 4, 3, 1, 2, 4, 4, 5,
    -- filter=237 channel=62
    8, 0, 1, -5, 0, -1, 7, -1, 5,
    -- filter=237 channel=63
    -9, 2, -5, 0, 8, -1, -5, 5, -1,
    -- filter=237 channel=64
    0, -8, 7, -11, -7, -5, 0, -5, -4,
    -- filter=237 channel=65
    4, 1, -6, 5, -4, 0, -3, -6, 5,
    -- filter=237 channel=66
    4, 1, 1, 0, -2, -10, 1, -7, -1,
    -- filter=237 channel=67
    2, -6, 3, -5, -7, -8, 0, -4, -2,
    -- filter=237 channel=68
    0, -3, 4, 5, -12, 2, 2, 2, 8,
    -- filter=237 channel=69
    4, -6, -5, -5, -1, 2, -2, -2, 0,
    -- filter=237 channel=70
    -9, -5, 1, -1, -1, 2, -8, -3, 0,
    -- filter=237 channel=71
    3, -7, -7, -1, -6, -1, -7, 4, 0,
    -- filter=237 channel=72
    -5, 1, 2, -5, -5, 2, -5, -9, 8,
    -- filter=237 channel=73
    -1, 1, 0, -3, -13, -6, 2, 1, 6,
    -- filter=237 channel=74
    -2, 0, -1, 2, 10, -6, 7, 3, -2,
    -- filter=237 channel=75
    -13, 17, -7, 5, 43, -9, -8, 10, -23,
    -- filter=237 channel=76
    3, -6, 4, -3, -23, -7, 11, 4, 15,
    -- filter=237 channel=77
    -6, 2, 1, -3, 3, 0, 0, -5, 4,
    -- filter=237 channel=78
    -2, 6, 0, 1, 12, 6, 0, 8, 1,
    -- filter=237 channel=79
    3, -7, 7, -5, -16, -9, 9, 6, 4,
    -- filter=237 channel=80
    -1, -1, 3, 0, 8, 9, 3, -6, 3,
    -- filter=237 channel=81
    -1, -6, 6, -3, 3, 2, 7, -1, -6,
    -- filter=237 channel=82
    -4, 1, 0, 6, -2, -4, -7, 3, -4,
    -- filter=237 channel=83
    -3, 1, 3, 0, 0, -2, -1, -2, -4,
    -- filter=237 channel=84
    -1, 6, 1, -5, 0, 0, 9, 8, 7,
    -- filter=237 channel=85
    -3, -3, 4, 3, 6, 6, 0, 1, 2,
    -- filter=237 channel=86
    -7, 3, -3, 2, 8, -2, -5, 1, -4,
    -- filter=237 channel=87
    2, -2, 4, -3, -8, -2, -4, 7, 2,
    -- filter=237 channel=88
    -3, -9, -3, -10, -15, 3, -5, -9, -3,
    -- filter=237 channel=89
    -2, 1, 14, -6, -19, 3, -5, -7, 13,
    -- filter=237 channel=90
    5, -6, 4, -10, -14, -3, -7, -1, 5,
    -- filter=237 channel=91
    -2, 0, 5, -10, -14, -3, -1, -1, 6,
    -- filter=237 channel=92
    0, -2, -2, -6, -3, 0, 3, 4, -1,
    -- filter=237 channel=93
    -5, 0, -5, 8, 35, 4, -8, 10, -12,
    -- filter=237 channel=94
    7, 2, -6, 2, -1, 4, -3, 0, 5,
    -- filter=237 channel=95
    -3, -1, 0, 4, 0, 0, -2, 0, 6,
    -- filter=237 channel=96
    -1, 2, 4, -4, -6, -2, 5, 6, -4,
    -- filter=237 channel=97
    -5, 1, 1, -7, -7, 0, -9, 6, -1,
    -- filter=237 channel=98
    -8, 1, -5, 0, 4, -3, 4, 9, 6,
    -- filter=237 channel=99
    0, 3, 7, -5, -17, 4, -1, -1, 6,
    -- filter=237 channel=100
    -1, -3, -4, -3, 3, -5, -2, -3, -10,
    -- filter=237 channel=101
    -5, -5, 9, 1, 3, 6, -1, 11, 3,
    -- filter=237 channel=102
    -7, -4, -3, -2, 4, 0, -2, -6, -2,
    -- filter=237 channel=103
    2, 2, 0, 12, 22, 4, -13, 4, -12,
    -- filter=237 channel=104
    6, 2, 4, 6, 4, 11, -6, -5, 2,
    -- filter=237 channel=105
    6, 7, -2, -5, -5, 0, 6, -5, 13,
    -- filter=237 channel=106
    0, -7, 3, -8, -7, -6, 4, -1, 4,
    -- filter=237 channel=107
    7, 2, -3, -9, -8, -1, 9, -4, 4,
    -- filter=237 channel=108
    0, 8, -4, 5, 1, -10, 5, -2, -6,
    -- filter=237 channel=109
    6, 6, 3, 7, -9, -4, 3, -3, 4,
    -- filter=237 channel=110
    0, -1, 6, -2, -3, 9, -6, -6, 12,
    -- filter=237 channel=111
    5, 0, 4, 11, 2, 0, 1, 7, -4,
    -- filter=237 channel=112
    0, -1, 7, 10, 9, -5, 6, 3, 0,
    -- filter=237 channel=113
    3, -3, -2, -4, -4, -4, -8, -8, 7,
    -- filter=237 channel=114
    -5, 7, -8, 17, 9, -12, 18, 18, 0,
    -- filter=237 channel=115
    -3, 0, 7, -7, 6, -6, 2, 4, 2,
    -- filter=237 channel=116
    -3, -7, 8, -4, -5, 9, 14, 0, 7,
    -- filter=237 channel=117
    7, -3, -5, 0, 0, 5, -1, -2, 0,
    -- filter=237 channel=118
    2, 7, -1, -5, -2, 2, 3, -7, -7,
    -- filter=237 channel=119
    6, 5, -8, 2, 8, -16, 5, -6, -7,
    -- filter=237 channel=120
    4, -1, 2, -6, -8, -9, 0, 9, 9,
    -- filter=237 channel=121
    8, -5, 2, -7, -1, 0, 0, 2, 6,
    -- filter=237 channel=122
    -9, -9, -8, 5, 22, 13, -19, -10, -1,
    -- filter=237 channel=123
    -2, -7, -6, 2, 0, -10, 2, 4, -4,
    -- filter=237 channel=124
    4, 4, 1, 5, -8, -3, 2, 1, -2,
    -- filter=237 channel=125
    10, 0, 4, 1, -6, 4, 8, 5, 11,
    -- filter=237 channel=126
    8, 6, -5, 0, -7, -4, -4, -8, -2,
    -- filter=237 channel=127
    5, 1, -2, 0, -7, -9, 5, 0, -9,
    -- filter=238 channel=0
    1, 0, -8, 5, -5, 0, 0, -4, 0,
    -- filter=238 channel=1
    1, -7, -11, 6, -7, -9, 4, -9, 3,
    -- filter=238 channel=2
    1, 7, 4, 2, 1, 2, -3, 2, 6,
    -- filter=238 channel=3
    -5, -10, 0, -13, -16, -6, 3, -13, -14,
    -- filter=238 channel=4
    0, -4, 0, -3, -9, 5, 0, 15, 1,
    -- filter=238 channel=5
    6, -6, -4, 7, -2, -3, 0, -5, -5,
    -- filter=238 channel=6
    -9, 7, 5, -7, 8, 9, 0, 3, 7,
    -- filter=238 channel=7
    2, -2, -5, 1, 2, 5, 2, -1, 0,
    -- filter=238 channel=8
    -3, 3, -1, 0, 5, 10, 7, 6, 2,
    -- filter=238 channel=9
    -6, 3, 0, -2, -1, 0, -3, 9, 2,
    -- filter=238 channel=10
    -5, -6, -6, -8, 3, -3, 1, -6, 2,
    -- filter=238 channel=11
    -4, 10, 7, -3, 15, 11, -2, 10, 7,
    -- filter=238 channel=12
    -1, 0, 8, 9, -4, 0, -3, 4, 6,
    -- filter=238 channel=13
    -5, -8, 0, 1, -7, 6, -5, 0, -4,
    -- filter=238 channel=14
    3, 3, 2, 0, 3, 1, -2, 0, 1,
    -- filter=238 channel=15
    -21, 0, 9, -5, 7, 15, -5, 0, 9,
    -- filter=238 channel=16
    -3, -8, -4, -1, -7, -8, -6, -3, 0,
    -- filter=238 channel=17
    4, 0, -3, 7, 3, 0, 1, 2, -6,
    -- filter=238 channel=18
    -19, -14, 12, -1, 0, 11, 3, 8, 12,
    -- filter=238 channel=19
    2, 4, 6, 3, -2, -1, 6, 5, 3,
    -- filter=238 channel=20
    -9, 7, 10, 1, 24, 17, -11, 0, 4,
    -- filter=238 channel=21
    1, -17, -5, -3, -9, -7, -8, -10, -6,
    -- filter=238 channel=22
    2, -5, 8, -9, 5, 9, 2, -1, 0,
    -- filter=238 channel=23
    -10, -4, 11, -9, 10, 7, -4, 0, 1,
    -- filter=238 channel=24
    5, 2, 6, -4, 6, 4, 0, -2, 6,
    -- filter=238 channel=25
    -10, -18, 3, -10, -15, 0, 4, 4, 11,
    -- filter=238 channel=26
    3, -3, 3, 0, 2, 0, -7, 3, 0,
    -- filter=238 channel=27
    -15, -8, 3, -7, 0, 5, -2, 14, 25,
    -- filter=238 channel=28
    5, 0, 1, -4, -1, -4, -5, -5, -1,
    -- filter=238 channel=29
    0, 8, 4, 4, 22, 17, -1, 3, 8,
    -- filter=238 channel=30
    -5, -9, -7, 2, -13, -1, 0, 2, 8,
    -- filter=238 channel=31
    1, -7, -12, -1, 0, 0, 0, -3, 3,
    -- filter=238 channel=32
    -18, -14, 3, -4, -4, 16, -7, 5, 15,
    -- filter=238 channel=33
    -12, -11, 2, -15, -10, 7, -4, -3, 9,
    -- filter=238 channel=34
    3, 12, 6, -3, 6, 4, -2, 5, 11,
    -- filter=238 channel=35
    -3, 0, 5, -2, -1, 0, -5, -3, 2,
    -- filter=238 channel=36
    -4, -4, -2, 4, -7, -4, -4, -5, -5,
    -- filter=238 channel=37
    6, -3, -10, -6, -17, -9, 0, -2, -10,
    -- filter=238 channel=38
    2, -3, 2, -2, 3, -3, -7, 5, 0,
    -- filter=238 channel=39
    3, 9, 8, -5, 5, 7, -3, -6, 2,
    -- filter=238 channel=40
    -5, -4, 4, 4, 1, -2, 0, 0, -3,
    -- filter=238 channel=41
    -4, 4, 9, 0, 0, 10, -2, 0, 12,
    -- filter=238 channel=42
    -4, -9, 6, -1, -7, -7, 4, 0, -3,
    -- filter=238 channel=43
    -13, -4, -7, -12, 4, 6, -12, -10, -7,
    -- filter=238 channel=44
    -8, -5, -12, -2, -8, -5, 7, -9, 2,
    -- filter=238 channel=45
    5, -4, 0, 7, -1, 0, -7, 4, -2,
    -- filter=238 channel=46
    3, -2, -3, 2, 7, 0, -1, -3, 3,
    -- filter=238 channel=47
    -5, -11, -16, -1, -19, -16, -1, -16, -4,
    -- filter=238 channel=48
    0, -17, -7, -11, -16, -5, 12, 0, 0,
    -- filter=238 channel=49
    -6, 1, 4, 5, 9, 8, 6, 11, 9,
    -- filter=238 channel=50
    -9, 2, -3, 1, -2, -1, 2, 7, 10,
    -- filter=238 channel=51
    4, 1, -1, -1, 4, 1, -2, -6, 5,
    -- filter=238 channel=52
    -3, 8, 2, 0, 0, -1, 3, -1, -1,
    -- filter=238 channel=53
    2, -5, 0, -6, 8, 11, 1, 5, 9,
    -- filter=238 channel=54
    3, 6, -5, 7, 1, -1, -4, -2, -5,
    -- filter=238 channel=55
    -8, -2, 4, -10, 7, 3, -9, -5, 6,
    -- filter=238 channel=56
    2, -3, 8, 4, 5, -2, 1, 4, 7,
    -- filter=238 channel=57
    -2, 5, -2, -5, -9, 2, 7, -4, 0,
    -- filter=238 channel=58
    -2, 0, 7, 8, -2, 6, -2, 2, 3,
    -- filter=238 channel=59
    -4, -9, -5, -5, -8, 5, 2, 0, 3,
    -- filter=238 channel=60
    3, 0, -5, -3, 3, -5, 5, -3, 2,
    -- filter=238 channel=61
    4, -4, 0, -5, 6, 0, -6, 5, -2,
    -- filter=238 channel=62
    1, -8, 0, -3, 4, 1, -2, -3, 6,
    -- filter=238 channel=63
    1, 2, 4, 3, -2, -2, -7, 3, -5,
    -- filter=238 channel=64
    -5, 4, -7, 1, 2, -7, -1, 3, -7,
    -- filter=238 channel=65
    0, 0, -5, 6, 2, -3, -6, -4, 2,
    -- filter=238 channel=66
    2, 4, 9, 0, 4, 7, 7, 6, 0,
    -- filter=238 channel=67
    0, 7, 2, -6, -2, 0, 6, -3, -1,
    -- filter=238 channel=68
    -7, -3, 0, 1, 4, 0, -5, -2, 4,
    -- filter=238 channel=69
    1, 2, -2, 2, -3, 3, -3, -4, -1,
    -- filter=238 channel=70
    -16, 3, -2, -1, 4, 8, 6, 2, 13,
    -- filter=238 channel=71
    3, -2, 1, 0, -7, -6, -5, 1, -3,
    -- filter=238 channel=72
    -8, -5, -6, -5, -4, 2, 5, -5, 5,
    -- filter=238 channel=73
    -15, -6, 0, -5, -2, 6, 0, 3, 9,
    -- filter=238 channel=74
    0, 6, 0, -5, 9, 5, -4, 2, 3,
    -- filter=238 channel=75
    3, -8, -7, -6, -18, -14, 6, -8, -2,
    -- filter=238 channel=76
    -3, 7, 3, 2, 9, 16, -14, -5, -4,
    -- filter=238 channel=77
    6, 5, -3, -2, 0, 0, 7, 3, -1,
    -- filter=238 channel=78
    5, 1, 2, 0, 4, 0, -3, -2, -6,
    -- filter=238 channel=79
    -15, -18, 1, -5, 3, 10, -7, 3, 6,
    -- filter=238 channel=80
    0, -17, -1, -11, -6, 0, -1, 3, 5,
    -- filter=238 channel=81
    0, 6, -5, 5, -4, 2, -3, 6, 6,
    -- filter=238 channel=82
    -2, -7, 4, 3, 5, 3, -6, 0, -2,
    -- filter=238 channel=83
    -2, 0, -2, -7, 1, 4, 5, 4, 9,
    -- filter=238 channel=84
    -11, 0, 4, 4, 0, 3, -1, 0, 7,
    -- filter=238 channel=85
    6, -2, 2, 6, 2, 1, 4, 2, -1,
    -- filter=238 channel=86
    4, 6, -4, 0, 0, -6, -1, 5, 2,
    -- filter=238 channel=87
    0, 9, 2, -3, 1, 4, -1, 3, -3,
    -- filter=238 channel=88
    0, 2, -5, 6, 4, -2, 2, 5, 4,
    -- filter=238 channel=89
    -6, -5, -3, -12, -6, -2, -4, 0, 10,
    -- filter=238 channel=90
    1, 5, -12, -4, 4, -5, -6, -6, 2,
    -- filter=238 channel=91
    -7, 0, 9, -4, 0, 13, 8, 11, 17,
    -- filter=238 channel=92
    0, -4, 2, 1, 1, 6, -1, -2, -6,
    -- filter=238 channel=93
    -3, -9, -8, -10, -16, -18, 0, -4, 2,
    -- filter=238 channel=94
    1, 5, -6, -2, -7, 5, 0, 2, 6,
    -- filter=238 channel=95
    -3, 0, 4, -6, 3, 6, 0, -7, -5,
    -- filter=238 channel=96
    -2, 0, 0, -8, -3, -3, 1, 0, 4,
    -- filter=238 channel=97
    -4, -3, -11, -9, -13, -9, -8, 0, -5,
    -- filter=238 channel=98
    -13, -1, 9, -8, 1, 0, -4, 9, 6,
    -- filter=238 channel=99
    -3, 3, 5, -1, 11, 4, -7, 10, 13,
    -- filter=238 channel=100
    2, -2, -2, 9, 6, 4, 8, 2, -1,
    -- filter=238 channel=101
    -5, 0, 5, -6, -12, -5, -2, 1, 9,
    -- filter=238 channel=102
    0, 2, 2, 7, 4, 0, 3, 6, -5,
    -- filter=238 channel=103
    -3, -17, -13, -1, -21, -13, -7, -9, -9,
    -- filter=238 channel=104
    -10, -6, -11, -12, -12, 2, 4, 3, 5,
    -- filter=238 channel=105
    -5, 10, 10, 7, 9, 0, -2, 5, 0,
    -- filter=238 channel=106
    1, 1, -3, -6, 2, -2, -9, -5, -3,
    -- filter=238 channel=107
    -3, 5, 1, -5, 13, 14, -4, 2, 7,
    -- filter=238 channel=108
    -3, 4, -3, 1, -5, 5, 7, -6, 6,
    -- filter=238 channel=109
    -10, -11, 2, -12, -4, 8, 3, 15, 24,
    -- filter=238 channel=110
    -7, -6, -4, 3, 0, -2, 0, 3, -3,
    -- filter=238 channel=111
    1, -1, 2, -4, -4, -3, -5, -1, -5,
    -- filter=238 channel=112
    -6, 2, 1, -1, -8, 9, 1, 3, 12,
    -- filter=238 channel=113
    -4, -6, -6, -6, 1, -6, -4, -1, 0,
    -- filter=238 channel=114
    -20, -7, 9, -10, 8, 18, 4, 9, 13,
    -- filter=238 channel=115
    1, 0, -5, -1, 2, -3, -2, 6, 7,
    -- filter=238 channel=116
    -8, -4, -2, 0, 0, 8, 5, 14, 13,
    -- filter=238 channel=117
    2, -8, -6, -4, 2, -6, -2, -5, -2,
    -- filter=238 channel=118
    7, 3, -1, -2, -3, 6, -5, -6, 4,
    -- filter=238 channel=119
    -4, 13, 1, 1, -1, 11, 6, 9, 8,
    -- filter=238 channel=120
    -9, 6, 15, 0, 4, 13, 1, 21, 15,
    -- filter=238 channel=121
    -6, -11, -1, -4, 2, 0, -3, -9, -3,
    -- filter=238 channel=122
    -6, -27, -19, -15, -28, -16, -9, -22, -17,
    -- filter=238 channel=123
    -3, 5, -3, -1, 7, 6, -8, -5, 6,
    -- filter=238 channel=124
    1, 5, 11, -6, 11, 10, -7, 0, 0,
    -- filter=238 channel=125
    0, -7, 0, -9, -6, -4, 3, 13, 15,
    -- filter=238 channel=126
    -12, -1, 2, -3, -7, 1, 1, 3, 6,
    -- filter=238 channel=127
    -2, 5, -4, 0, -6, -6, 6, -2, 5,
    -- filter=239 channel=0
    -2, -7, -15, -1, 8, 5, -18, 11, 1,
    -- filter=239 channel=1
    -3, -8, -13, 9, 12, -6, -21, 12, 1,
    -- filter=239 channel=2
    -5, -2, -1, -6, 5, -8, -7, 4, -5,
    -- filter=239 channel=3
    -4, 7, -4, -1, -10, 2, 0, 3, 2,
    -- filter=239 channel=4
    7, -2, 1, -2, 1, -8, -14, 5, 0,
    -- filter=239 channel=5
    -6, 8, -5, 1, 20, 3, -8, 16, 8,
    -- filter=239 channel=6
    6, 0, -3, 8, -4, 6, 9, 1, 6,
    -- filter=239 channel=7
    -4, 0, -1, 2, 6, 0, -3, 0, 5,
    -- filter=239 channel=8
    -11, 5, -4, -4, 2, -3, 2, -9, 1,
    -- filter=239 channel=9
    -5, -2, 6, 0, -5, 2, -3, -2, -7,
    -- filter=239 channel=10
    -10, -4, 4, -1, -13, 2, 7, -2, 0,
    -- filter=239 channel=11
    2, -4, 3, 4, -15, 1, 1, -3, 0,
    -- filter=239 channel=12
    1, -9, 8, 4, -2, 10, -6, -5, -2,
    -- filter=239 channel=13
    1, -23, 11, 17, -25, 0, 0, 10, -2,
    -- filter=239 channel=14
    -3, -2, 6, 1, -2, -3, -2, 1, 0,
    -- filter=239 channel=15
    -5, -18, 1, 14, -23, -1, 4, -6, 0,
    -- filter=239 channel=16
    -7, 11, 4, 6, 2, 6, -1, 0, 4,
    -- filter=239 channel=17
    -6, -6, 0, 0, 1, -1, -4, -2, 5,
    -- filter=239 channel=18
    7, -25, 3, 15, -17, 0, 1, 13, -8,
    -- filter=239 channel=19
    -1, -5, 1, -3, 7, 4, 4, 5, -2,
    -- filter=239 channel=20
    -7, -7, 2, 15, -20, 1, 20, -4, 3,
    -- filter=239 channel=21
    -2, 1, 3, -1, 3, -1, -8, -2, 1,
    -- filter=239 channel=22
    -13, 5, -3, 7, -6, 8, 4, -1, -7,
    -- filter=239 channel=23
    -13, 2, 13, 9, -31, 16, 26, -15, 0,
    -- filter=239 channel=24
    7, -2, 5, 2, 5, -5, -6, 3, -5,
    -- filter=239 channel=25
    -1, -17, 0, 25, -6, 4, 0, 14, -13,
    -- filter=239 channel=26
    0, 1, -7, -9, 4, 5, -16, 9, 8,
    -- filter=239 channel=27
    -15, -8, 7, 25, -26, 4, 11, 2, -16,
    -- filter=239 channel=28
    -7, -5, -2, -2, 3, 2, -5, 3, 1,
    -- filter=239 channel=29
    3, -5, 15, 13, -14, 6, 9, -5, 1,
    -- filter=239 channel=30
    0, 3, 3, 3, -8, 0, -10, 15, 4,
    -- filter=239 channel=31
    -24, 0, 5, 6, -17, 12, 9, 1, -10,
    -- filter=239 channel=32
    1, -13, 7, 23, -15, 0, 0, 15, -10,
    -- filter=239 channel=33
    -4, -4, 9, 2, -13, -1, 12, 0, -9,
    -- filter=239 channel=34
    -6, 28, 4, 0, 9, 18, 16, -8, 6,
    -- filter=239 channel=35
    -1, 0, 1, 4, 2, 0, 0, -3, 4,
    -- filter=239 channel=36
    4, -3, 1, -6, -9, -1, 1, 0, 6,
    -- filter=239 channel=37
    -10, -5, -8, -2, 7, -1, -24, 2, 1,
    -- filter=239 channel=38
    -11, -6, 5, 0, -8, 3, 5, -4, -1,
    -- filter=239 channel=39
    1, -7, 3, 0, -4, 7, 1, -1, 7,
    -- filter=239 channel=40
    -7, -11, -6, -2, -8, 4, 4, -8, -5,
    -- filter=239 channel=41
    18, -15, -3, 16, 10, -4, -17, 13, -11,
    -- filter=239 channel=42
    -2, 2, -6, 0, 3, 8, -7, 2, 4,
    -- filter=239 channel=43
    -4, -2, 0, 1, -5, 2, 16, -8, -2,
    -- filter=239 channel=44
    0, 3, 0, 2, 1, 7, -4, 7, -2,
    -- filter=239 channel=45
    -12, -3, 3, 1, -5, -7, -5, 3, -2,
    -- filter=239 channel=46
    9, 0, 0, -3, 0, -1, 2, -1, -3,
    -- filter=239 channel=47
    -8, 12, -6, -1, 17, -5, -16, 15, -7,
    -- filter=239 channel=48
    7, -8, 0, 0, 6, -4, -11, 11, -8,
    -- filter=239 channel=49
    -1, -14, 12, 11, -6, 1, -2, 7, -5,
    -- filter=239 channel=50
    -11, -4, 1, 13, -21, -3, -2, -3, -3,
    -- filter=239 channel=51
    -7, 0, 4, 5, 5, -1, -6, -4, -5,
    -- filter=239 channel=52
    -12, 6, -3, 6, -14, 10, 1, 2, -3,
    -- filter=239 channel=53
    0, 3, 11, 5, -10, 10, 6, 4, -1,
    -- filter=239 channel=54
    -1, 1, -2, -1, 0, 6, 0, -4, 1,
    -- filter=239 channel=55
    -2, -13, 17, 15, -31, -1, 6, -2, -1,
    -- filter=239 channel=56
    3, 6, 0, -4, -5, -6, 7, -5, -2,
    -- filter=239 channel=57
    12, -6, 0, 2, 11, 5, 2, 7, 4,
    -- filter=239 channel=58
    0, 11, 0, 1, 16, 7, -11, 10, 3,
    -- filter=239 channel=59
    11, -12, 9, 16, -1, -6, -11, 14, -4,
    -- filter=239 channel=60
    3, -2, -2, -4, -3, -2, 6, 4, 6,
    -- filter=239 channel=61
    6, 0, 4, 9, 3, 0, 1, 2, 1,
    -- filter=239 channel=62
    -6, 4, -1, -6, -3, 0, 4, -5, -2,
    -- filter=239 channel=63
    -3, 10, -10, 2, 17, 11, -11, 4, -1,
    -- filter=239 channel=64
    2, -7, 2, 3, 0, -1, -5, -2, 0,
    -- filter=239 channel=65
    -7, 4, -5, -7, 6, 3, -1, 0, 5,
    -- filter=239 channel=66
    2, -2, 8, 11, -1, 9, 0, 15, -8,
    -- filter=239 channel=67
    -6, -6, -3, -8, -2, -6, -5, -4, 3,
    -- filter=239 channel=68
    4, -5, 4, 6, -5, 0, -6, -5, 4,
    -- filter=239 channel=69
    -4, -6, 0, 7, 0, -6, -3, -2, 1,
    -- filter=239 channel=70
    -14, 0, 8, 5, -25, 0, 13, -6, -3,
    -- filter=239 channel=71
    -8, 7, 0, -8, -5, 6, -3, -2, -8,
    -- filter=239 channel=72
    -7, -7, 6, 15, -5, 3, 1, 3, -9,
    -- filter=239 channel=73
    1, -8, 9, 4, -3, -7, 9, 7, 6,
    -- filter=239 channel=74
    -16, -3, 7, 6, -13, 5, 14, -14, -10,
    -- filter=239 channel=75
    -10, 8, -4, 6, 5, 5, -9, 1, -2,
    -- filter=239 channel=76
    0, -8, 7, 2, -23, -4, 10, -5, -5,
    -- filter=239 channel=77
    4, 4, 0, -4, -3, -2, -1, 0, -5,
    -- filter=239 channel=78
    -10, 4, -2, -12, 8, 4, 3, -4, 10,
    -- filter=239 channel=79
    -4, -22, 11, 30, -36, 10, 1, 8, -9,
    -- filter=239 channel=80
    5, -7, 17, 14, -10, 0, 0, 14, -9,
    -- filter=239 channel=81
    6, -7, -5, 3, 1, 0, 5, -3, -3,
    -- filter=239 channel=82
    2, 8, 0, -4, 5, 0, -4, -4, 0,
    -- filter=239 channel=83
    -6, -8, 1, -4, 0, -5, -5, 10, -6,
    -- filter=239 channel=84
    0, -17, 11, 10, -14, -1, -1, 10, -4,
    -- filter=239 channel=85
    3, 2, -4, 4, -1, -1, -3, -2, 0,
    -- filter=239 channel=86
    -5, 7, 9, 6, -5, 8, 5, 7, -1,
    -- filter=239 channel=87
    -8, 6, 7, 6, -9, 5, 9, 3, 6,
    -- filter=239 channel=88
    -6, 4, -7, 1, -7, 0, -2, 1, -3,
    -- filter=239 channel=89
    3, -20, 18, 8, -29, 9, 2, -4, -12,
    -- filter=239 channel=90
    -6, 10, 4, -13, -10, 8, 0, -10, -2,
    -- filter=239 channel=91
    2, -17, 14, 18, -25, 0, 7, 9, -7,
    -- filter=239 channel=92
    -4, 6, 2, 6, 7, 5, 7, 3, 3,
    -- filter=239 channel=93
    -4, 8, -10, -3, 15, 4, -14, 6, 4,
    -- filter=239 channel=94
    -4, -6, -2, 0, -4, -5, 2, -6, 3,
    -- filter=239 channel=95
    0, 4, -6, -4, -6, 7, 7, -10, 3,
    -- filter=239 channel=96
    5, -1, -4, -4, -7, 0, 0, 0, 5,
    -- filter=239 channel=97
    -4, -2, 6, -14, -1, 7, 0, -4, -5,
    -- filter=239 channel=98
    -5, -12, 7, 7, -20, 8, 5, 4, 0,
    -- filter=239 channel=99
    -15, 1, 17, 14, -23, 10, 27, 0, -4,
    -- filter=239 channel=100
    6, 8, -4, 4, 10, -1, -4, -2, 9,
    -- filter=239 channel=101
    4, -12, 5, -2, 0, -5, -6, 10, -3,
    -- filter=239 channel=102
    -2, -6, 7, 0, 2, 5, -3, -3, -3,
    -- filter=239 channel=103
    -13, 17, -1, -10, 7, -2, 2, 9, -2,
    -- filter=239 channel=104
    0, -8, 1, 7, 2, -7, -4, 10, -6,
    -- filter=239 channel=105
    4, 2, 9, 3, -9, 7, 3, -2, 0,
    -- filter=239 channel=106
    9, -11, -8, 2, 0, -8, 3, -5, 3,
    -- filter=239 channel=107
    -9, -10, 7, 0, -19, 7, 11, -15, 4,
    -- filter=239 channel=108
    2, 5, 0, 8, 14, 0, -7, 2, 7,
    -- filter=239 channel=109
    8, -11, 13, 23, -19, 6, 7, 17, -12,
    -- filter=239 channel=110
    -8, -2, 15, 8, -9, 19, 2, -2, 9,
    -- filter=239 channel=111
    4, 1, 0, 8, 10, -6, 0, 0, 2,
    -- filter=239 channel=112
    -20, 2, -2, 0, -13, 0, -1, -2, -9,
    -- filter=239 channel=113
    -4, 1, 11, 7, -15, 1, 5, 3, -3,
    -- filter=239 channel=114
    3, -24, 1, 17, -6, 1, 3, 21, -3,
    -- filter=239 channel=115
    -6, 6, -5, 8, -6, -2, 3, 0, -6,
    -- filter=239 channel=116
    11, -8, 13, 24, -9, -2, -5, 19, 0,
    -- filter=239 channel=117
    -4, -11, 6, 7, 0, 2, -6, 2, 0,
    -- filter=239 channel=118
    2, 2, 0, -5, 0, -3, -3, -5, -2,
    -- filter=239 channel=119
    -7, 22, 2, 3, 10, -3, 16, -9, 1,
    -- filter=239 channel=120
    -20, -9, 7, -3, -40, 8, 16, -15, 1,
    -- filter=239 channel=121
    -1, -11, 1, 5, -11, -2, 4, 1, 0,
    -- filter=239 channel=122
    0, 17, -11, 2, 12, 7, -17, 4, -4,
    -- filter=239 channel=123
    -7, 7, 7, 1, 10, 9, 14, -8, 5,
    -- filter=239 channel=124
    0, -3, 4, 9, -3, 3, 6, -7, 0,
    -- filter=239 channel=125
    5, -9, 6, 20, -20, 5, 7, 6, 0,
    -- filter=239 channel=126
    -2, -8, 2, 9, -4, -4, -7, -3, -10,
    -- filter=239 channel=127
    0, -8, -6, 1, 1, -3, -5, -3, -1,
    -- filter=240 channel=0
    3, -9, -17, -5, -2, -5, 14, -4, -9,
    -- filter=240 channel=1
    4, 6, -13, -4, 1, -1, 17, 10, -4,
    -- filter=240 channel=2
    -2, 4, -2, 0, -3, 4, -2, 3, 6,
    -- filter=240 channel=3
    -9, -13, 0, -9, -17, -1, -4, -4, -2,
    -- filter=240 channel=4
    -4, -8, 0, 4, -13, 3, -3, -17, 2,
    -- filter=240 channel=5
    1, 4, -1, 5, 7, -5, 2, 6, -11,
    -- filter=240 channel=6
    -2, 8, 5, 1, -3, -2, -2, 5, -4,
    -- filter=240 channel=7
    3, -1, 0, -2, 0, -2, -2, -6, 5,
    -- filter=240 channel=8
    -7, 3, -3, 7, -2, -2, 2, 0, -5,
    -- filter=240 channel=9
    -1, 1, -8, -5, 4, 4, -3, -6, -8,
    -- filter=240 channel=10
    -3, 8, 5, -15, 16, 3, 0, -3, 2,
    -- filter=240 channel=11
    0, -5, 8, -2, -6, -3, -2, -11, 1,
    -- filter=240 channel=12
    3, 10, -4, 10, 9, 3, 17, 11, 2,
    -- filter=240 channel=13
    -9, 12, -2, -1, 11, -2, 0, 0, 1,
    -- filter=240 channel=14
    -3, 0, -3, -5, -4, 0, -4, 6, -6,
    -- filter=240 channel=15
    -3, 0, -2, -4, 1, -12, 5, 3, 2,
    -- filter=240 channel=16
    4, 8, 3, -6, 13, 4, -9, 6, -3,
    -- filter=240 channel=17
    2, 6, 4, 3, -4, 6, 5, 5, -3,
    -- filter=240 channel=18
    0, 12, -5, 3, 15, -12, 16, 0, 0,
    -- filter=240 channel=19
    -4, -1, 3, 6, -6, 6, 3, 5, -6,
    -- filter=240 channel=20
    1, 2, -4, -4, -5, 0, -1, -1, 4,
    -- filter=240 channel=21
    -9, 15, 9, -15, 19, 4, -7, 7, 1,
    -- filter=240 channel=22
    6, 1, -8, 2, 0, -1, 9, 7, -1,
    -- filter=240 channel=23
    0, 8, 5, -8, 18, -10, -15, 10, -12,
    -- filter=240 channel=24
    -5, -6, -2, 5, 6, -1, -2, 0, 4,
    -- filter=240 channel=25
    -14, 27, -11, -19, 26, -12, 3, 14, -2,
    -- filter=240 channel=26
    -2, 10, 0, -7, 4, 4, 0, 0, 1,
    -- filter=240 channel=27
    -11, 22, -16, -14, 35, -7, -2, 13, 0,
    -- filter=240 channel=28
    7, 2, 3, 0, -2, 5, 4, -6, 4,
    -- filter=240 channel=29
    0, -1, 0, 2, -7, 5, 7, -6, -4,
    -- filter=240 channel=30
    -10, 4, 0, -6, 17, -3, 0, -3, -5,
    -- filter=240 channel=31
    -15, 14, -2, -32, 29, -5, -32, 0, -11,
    -- filter=240 channel=32
    -3, 12, -13, -6, 25, -2, 3, -1, -12,
    -- filter=240 channel=33
    -7, 5, -11, -10, 14, -2, 0, 9, 0,
    -- filter=240 channel=34
    13, 6, -3, 21, 24, -6, -2, 10, -10,
    -- filter=240 channel=35
    -6, 5, 3, 0, 6, 1, 2, 0, -1,
    -- filter=240 channel=36
    -2, 3, -4, -6, 4, 0, 6, -3, -3,
    -- filter=240 channel=37
    7, -7, -7, 4, 11, -10, 12, 1, -10,
    -- filter=240 channel=38
    -10, 4, -2, -8, 14, 1, -2, -4, -1,
    -- filter=240 channel=39
    6, -4, -4, -6, -10, -4, 0, 0, -4,
    -- filter=240 channel=40
    4, -6, -2, -3, 1, 0, -6, 4, 1,
    -- filter=240 channel=41
    11, 21, -17, 27, 12, 0, 26, 11, -10,
    -- filter=240 channel=42
    3, 0, 9, -3, -3, 10, 0, 0, 8,
    -- filter=240 channel=43
    -3, -9, -9, -6, -3, 1, -1, -6, -9,
    -- filter=240 channel=44
    -5, 8, -8, -7, 17, -7, -3, 3, -11,
    -- filter=240 channel=45
    -4, 5, -1, -4, -6, -5, -6, 0, 0,
    -- filter=240 channel=46
    -3, -6, 4, 3, 2, -6, -2, 2, -5,
    -- filter=240 channel=47
    -7, 12, -1, -9, 24, -3, -6, 2, 1,
    -- filter=240 channel=48
    -12, 17, 4, -22, 22, -6, -1, -3, 6,
    -- filter=240 channel=49
    -8, -1, 2, 2, -8, 2, 1, 0, -1,
    -- filter=240 channel=50
    -6, 8, -5, -12, 14, -7, -12, 8, -7,
    -- filter=240 channel=51
    1, 3, 2, 3, -6, 2, -3, 5, 2,
    -- filter=240 channel=52
    0, 14, -9, 6, 10, 1, 0, 1, 0,
    -- filter=240 channel=53
    -6, 0, 0, -4, 1, -1, -4, 0, 5,
    -- filter=240 channel=54
    1, -5, 2, -2, 0, 3, -6, -1, -2,
    -- filter=240 channel=55
    -7, 9, 0, -11, 11, -2, 3, -2, -8,
    -- filter=240 channel=56
    1, 4, 8, 5, 11, 0, 6, 7, -7,
    -- filter=240 channel=57
    5, 8, -1, 9, -6, 7, 8, 7, 1,
    -- filter=240 channel=58
    9, -5, 4, -2, 0, -5, 9, -1, 6,
    -- filter=240 channel=59
    -13, 19, 1, -23, 26, 1, -6, 1, -2,
    -- filter=240 channel=60
    1, 4, 0, -6, -7, -7, 6, 3, 6,
    -- filter=240 channel=61
    7, 12, -8, -5, 17, 5, 2, 5, 6,
    -- filter=240 channel=62
    0, -3, 0, 4, 3, -5, -3, -4, 0,
    -- filter=240 channel=63
    4, 5, -4, -4, 3, 4, 7, -1, -7,
    -- filter=240 channel=64
    6, 7, 4, -2, 3, 5, -4, -3, -7,
    -- filter=240 channel=65
    1, 3, -5, 0, 2, -2, 1, -2, 1,
    -- filter=240 channel=66
    9, 24, -18, 13, 26, 0, 19, 23, -2,
    -- filter=240 channel=67
    6, 3, -6, 0, 4, 2, 0, -4, 1,
    -- filter=240 channel=68
    2, -6, -4, -2, 0, 4, -5, 0, 5,
    -- filter=240 channel=69
    1, -1, -2, -2, 7, -1, 2, -3, 0,
    -- filter=240 channel=70
    8, -2, 0, -9, 8, -7, 4, 0, 0,
    -- filter=240 channel=71
    0, -11, 5, -11, -1, -2, -6, -1, 2,
    -- filter=240 channel=72
    -11, 9, 3, -17, 16, -1, -13, -2, -3,
    -- filter=240 channel=73
    -4, 9, -5, -11, 5, -1, -2, 5, -4,
    -- filter=240 channel=74
    -1, 12, -11, 1, 31, -22, -3, 14, -17,
    -- filter=240 channel=75
    6, 0, -14, 1, 3, -10, 9, 2, -4,
    -- filter=240 channel=76
    0, -6, -7, 5, -10, 0, 5, -9, 3,
    -- filter=240 channel=77
    -4, 1, 6, 1, 1, -1, 0, 7, -7,
    -- filter=240 channel=78
    8, -4, -7, 2, 2, 3, 4, 3, 0,
    -- filter=240 channel=79
    -12, 23, -12, -16, 24, -10, 2, 12, -2,
    -- filter=240 channel=80
    -23, 27, -3, -36, 34, 5, -17, 6, -6,
    -- filter=240 channel=81
    -5, 1, 0, 7, 7, 1, -2, -3, -6,
    -- filter=240 channel=82
    7, -3, -5, 1, -4, 6, -6, 2, -8,
    -- filter=240 channel=83
    -13, 9, 0, -12, 7, 0, -6, 1, 3,
    -- filter=240 channel=84
    1, 15, 0, 4, 16, -5, 2, -1, -6,
    -- filter=240 channel=85
    7, -2, 6, -2, -6, 5, 2, 3, 2,
    -- filter=240 channel=86
    5, 10, -12, -8, 11, -1, 2, 9, 0,
    -- filter=240 channel=87
    5, 10, 0, 1, 5, -6, -1, 4, -2,
    -- filter=240 channel=88
    -8, -1, 3, 1, 16, -2, -1, 6, -6,
    -- filter=240 channel=89
    -4, 10, -4, -25, 11, -1, 0, -3, 0,
    -- filter=240 channel=90
    1, 5, 0, -8, 16, -1, -17, -2, -8,
    -- filter=240 channel=91
    -14, 11, -7, -16, 8, 2, 4, 4, 0,
    -- filter=240 channel=92
    5, -7, 0, 9, 3, -6, 3, -2, -2,
    -- filter=240 channel=93
    -5, 7, -9, -5, 9, -5, 7, 0, -8,
    -- filter=240 channel=94
    -6, -3, 2, 0, -2, -2, 5, -1, 5,
    -- filter=240 channel=95
    1, 3, 6, 0, 5, 0, 3, 2, -2,
    -- filter=240 channel=96
    -4, -4, -5, -7, -4, -2, -1, -7, 2,
    -- filter=240 channel=97
    -8, -4, -3, -2, 1, -2, -3, 4, 4,
    -- filter=240 channel=98
    -15, 23, -1, -25, 26, -13, -1, 14, -11,
    -- filter=240 channel=99
    -10, 23, -11, -17, 37, -18, -20, 7, -7,
    -- filter=240 channel=100
    10, 0, -4, 11, 10, 1, 10, 4, 0,
    -- filter=240 channel=101
    -9, 0, 4, 0, -15, 0, 3, -1, -8,
    -- filter=240 channel=102
    -7, 6, -6, -6, -4, -4, 1, 7, 0,
    -- filter=240 channel=103
    -7, 2, -7, -8, 21, 3, -6, 0, -2,
    -- filter=240 channel=104
    -11, 22, -5, -27, 21, -2, -11, 8, 6,
    -- filter=240 channel=105
    8, 1, 6, -2, -1, 8, 1, 6, -6,
    -- filter=240 channel=106
    7, -5, 1, 10, -5, -3, -5, 1, -5,
    -- filter=240 channel=107
    13, 0, -8, 6, 3, -11, 10, 6, -6,
    -- filter=240 channel=108
    1, 4, -11, 7, 1, -7, 5, -2, -3,
    -- filter=240 channel=109
    -6, 17, -7, -17, 26, -7, 8, 10, 0,
    -- filter=240 channel=110
    -6, 4, 2, -14, 13, -2, -8, -2, -1,
    -- filter=240 channel=111
    0, 4, -5, 3, 5, -6, 9, 6, 0,
    -- filter=240 channel=112
    0, 8, -3, -4, 4, -16, -10, 7, 0,
    -- filter=240 channel=113
    -3, 9, 5, -14, 20, 3, 0, 1, -2,
    -- filter=240 channel=114
    5, 9, -10, -5, 6, -17, 8, 11, -11,
    -- filter=240 channel=115
    1, -3, -1, 4, -4, -1, -5, 5, 1,
    -- filter=240 channel=116
    -16, 13, -1, -20, 8, 6, -1, 4, -2,
    -- filter=240 channel=117
    -8, 7, 2, -8, 1, -1, 0, -4, 0,
    -- filter=240 channel=118
    5, 7, -5, -1, 0, -3, 5, 0, 0,
    -- filter=240 channel=119
    19, 1, -3, 13, 11, 7, 9, 18, -10,
    -- filter=240 channel=120
    -9, 14, -15, -17, 16, -20, -3, 2, -9,
    -- filter=240 channel=121
    0, 16, -3, 0, 15, 4, 2, 6, 3,
    -- filter=240 channel=122
    -10, 26, -3, -24, 32, 5, -11, 3, 2,
    -- filter=240 channel=123
    15, 8, -2, 0, 4, 6, 2, 4, 1,
    -- filter=240 channel=124
    -1, 2, 6, -5, 6, 5, -6, -7, 2,
    -- filter=240 channel=125
    -9, 29, -9, -23, 24, -2, -13, 8, -2,
    -- filter=240 channel=126
    -9, 9, 0, -9, 2, 2, -5, -5, -6,
    -- filter=240 channel=127
    0, -1, 3, 8, 1, 2, 7, 3, 1,
    -- filter=241 channel=0
    -2, 3, 5, -8, -8, 10, -6, -6, 14,
    -- filter=241 channel=1
    1, -6, 8, -19, -8, 12, -6, -5, 4,
    -- filter=241 channel=2
    0, -1, 3, -1, -1, 7, 2, 3, -3,
    -- filter=241 channel=3
    1, 1, 2, -8, -6, -2, -6, 0, 4,
    -- filter=241 channel=4
    0, -2, 0, -3, -3, 8, 4, -10, -2,
    -- filter=241 channel=5
    -4, -4, 5, -9, -14, 12, 0, 7, 8,
    -- filter=241 channel=6
    1, 5, -3, 13, 0, 5, 5, -2, -3,
    -- filter=241 channel=7
    -5, -6, 2, -5, -6, 6, -1, 2, 0,
    -- filter=241 channel=8
    3, 4, 3, -3, -3, 5, -2, 3, -3,
    -- filter=241 channel=9
    0, 4, 0, -11, -3, 0, 0, 7, 1,
    -- filter=241 channel=10
    2, 0, 4, 4, 5, -5, 1, -9, -3,
    -- filter=241 channel=11
    -7, 2, -10, 6, 8, 0, -5, 0, -9,
    -- filter=241 channel=12
    0, 0, -2, 11, 1, 0, 8, -2, 1,
    -- filter=241 channel=13
    3, -4, -1, 6, 2, -7, 8, -8, 1,
    -- filter=241 channel=14
    0, 5, -5, -2, -1, -7, 0, 1, -7,
    -- filter=241 channel=15
    -3, -4, -5, 10, 15, -1, 6, 5, -14,
    -- filter=241 channel=16
    5, -1, 4, -9, -6, 6, -8, -4, 4,
    -- filter=241 channel=17
    2, 5, -4, 4, 1, 0, 3, -4, -4,
    -- filter=241 channel=18
    -8, 0, -2, 6, 21, -1, 5, 6, -3,
    -- filter=241 channel=19
    -3, -2, 1, 5, -2, 0, 2, 3, 5,
    -- filter=241 channel=20
    2, -2, -2, 16, 18, -12, 0, 8, -17,
    -- filter=241 channel=21
    -6, -6, 12, -15, -9, 14, -2, -7, 10,
    -- filter=241 channel=22
    -7, 1, 4, -6, 3, 0, -4, 10, -2,
    -- filter=241 channel=23
    2, 0, -9, 9, 9, -10, 7, 11, -13,
    -- filter=241 channel=24
    -3, -3, -7, 0, -1, -7, 1, 1, -6,
    -- filter=241 channel=25
    -2, -2, 3, -9, 6, 10, 2, -1, 10,
    -- filter=241 channel=26
    1, -2, 0, -10, -1, 0, -3, 4, 6,
    -- filter=241 channel=27
    -5, 2, -7, -11, 8, 3, 0, 5, 5,
    -- filter=241 channel=28
    2, 0, 3, -2, 2, 4, 6, -3, 0,
    -- filter=241 channel=29
    -3, 6, -6, 4, 19, -2, -1, -1, -4,
    -- filter=241 channel=30
    2, -4, 2, -13, -7, 3, -11, 4, 10,
    -- filter=241 channel=31
    1, -1, 0, -22, -6, 3, -7, -5, 5,
    -- filter=241 channel=32
    -9, -6, -5, -1, 14, 5, 0, 8, 2,
    -- filter=241 channel=33
    2, -8, 4, -6, 3, 5, -6, 5, 3,
    -- filter=241 channel=34
    4, 2, 0, 10, 9, -8, 0, 11, 2,
    -- filter=241 channel=35
    5, -1, 6, 0, 2, -7, -2, -3, -2,
    -- filter=241 channel=36
    2, 4, 6, -6, -3, -1, 5, 1, 0,
    -- filter=241 channel=37
    -10, -11, 4, -8, -17, 8, -2, -12, 15,
    -- filter=241 channel=38
    0, 5, 6, -10, -2, 1, -5, 6, 2,
    -- filter=241 channel=39
    -8, 2, 3, 6, 0, -2, 1, 1, -4,
    -- filter=241 channel=40
    -9, -7, -5, 0, 8, -7, -2, 7, -11,
    -- filter=241 channel=41
    0, -1, 13, 6, 1, 3, 0, -5, -1,
    -- filter=241 channel=42
    -8, -3, 7, 0, -9, 7, -6, -5, 7,
    -- filter=241 channel=43
    -3, 0, 0, 9, -4, -8, 4, 8, 1,
    -- filter=241 channel=44
    -3, -4, 6, -21, -5, 0, -14, -10, 0,
    -- filter=241 channel=45
    3, -2, 0, 3, -5, -4, -7, 2, -2,
    -- filter=241 channel=46
    0, -3, 3, 5, 7, -4, 2, -1, 0,
    -- filter=241 channel=47
    1, -4, 11, -23, -16, 5, -13, -7, 11,
    -- filter=241 channel=48
    -3, 2, 12, -17, -4, 10, -12, -4, 5,
    -- filter=241 channel=49
    -1, 2, -10, 5, 1, 4, 0, -3, 0,
    -- filter=241 channel=50
    0, -4, -1, -3, -2, 7, 0, -5, 8,
    -- filter=241 channel=51
    -4, -4, -5, 2, -2, 2, -1, -7, -7,
    -- filter=241 channel=52
    -4, 3, -5, -2, 9, 4, 1, 4, -4,
    -- filter=241 channel=53
    -5, -3, -8, 2, 3, -1, 6, 3, -10,
    -- filter=241 channel=54
    3, -4, 2, 3, -6, 1, -3, 3, 6,
    -- filter=241 channel=55
    1, -4, -5, 0, 16, -13, 0, -1, -17,
    -- filter=241 channel=56
    2, 7, -1, 3, 4, -5, 7, 1, 0,
    -- filter=241 channel=57
    -3, -7, 7, 0, -5, -2, 1, 3, 0,
    -- filter=241 channel=58
    4, -4, 3, -8, -3, -3, -4, 4, 5,
    -- filter=241 channel=59
    -7, 0, 3, -7, -1, 7, -5, -9, 10,
    -- filter=241 channel=60
    2, 1, -4, -7, 7, -5, -6, 6, -1,
    -- filter=241 channel=61
    6, 6, -2, 7, -2, 0, 5, -2, -5,
    -- filter=241 channel=62
    3, 1, 1, 6, 1, -6, 4, -4, 6,
    -- filter=241 channel=63
    2, 8, 10, -1, -4, 2, -5, -6, 6,
    -- filter=241 channel=64
    0, -7, 4, -4, 6, 5, -2, 4, -3,
    -- filter=241 channel=65
    0, 0, 0, -2, -2, 5, 7, 4, -3,
    -- filter=241 channel=66
    6, 5, 7, 0, -2, 7, 5, -1, 7,
    -- filter=241 channel=67
    -2, 0, 3, -5, -4, -1, 3, 6, 2,
    -- filter=241 channel=68
    1, -6, -3, -2, 6, 3, 0, -4, -9,
    -- filter=241 channel=69
    -5, -2, 5, 1, -2, 7, 0, -5, 0,
    -- filter=241 channel=70
    -7, 5, -8, 0, 2, -1, -4, 6, -9,
    -- filter=241 channel=71
    -3, 1, 0, -4, -7, 4, -1, -3, 0,
    -- filter=241 channel=72
    -4, -10, -3, -8, -10, -1, -1, -2, 3,
    -- filter=241 channel=73
    3, 1, 2, 5, 3, 5, -1, -2, -12,
    -- filter=241 channel=74
    2, -2, -3, -9, 0, 0, 1, -8, 0,
    -- filter=241 channel=75
    -9, -4, 11, -24, -16, -1, -1, 0, 23,
    -- filter=241 channel=76
    -7, -1, -7, 10, 7, -12, 8, 0, -11,
    -- filter=241 channel=77
    1, -1, 4, 0, -4, 7, 2, 0, -1,
    -- filter=241 channel=78
    -2, 0, 3, -8, 1, 0, -7, -4, 9,
    -- filter=241 channel=79
    3, -9, -12, 0, 5, -5, -7, 2, -13,
    -- filter=241 channel=80
    1, -3, 8, -9, -14, 12, -5, 0, 4,
    -- filter=241 channel=81
    4, -2, 1, 3, -3, -2, 0, 7, -2,
    -- filter=241 channel=82
    0, -8, 3, 4, 2, -8, 0, 2, 6,
    -- filter=241 channel=83
    1, -4, -1, -5, 3, 2, 2, -4, 9,
    -- filter=241 channel=84
    -2, -6, -2, 6, 2, -4, 3, 5, 2,
    -- filter=241 channel=85
    3, -2, 4, -6, 1, 0, -5, -7, -6,
    -- filter=241 channel=86
    0, 0, 4, -4, 1, 5, -4, -6, -1,
    -- filter=241 channel=87
    4, 1, -6, 11, 5, 0, -4, -4, 0,
    -- filter=241 channel=88
    -2, 3, -1, -4, 1, 5, 3, -3, 5,
    -- filter=241 channel=89
    5, -13, -8, 6, 4, -1, 9, 0, -5,
    -- filter=241 channel=90
    1, 2, 3, 2, 1, 6, 1, -6, -4,
    -- filter=241 channel=91
    4, -6, 0, -2, 8, -6, 5, 0, -5,
    -- filter=241 channel=92
    -1, 4, 5, 4, -5, -6, 1, 6, -3,
    -- filter=241 channel=93
    -8, -3, 2, -16, -6, 5, -6, 0, 11,
    -- filter=241 channel=94
    -5, 0, 0, -4, 5, 2, 2, 6, -1,
    -- filter=241 channel=95
    -4, 3, 0, 2, 5, 6, 1, 0, -1,
    -- filter=241 channel=96
    4, 0, -6, 5, -6, 2, 5, 2, 0,
    -- filter=241 channel=97
    -9, -7, -1, -4, 0, 7, 3, 0, 4,
    -- filter=241 channel=98
    -4, -5, 4, -17, 5, 2, -10, 0, 10,
    -- filter=241 channel=99
    -1, -3, 1, 0, -1, 7, -5, -3, 0,
    -- filter=241 channel=100
    4, -1, 3, -3, 1, 5, -2, 4, 2,
    -- filter=241 channel=101
    3, -6, -5, -8, 6, 0, 0, 0, 1,
    -- filter=241 channel=102
    6, -3, 4, -4, 2, 1, -3, -4, 6,
    -- filter=241 channel=103
    0, -6, 11, -10, -6, 8, -8, -7, 18,
    -- filter=241 channel=104
    -5, 3, 9, -13, -1, 10, -6, 0, 0,
    -- filter=241 channel=105
    -8, -2, -7, 13, 3, -6, 9, 4, -2,
    -- filter=241 channel=106
    -3, -5, 1, 6, 3, -3, 0, -3, -1,
    -- filter=241 channel=107
    -4, 0, 1, 11, 15, 1, 3, 6, -2,
    -- filter=241 channel=108
    3, 0, 0, 0, -7, 4, -1, -2, 0,
    -- filter=241 channel=109
    3, 7, 2, -3, 14, 0, 3, 10, 0,
    -- filter=241 channel=110
    -6, 0, -4, -4, -12, 1, 0, -6, 6,
    -- filter=241 channel=111
    -2, 0, 5, -4, -1, -2, -2, 5, -1,
    -- filter=241 channel=112
    1, 6, 0, -8, -4, 1, 2, -1, -1,
    -- filter=241 channel=113
    3, 3, 5, -3, -5, 0, 0, 5, 0,
    -- filter=241 channel=114
    -10, 11, -1, 3, 8, 4, 1, -1, -3,
    -- filter=241 channel=115
    7, -5, -4, 5, -5, -6, 2, -7, 3,
    -- filter=241 channel=116
    -1, 2, 0, -5, 0, -2, -3, -7, 0,
    -- filter=241 channel=117
    -2, -4, -3, -7, -6, -2, 0, -7, -3,
    -- filter=241 channel=118
    -3, -3, -6, 4, 6, 0, -4, 2, -2,
    -- filter=241 channel=119
    0, 5, -3, 14, 10, 8, 1, 13, 6,
    -- filter=241 channel=120
    -8, -4, 2, 1, 10, -2, -11, -8, 0,
    -- filter=241 channel=121
    -6, 0, 5, -3, -6, 0, -4, 5, 6,
    -- filter=241 channel=122
    -5, -9, 8, -24, -21, 12, -24, -6, 12,
    -- filter=241 channel=123
    0, -5, 2, 2, 10, 6, -1, 7, 0,
    -- filter=241 channel=124
    1, -3, -7, 2, -1, -9, -3, -2, -3,
    -- filter=241 channel=125
    -1, -9, 5, -3, 1, 3, 2, -2, 3,
    -- filter=241 channel=126
    5, -4, 3, -5, 0, 2, -4, 5, 4,
    -- filter=241 channel=127
    3, 1, 7, -7, 2, 2, -2, 5, 6,
    -- filter=242 channel=0
    13, -3, -7, -6, -24, -14, 2, -15, -20,
    -- filter=242 channel=1
    1, -13, -9, -2, -29, -18, -13, -22, -12,
    -- filter=242 channel=2
    -6, 2, 1, 0, 1, -5, 3, 0, -6,
    -- filter=242 channel=3
    6, 9, 2, -5, 3, -6, 1, 3, 2,
    -- filter=242 channel=4
    -10, -16, -11, -20, -15, -7, -8, -4, -7,
    -- filter=242 channel=5
    7, -4, 5, 1, -9, -10, -10, -9, -5,
    -- filter=242 channel=6
    -11, -11, -7, -8, 1, -3, 2, 11, 8,
    -- filter=242 channel=7
    -5, 4, 3, 4, -2, 2, 7, 4, 0,
    -- filter=242 channel=8
    -10, 0, 5, -6, -1, 2, 0, -3, 2,
    -- filter=242 channel=9
    0, 2, 5, -5, 4, -4, 0, -7, -6,
    -- filter=242 channel=10
    7, 15, 9, 7, 8, 7, -6, 0, 7,
    -- filter=242 channel=11
    -4, -2, -3, 2, 14, 8, 6, 10, 5,
    -- filter=242 channel=12
    -6, -4, -3, -2, 0, 7, -2, -1, -3,
    -- filter=242 channel=13
    6, -2, 7, 3, 0, 4, 3, -8, 1,
    -- filter=242 channel=14
    3, -2, -3, 3, 6, 0, -7, -7, -2,
    -- filter=242 channel=15
    -1, -8, -4, 0, -4, 0, 0, 11, 6,
    -- filter=242 channel=16
    4, 6, 1, 0, 4, -1, -13, -14, -10,
    -- filter=242 channel=17
    4, -5, -7, -6, -5, 1, -2, 6, 3,
    -- filter=242 channel=18
    4, -10, -13, 2, -14, 5, 7, 4, 10,
    -- filter=242 channel=19
    -1, -2, -5, 3, 5, -3, 3, -6, 4,
    -- filter=242 channel=20
    -14, -15, -4, -2, 20, 19, 4, 30, 27,
    -- filter=242 channel=21
    8, 14, 14, 0, 9, -3, -11, -16, -10,
    -- filter=242 channel=22
    1, -7, -10, -6, 1, -3, 3, -7, 3,
    -- filter=242 channel=23
    3, 3, 0, -8, 8, 5, -1, 6, 8,
    -- filter=242 channel=24
    5, 1, -2, -5, -3, -2, 2, -6, 5,
    -- filter=242 channel=25
    1, 4, 0, 2, -10, 4, -12, -12, -9,
    -- filter=242 channel=26
    4, 6, 10, -5, -3, 1, 0, 0, -6,
    -- filter=242 channel=27
    15, 0, -11, -7, -12, -5, -5, -10, -10,
    -- filter=242 channel=28
    1, 5, -2, -2, 0, -5, -3, -3, 1,
    -- filter=242 channel=29
    -4, -12, -9, 5, 9, 20, 0, 15, 15,
    -- filter=242 channel=30
    9, 7, -5, 0, -9, -2, -4, -13, -9,
    -- filter=242 channel=31
    17, 31, 8, 3, 14, -4, -7, -9, -2,
    -- filter=242 channel=32
    -2, -13, -9, 0, -15, 7, -2, 1, -1,
    -- filter=242 channel=33
    19, 4, 7, 6, -9, -5, -2, -16, 2,
    -- filter=242 channel=34
    -4, -10, 4, -5, -6, -9, -17, -3, 4,
    -- filter=242 channel=35
    -2, 5, -1, -3, -1, 5, -1, -5, 0,
    -- filter=242 channel=36
    0, -7, 5, 0, 0, 5, -5, 10, 1,
    -- filter=242 channel=37
    -4, -7, 1, -14, -16, -18, -9, -25, -23,
    -- filter=242 channel=38
    10, 4, 8, 3, 7, -4, -8, 3, 0,
    -- filter=242 channel=39
    -11, -11, -2, 0, 2, 12, -1, 7, 10,
    -- filter=242 channel=40
    -10, -10, -7, 7, 4, 4, -6, 10, 6,
    -- filter=242 channel=41
    -3, -16, 9, 1, -12, -1, 4, -4, 8,
    -- filter=242 channel=42
    4, 6, 4, -7, -9, -5, -4, -5, -10,
    -- filter=242 channel=43
    13, -2, 1, 8, 5, -7, -3, 3, 3,
    -- filter=242 channel=44
    4, 5, 0, -2, -5, -13, -6, -6, -4,
    -- filter=242 channel=45
    -7, 2, 1, 2, 3, 4, -2, -7, -5,
    -- filter=242 channel=46
    2, 3, 5, -2, 0, -9, -1, -6, 0,
    -- filter=242 channel=47
    15, 8, 13, -6, -13, 0, -7, -18, -18,
    -- filter=242 channel=48
    0, -2, 0, 1, -10, -14, -10, -14, -13,
    -- filter=242 channel=49
    -9, -13, -12, -4, -5, 1, -4, 6, -6,
    -- filter=242 channel=50
    4, 4, 0, 6, 5, -1, -1, 3, -6,
    -- filter=242 channel=51
    1, -6, 0, 3, -3, -2, -4, -2, 0,
    -- filter=242 channel=52
    0, -4, 2, -4, -8, 5, -3, 7, 1,
    -- filter=242 channel=53
    -6, -7, -7, -3, -2, 4, 3, 11, 5,
    -- filter=242 channel=54
    0, -4, 4, -6, -6, -6, -5, -5, 0,
    -- filter=242 channel=55
    -1, 2, -4, 1, 1, 11, 10, 14, 18,
    -- filter=242 channel=56
    3, 3, 4, -8, 2, -1, 0, 8, -7,
    -- filter=242 channel=57
    3, 0, 0, -3, -2, 3, 6, 5, -3,
    -- filter=242 channel=58
    -5, -6, -5, 0, -11, -8, 2, 0, 0,
    -- filter=242 channel=59
    5, 14, 2, 8, -2, -8, -2, -13, -10,
    -- filter=242 channel=60
    -4, -6, 1, -5, 4, 5, 0, 5, -6,
    -- filter=242 channel=61
    -3, -1, -4, 0, 4, 8, -5, -2, 0,
    -- filter=242 channel=62
    0, 0, 7, -4, 4, -1, 5, 8, 3,
    -- filter=242 channel=63
    0, 7, 10, -1, -3, -3, -4, -5, -8,
    -- filter=242 channel=64
    0, 0, 3, -2, 9, 3, 4, 8, -5,
    -- filter=242 channel=65
    7, 5, -4, 5, 0, 3, -6, 5, -3,
    -- filter=242 channel=66
    1, -3, 2, 0, 0, 5, 9, 0, 8,
    -- filter=242 channel=67
    -1, -3, -2, 0, 2, -5, 7, 3, -7,
    -- filter=242 channel=68
    -9, 0, -5, 6, 0, 0, -6, 6, -3,
    -- filter=242 channel=69
    1, 5, 2, 6, -4, 3, 7, -4, 3,
    -- filter=242 channel=70
    7, 5, 0, -3, -14, -2, -17, -6, -8,
    -- filter=242 channel=71
    3, 8, 5, 4, -3, 6, -2, -1, -3,
    -- filter=242 channel=72
    15, 21, 13, 11, 12, 2, 1, 4, -1,
    -- filter=242 channel=73
    -5, -1, -6, -8, 0, 5, 0, 3, -6,
    -- filter=242 channel=74
    -5, -2, 4, -2, 0, 2, -1, 1, 0,
    -- filter=242 channel=75
    3, 8, 1, -6, -11, -14, -6, -29, -6,
    -- filter=242 channel=76
    -5, -16, -5, 6, 12, 9, 10, 16, 11,
    -- filter=242 channel=77
    -4, -6, 4, -4, 2, 0, 0, 4, -6,
    -- filter=242 channel=78
    2, -1, 4, 0, 2, -6, 0, 0, 2,
    -- filter=242 channel=79
    8, -5, 2, 0, -12, 2, 5, -13, 7,
    -- filter=242 channel=80
    17, 28, 18, 8, -1, 1, 1, -18, 0,
    -- filter=242 channel=81
    6, -6, -5, -6, -3, 5, 0, -4, -1,
    -- filter=242 channel=82
    -3, 7, 0, 5, 8, 5, -4, 7, 3,
    -- filter=242 channel=83
    10, 7, 0, 2, 1, -1, 4, 1, 1,
    -- filter=242 channel=84
    -2, -5, -1, -5, -7, -1, -5, -10, -9,
    -- filter=242 channel=85
    -1, 3, 4, 7, 0, 2, 0, -5, 2,
    -- filter=242 channel=86
    -11, 0, 3, -11, -12, -4, -5, -1, 5,
    -- filter=242 channel=87
    -4, -11, 2, -1, 6, 0, -8, 4, 4,
    -- filter=242 channel=88
    2, -4, 4, 0, 6, -1, -7, 12, -1,
    -- filter=242 channel=89
    20, 8, -1, 2, 5, -3, 0, -7, 6,
    -- filter=242 channel=90
    0, 5, 1, -1, 3, -6, -2, 10, 2,
    -- filter=242 channel=91
    -7, -6, -14, -8, -13, -4, -9, 2, -11,
    -- filter=242 channel=92
    4, 4, 4, -1, 0, -3, 0, 5, -7,
    -- filter=242 channel=93
    1, 2, 0, -10, -14, -12, -19, -20, -10,
    -- filter=242 channel=94
    4, -7, -4, -5, -3, -6, 0, 1, -7,
    -- filter=242 channel=95
    7, 3, 3, 0, 0, 6, 0, -7, 3,
    -- filter=242 channel=96
    6, 0, -4, 5, 6, -6, 2, 2, 5,
    -- filter=242 channel=97
    11, 3, 3, 2, -1, -9, -6, 2, 3,
    -- filter=242 channel=98
    21, 18, 12, 4, -6, 0, -7, -12, -5,
    -- filter=242 channel=99
    6, 7, 4, -5, 6, 6, -14, 8, 7,
    -- filter=242 channel=100
    1, -8, 2, 4, 5, -3, -3, 8, -1,
    -- filter=242 channel=101
    -8, -11, -3, -10, -8, -7, -7, 7, 4,
    -- filter=242 channel=102
    -6, 2, 7, 2, -6, 5, 0, -3, 1,
    -- filter=242 channel=103
    16, 14, 9, 0, -10, -1, -13, -14, -11,
    -- filter=242 channel=104
    20, 17, 11, 1, 5, 3, -8, -6, 0,
    -- filter=242 channel=105
    -4, -16, -1, 6, 11, 0, 11, 22, 21,
    -- filter=242 channel=106
    2, 0, 2, 5, 2, 6, 7, 13, 5,
    -- filter=242 channel=107
    -13, -8, -19, 2, 1, 0, 2, 5, 10,
    -- filter=242 channel=108
    -9, -8, -2, -5, -5, 7, 6, -3, 1,
    -- filter=242 channel=109
    13, -6, 2, -9, -9, -5, -12, -12, 1,
    -- filter=242 channel=110
    8, 8, 6, 7, 3, 9, 0, 5, 3,
    -- filter=242 channel=111
    -7, 3, -1, -5, -5, 0, 6, -1, 7,
    -- filter=242 channel=112
    9, -4, 3, -5, -7, -5, -11, 0, -11,
    -- filter=242 channel=113
    19, 16, 15, 2, 0, 5, -5, -4, -5,
    -- filter=242 channel=114
    -4, -15, -12, 0, -25, -10, -6, -7, -10,
    -- filter=242 channel=115
    -8, -3, -7, -6, -2, -4, -2, 1, 1,
    -- filter=242 channel=116
    4, -5, 1, 7, 0, -5, 0, -1, 7,
    -- filter=242 channel=117
    7, 1, -4, -5, 4, 2, -2, -1, 1,
    -- filter=242 channel=118
    1, 1, 0, 2, 1, 6, 7, 1, -5,
    -- filter=242 channel=119
    2, -9, -4, 0, 3, -1, -12, 13, -13,
    -- filter=242 channel=120
    0, -3, -4, -12, -4, -5, -11, 15, -8,
    -- filter=242 channel=121
    11, 6, 12, -2, 1, 3, 5, -10, -4,
    -- filter=242 channel=122
    12, 20, 12, 5, -2, -13, -14, -30, -10,
    -- filter=242 channel=123
    6, 2, 2, 0, 1, 4, 2, 2, -2,
    -- filter=242 channel=124
    -13, -9, -2, 2, 6, 8, 8, 15, 3,
    -- filter=242 channel=125
    2, 12, 7, 6, 8, 3, 1, 0, 3,
    -- filter=242 channel=126
    12, 0, 9, 3, 4, 3, 8, -2, 8,
    -- filter=242 channel=127
    -7, -3, -4, -5, 1, -1, 0, -6, 1,
    -- filter=243 channel=0
    5, -3, -5, -2, -5, 3, 1, 6, -5,
    -- filter=243 channel=1
    4, -7, 2, 1, 5, 0, -3, -5, 5,
    -- filter=243 channel=2
    -5, 5, -7, -5, 4, 5, 5, 5, -5,
    -- filter=243 channel=3
    -2, -8, 2, -5, 3, 2, 1, -2, 7,
    -- filter=243 channel=4
    -4, 3, 0, 6, 3, -2, -6, -2, -6,
    -- filter=243 channel=5
    5, -4, -6, 4, 5, -5, 0, 4, -3,
    -- filter=243 channel=6
    0, -1, 4, 0, 3, 4, -7, 3, 2,
    -- filter=243 channel=7
    5, -6, 6, 3, 5, -4, 6, 1, 0,
    -- filter=243 channel=8
    0, -6, -3, -1, -2, -3, 3, 0, 0,
    -- filter=243 channel=9
    -5, -3, 5, -2, -5, -6, 6, -7, -2,
    -- filter=243 channel=10
    -4, -6, 7, -1, -6, 0, 2, -6, -2,
    -- filter=243 channel=11
    -2, 5, 2, -4, 0, 0, 0, 5, 4,
    -- filter=243 channel=12
    3, 7, 3, 3, 1, 2, 1, 2, -2,
    -- filter=243 channel=13
    -2, -1, -2, 7, 4, 6, -2, 1, 0,
    -- filter=243 channel=14
    4, -5, 0, 6, -5, -1, -2, -1, 5,
    -- filter=243 channel=15
    -6, -7, -5, 5, 0, 4, 1, -7, 0,
    -- filter=243 channel=16
    -3, -2, -2, -3, 3, -5, 0, 4, -4,
    -- filter=243 channel=17
    1, -6, 6, 5, 2, 6, -3, 3, -4,
    -- filter=243 channel=18
    5, -6, -4, 7, 1, 2, 4, -3, -10,
    -- filter=243 channel=19
    -6, -1, 0, 3, -7, 4, 3, 3, -3,
    -- filter=243 channel=20
    7, 0, -5, -1, 5, 3, 7, 0, -6,
    -- filter=243 channel=21
    3, 0, -2, 6, -7, -4, -7, 0, 6,
    -- filter=243 channel=22
    -1, -6, -3, -4, -6, 0, -6, 6, -5,
    -- filter=243 channel=23
    0, 2, -2, 4, 0, -5, -6, -3, -2,
    -- filter=243 channel=24
    4, 5, -6, -4, -1, 6, -4, -5, 2,
    -- filter=243 channel=25
    5, -2, -3, 0, -3, 4, -2, -1, 4,
    -- filter=243 channel=26
    -3, 7, -5, 1, 4, 6, 6, 3, 4,
    -- filter=243 channel=27
    -3, -6, 4, 6, -6, 5, 3, -2, 1,
    -- filter=243 channel=28
    -5, 6, 6, 3, -6, 7, 3, 6, -4,
    -- filter=243 channel=29
    2, -5, 7, 1, -2, -5, -4, 4, -8,
    -- filter=243 channel=30
    1, 1, -2, 0, -2, 6, 6, 0, -1,
    -- filter=243 channel=31
    -6, 3, 7, -1, -1, 3, -6, -1, 0,
    -- filter=243 channel=32
    7, 3, 2, 1, -8, 5, -5, -8, -6,
    -- filter=243 channel=33
    -1, -4, 1, 2, -5, -4, 0, 0, -5,
    -- filter=243 channel=34
    6, 2, 0, 1, 5, -5, -3, -5, 2,
    -- filter=243 channel=35
    2, 1, 0, 4, -1, 0, -6, -2, -2,
    -- filter=243 channel=36
    7, 6, 2, 0, 7, -3, 8, 4, 0,
    -- filter=243 channel=37
    -7, -3, 7, 2, -6, -2, 0, 2, -1,
    -- filter=243 channel=38
    5, 0, 1, -5, -5, -1, 4, 5, 3,
    -- filter=243 channel=39
    1, -3, -1, 3, 5, -6, -3, -5, 4,
    -- filter=243 channel=40
    -4, -1, 5, 6, -6, 5, 5, -6, 0,
    -- filter=243 channel=41
    5, -7, 7, -5, -1, -2, -1, 2, -7,
    -- filter=243 channel=42
    6, 7, -2, 2, -5, 0, 5, 7, 0,
    -- filter=243 channel=43
    0, 0, -3, 7, -3, -3, 0, 5, -7,
    -- filter=243 channel=44
    -2, 6, -3, -3, 4, 0, -7, 0, 5,
    -- filter=243 channel=45
    0, 5, 5, 1, -4, 0, 1, 5, -6,
    -- filter=243 channel=46
    -1, 1, 0, -5, 7, 2, 2, 4, 0,
    -- filter=243 channel=47
    -3, -6, -5, 0, 1, 8, -3, -2, -4,
    -- filter=243 channel=48
    -6, 0, -1, -7, -1, 8, 1, 2, 4,
    -- filter=243 channel=49
    -7, -3, 6, 5, -8, 2, -7, 0, -1,
    -- filter=243 channel=50
    -7, 5, 2, 3, 3, -2, -4, 0, 7,
    -- filter=243 channel=51
    -4, -4, 5, 4, 2, -3, -4, -6, 5,
    -- filter=243 channel=52
    2, -1, -1, 5, 5, -1, 0, -3, 0,
    -- filter=243 channel=53
    -4, 2, -1, -1, 6, 2, 6, 4, 5,
    -- filter=243 channel=54
    -3, -4, 2, 3, 0, -6, 0, -2, 0,
    -- filter=243 channel=55
    5, -6, -1, 3, 0, 5, 4, -6, -7,
    -- filter=243 channel=56
    2, 5, -4, 1, 0, 7, 5, 2, 0,
    -- filter=243 channel=57
    2, -3, -6, -4, -6, -1, 1, 6, 6,
    -- filter=243 channel=58
    3, -4, -5, 3, -3, -5, 4, 1, -6,
    -- filter=243 channel=59
    -1, 0, 2, 8, -3, 5, -6, -4, 6,
    -- filter=243 channel=60
    1, -6, -5, -6, 1, -3, 0, -4, -1,
    -- filter=243 channel=61
    0, 0, -4, -4, -3, 3, -3, -6, -6,
    -- filter=243 channel=62
    -7, 0, -2, 4, 3, -2, -3, -4, 2,
    -- filter=243 channel=63
    -1, -2, -2, 7, -4, 4, -2, 7, 2,
    -- filter=243 channel=64
    3, -2, 0, 4, -6, 0, -3, -7, 3,
    -- filter=243 channel=65
    -6, -5, 2, 3, 1, -6, -5, 1, 0,
    -- filter=243 channel=66
    3, -2, 0, -4, 2, -4, 3, 2, 2,
    -- filter=243 channel=67
    -7, 6, -2, 1, -3, 5, -4, -5, 1,
    -- filter=243 channel=68
    7, -1, -6, 1, 3, -6, 3, 6, 6,
    -- filter=243 channel=69
    3, -4, 1, 4, 0, 6, 8, -2, -2,
    -- filter=243 channel=70
    -5, -1, 0, -7, 3, 5, -3, 0, 1,
    -- filter=243 channel=71
    6, -3, -2, -4, -2, 0, 6, -3, -5,
    -- filter=243 channel=72
    -5, 0, 0, -1, 4, 0, -7, 3, -4,
    -- filter=243 channel=73
    3, 4, -6, 0, -4, -8, 0, -5, 5,
    -- filter=243 channel=74
    -2, 0, -5, 2, 3, 0, -2, 0, 1,
    -- filter=243 channel=75
    -5, -3, -7, -5, -6, 6, -6, -5, 1,
    -- filter=243 channel=76
    4, 1, 8, -3, 3, 4, 9, 3, -7,
    -- filter=243 channel=77
    -3, 6, -1, 3, 2, 3, -4, 5, 4,
    -- filter=243 channel=78
    7, -2, 3, 0, 0, 2, 3, -1, 2,
    -- filter=243 channel=79
    1, 4, 1, 10, 5, -1, 8, -2, -5,
    -- filter=243 channel=80
    0, -2, -7, -1, -5, 0, -1, -6, 3,
    -- filter=243 channel=81
    6, -3, 4, -3, 5, 1, 4, 0, 4,
    -- filter=243 channel=82
    5, -6, -5, -2, 3, 0, -2, -2, -5,
    -- filter=243 channel=83
    4, -2, -2, -7, -4, -1, 3, -1, -2,
    -- filter=243 channel=84
    6, 2, -2, 2, -7, 6, -5, -6, -5,
    -- filter=243 channel=85
    -1, 0, -1, 2, -6, 0, -2, -5, -5,
    -- filter=243 channel=86
    6, -2, -6, 6, 1, -3, -3, 0, -2,
    -- filter=243 channel=87
    -6, -2, 4, 5, -1, -2, -6, -3, 4,
    -- filter=243 channel=88
    -5, 5, 0, 5, 2, -2, 0, 4, 7,
    -- filter=243 channel=89
    6, 0, -3, 5, -5, 2, -2, -1, 4,
    -- filter=243 channel=90
    0, 3, 0, 3, 4, 9, -6, -4, 8,
    -- filter=243 channel=91
    -4, -6, 0, 1, -5, 3, -3, 4, -7,
    -- filter=243 channel=92
    -2, -2, 1, -3, 6, 0, 0, -6, 8,
    -- filter=243 channel=93
    -3, -1, -4, -6, -7, -5, 0, 5, 7,
    -- filter=243 channel=94
    2, -3, -5, 5, 2, 4, 5, 1, -6,
    -- filter=243 channel=95
    -3, -5, -2, 0, -3, -1, 7, 6, -3,
    -- filter=243 channel=96
    7, 5, 4, -5, -2, 4, 1, -1, 0,
    -- filter=243 channel=97
    2, 1, 2, -3, -2, 4, -1, 2, -5,
    -- filter=243 channel=98
    4, -4, -8, 1, -8, 1, 8, -7, 2,
    -- filter=243 channel=99
    5, -4, -4, 0, 3, 4, -6, -6, 0,
    -- filter=243 channel=100
    1, 3, -1, -2, 1, 1, -4, 2, 0,
    -- filter=243 channel=101
    3, -4, 5, 5, 0, -2, 3, 0, -1,
    -- filter=243 channel=102
    -3, -6, 0, 5, 4, -3, 0, -7, 5,
    -- filter=243 channel=103
    1, 3, -4, -1, -8, 3, 0, -6, 6,
    -- filter=243 channel=104
    -3, 1, 3, -7, -5, -4, -3, 1, 5,
    -- filter=243 channel=105
    0, -4, -1, 1, -5, -4, 3, 3, 2,
    -- filter=243 channel=106
    6, 3, -6, 4, -1, 0, 2, 4, -2,
    -- filter=243 channel=107
    5, -2, 7, -1, 3, -6, 7, 2, -6,
    -- filter=243 channel=108
    7, 3, -5, 6, 3, 4, 4, 5, -7,
    -- filter=243 channel=109
    3, 2, -7, 7, 4, -6, 6, 0, -7,
    -- filter=243 channel=110
    0, -5, 1, -4, 0, -1, -3, -7, 0,
    -- filter=243 channel=111
    -1, 6, 2, 3, 6, -6, 3, 4, -7,
    -- filter=243 channel=112
    0, 6, -7, -6, 3, 2, 4, 0, -1,
    -- filter=243 channel=113
    -2, -3, -6, 2, -7, -5, 1, -2, 0,
    -- filter=243 channel=114
    -2, -6, -3, 7, -6, 3, 0, 3, -5,
    -- filter=243 channel=115
    1, -4, -4, 3, -2, -4, 0, 0, 4,
    -- filter=243 channel=116
    -2, 4, -5, 2, -6, 2, -4, 2, 0,
    -- filter=243 channel=117
    -4, 1, 0, 3, 5, -4, 1, -5, -4,
    -- filter=243 channel=118
    7, 7, -6, -5, -5, 7, 5, -1, 3,
    -- filter=243 channel=119
    -5, 6, 5, 4, -3, 0, -2, 6, 1,
    -- filter=243 channel=120
    -3, -5, -4, 2, -9, -6, 0, -7, -3,
    -- filter=243 channel=121
    -1, 1, -2, 0, -2, -5, 2, 5, 6,
    -- filter=243 channel=122
    -3, 1, -2, 3, 1, 7, -4, 7, -2,
    -- filter=243 channel=123
    -4, -3, 3, -5, -7, -2, 4, 7, -1,
    -- filter=243 channel=124
    4, 5, 7, 3, 4, -4, -4, -7, -1,
    -- filter=243 channel=125
    2, -5, -5, 4, -9, -2, 2, 5, -1,
    -- filter=243 channel=126
    -4, -5, 6, 1, 0, 4, 4, 5, 0,
    -- filter=243 channel=127
    -2, -2, 0, 3, 0, 5, -5, 5, -5,
    -- filter=244 channel=0
    5, 5, -1, 2, 0, -3, 3, 5, -7,
    -- filter=244 channel=1
    5, 2, -4, 3, -6, -1, -4, 3, -6,
    -- filter=244 channel=2
    3, 6, 2, 0, -6, 1, 1, 0, 3,
    -- filter=244 channel=3
    -1, -3, -2, -5, 2, 0, -1, -6, 4,
    -- filter=244 channel=4
    -4, 0, -3, -3, 8, 3, -5, 9, 0,
    -- filter=244 channel=5
    -1, 1, -2, 5, 5, -1, -5, 1, -3,
    -- filter=244 channel=6
    -2, 0, -5, -5, -6, 3, -3, 6, 0,
    -- filter=244 channel=7
    -7, -5, 5, 2, 6, -4, -2, 5, 0,
    -- filter=244 channel=8
    1, -6, 0, 1, 2, 6, -2, -3, -4,
    -- filter=244 channel=9
    -4, 1, 4, 3, -7, -6, 5, 5, 0,
    -- filter=244 channel=10
    5, -6, 0, 1, -4, -3, 9, 5, 7,
    -- filter=244 channel=11
    -5, -5, 6, -6, 6, -1, 0, 3, 0,
    -- filter=244 channel=12
    1, -3, -7, 1, 0, 0, 0, 6, 1,
    -- filter=244 channel=13
    -4, -2, -6, 2, -2, -8, 3, -6, 0,
    -- filter=244 channel=14
    3, -2, -4, 3, -4, 0, -1, 2, 0,
    -- filter=244 channel=15
    -5, -7, -1, 5, -7, -2, 0, 2, -3,
    -- filter=244 channel=16
    4, -2, -5, 8, -1, -3, 4, -7, 3,
    -- filter=244 channel=17
    1, 7, 5, 1, 2, -1, 5, -3, 5,
    -- filter=244 channel=18
    -5, -2, 0, -3, 3, -6, -7, 3, -4,
    -- filter=244 channel=19
    3, 1, 0, 2, 5, 0, 0, 0, 2,
    -- filter=244 channel=20
    2, 3, 1, 2, 2, 0, 9, 0, -2,
    -- filter=244 channel=21
    4, -6, -4, 9, -5, -5, 1, 1, -2,
    -- filter=244 channel=22
    -6, -5, -1, -3, 5, -6, 0, 1, -6,
    -- filter=244 channel=23
    -1, 4, 5, -7, -10, -7, -6, 3, -2,
    -- filter=244 channel=24
    -7, 0, 5, 6, 7, -3, 4, 0, 4,
    -- filter=244 channel=25
    -4, -1, -4, -3, -3, -3, -4, -1, -7,
    -- filter=244 channel=26
    3, 0, -5, 2, 2, 0, 6, -5, 1,
    -- filter=244 channel=27
    4, -7, -6, 4, 0, -1, 3, 1, -5,
    -- filter=244 channel=28
    -3, -6, -1, -1, 6, 3, -3, 4, 0,
    -- filter=244 channel=29
    5, 0, 2, 3, 7, -5, -4, 6, 3,
    -- filter=244 channel=30
    5, -6, -8, -5, 3, 5, -6, -5, 4,
    -- filter=244 channel=31
    2, 1, -5, -2, -9, -7, 10, 0, 0,
    -- filter=244 channel=32
    -6, -3, -1, 2, -5, -3, -4, 0, 1,
    -- filter=244 channel=33
    -3, 4, 3, -4, -9, 4, 0, -1, 4,
    -- filter=244 channel=34
    2, 1, 2, -5, 4, -3, 1, 5, 3,
    -- filter=244 channel=35
    -6, 0, -5, 0, 2, -6, -4, 3, -4,
    -- filter=244 channel=36
    0, 5, -5, -5, 6, 3, 9, -1, 9,
    -- filter=244 channel=37
    -5, 3, -6, -5, 5, 2, 4, -6, -1,
    -- filter=244 channel=38
    0, 0, 0, -4, -7, 0, -4, 1, 5,
    -- filter=244 channel=39
    2, -4, -4, 2, 8, 4, 1, 5, 8,
    -- filter=244 channel=40
    5, 2, -5, -6, 7, 3, 0, -3, 4,
    -- filter=244 channel=41
    -7, 1, 0, 6, -3, -4, -4, -5, 0,
    -- filter=244 channel=42
    -6, 4, 5, -5, 1, 1, 6, 2, -1,
    -- filter=244 channel=43
    -6, -1, 7, -6, -2, -3, 4, 3, -6,
    -- filter=244 channel=44
    -3, -2, -10, -7, -5, 4, -1, -5, 3,
    -- filter=244 channel=45
    0, 6, -5, 4, 1, 2, 7, -2, -6,
    -- filter=244 channel=46
    -5, -6, 0, 1, 7, -4, -1, 4, -3,
    -- filter=244 channel=47
    -5, 2, -2, 7, -1, -5, 6, -5, 2,
    -- filter=244 channel=48
    3, -5, 2, 5, -6, 5, 4, 4, 6,
    -- filter=244 channel=49
    -2, -5, -1, 0, -4, -7, -4, 4, -4,
    -- filter=244 channel=50
    1, 1, 2, 2, 1, -3, 7, 4, -5,
    -- filter=244 channel=51
    4, 4, 0, 3, 5, 0, -3, 0, -5,
    -- filter=244 channel=52
    -2, -5, 7, -7, 7, 6, 4, -1, -4,
    -- filter=244 channel=53
    1, 0, -3, 2, 1, -2, 7, -1, -4,
    -- filter=244 channel=54
    -6, 3, 0, 7, 7, -1, -3, -6, 0,
    -- filter=244 channel=55
    -5, -4, 2, 1, 2, -1, 0, -6, 6,
    -- filter=244 channel=56
    1, 0, 0, 6, -7, 7, 0, 1, -7,
    -- filter=244 channel=57
    -3, -4, -2, 5, -1, -6, -1, 4, -1,
    -- filter=244 channel=58
    -3, 3, -4, -6, 7, 0, -7, 4, 0,
    -- filter=244 channel=59
    0, 2, -9, 7, -8, 3, -4, 4, -1,
    -- filter=244 channel=60
    0, 4, 5, -2, -1, -6, -4, -1, 7,
    -- filter=244 channel=61
    3, -2, 2, -2, 6, -4, -5, 1, 1,
    -- filter=244 channel=62
    -3, -5, -5, -3, -5, -3, -2, -6, -6,
    -- filter=244 channel=63
    4, -2, 6, 4, -4, 0, 1, 3, 0,
    -- filter=244 channel=64
    -3, 0, 1, 1, 4, 3, 5, -5, 0,
    -- filter=244 channel=65
    -1, 1, 4, -7, -6, 2, -6, -3, 5,
    -- filter=244 channel=66
    -3, -1, 4, 5, -2, -2, -2, 3, -6,
    -- filter=244 channel=67
    -4, 1, -2, 0, -2, 0, 0, 0, 0,
    -- filter=244 channel=68
    -5, -5, -6, 3, -4, 5, 6, 4, -2,
    -- filter=244 channel=69
    0, 5, 1, 0, 6, 2, 3, 1, 6,
    -- filter=244 channel=70
    0, 2, 3, -2, -9, -7, -7, -7, -6,
    -- filter=244 channel=71
    7, 0, -6, 0, 4, 5, 7, 6, -4,
    -- filter=244 channel=72
    6, -8, 0, -3, 4, 3, 7, 0, 2,
    -- filter=244 channel=73
    5, -7, 2, 4, -2, -3, -5, 2, 3,
    -- filter=244 channel=74
    -7, -6, 2, -5, -9, -5, -7, -6, 0,
    -- filter=244 channel=75
    -6, 4, 5, -3, -2, -8, -2, 3, -6,
    -- filter=244 channel=76
    8, -4, 4, 7, 0, 9, 7, 9, 5,
    -- filter=244 channel=77
    6, 0, 4, -2, 2, 0, 0, -5, -1,
    -- filter=244 channel=78
    -2, 5, -4, -6, -2, -1, -6, -3, -1,
    -- filter=244 channel=79
    -1, -3, -7, 6, 2, -5, -5, -2, -6,
    -- filter=244 channel=80
    -4, 3, -3, -1, -2, 0, 3, 4, 4,
    -- filter=244 channel=81
    0, -5, 3, -2, 6, 0, -2, 2, 4,
    -- filter=244 channel=82
    0, -4, -6, 5, -1, 0, 4, -2, -1,
    -- filter=244 channel=83
    1, 0, 2, 2, 3, -3, 6, 4, -3,
    -- filter=244 channel=84
    0, 3, 5, -5, -6, 1, -6, -6, 0,
    -- filter=244 channel=85
    -4, -3, 2, 3, 0, 0, 1, 4, 7,
    -- filter=244 channel=86
    1, 3, -3, 4, -3, -3, -5, 2, -4,
    -- filter=244 channel=87
    -5, 7, -3, 0, 4, -1, 6, 3, -1,
    -- filter=244 channel=88
    -6, 2, -3, 5, -2, 2, 9, 6, 6,
    -- filter=244 channel=89
    2, -8, -4, 0, -8, 1, 5, -1, -1,
    -- filter=244 channel=90
    -3, -5, -2, 5, 7, 0, 1, 8, 6,
    -- filter=244 channel=91
    0, -6, -8, 3, -3, 0, 0, 0, 0,
    -- filter=244 channel=92
    -7, -3, -5, -2, -4, -1, 0, -5, -5,
    -- filter=244 channel=93
    2, -1, 4, -2, -3, 3, 3, -1, 0,
    -- filter=244 channel=94
    0, 1, 6, 0, 5, -4, 5, 5, 6,
    -- filter=244 channel=95
    0, -2, -3, 3, -4, -6, 3, -5, 6,
    -- filter=244 channel=96
    0, 4, 0, -5, 0, 1, -1, -1, 0,
    -- filter=244 channel=97
    5, 0, 0, 5, -3, 2, 4, 0, -7,
    -- filter=244 channel=98
    8, -4, -5, -1, -1, -2, -3, 6, -5,
    -- filter=244 channel=99
    2, 0, -7, -5, 0, -1, 8, 2, -3,
    -- filter=244 channel=100
    6, 3, 1, 6, -7, 0, 1, 2, -3,
    -- filter=244 channel=101
    -2, 0, 2, -6, -3, -4, 2, 0, 8,
    -- filter=244 channel=102
    2, -1, -2, 7, -6, -6, -5, 5, 1,
    -- filter=244 channel=103
    2, -6, -8, 0, -4, -5, 0, 4, 1,
    -- filter=244 channel=104
    7, -5, -9, 4, 1, 2, 9, 4, -1,
    -- filter=244 channel=105
    1, 0, 0, -2, 5, 7, -5, 5, 0,
    -- filter=244 channel=106
    3, 8, 6, -2, 8, -2, 1, 0, 0,
    -- filter=244 channel=107
    5, -1, 8, 2, 5, -2, 5, -6, -3,
    -- filter=244 channel=108
    5, -3, -1, 3, -1, 0, 0, -4, -6,
    -- filter=244 channel=109
    3, -8, 0, -3, -3, 4, 5, 2, 0,
    -- filter=244 channel=110
    3, -5, 4, 0, 0, 3, 3, -1, -5,
    -- filter=244 channel=111
    -2, -6, 1, 5, -3, 5, -2, -6, 0,
    -- filter=244 channel=112
    2, -6, -1, 0, -3, 6, -7, -4, 1,
    -- filter=244 channel=113
    0, 3, -6, 1, 1, -5, 4, -5, 5,
    -- filter=244 channel=114
    -6, -1, -7, -5, -7, 2, -4, -2, -7,
    -- filter=244 channel=115
    -5, 1, 3, 0, 3, -2, -4, 0, -6,
    -- filter=244 channel=116
    7, 3, -10, 4, -4, -7, 0, -3, 5,
    -- filter=244 channel=117
    -1, 0, -7, 7, 7, 1, 5, -2, -3,
    -- filter=244 channel=118
    -7, 1, -1, -4, -6, -3, -2, 7, 1,
    -- filter=244 channel=119
    -5, 0, 0, -8, -6, -5, -7, -3, 0,
    -- filter=244 channel=120
    -4, -3, 1, -2, -5, 7, -2, 1, 6,
    -- filter=244 channel=121
    -1, 2, -5, -7, 0, -1, 1, -4, 0,
    -- filter=244 channel=122
    6, 1, -3, 5, 1, -6, 10, 5, -2,
    -- filter=244 channel=123
    -7, 0, 2, -7, 0, -3, 0, -2, 7,
    -- filter=244 channel=124
    6, -6, 0, 2, 3, -4, 7, -2, -3,
    -- filter=244 channel=125
    7, -2, 0, 2, -5, -2, -3, 5, 5,
    -- filter=244 channel=126
    3, -4, 6, -2, -6, 0, 0, -7, 3,
    -- filter=244 channel=127
    0, 4, 2, -3, 4, 5, 6, -5, 3,
    -- filter=245 channel=0
    -6, 7, 36, -21, -14, 24, -15, -18, 14,
    -- filter=245 channel=1
    -6, 4, 22, -17, -10, 22, -18, -21, 12,
    -- filter=245 channel=2
    -7, 3, 1, 3, -5, 1, -5, -1, -10,
    -- filter=245 channel=3
    -11, -14, 1, -17, -16, -9, -14, -17, -3,
    -- filter=245 channel=4
    -3, -6, 0, -5, -11, -2, -7, -12, -11,
    -- filter=245 channel=5
    -19, 14, 20, -27, -6, 22, -17, -2, 15,
    -- filter=245 channel=6
    -4, -3, -2, 5, 1, 4, -6, 7, 6,
    -- filter=245 channel=7
    3, 3, 0, -3, -1, 3, -3, -5, -5,
    -- filter=245 channel=8
    -1, -4, -8, -5, 0, -9, -6, 3, -9,
    -- filter=245 channel=9
    -7, 0, 10, 1, -1, 6, -8, 2, 2,
    -- filter=245 channel=10
    7, -7, -12, 3, 1, 0, -1, 5, 2,
    -- filter=245 channel=11
    -1, 6, -8, 8, 13, -14, 11, 8, 1,
    -- filter=245 channel=12
    2, 1, 1, 4, -7, -5, 6, -11, -2,
    -- filter=245 channel=13
    12, -4, -16, 8, -5, -2, 3, -6, 4,
    -- filter=245 channel=14
    1, 4, 1, -7, 4, -3, -2, -1, -6,
    -- filter=245 channel=15
    0, 1, -4, 2, -3, -5, 9, 10, -5,
    -- filter=245 channel=16
    -12, 6, 3, -12, 4, 11, -11, 0, 11,
    -- filter=245 channel=17
    0, -7, 3, 0, -4, 5, 2, -5, 0,
    -- filter=245 channel=18
    -7, -5, -3, -1, 0, 7, -5, 3, 1,
    -- filter=245 channel=19
    -3, -2, -7, -6, 3, 0, 3, 0, 6,
    -- filter=245 channel=20
    -6, -4, -11, 15, 13, -21, 8, 24, -3,
    -- filter=245 channel=21
    -2, 4, 4, 6, -5, 0, 8, -5, 7,
    -- filter=245 channel=22
    -11, -1, -4, -2, 9, 0, -12, 6, 8,
    -- filter=245 channel=23
    4, -12, -23, 7, 8, -22, 6, 11, 0,
    -- filter=245 channel=24
    -2, 3, 0, 3, 5, -1, -7, 0, 0,
    -- filter=245 channel=25
    6, 0, 11, 5, 0, 2, 3, -14, 8,
    -- filter=245 channel=26
    -11, 3, 10, -7, 6, 7, -13, -7, -3,
    -- filter=245 channel=27
    9, 0, 4, -10, 4, 1, -3, -5, 0,
    -- filter=245 channel=28
    3, 4, 3, -6, -2, -5, 0, -1, 3,
    -- filter=245 channel=29
    0, -1, -21, 11, 12, -7, 14, 13, 6,
    -- filter=245 channel=30
    2, 11, 17, -12, 3, 7, -12, -7, 14,
    -- filter=245 channel=31
    1, 0, -15, 5, 1, -8, 7, -1, 1,
    -- filter=245 channel=32
    7, -7, -6, -3, -8, -2, -5, 0, 12,
    -- filter=245 channel=33
    -3, -4, -1, -4, 1, 2, -5, -10, 5,
    -- filter=245 channel=34
    1, -3, 0, -14, 14, 4, -15, -7, 4,
    -- filter=245 channel=35
    0, -1, 0, 7, -5, -7, 1, -2, -5,
    -- filter=245 channel=36
    4, -3, -18, 9, 1, -20, 8, 8, -12,
    -- filter=245 channel=37
    -18, -2, 29, -22, -11, 22, -22, -26, 14,
    -- filter=245 channel=38
    -3, 6, -7, 5, 7, 0, -3, 7, 2,
    -- filter=245 channel=39
    1, -3, -10, 2, -4, -4, 10, 9, -4,
    -- filter=245 channel=40
    -3, 0, -5, 6, 7, -9, -1, 6, -7,
    -- filter=245 channel=41
    -1, -12, 1, -5, -4, 8, -2, -10, 1,
    -- filter=245 channel=42
    -4, 3, 10, -2, -7, 14, 4, -5, 6,
    -- filter=245 channel=43
    -2, -6, -6, -1, -9, -5, -11, 0, -7,
    -- filter=245 channel=44
    -6, 2, 22, -21, -6, 10, -6, -1, 12,
    -- filter=245 channel=45
    -4, 2, 0, -1, -5, 9, -1, 0, 6,
    -- filter=245 channel=46
    -4, 6, -3, -4, -5, 6, -9, -7, 0,
    -- filter=245 channel=47
    -13, -6, 14, -8, 3, 20, -1, 1, 9,
    -- filter=245 channel=48
    1, 4, 19, -4, -8, 14, -7, -11, 8,
    -- filter=245 channel=49
    -6, 4, 4, 1, -2, -10, 1, -3, -2,
    -- filter=245 channel=50
    1, 7, 3, 3, -4, 4, -2, 5, -2,
    -- filter=245 channel=51
    -4, 1, -6, -4, -3, -5, 2, 7, 1,
    -- filter=245 channel=52
    0, -9, -12, 2, 0, -11, -5, -3, -1,
    -- filter=245 channel=53
    6, -4, -11, 12, -3, -7, 8, 14, -4,
    -- filter=245 channel=54
    6, -4, -2, 2, -5, -3, 0, 6, 6,
    -- filter=245 channel=55
    6, 0, -19, 14, 13, -14, 8, 14, -7,
    -- filter=245 channel=56
    4, 2, -4, 1, 5, 2, -7, 9, -3,
    -- filter=245 channel=57
    4, -4, 1, -3, 5, 6, 0, 3, -1,
    -- filter=245 channel=58
    -14, 0, 12, -11, 0, 10, -2, -3, 5,
    -- filter=245 channel=59
    4, 5, 8, 8, 0, 6, 4, -5, 4,
    -- filter=245 channel=60
    -2, -7, -5, 2, 2, 5, 1, -4, -1,
    -- filter=245 channel=61
    -6, 0, -5, -6, -2, -4, -2, -3, -1,
    -- filter=245 channel=62
    0, -3, -3, -1, 4, -7, 5, 5, 1,
    -- filter=245 channel=63
    -3, 0, 8, -4, -1, 7, -11, -5, 10,
    -- filter=245 channel=64
    -5, -3, -14, 2, 3, -1, 7, 2, -8,
    -- filter=245 channel=65
    -2, -1, 0, 0, -4, 7, 7, 0, 6,
    -- filter=245 channel=66
    6, -1, 3, 6, -9, 7, 5, -7, 7,
    -- filter=245 channel=67
    2, 0, -2, 3, 0, -8, 1, 6, 2,
    -- filter=245 channel=68
    5, -8, 3, 6, -5, -8, -2, -5, 1,
    -- filter=245 channel=69
    -1, -1, 2, 5, -5, 7, 4, 1, 8,
    -- filter=245 channel=70
    3, -3, 2, 6, 3, -11, -6, 1, 0,
    -- filter=245 channel=71
    -3, -2, -8, 3, 0, 0, 1, -8, -7,
    -- filter=245 channel=72
    3, -7, -6, 19, 0, -2, 17, -4, -6,
    -- filter=245 channel=73
    4, -5, -2, 0, 3, -4, 7, 3, -11,
    -- filter=245 channel=74
    -5, 4, 0, -3, 5, 5, -14, 4, -1,
    -- filter=245 channel=75
    -7, -8, 22, -24, -11, 23, -17, -17, 11,
    -- filter=245 channel=76
    3, -2, -14, 14, 8, -6, 13, 21, -5,
    -- filter=245 channel=77
    -1, -4, 3, 0, 0, 5, -2, -3, 0,
    -- filter=245 channel=78
    -10, 6, 1, -6, -1, 2, 2, 3, 10,
    -- filter=245 channel=79
    7, -3, 0, 8, -7, 11, 0, -3, 12,
    -- filter=245 channel=80
    16, -3, -4, 14, -5, 5, 12, 1, 3,
    -- filter=245 channel=81
    -3, 2, 2, 2, -1, 6, 0, -2, 0,
    -- filter=245 channel=82
    -1, 3, 0, 3, -2, 5, -4, 4, -2,
    -- filter=245 channel=83
    3, 8, 7, -7, -1, 10, 4, 5, 1,
    -- filter=245 channel=84
    -2, 4, 3, 2, 2, 7, -2, -9, 3,
    -- filter=245 channel=85
    -5, -5, -2, -6, 6, -3, -4, 2, -4,
    -- filter=245 channel=86
    -7, 2, 11, 0, 3, 3, -8, -5, 0,
    -- filter=245 channel=87
    -5, 0, -2, 3, 0, 0, -5, 10, 2,
    -- filter=245 channel=88
    -4, -1, -5, 2, -1, -19, -3, 7, -8,
    -- filter=245 channel=89
    10, -17, -10, 15, -1, -5, 11, -5, -7,
    -- filter=245 channel=90
    -7, -5, -13, 0, 6, -20, 3, 12, -5,
    -- filter=245 channel=91
    8, -4, -12, 3, 0, -5, 0, -4, -1,
    -- filter=245 channel=92
    1, 0, 3, -6, 6, -3, -8, 1, 5,
    -- filter=245 channel=93
    -11, 4, 21, -15, -13, 17, -4, -2, 3,
    -- filter=245 channel=94
    6, 6, 0, 4, -4, 4, -2, -6, -3,
    -- filter=245 channel=95
    -6, 0, -8, 4, 3, -1, 0, -4, -3,
    -- filter=245 channel=96
    -4, -8, 1, -3, 0, -1, -2, 4, 1,
    -- filter=245 channel=97
    4, -12, -5, 0, 2, 3, -10, -3, 0,
    -- filter=245 channel=98
    11, -8, -2, 1, -9, 9, -7, -12, 9,
    -- filter=245 channel=99
    -3, 0, -18, 7, 10, -24, -2, 9, -11,
    -- filter=245 channel=100
    5, 5, -4, 1, 4, -3, 0, 3, -5,
    -- filter=245 channel=101
    -6, -9, -11, -8, -7, -6, -6, -14, -2,
    -- filter=245 channel=102
    -4, -7, -5, -5, 5, 7, 0, -2, -5,
    -- filter=245 channel=103
    -6, 5, 7, -8, 0, 13, 1, -8, 6,
    -- filter=245 channel=104
    4, 2, -5, 3, -5, 1, 3, -2, -2,
    -- filter=245 channel=105
    -8, -9, -6, 4, 3, -7, 4, 6, -5,
    -- filter=245 channel=106
    4, -2, 0, -2, 0, -11, -2, 10, 4,
    -- filter=245 channel=107
    -11, -7, -3, -5, -2, 0, 0, -1, 3,
    -- filter=245 channel=108
    -7, 0, 7, -9, -6, -1, -7, -7, -1,
    -- filter=245 channel=109
    1, 4, 5, -4, 8, 5, -11, -2, 1,
    -- filter=245 channel=110
    -1, -1, -6, 4, -7, -9, 0, 3, -10,
    -- filter=245 channel=111
    2, 2, -6, -5, 0, -2, 0, 4, 2,
    -- filter=245 channel=112
    -8, 5, 2, -11, -2, 9, -11, -8, 8,
    -- filter=245 channel=113
    8, 0, -3, 0, -3, 4, 1, 1, 5,
    -- filter=245 channel=114
    -3, 8, 21, -9, -7, 20, -7, -13, 1,
    -- filter=245 channel=115
    -2, 5, -3, 2, 7, -3, 0, 5, 1,
    -- filter=245 channel=116
    11, 1, -1, 8, -2, -7, 11, 4, -6,
    -- filter=245 channel=117
    -1, 4, 1, 9, 0, 0, 3, 0, -5,
    -- filter=245 channel=118
    -8, -5, 2, 2, -2, -4, 6, 3, -4,
    -- filter=245 channel=119
    -3, -1, 6, -2, 9, -4, -11, 6, 0,
    -- filter=245 channel=120
    -12, -3, -7, 4, 2, -8, -1, 7, 2,
    -- filter=245 channel=121
    2, -10, -9, 2, -9, -1, 0, -2, 5,
    -- filter=245 channel=122
    -19, -2, 10, -17, 1, 4, -8, 3, 2,
    -- filter=245 channel=123
    2, -8, 0, 1, -3, -4, 2, -3, -6,
    -- filter=245 channel=124
    3, -6, -10, 4, 5, -3, -4, 13, 6,
    -- filter=245 channel=125
    0, 1, -4, 6, 0, 2, 8, 8, 3,
    -- filter=245 channel=126
    0, 0, -4, 2, -10, 7, 1, -1, 8,
    -- filter=245 channel=127
    3, -3, -2, -1, -1, -3, 0, 3, 7,
    -- filter=246 channel=0
    6, -3, 3, -5, -3, -5, 1, -7, 3,
    -- filter=246 channel=1
    4, -2, 0, -4, -2, -2, 0, 4, 5,
    -- filter=246 channel=2
    -6, 4, -1, -6, 0, 6, -7, -2, -1,
    -- filter=246 channel=3
    -5, -5, -4, 6, 4, 1, 4, 0, 0,
    -- filter=246 channel=4
    -2, -4, 2, 0, -5, 5, -4, -6, -1,
    -- filter=246 channel=5
    -6, -5, 6, 1, -3, 4, 3, -6, 2,
    -- filter=246 channel=6
    2, 6, -6, 2, -4, 0, -5, -6, 1,
    -- filter=246 channel=7
    -6, 4, -1, -4, -5, -6, 3, -3, 4,
    -- filter=246 channel=8
    6, 0, -5, 6, 6, -5, -2, 1, -3,
    -- filter=246 channel=9
    -2, -3, -1, 3, 0, 1, 1, -1, 7,
    -- filter=246 channel=10
    2, 4, 5, -5, 3, -6, -6, 4, -2,
    -- filter=246 channel=11
    1, -2, -2, 7, 4, 5, -2, 0, 5,
    -- filter=246 channel=12
    -1, 3, -1, 0, 1, 0, 6, -4, 0,
    -- filter=246 channel=13
    -2, -3, 6, 5, -4, -2, 2, -1, -2,
    -- filter=246 channel=14
    4, 5, 1, 2, -6, -6, 7, -5, 2,
    -- filter=246 channel=15
    3, -6, 1, -5, 0, 1, -7, -6, 3,
    -- filter=246 channel=16
    4, 4, -5, -6, 6, 3, -3, 5, 6,
    -- filter=246 channel=17
    -1, 1, -3, 2, 2, -2, 0, 0, -6,
    -- filter=246 channel=18
    6, 2, 1, -3, -2, 3, 6, -3, -5,
    -- filter=246 channel=19
    1, 2, 5, 2, 6, 6, 5, -3, 2,
    -- filter=246 channel=20
    -4, 2, 0, 0, 0, 4, 3, -6, 3,
    -- filter=246 channel=21
    1, -5, 0, 3, -6, -6, 0, -3, 6,
    -- filter=246 channel=22
    1, 3, -2, -1, -6, 0, -2, -2, -4,
    -- filter=246 channel=23
    -1, 1, 0, 1, 5, 6, -6, 7, 1,
    -- filter=246 channel=24
    4, 4, 3, -2, -4, -1, 6, -1, -6,
    -- filter=246 channel=25
    3, 2, -7, -6, -5, 4, -1, 1, 0,
    -- filter=246 channel=26
    -5, -7, 0, -5, 0, 6, -6, 2, 6,
    -- filter=246 channel=27
    -1, 7, -1, 1, -1, 0, 1, 6, -6,
    -- filter=246 channel=28
    -1, -4, 1, 3, -1, 4, -5, -7, -4,
    -- filter=246 channel=29
    -6, 1, -1, 2, -2, -6, 1, -3, 2,
    -- filter=246 channel=30
    -3, 1, 0, 1, 3, 3, -5, -4, -4,
    -- filter=246 channel=31
    -7, 4, 2, -7, 0, -4, 5, -2, -2,
    -- filter=246 channel=32
    -1, 3, -6, -1, -2, 4, 2, -1, 0,
    -- filter=246 channel=33
    -5, 3, 2, -7, 4, -1, 4, 2, -6,
    -- filter=246 channel=34
    0, -5, -1, 3, 1, 1, 1, 4, -5,
    -- filter=246 channel=35
    5, -6, 0, 3, -5, -2, 1, -1, 0,
    -- filter=246 channel=36
    -7, 2, -7, -4, 0, 2, 0, -4, 5,
    -- filter=246 channel=37
    -4, 2, -3, 3, 3, -7, 4, 6, 4,
    -- filter=246 channel=38
    1, 4, -1, 1, 2, -4, -7, 4, 7,
    -- filter=246 channel=39
    -5, -3, 0, -4, 2, -5, 5, -5, 0,
    -- filter=246 channel=40
    2, 2, 1, -7, -2, -4, 2, 2, 6,
    -- filter=246 channel=41
    5, 3, -2, -1, -7, 2, 3, -5, 5,
    -- filter=246 channel=42
    6, 3, 5, 2, -1, -5, 2, 0, 5,
    -- filter=246 channel=43
    -1, 4, -3, 0, -3, 6, 0, 7, -1,
    -- filter=246 channel=44
    7, -4, 2, 7, -5, 4, 3, 5, -2,
    -- filter=246 channel=45
    -4, 1, -3, -1, 1, 7, 0, 1, 5,
    -- filter=246 channel=46
    3, 2, 1, 3, -5, 2, 0, -6, 6,
    -- filter=246 channel=47
    0, 0, -6, 5, -2, 0, 1, -1, -2,
    -- filter=246 channel=48
    -2, -6, -5, 3, 2, -4, 3, -4, 1,
    -- filter=246 channel=49
    -3, 3, 3, 4, 2, 3, -3, -4, 3,
    -- filter=246 channel=50
    -7, 3, 4, 3, 5, 1, 5, 7, -5,
    -- filter=246 channel=51
    6, 0, 0, 5, 4, -4, -3, 1, 0,
    -- filter=246 channel=52
    2, -4, 1, 0, 0, -4, -3, -5, 1,
    -- filter=246 channel=53
    -3, 4, 4, -5, 4, 2, 5, 0, 1,
    -- filter=246 channel=54
    1, 4, -3, -2, 2, -1, 3, -4, 1,
    -- filter=246 channel=55
    2, 4, -2, -1, 5, -2, 6, 0, 6,
    -- filter=246 channel=56
    6, -2, 1, 3, 6, -6, -6, -4, 0,
    -- filter=246 channel=57
    -2, 6, 3, -3, 0, 0, -7, 4, 5,
    -- filter=246 channel=58
    0, 2, 3, -6, 5, -5, -2, 0, 1,
    -- filter=246 channel=59
    0, -1, -6, -2, 0, 3, 5, 6, 2,
    -- filter=246 channel=60
    3, -2, 3, -4, 4, 6, -7, -4, -1,
    -- filter=246 channel=61
    1, -7, -2, 6, -6, 4, 0, 2, -2,
    -- filter=246 channel=62
    0, -2, -3, -7, 3, 5, -5, -1, -5,
    -- filter=246 channel=63
    0, -3, 6, 0, 6, 0, 0, 5, -6,
    -- filter=246 channel=64
    -6, -1, -2, 3, -4, 4, 5, -6, 5,
    -- filter=246 channel=65
    -1, -6, -3, 0, 1, -4, 4, 1, -3,
    -- filter=246 channel=66
    0, 0, -2, -6, 3, -5, 0, -5, 3,
    -- filter=246 channel=67
    -2, 0, -3, 5, 6, 6, 3, 7, -1,
    -- filter=246 channel=68
    7, 4, 4, 2, 0, -3, -3, -4, 6,
    -- filter=246 channel=69
    5, -5, -6, 6, 1, -3, 0, 6, 3,
    -- filter=246 channel=70
    0, -2, 3, -3, 2, -3, -2, 1, 7,
    -- filter=246 channel=71
    4, 6, -2, -4, -3, 2, -6, 6, -5,
    -- filter=246 channel=72
    -7, 7, -2, 4, 6, 6, -6, 5, 0,
    -- filter=246 channel=73
    2, -2, 6, -4, -1, -6, -5, 2, 3,
    -- filter=246 channel=74
    -3, -6, 0, -3, -6, -4, -2, -5, -6,
    -- filter=246 channel=75
    0, -5, -1, 1, 1, 2, -4, 5, 2,
    -- filter=246 channel=76
    -2, -6, 0, 1, 0, 1, 6, -4, -4,
    -- filter=246 channel=77
    3, -7, 5, 1, 5, -3, -2, -4, 2,
    -- filter=246 channel=78
    3, -4, -1, -5, -2, 2, -2, 3, 1,
    -- filter=246 channel=79
    -4, -1, 0, 0, -2, -6, 3, -5, -6,
    -- filter=246 channel=80
    -2, -6, 2, 0, 0, 0, 3, -2, -5,
    -- filter=246 channel=81
    -4, 1, -3, 3, -5, -7, -7, 6, 0,
    -- filter=246 channel=82
    -1, 2, 2, 5, 0, -5, 0, 3, 1,
    -- filter=246 channel=83
    4, -1, 2, 0, 1, -3, -4, 2, 3,
    -- filter=246 channel=84
    5, 1, 3, 2, -6, 1, -7, -6, 1,
    -- filter=246 channel=85
    6, 0, -6, -1, -1, -3, -5, -1, 0,
    -- filter=246 channel=86
    -3, 7, 3, 6, -6, 1, 4, 7, -1,
    -- filter=246 channel=87
    5, 0, -6, 2, 0, -2, 5, -5, 4,
    -- filter=246 channel=88
    7, 2, -6, -5, -1, -2, -1, 0, 4,
    -- filter=246 channel=89
    -2, 4, -6, 1, -5, -3, 0, -4, -2,
    -- filter=246 channel=90
    0, 2, -4, -5, -2, -5, 1, -5, 6,
    -- filter=246 channel=91
    6, -2, 2, 2, -4, 2, 4, 5, 2,
    -- filter=246 channel=92
    5, 4, -6, -2, 0, -2, -3, 0, -4,
    -- filter=246 channel=93
    7, -5, -7, -2, -5, 7, -3, -2, -3,
    -- filter=246 channel=94
    6, 0, -4, -6, -1, 6, 0, -4, 2,
    -- filter=246 channel=95
    -2, -4, 3, -1, 2, 7, 4, -2, -5,
    -- filter=246 channel=96
    -1, 0, 0, -5, 7, 4, 5, 3, -2,
    -- filter=246 channel=97
    -4, 0, 1, 4, -5, 0, -3, 3, 4,
    -- filter=246 channel=98
    -4, 0, 0, 0, 5, -6, -5, 5, 2,
    -- filter=246 channel=99
    -1, -5, -2, -7, 1, -6, 4, -1, -6,
    -- filter=246 channel=100
    -7, 1, -5, 0, 4, -1, -2, -5, -2,
    -- filter=246 channel=101
    0, -7, 6, -7, -4, 1, 6, -6, -4,
    -- filter=246 channel=102
    6, 4, 3, 3, -2, -7, 1, 1, -4,
    -- filter=246 channel=103
    -5, 4, 0, -6, 6, 0, -7, -2, 1,
    -- filter=246 channel=104
    -3, 0, 4, -2, -3, -6, 6, 5, -7,
    -- filter=246 channel=105
    3, 3, -4, 2, -5, 1, -5, 6, 5,
    -- filter=246 channel=106
    1, 4, 1, -3, 3, -3, -7, -4, 6,
    -- filter=246 channel=107
    -1, 4, -6, -7, 2, -6, 1, -5, -6,
    -- filter=246 channel=108
    0, -7, 3, -7, 4, -5, 3, -4, -7,
    -- filter=246 channel=109
    5, -6, 6, 3, 0, -4, -5, -4, 2,
    -- filter=246 channel=110
    -5, 3, -4, -4, -4, 6, 2, 2, -6,
    -- filter=246 channel=111
    -2, -3, 4, 2, -3, -3, 1, 4, -3,
    -- filter=246 channel=112
    7, -3, 0, -3, -3, -3, -3, -5, -2,
    -- filter=246 channel=113
    -4, -6, 0, -3, -3, 0, -2, 6, -1,
    -- filter=246 channel=114
    -4, -6, -6, 0, 0, -3, -2, 1, 5,
    -- filter=246 channel=115
    0, -4, -6, -6, 2, -6, 1, -4, -4,
    -- filter=246 channel=116
    -3, -3, -1, 4, 4, 1, 0, -1, -6,
    -- filter=246 channel=117
    5, 0, 4, 3, -5, 3, 4, 0, 3,
    -- filter=246 channel=118
    -5, 0, 5, 4, 6, 0, 6, -2, -5,
    -- filter=246 channel=119
    -1, -3, -6, -2, 5, -4, 6, -2, -5,
    -- filter=246 channel=120
    0, 1, 5, 1, -4, -2, 2, -1, -7,
    -- filter=246 channel=121
    1, 0, -6, 2, -4, -1, -7, -1, -7,
    -- filter=246 channel=122
    5, -3, -6, 2, 5, 5, -7, 6, 5,
    -- filter=246 channel=123
    0, 0, 0, 3, 0, 4, 3, 6, -5,
    -- filter=246 channel=124
    0, 2, 0, 0, -6, -7, 7, -4, 4,
    -- filter=246 channel=125
    -7, -2, 0, 4, 3, 4, 0, 0, -4,
    -- filter=246 channel=126
    -2, -1, 4, -5, 1, 5, -1, 5, -7,
    -- filter=246 channel=127
    -3, 3, -5, 3, -7, 2, 7, 7, -6,
    -- filter=247 channel=0
    -2, -7, 0, 4, -10, -3, 9, 0, 7,
    -- filter=247 channel=1
    0, 3, -4, -5, -8, 1, 14, 9, 6,
    -- filter=247 channel=2
    5, 6, -3, 2, -1, 6, 13, 9, -7,
    -- filter=247 channel=3
    -1, 17, 9, 5, 9, -3, -3, 17, 19,
    -- filter=247 channel=4
    -2, -1, 0, 0, 8, 8, 25, 24, -2,
    -- filter=247 channel=5
    0, -5, -11, 5, -10, -5, -4, 6, 6,
    -- filter=247 channel=6
    3, -7, 6, 0, 1, 7, 6, 8, 1,
    -- filter=247 channel=7
    -4, 3, 3, 1, -6, 5, 2, 0, 3,
    -- filter=247 channel=8
    0, -8, 4, 0, 3, 7, 4, -1, 5,
    -- filter=247 channel=9
    -1, 5, 0, 0, -2, -7, 6, 0, 2,
    -- filter=247 channel=10
    -1, 12, -9, 2, -7, -10, -12, 1, 5,
    -- filter=247 channel=11
    3, 4, 3, 0, -3, -2, -1, -1, 3,
    -- filter=247 channel=12
    0, 7, 6, 7, -8, 2, -3, -4, 9,
    -- filter=247 channel=13
    0, 5, -4, -2, -13, 0, 0, 5, 10,
    -- filter=247 channel=14
    7, 0, -5, -3, -3, -2, 0, -2, -7,
    -- filter=247 channel=15
    -7, -1, 6, -4, -11, 0, 0, 8, 7,
    -- filter=247 channel=16
    4, 12, -6, 9, 4, 5, -8, -2, 8,
    -- filter=247 channel=17
    4, -2, 1, -3, -3, 0, -2, -3, -2,
    -- filter=247 channel=18
    1, -13, -2, -5, -25, 0, 1, -3, 11,
    -- filter=247 channel=19
    -5, 0, -2, 0, -6, 2, -2, 6, 2,
    -- filter=247 channel=20
    -6, -9, 7, -7, -8, 11, 0, 0, 1,
    -- filter=247 channel=21
    12, 14, -4, -2, -5, -10, -8, -7, 1,
    -- filter=247 channel=22
    1, 1, -4, -6, -4, 5, 0, -4, 2,
    -- filter=247 channel=23
    -3, -9, 0, -16, -9, 1, -10, -2, 6,
    -- filter=247 channel=24
    6, -5, 4, 6, -3, 2, 0, -1, 3,
    -- filter=247 channel=25
    5, 2, -10, -9, -9, 8, 0, 13, 6,
    -- filter=247 channel=26
    3, -6, -2, 0, 6, 9, 5, -4, 0,
    -- filter=247 channel=27
    0, -8, -5, -21, -22, 5, 14, 17, 6,
    -- filter=247 channel=28
    6, -3, 6, 6, -6, -6, 5, 5, -4,
    -- filter=247 channel=29
    3, -1, 14, -15, 0, 4, -10, 5, 1,
    -- filter=247 channel=30
    0, -7, -8, -8, -11, -4, 0, 12, -6,
    -- filter=247 channel=31
    9, 3, -3, -3, -1, 0, -4, 5, -1,
    -- filter=247 channel=32
    7, -7, 0, -6, -13, 3, 2, 2, 11,
    -- filter=247 channel=33
    -4, -2, 2, -8, -10, 1, -2, 4, 13,
    -- filter=247 channel=34
    -13, -4, 11, 0, -5, 6, 12, 7, -7,
    -- filter=247 channel=35
    -7, 0, 3, 7, 3, 5, 0, 0, -1,
    -- filter=247 channel=36
    3, 3, -3, -9, 0, -5, 0, 3, 1,
    -- filter=247 channel=37
    1, -2, -13, 0, 0, 6, 2, 6, -4,
    -- filter=247 channel=38
    -1, 1, -2, -4, -6, 5, -5, 4, 8,
    -- filter=247 channel=39
    5, -1, 10, 2, -8, -2, 2, 0, -3,
    -- filter=247 channel=40
    -1, -6, -2, -2, 0, -3, -8, -3, 1,
    -- filter=247 channel=41
    -3, -5, -1, 7, -2, -13, 9, 0, 1,
    -- filter=247 channel=42
    -8, 6, 0, -3, -5, 4, 5, 1, -5,
    -- filter=247 channel=43
    3, 0, -2, 4, -4, 0, -5, 2, 6,
    -- filter=247 channel=44
    -3, -9, -12, 2, -6, 8, 9, 10, -2,
    -- filter=247 channel=45
    6, -6, -7, -1, -6, 6, -2, -2, -5,
    -- filter=247 channel=46
    5, 1, 2, -7, 0, -2, 0, 4, 3,
    -- filter=247 channel=47
    6, 11, -6, -5, 4, -10, -4, 7, -3,
    -- filter=247 channel=48
    4, -7, -16, -5, 0, 1, 1, 14, -1,
    -- filter=247 channel=49
    -3, -14, 4, -14, -2, 12, 8, 2, -2,
    -- filter=247 channel=50
    10, 0, 0, -2, -10, 3, 1, -3, 4,
    -- filter=247 channel=51
    -1, 2, 7, 6, 1, 0, -1, -2, 0,
    -- filter=247 channel=52
    2, 0, 6, 0, 7, -2, 8, 0, -5,
    -- filter=247 channel=53
    0, -5, 2, -11, 3, -2, 0, 5, -2,
    -- filter=247 channel=54
    6, 3, 1, -5, 1, -7, -2, -6, 4,
    -- filter=247 channel=55
    11, -10, 0, -6, -12, 6, -7, -6, 3,
    -- filter=247 channel=56
    -2, -6, 13, -6, 6, 1, 6, 6, 0,
    -- filter=247 channel=57
    0, 0, -3, 2, -8, -4, 2, 2, -8,
    -- filter=247 channel=58
    -4, 2, 0, 3, -5, -3, 0, 5, 8,
    -- filter=247 channel=59
    1, 2, -14, 0, -18, -5, -2, 0, 8,
    -- filter=247 channel=60
    -3, -7, 2, 0, 4, 0, -4, -4, 5,
    -- filter=247 channel=61
    1, 3, 7, 0, 3, 2, 3, -7, 0,
    -- filter=247 channel=62
    0, -2, -2, -1, 0, -2, -3, 0, 6,
    -- filter=247 channel=63
    -4, 2, -3, 5, 1, -6, -8, -3, 1,
    -- filter=247 channel=64
    0, -5, 3, 0, 0, 2, 5, -6, -6,
    -- filter=247 channel=65
    7, -5, -3, 0, -2, -4, 5, 0, -1,
    -- filter=247 channel=66
    -3, 6, -3, 0, 0, 4, 6, -7, -1,
    -- filter=247 channel=67
    4, 5, -2, -6, 4, 3, 1, 6, -4,
    -- filter=247 channel=68
    5, 1, 4, -2, -5, 8, 8, 1, -3,
    -- filter=247 channel=69
    -7, -3, 6, 0, 4, -5, -5, -6, -3,
    -- filter=247 channel=70
    -3, -12, 4, -17, -4, -1, -4, 0, -1,
    -- filter=247 channel=71
    8, 2, -1, 5, 5, -1, -2, -3, 9,
    -- filter=247 channel=72
    12, 9, -4, 0, -15, 2, -9, 3, 0,
    -- filter=247 channel=73
    1, 2, -1, -18, -1, 11, 9, 14, 1,
    -- filter=247 channel=74
    2, -17, 5, -2, -2, 7, 4, 8, -9,
    -- filter=247 channel=75
    4, 10, -11, -3, -10, -6, -3, 8, 19,
    -- filter=247 channel=76
    6, 5, 8, -8, -13, 5, -2, 0, 8,
    -- filter=247 channel=77
    3, 4, -1, 1, 0, 5, -1, 3, 1,
    -- filter=247 channel=78
    0, -4, -7, 0, -3, -5, 5, -4, -3,
    -- filter=247 channel=79
    0, -1, -8, -13, -22, 10, -6, 3, 15,
    -- filter=247 channel=80
    7, 5, -8, -5, -14, -7, -3, -1, 1,
    -- filter=247 channel=81
    0, -4, 3, 0, 4, 0, 0, -2, 5,
    -- filter=247 channel=82
    6, 1, 5, -2, 6, 5, -8, -4, -7,
    -- filter=247 channel=83
    8, 1, 0, -4, 2, -7, -2, 4, 0,
    -- filter=247 channel=84
    4, -1, 6, -11, -8, 2, 0, 10, -3,
    -- filter=247 channel=85
    1, 2, -3, 2, 2, -5, 6, 0, -1,
    -- filter=247 channel=86
    -5, -4, 5, -2, 4, 9, 11, 4, -3,
    -- filter=247 channel=87
    0, 0, 5, -7, 0, 12, 8, -2, -2,
    -- filter=247 channel=88
    3, 1, 0, -4, -3, 6, 0, 2, -8,
    -- filter=247 channel=89
    6, 11, -5, 0, -21, 5, -9, 4, 17,
    -- filter=247 channel=90
    -4, 4, 0, 7, -1, 1, -5, 1, -13,
    -- filter=247 channel=91
    6, -12, 6, -16, -10, 2, 16, 12, -8,
    -- filter=247 channel=92
    0, 2, -7, 2, 0, -1, -4, -8, 0,
    -- filter=247 channel=93
    6, -7, 0, -9, -4, 8, 12, 11, -7,
    -- filter=247 channel=94
    -1, 0, -1, -3, -5, 4, 5, -4, 4,
    -- filter=247 channel=95
    3, -1, 3, 0, 0, -1, -5, 0, 8,
    -- filter=247 channel=96
    0, 7, -1, 5, 4, -3, -8, 0, 4,
    -- filter=247 channel=97
    6, 13, 0, 14, 2, -1, 0, 1, 1,
    -- filter=247 channel=98
    6, 8, -9, -9, -9, -4, -5, 12, 10,
    -- filter=247 channel=99
    11, -4, 1, -14, -10, 11, -1, 2, -4,
    -- filter=247 channel=100
    5, -4, 2, -8, 1, 5, -4, 5, 6,
    -- filter=247 channel=101
    0, 3, -4, 0, 8, 5, 9, 4, 1,
    -- filter=247 channel=102
    2, 5, 6, 1, 3, 5, -4, 5, 1,
    -- filter=247 channel=103
    12, 12, -3, 4, -5, -11, -5, 5, 6,
    -- filter=247 channel=104
    15, 7, -6, -7, -7, -7, -6, 2, 2,
    -- filter=247 channel=105
    5, 3, 7, -8, -2, 4, -11, 2, 10,
    -- filter=247 channel=106
    5, -8, -2, -6, -3, 2, -2, 0, -3,
    -- filter=247 channel=107
    -1, -8, 10, -1, -1, 11, -6, 0, 10,
    -- filter=247 channel=108
    1, 0, 0, -2, -4, -2, 3, -2, 10,
    -- filter=247 channel=109
    8, -14, 0, -20, -10, 8, 5, 9, 8,
    -- filter=247 channel=110
    7, 9, -2, 4, -1, -6, -4, 3, 0,
    -- filter=247 channel=111
    0, 0, 1, 2, 3, 6, -3, 3, -4,
    -- filter=247 channel=112
    0, -1, -4, -10, -6, 3, 1, -3, 0,
    -- filter=247 channel=113
    9, 0, -1, 2, -15, 1, 1, 0, 4,
    -- filter=247 channel=114
    1, -8, -2, -22, -23, 14, 1, 20, 14,
    -- filter=247 channel=115
    1, 5, -5, 1, 0, -2, -3, 7, 1,
    -- filter=247 channel=116
    9, -5, 2, -15, -16, 0, -1, 7, -7,
    -- filter=247 channel=117
    -2, 7, -3, 0, -9, 0, 7, 5, -6,
    -- filter=247 channel=118
    6, 5, 5, 2, 4, -7, -2, 3, -5,
    -- filter=247 channel=119
    0, -3, 12, -8, 2, 3, 6, 7, -1,
    -- filter=247 channel=120
    -1, -19, 9, -28, 1, 23, 18, 18, -9,
    -- filter=247 channel=121
    5, -2, 0, -2, -11, 3, 2, 2, 6,
    -- filter=247 channel=122
    9, 9, -10, 0, 2, -8, 1, -4, -7,
    -- filter=247 channel=123
    3, -4, 2, -6, 6, 3, -5, 0, 3,
    -- filter=247 channel=124
    4, 1, 3, 0, 5, 1, -9, 2, 4,
    -- filter=247 channel=125
    10, 1, -11, -15, -3, 6, -1, -1, -1,
    -- filter=247 channel=126
    -2, 1, 4, 5, -14, -7, -10, 0, 15,
    -- filter=247 channel=127
    -6, 7, -6, -2, 1, 0, 0, 3, -2,
    -- filter=248 channel=0
    11, 11, 0, 12, -14, -14, 5, -10, -15,
    -- filter=248 channel=1
    5, 0, 2, 8, -7, -9, 14, -14, 1,
    -- filter=248 channel=2
    4, 0, 0, 3, -5, 7, -6, -2, -2,
    -- filter=248 channel=3
    5, 0, 1, -5, -5, -8, -7, -3, -4,
    -- filter=248 channel=4
    -7, 2, -9, -2, -8, -4, -6, 3, 0,
    -- filter=248 channel=5
    5, 2, 1, 8, -6, -1, -5, -9, -5,
    -- filter=248 channel=6
    9, 0, 0, 6, 5, 0, -1, 1, -2,
    -- filter=248 channel=7
    -7, -7, -2, -3, 0, -3, -5, 1, -2,
    -- filter=248 channel=8
    0, 11, 6, 10, 0, 4, -2, 5, 0,
    -- filter=248 channel=9
    -7, -6, 0, 0, 2, -6, -3, 3, 6,
    -- filter=248 channel=10
    6, 6, -1, 9, -2, -5, 0, 5, 3,
    -- filter=248 channel=11
    7, -6, 0, -2, -10, 4, -6, -7, 5,
    -- filter=248 channel=12
    7, 13, 0, 3, -3, 9, 13, 6, 5,
    -- filter=248 channel=13
    8, -2, 2, 15, 0, -5, 9, -7, 2,
    -- filter=248 channel=14
    -2, -3, 5, -1, -7, 6, 4, -3, 4,
    -- filter=248 channel=15
    12, -2, -4, 4, -15, -5, -2, -11, 2,
    -- filter=248 channel=16
    6, 3, 0, 4, -1, -1, 1, 9, 0,
    -- filter=248 channel=17
    1, 1, -5, 3, 4, -3, -4, -6, -2,
    -- filter=248 channel=18
    17, -3, -6, 17, -4, -16, 20, -23, 0,
    -- filter=248 channel=19
    0, 2, -4, 2, 0, 4, 3, 0, -5,
    -- filter=248 channel=20
    10, -7, -9, 10, -11, 0, 3, -10, -4,
    -- filter=248 channel=21
    2, -3, -6, -10, -6, 0, -1, 6, 5,
    -- filter=248 channel=22
    0, 4, -5, 4, -10, 4, 1, -5, -1,
    -- filter=248 channel=23
    3, -3, -7, 6, -6, -1, -6, 0, 3,
    -- filter=248 channel=24
    3, 1, 2, 7, 6, -6, -3, 3, 0,
    -- filter=248 channel=25
    -3, 8, 0, 6, -12, -8, 3, -10, 1,
    -- filter=248 channel=26
    0, -3, 0, -8, 4, 5, -2, 0, 0,
    -- filter=248 channel=27
    4, 7, -11, 16, -18, -6, 1, -5, 1,
    -- filter=248 channel=28
    5, 2, 1, 6, -6, 7, -6, -2, 3,
    -- filter=248 channel=29
    9, 3, -10, 5, -10, -7, 2, -19, -7,
    -- filter=248 channel=30
    8, -5, 1, -3, -3, -4, -7, -8, 0,
    -- filter=248 channel=31
    -7, -6, -12, -2, 0, 5, -13, 15, 14,
    -- filter=248 channel=32
    11, 2, 2, 13, -15, -3, 9, -19, 5,
    -- filter=248 channel=33
    -1, 9, 5, 9, -7, 0, 7, -7, -4,
    -- filter=248 channel=34
    14, 12, 4, 13, 3, -6, 6, 16, -1,
    -- filter=248 channel=35
    2, 0, 0, -4, 6, -2, -7, 2, -2,
    -- filter=248 channel=36
    1, 3, 3, 0, 6, 6, -2, 2, 15,
    -- filter=248 channel=37
    7, 9, -3, 3, -5, -1, 8, -1, -4,
    -- filter=248 channel=38
    3, 0, -2, -6, -8, 0, -6, -5, 2,
    -- filter=248 channel=39
    -7, -5, -9, -1, -5, -8, -2, -2, 7,
    -- filter=248 channel=40
    -2, 6, -1, -3, 7, 7, 2, -7, 1,
    -- filter=248 channel=41
    14, -2, 12, 29, 20, -9, 44, -1, 5,
    -- filter=248 channel=42
    -4, 1, 0, 4, 3, 1, 3, -9, -1,
    -- filter=248 channel=43
    -3, -1, 4, 8, -3, -7, 0, -4, 0,
    -- filter=248 channel=44
    7, 7, 1, -4, -10, 0, -7, 0, 9,
    -- filter=248 channel=45
    -3, -3, -3, -3, -9, -1, -4, 4, 5,
    -- filter=248 channel=46
    3, 0, 1, 10, 2, -4, 7, 6, 4,
    -- filter=248 channel=47
    -11, -3, -9, -8, -4, 1, 5, 10, 5,
    -- filter=248 channel=48
    3, -3, -13, 5, -14, -2, -2, -8, 8,
    -- filter=248 channel=49
    10, 0, -6, 3, -16, 1, 2, -5, -3,
    -- filter=248 channel=50
    -8, -1, -10, 5, -12, -3, -1, -4, 0,
    -- filter=248 channel=51
    -5, 1, 0, 0, 0, 6, -6, 3, -3,
    -- filter=248 channel=52
    12, 11, 3, 14, 1, 5, 2, 9, -2,
    -- filter=248 channel=53
    8, -1, 0, 1, 2, 2, 1, -7, 4,
    -- filter=248 channel=54
    3, 6, 1, 2, -5, -1, -3, -3, 2,
    -- filter=248 channel=55
    1, -5, -7, 17, -3, -2, 2, -10, 3,
    -- filter=248 channel=56
    4, -1, -1, 7, 8, 7, -1, 11, 2,
    -- filter=248 channel=57
    -5, 0, -3, 2, -7, 5, 10, -8, -6,
    -- filter=248 channel=58
    9, 0, -5, -3, -5, -2, -1, 2, -11,
    -- filter=248 channel=59
    6, -7, -6, 10, -3, 0, 9, -6, 1,
    -- filter=248 channel=60
    1, 3, -4, 3, -3, -2, 4, 4, 0,
    -- filter=248 channel=61
    9, 0, -6, 1, 5, -1, 0, 10, -1,
    -- filter=248 channel=62
    -3, 0, 2, 0, 1, -5, -2, -7, -3,
    -- filter=248 channel=63
    0, -2, -1, 0, 8, -7, 1, 2, 4,
    -- filter=248 channel=64
    7, 6, -2, -1, 4, 0, 0, 10, 2,
    -- filter=248 channel=65
    -4, -4, 5, -6, -3, -4, 3, -4, 4,
    -- filter=248 channel=66
    8, 4, 2, 15, 1, -5, 12, 4, 0,
    -- filter=248 channel=67
    -6, -1, -3, -1, 3, -3, 6, 7, 3,
    -- filter=248 channel=68
    -3, 0, -4, -1, -5, -6, -3, -4, 4,
    -- filter=248 channel=69
    -4, 4, -5, -3, -3, 0, -1, 3, 1,
    -- filter=248 channel=70
    0, 8, 2, -1, -8, -2, -5, -8, 13,
    -- filter=248 channel=71
    4, 1, 9, -8, -4, 4, 2, -6, -7,
    -- filter=248 channel=72
    5, -5, -4, -5, 0, 5, 1, 2, 12,
    -- filter=248 channel=73
    6, 6, -10, 12, -12, -8, -4, -13, 10,
    -- filter=248 channel=74
    9, 10, -7, 4, -9, 7, -2, 0, 8,
    -- filter=248 channel=75
    11, 2, 4, 8, -10, -11, 10, -13, -9,
    -- filter=248 channel=76
    8, -4, -3, 13, 1, -7, 6, 0, -5,
    -- filter=248 channel=77
    -6, 1, 0, 8, 5, -1, 7, 6, 0,
    -- filter=248 channel=78
    4, -2, -10, -5, -7, 0, -3, 7, -7,
    -- filter=248 channel=79
    16, 4, 7, 10, -10, -13, 14, -23, -6,
    -- filter=248 channel=80
    -3, -6, -5, -10, -2, -9, 0, 3, 4,
    -- filter=248 channel=81
    3, -2, -3, 2, 3, -2, 0, -6, 3,
    -- filter=248 channel=82
    5, 5, -1, -2, 5, -6, -3, -2, 2,
    -- filter=248 channel=83
    0, -1, -8, -10, -10, 3, -12, -1, 0,
    -- filter=248 channel=84
    0, -3, -6, 10, -15, -9, 6, 2, 9,
    -- filter=248 channel=85
    -1, -2, 4, 6, -6, 1, -7, 1, -1,
    -- filter=248 channel=86
    8, 12, 3, 18, 5, 3, 11, 3, -5,
    -- filter=248 channel=87
    11, 0, 1, 5, 3, 5, 1, -4, 0,
    -- filter=248 channel=88
    4, 5, 0, -4, 11, 10, -7, 17, 5,
    -- filter=248 channel=89
    0, 6, 1, 1, 1, -6, 9, -9, 9,
    -- filter=248 channel=90
    -2, -1, -4, -1, 6, 2, -6, 9, 9,
    -- filter=248 channel=91
    8, 6, -8, 0, -15, -4, -8, -9, 14,
    -- filter=248 channel=92
    -4, -5, -9, 5, 1, -8, 1, -2, 5,
    -- filter=248 channel=93
    7, 6, -9, -1, -14, 0, -4, 0, 1,
    -- filter=248 channel=94
    -6, 6, 4, 0, 0, 2, 1, -3, -5,
    -- filter=248 channel=95
    2, -1, 5, 3, 0, 8, 2, 6, -3,
    -- filter=248 channel=96
    -5, 0, 6, 1, 5, 1, 6, 3, -8,
    -- filter=248 channel=97
    -5, 0, 0, -11, 4, -2, -5, 4, -1,
    -- filter=248 channel=98
    -7, -2, -3, 2, -13, -12, 1, -9, -5,
    -- filter=248 channel=99
    9, 4, -13, 8, -12, -6, -15, 3, 0,
    -- filter=248 channel=100
    5, 5, 3, 1, 0, 0, 1, -1, 6,
    -- filter=248 channel=101
    -8, 0, -5, -9, 0, -1, -7, -3, 9,
    -- filter=248 channel=102
    0, 3, 6, 5, 1, -1, -3, 4, 4,
    -- filter=248 channel=103
    -9, 3, -1, -7, -8, 0, -7, 4, 0,
    -- filter=248 channel=104
    -1, 3, -10, -8, 3, -3, -10, 10, 13,
    -- filter=248 channel=105
    5, -3, 2, -2, -7, 0, 0, -11, -8,
    -- filter=248 channel=106
    6, 0, -3, 6, -2, -1, 9, 5, -2,
    -- filter=248 channel=107
    2, -2, 1, 13, -5, -4, 6, -10, -6,
    -- filter=248 channel=108
    11, -7, 0, 3, 4, -2, 8, -6, 4,
    -- filter=248 channel=109
    2, 0, -1, 10, -21, 0, 1, -15, 2,
    -- filter=248 channel=110
    -6, 5, 3, -2, 1, -2, 0, 3, 0,
    -- filter=248 channel=111
    9, -3, 10, 12, 7, -6, 0, 3, 5,
    -- filter=248 channel=112
    -2, 5, 3, -7, -1, 3, -1, -3, 5,
    -- filter=248 channel=113
    3, 11, -2, 4, -7, 0, 1, -3, -3,
    -- filter=248 channel=114
    21, 7, 1, 14, -19, -12, 7, -26, -6,
    -- filter=248 channel=115
    -5, -1, 6, 0, -1, 6, -5, 7, -6,
    -- filter=248 channel=116
    1, -2, 0, 5, -13, 0, 0, -8, 8,
    -- filter=248 channel=117
    5, 0, -4, 5, -2, 6, 0, 6, 9,
    -- filter=248 channel=118
    0, 0, 0, 0, -6, 0, 6, 5, 5,
    -- filter=248 channel=119
    13, 4, -6, 7, 6, -8, 0, 10, 2,
    -- filter=248 channel=120
    1, 2, -4, 9, -25, -2, -10, -13, 7,
    -- filter=248 channel=121
    8, 6, 0, 4, 0, -4, 7, -2, 3,
    -- filter=248 channel=122
    2, 0, 0, -13, -5, 9, -1, 16, 6,
    -- filter=248 channel=123
    3, -1, -5, 7, 6, -1, -1, 2, -1,
    -- filter=248 channel=124
    0, -5, -4, -2, 2, -4, 4, 0, -3,
    -- filter=248 channel=125
    0, 2, -13, 0, 0, 3, -7, 1, 12,
    -- filter=248 channel=126
    4, -6, 1, 13, 8, -1, 15, -2, -8,
    -- filter=248 channel=127
    9, 0, 0, 13, 3, -5, 9, 0, 6,
    -- filter=249 channel=0
    -15, -10, 2, -4, 0, 16, -10, 2, 10,
    -- filter=249 channel=1
    -10, -5, -8, -13, -8, 2, -5, 1, 7,
    -- filter=249 channel=2
    1, -1, 1, -6, -3, -7, -4, -2, -6,
    -- filter=249 channel=3
    -1, -3, 1, -2, -4, 11, -2, -7, -4,
    -- filter=249 channel=4
    -4, 1, -5, -1, -11, 7, -3, -14, -1,
    -- filter=249 channel=5
    0, -9, 0, -1, -1, -5, -10, 2, 5,
    -- filter=249 channel=6
    -4, -1, 7, -9, -8, 6, -1, 5, 1,
    -- filter=249 channel=7
    -1, 6, 3, 2, -5, 6, 2, -3, 0,
    -- filter=249 channel=8
    0, 7, 5, 1, 2, -2, -3, 6, -1,
    -- filter=249 channel=9
    6, 0, -2, 0, 3, -2, 0, -6, -6,
    -- filter=249 channel=10
    4, 4, 4, -4, 11, -4, 1, -4, -9,
    -- filter=249 channel=11
    6, 9, 9, -7, 4, 0, 0, -8, -6,
    -- filter=249 channel=12
    3, 0, 2, -7, -2, -4, -5, -6, 3,
    -- filter=249 channel=13
    -15, 12, 7, -8, 9, 5, -16, 0, 3,
    -- filter=249 channel=14
    5, 1, 0, 4, -3, -5, 5, 5, -6,
    -- filter=249 channel=15
    -16, 1, 15, -22, 3, 12, -11, -2, 8,
    -- filter=249 channel=16
    6, -9, -14, 5, 4, -3, -2, 1, -2,
    -- filter=249 channel=17
    -4, 6, -6, -2, -7, 2, 7, 5, 1,
    -- filter=249 channel=18
    -18, 0, 11, -27, 0, 20, -12, 7, 7,
    -- filter=249 channel=19
    4, 7, -6, 5, 1, -1, 3, -7, 0,
    -- filter=249 channel=20
    -3, 2, 12, -2, -8, 2, -11, -9, -3,
    -- filter=249 channel=21
    17, -2, -5, 17, 9, -11, -1, -3, -11,
    -- filter=249 channel=22
    -10, 3, 0, -11, -6, 12, -5, 5, -1,
    -- filter=249 channel=23
    0, 13, 19, -10, 14, 0, -9, 11, -9,
    -- filter=249 channel=24
    -5, 3, 1, 4, -4, -6, -3, -2, 6,
    -- filter=249 channel=25
    -10, 7, 1, -16, -4, 4, -13, -1, 0,
    -- filter=249 channel=26
    8, -2, 0, 8, 4, -2, -5, -8, -1,
    -- filter=249 channel=27
    -13, 2, 5, -21, 7, 7, -9, 13, 12,
    -- filter=249 channel=28
    6, -2, -5, -4, -2, -5, 3, 1, -6,
    -- filter=249 channel=29
    -9, 2, 6, -12, -6, -7, -2, 0, -1,
    -- filter=249 channel=30
    -2, -5, 8, -1, -1, 0, 4, 5, 3,
    -- filter=249 channel=31
    26, 21, -2, 15, 16, -13, 10, 6, -14,
    -- filter=249 channel=32
    -22, -1, 15, -23, -3, 7, -18, -1, 12,
    -- filter=249 channel=33
    -17, 0, 13, -9, 8, 0, -6, 7, 12,
    -- filter=249 channel=34
    -4, -3, 0, -14, 0, 5, -4, 3, -1,
    -- filter=249 channel=35
    0, 0, -6, -6, -3, 6, 4, 4, 0,
    -- filter=249 channel=36
    8, 15, -5, 16, 9, -5, 0, -3, -4,
    -- filter=249 channel=37
    -7, -10, -9, -11, 2, 9, -2, 3, 0,
    -- filter=249 channel=38
    -7, 7, 7, -1, -3, 4, 3, 0, 7,
    -- filter=249 channel=39
    0, -3, 7, 5, -2, 0, 6, -6, -4,
    -- filter=249 channel=40
    9, 10, 11, -4, 10, 0, 6, 0, 5,
    -- filter=249 channel=41
    -28, -16, 6, -25, -9, -14, -14, -7, 6,
    -- filter=249 channel=42
    -4, -7, 3, 1, -3, 4, -7, 7, 0,
    -- filter=249 channel=43
    -6, -3, -2, -15, -5, 13, 0, -6, -2,
    -- filter=249 channel=44
    -4, 2, -9, 0, 1, -5, -7, -5, 1,
    -- filter=249 channel=45
    8, 8, -4, 4, 0, 9, 7, 0, 2,
    -- filter=249 channel=46
    3, -1, -5, -4, -4, -4, -2, 2, 7,
    -- filter=249 channel=47
    10, 0, -16, 10, 2, -15, 1, -5, -7,
    -- filter=249 channel=48
    8, 0, 1, -4, -2, -9, -8, 0, 2,
    -- filter=249 channel=49
    -12, 8, 7, -13, -7, -1, -2, -4, 5,
    -- filter=249 channel=50
    -2, 11, 0, 1, 3, 0, 6, 8, 7,
    -- filter=249 channel=51
    3, 6, 0, 4, -6, -1, -6, 0, 1,
    -- filter=249 channel=52
    0, 10, 4, -5, 7, 4, -7, 0, 2,
    -- filter=249 channel=53
    4, 7, 9, 0, -4, 5, -3, 3, 0,
    -- filter=249 channel=54
    0, 3, 5, 2, 0, -3, -1, -4, -4,
    -- filter=249 channel=55
    -3, 1, 11, -6, 5, 0, -10, 8, -4,
    -- filter=249 channel=56
    -4, 7, 4, 3, 5, 0, 6, -7, -1,
    -- filter=249 channel=57
    -5, -3, -1, -10, -9, 0, -6, -8, -2,
    -- filter=249 channel=58
    3, 0, -9, -1, -5, -1, 1, -7, -3,
    -- filter=249 channel=59
    2, 2, -6, -4, 5, 4, -15, 4, -3,
    -- filter=249 channel=60
    -2, -4, -3, 5, 3, -2, -7, -2, 0,
    -- filter=249 channel=61
    8, 9, -5, -1, -1, -8, -7, -1, -10,
    -- filter=249 channel=62
    0, 3, 0, 6, -4, 1, -5, 6, 3,
    -- filter=249 channel=63
    -3, -5, -10, 10, -5, -8, 0, 0, -8,
    -- filter=249 channel=64
    -2, 7, 4, 11, 2, -5, 8, 0, 0,
    -- filter=249 channel=65
    6, 0, 2, 1, -2, 4, 0, 7, -5,
    -- filter=249 channel=66
    -12, -6, -10, -7, 0, 3, -2, -2, 7,
    -- filter=249 channel=67
    6, -6, -6, -4, -1, -3, 0, -6, -2,
    -- filter=249 channel=68
    3, 1, 2, 7, -7, -2, 7, -6, -6,
    -- filter=249 channel=69
    4, 3, 0, 2, -6, 2, 4, -5, 4,
    -- filter=249 channel=70
    -11, 9, 18, -6, 7, 5, -8, 7, 10,
    -- filter=249 channel=71
    -1, 0, 0, 4, 0, -4, 0, -5, 4,
    -- filter=249 channel=72
    14, 4, -6, 12, 12, -7, 1, 0, -9,
    -- filter=249 channel=73
    -7, 1, 7, -9, -5, -4, -12, 1, 0,
    -- filter=249 channel=74
    5, 14, -2, 0, 14, -2, 5, 10, 4,
    -- filter=249 channel=75
    -15, -3, 7, -10, -9, 0, -3, 3, 9,
    -- filter=249 channel=76
    -1, 9, 1, -8, 4, -3, -9, 0, -1,
    -- filter=249 channel=77
    -1, 5, 0, 2, -3, 0, 0, -3, 2,
    -- filter=249 channel=78
    -3, -2, -2, 4, 0, 0, 1, -3, 4,
    -- filter=249 channel=79
    -26, 0, 16, -35, 9, 17, -12, 10, 19,
    -- filter=249 channel=80
    16, 13, -9, 9, 3, -21, -11, 5, -8,
    -- filter=249 channel=81
    0, -5, -1, 2, -4, -5, 0, -2, 5,
    -- filter=249 channel=82
    3, 5, 6, -3, 0, -2, 2, 5, -4,
    -- filter=249 channel=83
    10, 8, -5, 4, -4, -6, 7, 2, 8,
    -- filter=249 channel=84
    -17, 8, 0, -7, -6, 2, -17, 5, 11,
    -- filter=249 channel=85
    0, 2, 0, -1, -4, -2, -4, -4, 1,
    -- filter=249 channel=86
    0, -3, -6, -8, 5, 1, -3, 10, 2,
    -- filter=249 channel=87
    -10, 1, 7, -10, -7, 1, -7, 2, 1,
    -- filter=249 channel=88
    12, 14, -3, 21, 0, -14, 1, -3, -8,
    -- filter=249 channel=89
    -8, 0, 0, -9, 9, -7, -17, 4, 4,
    -- filter=249 channel=90
    19, 12, 1, 20, 1, -8, 1, 6, -9,
    -- filter=249 channel=91
    -9, 6, 9, -18, 7, 0, -10, 14, 11,
    -- filter=249 channel=92
    -8, -1, 1, 1, -4, 7, 0, -3, 2,
    -- filter=249 channel=93
    1, -4, -5, 1, -12, -10, -5, -8, -6,
    -- filter=249 channel=94
    2, 0, 7, -6, 3, 1, -3, -3, 4,
    -- filter=249 channel=95
    -2, -1, -6, -5, -2, 3, -8, -1, -6,
    -- filter=249 channel=96
    -7, -7, 6, -5, -3, 6, 1, -2, 4,
    -- filter=249 channel=97
    6, 5, 1, 3, -4, -4, -2, -1, 5,
    -- filter=249 channel=98
    -15, -1, 4, -12, 6, -8, -16, 11, -3,
    -- filter=249 channel=99
    9, 12, 8, 12, 0, -5, -4, -1, -10,
    -- filter=249 channel=100
    -6, 0, 5, -6, -5, -4, 4, 0, 0,
    -- filter=249 channel=101
    4, -3, 5, -2, -1, 0, -9, -8, 1,
    -- filter=249 channel=102
    -1, -1, 2, -4, 6, -2, -5, 1, 4,
    -- filter=249 channel=103
    8, -6, -3, 5, -8, -7, -7, -5, -6,
    -- filter=249 channel=104
    18, 10, -9, 10, 10, -10, 0, -1, -13,
    -- filter=249 channel=105
    0, -7, 0, -3, -5, 2, -8, -6, -6,
    -- filter=249 channel=106
    5, 4, 3, 0, 1, 0, 6, 0, 3,
    -- filter=249 channel=107
    -19, 6, 10, -19, 0, 2, -2, 8, 0,
    -- filter=249 channel=108
    -7, -13, 5, -4, -4, -8, -9, -2, -8,
    -- filter=249 channel=109
    -18, 8, 14, -14, 1, 11, -18, 2, 3,
    -- filter=249 channel=110
    3, 9, -4, 5, -3, -12, 0, 5, -8,
    -- filter=249 channel=111
    3, -8, -2, -1, -5, -7, 5, 4, 6,
    -- filter=249 channel=112
    0, -2, 3, 1, 2, -1, 4, 13, -3,
    -- filter=249 channel=113
    0, 0, 6, -1, 8, 0, -7, 8, -7,
    -- filter=249 channel=114
    -34, 1, 13, -34, 4, 10, -23, 7, 14,
    -- filter=249 channel=115
    -5, -6, -6, -8, 4, 3, 0, -3, 4,
    -- filter=249 channel=116
    -7, 2, 2, 1, 5, -3, -3, -2, 3,
    -- filter=249 channel=117
    7, 10, -2, 7, 8, 1, 5, 3, -2,
    -- filter=249 channel=118
    3, -1, -1, -4, 1, 1, -1, 1, 3,
    -- filter=249 channel=119
    -10, -5, 3, 0, -9, 4, -2, -3, 10,
    -- filter=249 channel=120
    -2, 8, 10, -19, 11, 0, -6, 15, 2,
    -- filter=249 channel=121
    -9, 0, -3, -9, 0, 1, -10, -1, 4,
    -- filter=249 channel=122
    15, 5, -21, 24, 0, -16, 9, -4, -7,
    -- filter=249 channel=123
    4, -4, -1, 5, -5, 3, 2, -6, -4,
    -- filter=249 channel=124
    -6, -6, 3, 0, 3, 2, 0, -2, -5,
    -- filter=249 channel=125
    7, 12, -6, 8, 15, -3, -2, 10, -3,
    -- filter=249 channel=126
    -18, -10, 5, -11, -2, 7, -8, -10, 5,
    -- filter=249 channel=127
    -2, -7, 4, -10, 0, -1, -3, -2, -6,
    -- filter=250 channel=0
    -17, -10, 1, -7, -1, 0, 8, 14, 0,
    -- filter=250 channel=1
    -3, 0, 2, 3, 3, -12, 0, -4, -2,
    -- filter=250 channel=2
    4, -6, -2, 9, 7, 5, -1, 3, -2,
    -- filter=250 channel=3
    -12, -12, -4, -14, -15, -12, 5, 14, 5,
    -- filter=250 channel=4
    2, -7, -9, 6, -6, -8, 12, 13, -3,
    -- filter=250 channel=5
    -7, 7, 3, -2, 3, -1, 8, 6, 0,
    -- filter=250 channel=6
    -10, -1, -3, -7, 2, 1, -1, 4, 10,
    -- filter=250 channel=7
    0, 3, -1, 5, 6, -5, 5, 0, 1,
    -- filter=250 channel=8
    -4, 5, -7, -4, -9, -1, -2, 0, -2,
    -- filter=250 channel=9
    2, 6, -1, 7, -7, 4, 5, 7, 5,
    -- filter=250 channel=10
    -6, -9, 0, 0, -9, -4, 4, 4, 1,
    -- filter=250 channel=11
    3, -7, -1, 6, 0, 12, -3, -3, 4,
    -- filter=250 channel=12
    7, -4, -2, 8, 2, -3, 1, 0, -3,
    -- filter=250 channel=13
    -6, -4, 2, 1, -2, -7, 2, 7, 7,
    -- filter=250 channel=14
    -3, 4, 5, -1, 1, 0, -3, 2, 2,
    -- filter=250 channel=15
    -4, -14, -9, -7, 2, 11, -2, 8, 14,
    -- filter=250 channel=16
    2, -4, -6, -3, -9, -7, 0, 0, 2,
    -- filter=250 channel=17
    1, -2, 2, 4, -3, -5, 5, 0, -1,
    -- filter=250 channel=18
    -10, -15, -8, 2, 10, 15, 7, 11, 14,
    -- filter=250 channel=19
    4, 0, 6, 3, -6, -6, -6, 1, 3,
    -- filter=250 channel=20
    0, -2, 0, -5, 1, 24, 0, 1, 9,
    -- filter=250 channel=21
    -7, -2, -9, -2, -4, -5, -9, -11, -13,
    -- filter=250 channel=22
    -2, 2, 3, -2, 6, -7, 3, 1, 0,
    -- filter=250 channel=23
    -2, -14, -7, -9, -3, 5, 9, 4, 12,
    -- filter=250 channel=24
    5, -2, 6, 1, -4, 0, 2, -5, -1,
    -- filter=250 channel=25
    -7, 5, 0, 4, -7, 0, 14, 2, -7,
    -- filter=250 channel=26
    -5, -4, 4, 7, 0, 5, -3, 3, -7,
    -- filter=250 channel=27
    -3, -5, -9, 2, -6, 2, 7, 0, -7,
    -- filter=250 channel=28
    -5, 4, 0, -6, 5, 5, -3, -3, 3,
    -- filter=250 channel=29
    0, -2, 4, -2, 15, 23, -3, -3, 14,
    -- filter=250 channel=30
    -1, -1, 3, 4, -7, 0, 12, 0, -6,
    -- filter=250 channel=31
    -10, 3, 0, -2, -8, -12, 1, -4, -9,
    -- filter=250 channel=32
    -14, -9, 1, -2, 3, 4, 2, 13, 9,
    -- filter=250 channel=33
    -3, -14, 0, -9, 0, 0, 1, 6, 2,
    -- filter=250 channel=34
    -3, 2, -8, -3, 8, -4, 0, 4, -2,
    -- filter=250 channel=35
    -3, -4, -2, -4, 0, 3, 1, -3, -5,
    -- filter=250 channel=36
    10, -6, 2, 2, 7, 6, 5, -3, -8,
    -- filter=250 channel=37
    -4, -13, 2, 6, -13, -5, 4, -5, -7,
    -- filter=250 channel=38
    3, 2, 0, 0, -1, 3, 9, 0, -2,
    -- filter=250 channel=39
    -2, 5, 9, 3, 9, 8, 3, 7, 10,
    -- filter=250 channel=40
    -2, 2, 5, -2, 5, 6, -9, -6, 6,
    -- filter=250 channel=41
    -8, 0, -1, 3, 14, -4, -2, 16, -5,
    -- filter=250 channel=42
    -7, -7, 0, 0, 4, -3, -1, 5, 1,
    -- filter=250 channel=43
    -1, -5, 1, -4, -1, 6, -2, 1, 4,
    -- filter=250 channel=44
    -13, -4, -2, -5, -11, -14, 10, -10, -8,
    -- filter=250 channel=45
    -3, -1, -3, 5, -3, -4, 6, 6, 3,
    -- filter=250 channel=46
    -3, 0, 2, -1, 6, -3, 0, -3, -4,
    -- filter=250 channel=47
    -8, -11, -5, -10, -7, -14, -1, 0, -8,
    -- filter=250 channel=48
    1, -4, -7, 2, -2, -20, 9, 0, -4,
    -- filter=250 channel=49
    -4, -6, -4, 8, 6, 6, 1, 8, 13,
    -- filter=250 channel=50
    -1, -4, -1, -4, -7, -1, 0, -1, 4,
    -- filter=250 channel=51
    -3, 3, -2, 2, 0, -3, -1, 6, 6,
    -- filter=250 channel=52
    -5, -6, -6, 3, -4, 2, -1, 0, -7,
    -- filter=250 channel=53
    -2, -6, 5, -5, -2, 12, -2, -4, 8,
    -- filter=250 channel=54
    0, -5, -6, 3, -2, 7, -1, 1, -7,
    -- filter=250 channel=55
    -7, -8, 0, 2, -1, 15, 0, 1, 11,
    -- filter=250 channel=56
    -7, 4, -7, -3, -2, -1, -7, 1, 4,
    -- filter=250 channel=57
    -5, 3, -1, -7, 5, -1, 3, 7, -4,
    -- filter=250 channel=58
    1, 6, 4, 6, 8, 3, 1, 3, 0,
    -- filter=250 channel=59
    -2, -8, -11, -7, 0, -11, 12, 6, -3,
    -- filter=250 channel=60
    -2, 3, 2, 7, -1, 0, 0, -7, -4,
    -- filter=250 channel=61
    4, 3, 2, -5, 5, 6, 0, -6, -5,
    -- filter=250 channel=62
    0, -5, 6, 1, 3, -2, -3, 2, 4,
    -- filter=250 channel=63
    0, 1, 0, -2, 8, 6, 9, 4, 0,
    -- filter=250 channel=64
    1, -6, -3, 6, -4, 6, -4, 1, -2,
    -- filter=250 channel=65
    1, 1, 1, 6, -7, 4, 2, -6, 7,
    -- filter=250 channel=66
    1, 5, 10, 2, 4, 7, 3, -1, 0,
    -- filter=250 channel=67
    2, 6, 5, 3, 5, 1, 0, 0, 1,
    -- filter=250 channel=68
    7, -5, 6, 6, -2, 2, 6, -4, -1,
    -- filter=250 channel=69
    2, 3, 4, 5, -5, 1, -5, 2, 7,
    -- filter=250 channel=70
    -4, -7, -5, -5, -2, -9, 11, 2, -1,
    -- filter=250 channel=71
    -3, -10, -5, -6, -6, 2, 1, 1, 4,
    -- filter=250 channel=72
    6, 0, -10, 2, -5, -6, 2, -3, -9,
    -- filter=250 channel=73
    0, 0, 0, -1, 7, 3, -3, 0, 9,
    -- filter=250 channel=74
    -1, 0, -4, -2, -7, 1, -5, 0, -9,
    -- filter=250 channel=75
    -11, -14, -4, -3, -5, -1, 2, 12, 6,
    -- filter=250 channel=76
    2, -6, 7, -8, 2, 19, 1, -2, 14,
    -- filter=250 channel=77
    -6, -6, 4, -4, -5, 5, 4, 1, -5,
    -- filter=250 channel=78
    4, 1, -4, -5, 0, 7, 1, 9, 5,
    -- filter=250 channel=79
    -18, -17, 4, -6, -4, 10, 4, 5, 16,
    -- filter=250 channel=80
    0, -6, 0, 2, -11, -8, 6, 1, -4,
    -- filter=250 channel=81
    1, 0, 4, 0, -5, -3, 4, -2, 4,
    -- filter=250 channel=82
    -7, -3, 4, 0, 2, -5, -4, -2, -4,
    -- filter=250 channel=83
    3, 0, -1, -4, 0, 3, 1, 6, -8,
    -- filter=250 channel=84
    -8, -4, 6, -4, 2, 8, -2, 10, 12,
    -- filter=250 channel=85
    4, 6, -1, -2, -3, -1, 5, 0, 7,
    -- filter=250 channel=86
    -6, 7, 5, -4, 2, 5, 0, 1, -6,
    -- filter=250 channel=87
    3, 3, 7, 4, -2, 2, 3, 2, 3,
    -- filter=250 channel=88
    10, 4, 0, 7, -1, -6, -8, -7, 0,
    -- filter=250 channel=89
    0, -16, -3, -5, -6, -6, 11, 8, 5,
    -- filter=250 channel=90
    4, 5, -2, -4, 1, -1, -9, -6, -12,
    -- filter=250 channel=91
    -11, -13, 0, 1, 1, -4, 11, 6, 2,
    -- filter=250 channel=92
    -7, 5, -7, -1, 0, 3, -1, 2, -4,
    -- filter=250 channel=93
    -5, -6, -9, -3, -6, -4, 5, -2, -11,
    -- filter=250 channel=94
    0, -4, 4, 6, 6, 4, -1, 3, 1,
    -- filter=250 channel=95
    3, 1, 3, 0, 0, 6, -4, 0, -2,
    -- filter=250 channel=96
    2, 1, 6, -2, 6, 4, 1, 3, -4,
    -- filter=250 channel=97
    -2, -6, -7, -4, -1, -7, 3, 2, -1,
    -- filter=250 channel=98
    -2, 1, -6, -4, -7, -2, 6, 0, -9,
    -- filter=250 channel=99
    -3, -3, 0, 9, -4, 1, 8, -3, 2,
    -- filter=250 channel=100
    2, -4, -2, 3, -3, 1, -3, 2, -3,
    -- filter=250 channel=101
    -3, 3, -9, 1, -7, 0, 7, 8, -4,
    -- filter=250 channel=102
    -3, -2, 0, -1, -5, -1, 4, 3, -4,
    -- filter=250 channel=103
    -10, -11, 0, -12, -1, -14, 0, -5, 0,
    -- filter=250 channel=104
    4, -7, 0, -4, -5, -3, 8, -3, -12,
    -- filter=250 channel=105
    -10, -5, 5, 3, 7, 12, -1, 6, 17,
    -- filter=250 channel=106
    1, 1, -6, -3, 6, 7, -2, 2, -1,
    -- filter=250 channel=107
    -12, -11, 2, 0, 3, 3, 1, 0, 14,
    -- filter=250 channel=108
    -8, 7, 5, 1, 0, 2, 0, 8, 9,
    -- filter=250 channel=109
    0, -6, 3, 8, -2, 3, 7, -2, 0,
    -- filter=250 channel=110
    -5, 0, 0, 6, -10, 0, 4, 2, 4,
    -- filter=250 channel=111
    1, 6, 2, -7, 8, 6, 0, -2, 1,
    -- filter=250 channel=112
    2, 5, 4, 4, -3, -2, -2, 2, -1,
    -- filter=250 channel=113
    1, -6, -13, -3, -4, -7, 1, 0, -6,
    -- filter=250 channel=114
    -10, -14, -3, -1, 13, 14, 12, 22, 22,
    -- filter=250 channel=115
    6, 0, 2, -5, 7, -6, -4, 1, 6,
    -- filter=250 channel=116
    -1, 5, -3, -1, 0, 0, 6, 10, 1,
    -- filter=250 channel=117
    6, -4, -2, 3, 0, -4, -1, -5, 6,
    -- filter=250 channel=118
    1, 0, 5, 0, -2, 4, 0, 4, 5,
    -- filter=250 channel=119
    4, 0, -6, 9, 0, 8, 2, 0, -5,
    -- filter=250 channel=120
    -8, -5, 2, -6, 0, 3, 1, -1, 10,
    -- filter=250 channel=121
    0, -4, -1, 1, -5, -9, 5, 0, 0,
    -- filter=250 channel=122
    -14, -12, -17, -3, -13, -12, -9, -3, -15,
    -- filter=250 channel=123
    4, 3, 2, -5, 0, -2, -3, -2, 0,
    -- filter=250 channel=124
    -7, -4, 11, -10, -1, 14, -1, 6, 8,
    -- filter=250 channel=125
    5, -3, -6, 2, 2, -8, 0, 4, 0,
    -- filter=250 channel=126
    -10, -10, -9, -1, 0, 7, 0, 9, 6,
    -- filter=250 channel=127
    0, 8, -1, 0, 0, -4, -7, 6, -6,
    -- filter=251 channel=0
    -8, -11, 1, -13, -29, -1, 0, -7, 4,
    -- filter=251 channel=1
    1, 0, 11, -5, -16, 7, -6, -4, -2,
    -- filter=251 channel=2
    2, -4, 3, 1, 3, 6, 0, 0, -4,
    -- filter=251 channel=3
    -7, -9, 6, -15, -15, 2, -8, -5, 0,
    -- filter=251 channel=4
    -3, -8, 3, 0, -15, 13, -4, -6, -6,
    -- filter=251 channel=5
    -11, -8, -3, -10, -2, 0, 2, -2, 3,
    -- filter=251 channel=6
    -1, -3, 0, -1, -10, 5, -2, 1, 3,
    -- filter=251 channel=7
    -1, 0, -7, 7, -3, 1, -2, -5, 3,
    -- filter=251 channel=8
    -4, 2, 9, 0, 0, 5, -6, 5, 6,
    -- filter=251 channel=9
    0, -1, 0, 6, 3, 5, -5, 3, -6,
    -- filter=251 channel=10
    -2, 7, -13, 0, 20, -9, 7, 13, 2,
    -- filter=251 channel=11
    5, -3, 0, 4, 3, -3, 1, 5, -1,
    -- filter=251 channel=12
    2, 3, -3, 11, 6, 6, 10, 6, -1,
    -- filter=251 channel=13
    6, -7, -4, -3, -2, -3, 3, -3, 2,
    -- filter=251 channel=14
    5, -4, 4, -3, 6, -4, 4, 0, 1,
    -- filter=251 channel=15
    6, -17, -3, -4, -7, 3, 7, -4, 15,
    -- filter=251 channel=16
    3, 6, -4, 4, 12, -2, -8, 5, 0,
    -- filter=251 channel=17
    -5, 6, 4, 0, -4, 2, -7, 4, -2,
    -- filter=251 channel=18
    -3, -17, 0, -15, -25, 0, -4, -10, 7,
    -- filter=251 channel=19
    -5, -6, 7, -4, 5, 0, -6, -2, -3,
    -- filter=251 channel=20
    0, -6, -8, 5, -2, 5, 4, 4, 7,
    -- filter=251 channel=21
    2, 18, -17, 10, 36, -10, 0, 5, -13,
    -- filter=251 channel=22
    -9, -6, 0, 0, -5, 4, 3, -2, 5,
    -- filter=251 channel=23
    -1, -5, -1, -6, -1, -7, -4, 0, 5,
    -- filter=251 channel=24
    -6, 0, 3, 6, 4, 3, 6, 3, 5,
    -- filter=251 channel=25
    -8, -5, -6, -2, -2, 2, -1, -2, -4,
    -- filter=251 channel=26
    -10, 1, -1, 2, 11, -5, 1, 0, -11,
    -- filter=251 channel=27
    -8, -10, 1, -10, -3, 16, -4, -10, 13,
    -- filter=251 channel=28
    -6, -7, -1, 6, 5, -6, -5, -6, 2,
    -- filter=251 channel=29
    4, 0, 0, 10, -2, 1, 12, 3, 3,
    -- filter=251 channel=30
    -4, 0, -1, -7, -8, 6, 6, -10, 7,
    -- filter=251 channel=31
    -7, 2, -23, 3, 36, -19, -2, 5, -10,
    -- filter=251 channel=32
    2, -3, 1, -13, -13, 4, 8, -10, 7,
    -- filter=251 channel=33
    -6, -11, 2, -10, -7, 12, 1, -10, 10,
    -- filter=251 channel=34
    8, -1, 2, 6, -1, -5, 11, -3, 12,
    -- filter=251 channel=35
    -1, 6, 2, 0, 0, 0, 4, 1, -5,
    -- filter=251 channel=36
    4, 10, -17, 5, 20, -2, 8, -1, -8,
    -- filter=251 channel=37
    -11, 4, 9, -4, -10, 12, -9, -8, -2,
    -- filter=251 channel=38
    1, -5, 1, -7, 3, 3, -7, -3, -6,
    -- filter=251 channel=39
    5, 0, 3, 0, -5, 3, 3, -5, 8,
    -- filter=251 channel=40
    2, -8, -8, -4, -4, -3, 1, -3, -1,
    -- filter=251 channel=41
    17, 12, 1, 14, -2, -6, 9, 1, -7,
    -- filter=251 channel=42
    -6, -8, 7, -8, 5, 1, -1, 0, 2,
    -- filter=251 channel=43
    -1, -14, 0, -9, -17, 3, -11, -3, 1,
    -- filter=251 channel=44
    -1, 7, 0, -7, 2, 6, -9, -5, -4,
    -- filter=251 channel=45
    -4, -10, 3, -6, -9, 1, 2, -12, -5,
    -- filter=251 channel=46
    0, 3, 0, -4, -2, -4, -1, -1, -5,
    -- filter=251 channel=47
    -10, 14, -11, 0, 23, -2, -7, 1, -15,
    -- filter=251 channel=48
    -8, 4, -15, 0, 12, 1, 3, 1, -12,
    -- filter=251 channel=49
    -9, -12, 0, -6, -7, 5, 2, -9, 3,
    -- filter=251 channel=50
    -5, -6, -2, 4, -2, -1, 0, -8, -5,
    -- filter=251 channel=51
    -5, 3, 3, -1, -5, -7, 1, -4, 1,
    -- filter=251 channel=52
    4, -2, 0, 0, 7, 7, 3, 2, 4,
    -- filter=251 channel=53
    -2, -8, -8, 5, -5, -2, 5, 3, -5,
    -- filter=251 channel=54
    -3, -5, 0, -4, -5, 6, 2, -1, 3,
    -- filter=251 channel=55
    2, -6, -14, 8, -3, -8, 16, 0, 5,
    -- filter=251 channel=56
    -2, -5, 0, 6, 10, 7, 0, -2, 10,
    -- filter=251 channel=57
    -7, 6, -4, 3, 1, -4, 4, 3, -7,
    -- filter=251 channel=58
    0, -1, 4, -1, 0, 0, -2, 5, 3,
    -- filter=251 channel=59
    -8, 7, -15, 2, 11, 5, 6, 6, -4,
    -- filter=251 channel=60
    1, -1, 6, 0, 6, -4, -2, 6, -4,
    -- filter=251 channel=61
    3, 0, -5, 11, 9, 0, 1, 10, 0,
    -- filter=251 channel=62
    2, -3, 7, 1, 4, 7, 4, 0, 4,
    -- filter=251 channel=63
    6, 0, -4, 2, 12, -1, 0, 4, -8,
    -- filter=251 channel=64
    7, -4, -5, 8, 2, -2, 1, 10, 2,
    -- filter=251 channel=65
    6, 0, 1, -5, -4, -4, -7, 2, 6,
    -- filter=251 channel=66
    7, 8, -5, 13, -7, -4, 5, -2, 8,
    -- filter=251 channel=67
    -6, -9, 1, -4, -5, 0, 0, 6, -6,
    -- filter=251 channel=68
    -1, -2, -2, -1, -5, -7, 3, -8, 3,
    -- filter=251 channel=69
    -5, -5, 0, 6, 4, -9, -6, -7, 0,
    -- filter=251 channel=70
    6, -12, 7, -11, -13, 0, 3, -4, 9,
    -- filter=251 channel=71
    3, 5, -4, 0, 0, -3, -8, -7, -3,
    -- filter=251 channel=72
    -4, 8, -28, 12, 21, -16, 10, 11, -6,
    -- filter=251 channel=73
    -7, -11, 1, 1, -7, 1, 6, -7, 8,
    -- filter=251 channel=74
    -1, 1, -8, 8, 7, 3, 1, 4, 3,
    -- filter=251 channel=75
    -4, -2, 5, -2, -4, 9, 1, -7, 0,
    -- filter=251 channel=76
    9, 0, -5, 1, -2, -2, 0, -4, 1,
    -- filter=251 channel=77
    -4, -4, 4, 2, -1, -1, 0, 3, -1,
    -- filter=251 channel=78
    -7, -1, -1, -1, -1, 6, -1, 0, 0,
    -- filter=251 channel=79
    -5, -11, 12, -25, -23, 12, -4, -12, 11,
    -- filter=251 channel=80
    2, 2, -22, 11, 25, -9, 11, 12, -16,
    -- filter=251 channel=81
    1, -5, -5, -2, 1, -6, 3, -4, -1,
    -- filter=251 channel=82
    4, 0, -1, 0, 3, 6, -3, -1, -1,
    -- filter=251 channel=83
    0, -3, -2, 7, 9, -1, 3, -4, -2,
    -- filter=251 channel=84
    -4, -8, -3, 0, -16, 10, 1, -12, 0,
    -- filter=251 channel=85
    -5, 2, -3, -5, -2, -2, 7, -6, 5,
    -- filter=251 channel=86
    -5, -1, 1, 2, -6, 0, 0, 3, 0,
    -- filter=251 channel=87
    6, -2, 9, 0, 0, 3, -2, -4, 2,
    -- filter=251 channel=88
    1, 7, -9, 17, 23, -14, -1, 4, -4,
    -- filter=251 channel=89
    6, -12, -21, 5, -5, -8, 3, 11, 0,
    -- filter=251 channel=90
    -2, 13, -14, 9, 14, 0, -3, 15, 0,
    -- filter=251 channel=91
    -10, 0, 3, -10, -13, 3, 4, -6, 4,
    -- filter=251 channel=92
    10, -7, 1, -3, -6, -5, -5, 1, 2,
    -- filter=251 channel=93
    -1, 12, -9, 0, 17, 0, -4, -7, -13,
    -- filter=251 channel=94
    1, -1, -3, 4, 5, 4, 5, -3, 1,
    -- filter=251 channel=95
    0, 6, -4, -7, -2, 7, -3, 5, -5,
    -- filter=251 channel=96
    0, 2, -8, 3, 3, 3, 1, -6, -1,
    -- filter=251 channel=97
    9, -3, -6, 0, 2, 6, -6, 4, -8,
    -- filter=251 channel=98
    1, -8, -12, -12, 0, 0, -2, -2, -3,
    -- filter=251 channel=99
    3, 2, -14, 4, 29, -8, 2, 2, 2,
    -- filter=251 channel=100
    3, 6, -4, 3, 10, -1, 9, 0, -2,
    -- filter=251 channel=101
    -5, -3, 4, 3, -5, -2, 6, -3, -4,
    -- filter=251 channel=102
    -2, 0, 0, 0, 6, 7, -3, -3, 5,
    -- filter=251 channel=103
    1, 8, -19, -1, 22, -3, -10, 8, -14,
    -- filter=251 channel=104
    -7, 4, -14, 14, 22, -1, -5, 6, -4,
    -- filter=251 channel=105
    6, -2, -2, 1, 1, -2, -1, 1, 3,
    -- filter=251 channel=106
    6, 3, -5, 0, 1, 4, 0, 3, 0,
    -- filter=251 channel=107
    -11, -12, 0, -17, -23, -4, -13, -14, 8,
    -- filter=251 channel=108
    1, -7, -6, 0, -7, -4, -5, 3, -6,
    -- filter=251 channel=109
    0, -3, -4, 3, 2, 11, 15, -3, 6,
    -- filter=251 channel=110
    5, -1, -8, 0, 13, -14, 3, 4, -6,
    -- filter=251 channel=111
    -4, 1, 6, 4, 1, 2, 0, -2, -4,
    -- filter=251 channel=112
    -8, -2, -5, -9, -8, -5, -9, -10, 0,
    -- filter=251 channel=113
    0, 0, 0, -3, 10, -1, 0, 0, 10,
    -- filter=251 channel=114
    -7, -28, 9, -27, -37, 4, -8, -20, 8,
    -- filter=251 channel=115
    -5, -3, -4, -5, 0, 1, 1, 1, 0,
    -- filter=251 channel=116
    -6, -2, -15, 9, 9, -1, 11, -3, -1,
    -- filter=251 channel=117
    0, 3, -2, -6, -3, 0, 0, -6, -3,
    -- filter=251 channel=118
    -7, 4, 2, -2, 1, 4, 2, -6, 6,
    -- filter=251 channel=119
    0, 7, 1, 8, 11, 0, 4, 9, 12,
    -- filter=251 channel=120
    -8, -9, -6, -3, 0, 6, -4, -2, 16,
    -- filter=251 channel=121
    15, 0, 0, 12, 8, -2, 10, -1, 0,
    -- filter=251 channel=122
    -3, 20, -26, 8, 49, -5, -8, 15, -25,
    -- filter=251 channel=123
    5, -4, 3, 12, -3, 2, 7, 6, -1,
    -- filter=251 channel=124
    4, 0, 4, -8, -7, 3, 0, 5, -4,
    -- filter=251 channel=125
    -10, 5, -19, 3, 23, 5, 4, 6, 0,
    -- filter=251 channel=126
    0, -8, 2, 1, -2, 5, 7, -1, 8,
    -- filter=251 channel=127
    5, -5, -1, 2, -4, 7, 9, 4, -6,
    -- filter=252 channel=0
    -6, 7, 13, -18, -6, 7, -15, -12, 15,
    -- filter=252 channel=1
    -2, -2, 6, -6, 5, 11, -14, -6, 8,
    -- filter=252 channel=2
    2, -8, 0, 1, -2, 4, -4, 0, 3,
    -- filter=252 channel=3
    3, 7, 3, 9, -6, -2, 0, -8, 8,
    -- filter=252 channel=4
    -9, -13, -15, 2, -8, 2, 1, -2, 1,
    -- filter=252 channel=5
    -4, -2, -3, 0, 8, 0, -13, 8, 6,
    -- filter=252 channel=6
    5, 6, -4, -7, -1, -4, 1, 0, -6,
    -- filter=252 channel=7
    7, -5, 1, 1, 0, 0, -1, 3, 2,
    -- filter=252 channel=8
    0, -4, -2, -7, -1, 11, -9, 2, 3,
    -- filter=252 channel=9
    -5, -4, -7, -6, 6, 0, -5, 1, -4,
    -- filter=252 channel=10
    6, 10, 2, 0, -6, -5, 0, 2, -2,
    -- filter=252 channel=11
    7, -7, 3, -5, -3, 0, 3, -12, 1,
    -- filter=252 channel=12
    -10, 0, 7, 0, 2, 5, -2, -1, 8,
    -- filter=252 channel=13
    0, 4, 4, -2, -3, -5, 0, -7, 0,
    -- filter=252 channel=14
    0, 0, 0, 4, -3, 5, 5, -2, 7,
    -- filter=252 channel=15
    8, 8, 5, -9, -9, 5, -8, -10, 7,
    -- filter=252 channel=16
    2, -4, -1, 6, 4, -1, -4, 0, 6,
    -- filter=252 channel=17
    1, 5, -1, 3, 0, 2, -7, -3, 3,
    -- filter=252 channel=18
    6, 14, 7, -1, -17, 7, -5, -22, -2,
    -- filter=252 channel=19
    -5, 1, 1, 6, 0, 5, 3, 3, 0,
    -- filter=252 channel=20
    -3, -5, 8, -2, -14, -2, 10, -7, -3,
    -- filter=252 channel=21
    -1, 3, -11, -3, 0, 3, -1, 4, -2,
    -- filter=252 channel=22
    -6, 7, 1, -1, -1, 10, -6, -5, 5,
    -- filter=252 channel=23
    8, 8, 8, -9, -1, 12, -3, -5, 19,
    -- filter=252 channel=24
    -3, -3, 0, -4, 5, 0, 1, 0, -4,
    -- filter=252 channel=25
    -6, 4, -6, 0, 3, 4, -1, -6, 6,
    -- filter=252 channel=26
    -9, -5, -4, 6, -5, -2, -8, 9, 7,
    -- filter=252 channel=27
    -7, -5, 6, -4, -4, 14, -13, -12, 16,
    -- filter=252 channel=28
    -1, 1, 7, 1, -2, 0, -5, -5, -1,
    -- filter=252 channel=29
    0, 0, 3, 0, -4, -8, 10, -16, -1,
    -- filter=252 channel=30
    1, -5, -9, -7, -10, 1, -2, -3, 4,
    -- filter=252 channel=31
    4, 0, -5, 1, -1, -2, 4, -2, 7,
    -- filter=252 channel=32
    0, 6, 14, -2, -13, 6, -12, -11, 2,
    -- filter=252 channel=33
    3, 10, 10, -6, -6, 6, -2, -5, 17,
    -- filter=252 channel=34
    4, -1, 5, -8, -2, 24, -10, 4, 23,
    -- filter=252 channel=35
    2, 5, 4, 3, -2, 4, 0, -5, 3,
    -- filter=252 channel=36
    -9, -10, 1, -1, 5, 7, 7, -3, -6,
    -- filter=252 channel=37
    -5, 0, 2, -11, -3, 15, -4, -3, 16,
    -- filter=252 channel=38
    -3, -1, 5, -5, 0, 6, 2, -9, 6,
    -- filter=252 channel=39
    3, -5, 3, 7, 0, -2, -2, -5, -4,
    -- filter=252 channel=40
    8, -4, 1, -7, -1, 0, 5, -8, -7,
    -- filter=252 channel=41
    -10, 10, 2, -13, 1, 1, -4, 2, -5,
    -- filter=252 channel=42
    2, 4, -8, 7, 0, -2, 0, -5, 1,
    -- filter=252 channel=43
    6, -2, -2, -2, -4, 0, -4, -2, -2,
    -- filter=252 channel=44
    -7, -9, -5, -3, -3, 14, -5, 1, 13,
    -- filter=252 channel=45
    1, 2, 2, -4, 5, -1, -3, -6, 1,
    -- filter=252 channel=46
    -1, -5, -5, -3, -4, 3, 4, 3, 1,
    -- filter=252 channel=47
    -5, 0, 1, -1, 6, 3, 1, -1, 12,
    -- filter=252 channel=48
    -5, -2, -4, -8, 0, 2, -5, -1, 7,
    -- filter=252 channel=49
    5, 0, 3, -7, -6, 1, -4, -7, 4,
    -- filter=252 channel=50
    4, 4, 0, 0, -1, 1, 0, -10, 1,
    -- filter=252 channel=51
    -4, 4, 0, 7, -3, -1, -7, 2, 0,
    -- filter=252 channel=52
    3, 2, 0, -5, -9, 6, -3, -3, 0,
    -- filter=252 channel=53
    -4, 0, 1, -2, 0, 3, 0, -10, 0,
    -- filter=252 channel=54
    1, 3, -7, -2, -6, -4, 7, 5, 2,
    -- filter=252 channel=55
    0, 0, 12, 2, -6, 0, -2, -19, 2,
    -- filter=252 channel=56
    0, 0, 2, -4, -1, 5, -10, 1, -1,
    -- filter=252 channel=57
    2, 1, -6, -6, -3, 7, 4, -1, -4,
    -- filter=252 channel=58
    4, -4, -2, -10, 0, -3, -10, -6, 6,
    -- filter=252 channel=59
    -6, 8, -2, -8, -3, 5, 1, -2, 0,
    -- filter=252 channel=60
    5, -7, -3, 3, -7, -2, 1, 6, 3,
    -- filter=252 channel=61
    -6, 0, -4, -8, 2, 1, 1, 4, -3,
    -- filter=252 channel=62
    6, 8, 2, -7, -4, 1, 0, 0, 2,
    -- filter=252 channel=63
    1, -7, -3, -1, -2, 2, -5, 6, -3,
    -- filter=252 channel=64
    1, -2, 2, 7, 6, -2, -3, -2, 0,
    -- filter=252 channel=65
    -4, 5, 2, -3, 2, 0, 3, -3, -1,
    -- filter=252 channel=66
    -10, 8, 7, -9, -3, 12, 3, -3, 13,
    -- filter=252 channel=67
    -2, -7, -4, -9, -8, -2, -8, 1, -1,
    -- filter=252 channel=68
    -6, 3, -10, -4, 0, 3, 6, -5, 1,
    -- filter=252 channel=69
    0, 5, 0, -8, 1, -4, 0, 1, 7,
    -- filter=252 channel=70
    4, -1, 7, -7, -3, 12, -14, -9, 14,
    -- filter=252 channel=71
    4, 3, 0, -4, 6, 0, 4, 0, -6,
    -- filter=252 channel=72
    0, -8, 0, -3, -6, -2, 8, -5, -3,
    -- filter=252 channel=73
    3, 4, 4, -1, -14, 5, -11, -15, 0,
    -- filter=252 channel=74
    -5, -9, -1, -3, -10, 24, -18, -5, 16,
    -- filter=252 channel=75
    1, 12, 1, -4, 4, 7, -15, 1, 4,
    -- filter=252 channel=76
    7, 1, 3, 0, -1, -13, 3, -17, 0,
    -- filter=252 channel=77
    -8, -1, -3, 3, 0, 0, 6, 0, -5,
    -- filter=252 channel=78
    0, 6, -3, 0, -2, 4, -1, 9, 6,
    -- filter=252 channel=79
    10, 3, 9, 0, -16, 5, -11, -22, 9,
    -- filter=252 channel=80
    3, 3, -4, 4, 2, 0, 1, -1, 9,
    -- filter=252 channel=81
    -4, 0, 0, 4, -4, -6, 0, -3, 4,
    -- filter=252 channel=82
    8, 3, -5, 5, 3, -2, 3, -5, 2,
    -- filter=252 channel=83
    2, -2, -1, -3, -6, -1, 4, 4, 0,
    -- filter=252 channel=84
    4, 3, 8, -8, -4, 1, 0, -11, 6,
    -- filter=252 channel=85
    -3, 5, -5, 2, 3, 5, 0, 5, 2,
    -- filter=252 channel=86
    -7, 6, 11, -4, -1, 5, -10, -4, 17,
    -- filter=252 channel=87
    4, 7, 0, -9, -10, 0, -8, 2, -2,
    -- filter=252 channel=88
    -12, -10, -7, -1, 5, -2, 7, 9, 0,
    -- filter=252 channel=89
    -3, 8, 5, -1, -12, -10, 5, -6, -2,
    -- filter=252 channel=90
    -2, -6, 1, -7, 0, 5, -6, 12, 0,
    -- filter=252 channel=91
    -2, 3, -3, -1, -12, 9, -9, -13, 10,
    -- filter=252 channel=92
    -1, -4, -1, -1, 1, -1, 2, 8, 10,
    -- filter=252 channel=93
    -13, -8, 0, -1, 1, 10, -1, 4, 10,
    -- filter=252 channel=94
    -2, -1, -1, 0, -1, -4, 0, 0, 6,
    -- filter=252 channel=95
    -6, 1, -4, 3, -3, 0, -3, 0, 3,
    -- filter=252 channel=96
    -6, 5, 5, -2, 0, 0, 6, 4, -1,
    -- filter=252 channel=97
    6, 5, 7, 2, 10, 5, 5, -4, 2,
    -- filter=252 channel=98
    1, 0, -5, 3, 2, 4, -8, -4, 13,
    -- filter=252 channel=99
    2, -4, -1, -3, -2, 9, -12, -3, 11,
    -- filter=252 channel=100
    -3, -4, 12, -2, 4, 6, 1, 1, -1,
    -- filter=252 channel=101
    2, -10, -7, 0, -2, 6, -5, -7, -1,
    -- filter=252 channel=102
    -3, 6, 0, 0, 1, 4, -1, -5, -3,
    -- filter=252 channel=103
    3, 2, -4, 2, 11, -1, 4, 2, -2,
    -- filter=252 channel=104
    3, -7, -6, 6, 5, 6, -3, 1, 4,
    -- filter=252 channel=105
    9, 6, 4, -6, -3, 4, -3, -14, -1,
    -- filter=252 channel=106
    -6, 1, -2, 6, -2, -1, 9, -9, -1,
    -- filter=252 channel=107
    10, 3, 12, -4, -6, 0, -5, -6, 4,
    -- filter=252 channel=108
    -4, 1, 2, -3, 5, 3, -7, -5, -6,
    -- filter=252 channel=109
    -6, -4, 1, -4, -10, 8, -4, -12, 19,
    -- filter=252 channel=110
    2, 0, 4, 1, 3, -6, 4, -2, 0,
    -- filter=252 channel=111
    4, -2, 4, -5, 6, -4, -3, -5, -4,
    -- filter=252 channel=112
    -5, -1, 3, -11, -6, 17, -11, 2, 15,
    -- filter=252 channel=113
    -1, 2, 10, 2, 0, 8, -8, -6, 10,
    -- filter=252 channel=114
    0, -1, 12, -14, -18, 3, -22, -26, 8,
    -- filter=252 channel=115
    -1, -7, -1, 5, 4, 3, 0, 6, -4,
    -- filter=252 channel=116
    -10, 1, -5, 0, -2, -3, -7, -12, 4,
    -- filter=252 channel=117
    4, 0, -5, -2, 3, -3, 4, 0, 1,
    -- filter=252 channel=118
    1, -1, -4, -4, 2, -1, -5, 1, -5,
    -- filter=252 channel=119
    -1, -5, 17, -7, 4, 19, -4, 9, 7,
    -- filter=252 channel=120
    -8, -6, 3, -10, -5, 17, -8, -13, 23,
    -- filter=252 channel=121
    -1, 7, 6, 4, 5, 2, 0, 5, -5,
    -- filter=252 channel=122
    -13, -8, -7, 4, 9, 6, 4, 19, 12,
    -- filter=252 channel=123
    0, 5, -1, -1, 3, 2, -10, 1, 11,
    -- filter=252 channel=124
    4, -2, -1, -4, -3, -5, -1, -11, 1,
    -- filter=252 channel=125
    -6, -6, 2, 3, -6, 3, -4, -7, 13,
    -- filter=252 channel=126
    -2, -2, 6, -3, -3, -7, 0, -9, 3,
    -- filter=252 channel=127
    0, 6, -1, 1, -5, -5, 2, -3, 1,
    -- filter=253 channel=0
    -8, -7, 12, -2, -10, 4, 1, -7, 7,
    -- filter=253 channel=1
    4, -5, 0, 8, -3, 2, 14, 2, 7,
    -- filter=253 channel=2
    -5, -4, -9, 4, 7, 0, 3, 2, 7,
    -- filter=253 channel=3
    -8, -14, -2, -4, -11, -1, -10, -14, 1,
    -- filter=253 channel=4
    -1, 0, 0, 0, -13, -4, -2, 9, 14,
    -- filter=253 channel=5
    -9, 3, 6, -3, -7, 4, 5, -5, 8,
    -- filter=253 channel=6
    6, 7, 9, 2, -6, 2, 0, 0, 5,
    -- filter=253 channel=7
    4, -7, -1, -5, -4, 3, 4, 2, -2,
    -- filter=253 channel=8
    -3, -10, -9, -2, 0, -8, -4, 0, -3,
    -- filter=253 channel=9
    -5, -5, -2, -2, -3, 9, 6, 10, 0,
    -- filter=253 channel=10
    -8, -6, -17, -3, -6, -12, 5, -3, 0,
    -- filter=253 channel=11
    1, 12, 5, -8, 0, 11, 0, -4, 4,
    -- filter=253 channel=12
    0, -2, -8, 1, -16, -16, -10, -7, -15,
    -- filter=253 channel=13
    -4, -8, -6, 3, -13, -8, 9, -8, -4,
    -- filter=253 channel=14
    1, 0, 7, -1, 0, 6, -4, 0, 1,
    -- filter=253 channel=15
    -4, 7, -1, -5, -12, 0, 12, 1, 2,
    -- filter=253 channel=16
    -10, -1, -1, 1, -5, 3, -5, 0, 7,
    -- filter=253 channel=17
    -2, 1, -4, -3, 3, 5, -5, -3, 0,
    -- filter=253 channel=18
    8, -3, 12, 0, -5, 3, 17, 6, 4,
    -- filter=253 channel=19
    4, 4, 2, 6, 3, -5, -1, -1, 5,
    -- filter=253 channel=20
    12, 17, 10, -1, -10, 4, 1, -7, 3,
    -- filter=253 channel=21
    -3, -9, -10, 11, 13, 2, 9, 16, 16,
    -- filter=253 channel=22
    -8, 4, 6, -7, -10, 2, 4, -8, 2,
    -- filter=253 channel=23
    0, 0, -7, -16, -3, -13, 5, -9, -12,
    -- filter=253 channel=24
    -1, 4, -4, 1, 0, 2, -1, 2, -1,
    -- filter=253 channel=25
    -5, -4, -3, 2, -12, 4, 7, 12, -3,
    -- filter=253 channel=26
    0, -5, 3, 1, 6, -2, 3, 0, 0,
    -- filter=253 channel=27
    -12, 1, -6, 1, -5, 0, 26, 4, 6,
    -- filter=253 channel=28
    4, 4, 4, 6, 4, 2, 0, -3, 0,
    -- filter=253 channel=29
    7, 14, 13, -10, 0, 0, 3, -1, 4,
    -- filter=253 channel=30
    0, -10, 1, 0, 0, 6, 14, 8, 1,
    -- filter=253 channel=31
    -8, -1, -11, 2, 5, 2, 9, 6, 5,
    -- filter=253 channel=32
    -5, 0, -4, 2, -12, -10, 11, 0, 0,
    -- filter=253 channel=33
    -6, -1, -6, 0, -2, -9, 11, -10, -10,
    -- filter=253 channel=34
    -16, -11, -10, -19, -15, -22, -14, -27, -18,
    -- filter=253 channel=35
    4, 7, 4, 6, -7, 5, 7, -1, -7,
    -- filter=253 channel=36
    7, -2, 0, 12, -2, -1, 10, 0, 3,
    -- filter=253 channel=37
    -3, -10, -2, 0, -1, 1, 4, 10, 12,
    -- filter=253 channel=38
    -8, -2, -8, -6, -3, 0, -6, -2, -2,
    -- filter=253 channel=39
    5, 6, 0, -2, 5, 0, 0, 3, 7,
    -- filter=253 channel=40
    -2, 14, 5, -3, 3, 8, -4, 1, 1,
    -- filter=253 channel=41
    -3, -18, -18, 1, -15, -28, 9, -3, -18,
    -- filter=253 channel=42
    -7, 0, 1, 9, -3, 4, 12, 7, -1,
    -- filter=253 channel=43
    0, -8, -8, -10, -9, 0, -1, -7, -11,
    -- filter=253 channel=44
    -18, -11, -11, 0, -3, -1, 8, 2, 12,
    -- filter=253 channel=45
    0, 0, 2, 0, 12, 13, 5, -2, 2,
    -- filter=253 channel=46
    5, -8, 5, 7, -5, 0, 5, -7, -3,
    -- filter=253 channel=47
    -17, -3, 0, -1, 6, -1, 6, 13, 12,
    -- filter=253 channel=48
    -5, -2, -12, 17, 4, -5, 12, 17, 10,
    -- filter=253 channel=49
    12, 0, 3, 5, 7, 4, 21, 10, 5,
    -- filter=253 channel=50
    3, 4, 6, 6, 4, 6, 17, 7, 7,
    -- filter=253 channel=51
    1, 1, 1, -3, -6, 4, 6, -2, -1,
    -- filter=253 channel=52
    5, -3, -7, -3, -17, -13, -2, -8, 0,
    -- filter=253 channel=53
    1, -1, -1, 0, -9, 1, 0, 5, -1,
    -- filter=253 channel=54
    3, 6, -5, 4, 0, -1, 4, -7, -2,
    -- filter=253 channel=55
    1, 7, -5, -8, -11, 0, 5, -3, 0,
    -- filter=253 channel=56
    -9, 0, -12, -11, -11, -2, 0, -11, 0,
    -- filter=253 channel=57
    -7, -5, 2, -6, -7, -3, -4, 6, 0,
    -- filter=253 channel=58
    -3, -9, 5, -3, 0, -1, 0, -7, 3,
    -- filter=253 channel=59
    -10, -8, -15, 12, 6, 2, 19, 10, 11,
    -- filter=253 channel=60
    7, 0, -5, 4, 7, 5, -2, -5, 5,
    -- filter=253 channel=61
    4, -8, -3, -1, -9, -6, 3, 4, -1,
    -- filter=253 channel=62
    0, 0, -1, -4, -5, 3, 2, -2, -7,
    -- filter=253 channel=63
    -1, 4, -3, 4, 3, 1, -4, 2, 5,
    -- filter=253 channel=64
    0, 3, 2, 6, 6, -2, 0, 4, 4,
    -- filter=253 channel=65
    3, -3, 3, -5, 3, -4, 2, -6, 0,
    -- filter=253 channel=66
    1, -6, -12, -7, -17, -10, -5, -5, -14,
    -- filter=253 channel=67
    6, -3, 4, 2, -4, -7, 0, 4, 1,
    -- filter=253 channel=68
    8, 10, -4, 5, 0, 2, 8, 7, 8,
    -- filter=253 channel=69
    -4, 0, -2, -5, -5, 5, -2, -5, -3,
    -- filter=253 channel=70
    5, 0, 0, 2, -5, -3, 5, -4, -1,
    -- filter=253 channel=71
    0, -1, 1, -7, -7, 1, -9, 2, 2,
    -- filter=253 channel=72
    -2, -1, -10, 2, 9, 0, 15, 9, 9,
    -- filter=253 channel=73
    -4, -4, 0, 6, -2, -8, 16, -3, -4,
    -- filter=253 channel=74
    -1, 0, -16, 3, -4, -6, 8, -11, -3,
    -- filter=253 channel=75
    -18, -7, 3, 3, -3, -6, 5, -7, 6,
    -- filter=253 channel=76
    13, 10, 5, -4, -8, 7, 1, 5, -6,
    -- filter=253 channel=77
    5, -4, 1, 7, -5, -6, 0, -5, -3,
    -- filter=253 channel=78
    -4, 6, 1, -3, 0, 1, -1, -1, 1,
    -- filter=253 channel=79
    0, -8, 8, 4, -16, 3, 11, 2, 0,
    -- filter=253 channel=80
    -10, -9, -5, 8, 0, -5, 10, 16, 1,
    -- filter=253 channel=81
    2, 2, 7, 0, 3, 4, -6, 0, -1,
    -- filter=253 channel=82
    -8, -3, -3, -5, -4, 5, 4, -1, -6,
    -- filter=253 channel=83
    -6, -4, -9, 3, 1, 3, 12, 13, 8,
    -- filter=253 channel=84
    9, 6, 9, 0, -7, 1, 5, 1, 6,
    -- filter=253 channel=85
    0, 1, 5, 1, 6, -5, -3, 6, 2,
    -- filter=253 channel=86
    -5, -3, -3, -6, -8, -8, -6, -11, -10,
    -- filter=253 channel=87
    5, 6, 5, -12, -16, -7, -5, -8, 0,
    -- filter=253 channel=88
    10, 5, -3, -1, 11, -7, 9, 11, 0,
    -- filter=253 channel=89
    2, -6, -3, 6, -1, -9, 16, 9, -6,
    -- filter=253 channel=90
    2, -2, -9, 0, -8, -1, -9, 4, -7,
    -- filter=253 channel=91
    -2, 1, 0, 0, -1, 0, 25, 13, 5,
    -- filter=253 channel=92
    -6, -3, -9, -12, -3, 0, -8, -3, -4,
    -- filter=253 channel=93
    -6, -17, -12, 9, 3, 5, 2, 9, 7,
    -- filter=253 channel=94
    -3, 6, 2, 1, -1, -3, 7, -1, -6,
    -- filter=253 channel=95
    0, -10, 2, 3, 3, 2, -7, 2, 4,
    -- filter=253 channel=96
    4, 5, 3, 5, 5, 4, 0, -1, -2,
    -- filter=253 channel=97
    0, -4, -7, 1, -4, 2, -4, -11, -5,
    -- filter=253 channel=98
    -6, -2, -13, -6, -11, -4, 12, -2, 0,
    -- filter=253 channel=99
    -9, -6, -1, -1, 7, -5, -2, -4, -5,
    -- filter=253 channel=100
    -4, -12, 0, -3, -6, -8, -6, -11, -5,
    -- filter=253 channel=101
    -3, -2, 3, 0, 3, 0, 0, 3, 9,
    -- filter=253 channel=102
    -2, 5, -1, 5, 6, -2, 0, -5, -5,
    -- filter=253 channel=103
    -9, -12, -3, 0, 9, 5, 9, 14, 1,
    -- filter=253 channel=104
    -11, -5, -5, 12, 4, 8, 17, 17, 7,
    -- filter=253 channel=105
    -2, 8, 12, -6, 1, 5, 1, -2, 1,
    -- filter=253 channel=106
    6, 12, 6, 3, 0, -1, -1, -2, 1,
    -- filter=253 channel=107
    2, 11, 10, -9, 1, 5, 5, -13, 0,
    -- filter=253 channel=108
    5, -8, 0, 2, -4, 0, -8, -7, -7,
    -- filter=253 channel=109
    0, -8, -6, 1, -10, -10, 24, 6, 12,
    -- filter=253 channel=110
    -8, 2, -2, -12, -3, -12, -3, -6, 0,
    -- filter=253 channel=111
    4, 2, 6, -6, 3, 3, -2, 5, 1,
    -- filter=253 channel=112
    -5, 3, -8, -6, -8, -5, 7, -2, 1,
    -- filter=253 channel=113
    0, -10, -12, -12, -3, -9, 0, -2, 0,
    -- filter=253 channel=114
    9, 9, 19, -2, -18, 3, 24, -6, 1,
    -- filter=253 channel=115
    5, -2, -4, 4, 1, 1, -4, -3, 6,
    -- filter=253 channel=116
    0, 0, -4, 11, 4, 3, 20, 18, 1,
    -- filter=253 channel=117
    7, 1, 2, 8, 6, 1, 3, 5, 7,
    -- filter=253 channel=118
    4, -4, 3, -2, -6, 4, 0, -1, 0,
    -- filter=253 channel=119
    -3, -14, -18, -5, -19, -15, -1, -8, -3,
    -- filter=253 channel=120
    0, 7, -3, 8, -8, 3, 11, 3, 6,
    -- filter=253 channel=121
    -9, -6, -1, -5, -10, -6, -3, 0, -3,
    -- filter=253 channel=122
    -13, -13, -10, 2, 16, 5, -2, 22, 12,
    -- filter=253 channel=123
    2, 0, -11, -2, -5, -9, -2, -9, -9,
    -- filter=253 channel=124
    -2, 10, 7, -6, -8, -8, -1, -3, -9,
    -- filter=253 channel=125
    1, -7, -6, 5, -1, 0, 13, 12, 10,
    -- filter=253 channel=126
    -1, -11, -6, -8, -5, -10, -3, -4, -5,
    -- filter=253 channel=127
    -3, -8, -4, 3, 1, 1, -4, 0, -5,
    -- filter=254 channel=0
    4, 0, 2, -1, -5, 0, -5, -7, -3,
    -- filter=254 channel=1
    -3, -1, -6, 0, 2, 4, 1, -1, 0,
    -- filter=254 channel=2
    5, -6, -6, 5, -2, 0, -3, 1, -2,
    -- filter=254 channel=3
    7, 8, 2, -6, 0, 2, -4, 1, 2,
    -- filter=254 channel=4
    1, 6, 1, -4, -1, -7, 5, 5, 6,
    -- filter=254 channel=5
    -1, 2, 0, -7, -1, 4, -5, 6, 4,
    -- filter=254 channel=6
    6, 5, -4, 5, 7, 1, -3, -6, 7,
    -- filter=254 channel=7
    -2, 3, -6, 6, 1, 4, 5, -3, -3,
    -- filter=254 channel=8
    1, 2, -1, 0, -5, -3, -5, 0, 7,
    -- filter=254 channel=9
    -7, -6, 4, 1, 0, 2, -6, 5, -5,
    -- filter=254 channel=10
    -4, 0, -2, 1, 4, -6, 5, -1, 2,
    -- filter=254 channel=11
    -6, 5, 4, 0, -3, 3, 0, 3, -5,
    -- filter=254 channel=12
    4, -3, 1, -4, -5, -1, 0, 0, -3,
    -- filter=254 channel=13
    -3, 2, -3, 5, -3, 4, 0, 1, -1,
    -- filter=254 channel=14
    -2, -6, 1, -2, 0, -2, 6, -6, 7,
    -- filter=254 channel=15
    0, -4, 6, 1, 0, 0, -4, 2, 3,
    -- filter=254 channel=16
    -1, 7, -6, 0, 0, -1, 7, -5, -5,
    -- filter=254 channel=17
    -1, 1, 4, -4, 0, -5, 6, 5, 6,
    -- filter=254 channel=18
    -4, 3, -6, -1, 1, 0, 4, -4, -4,
    -- filter=254 channel=19
    -5, 0, 2, -1, 2, -5, -1, 0, 3,
    -- filter=254 channel=20
    4, 0, -5, 0, 1, -3, -2, 3, -2,
    -- filter=254 channel=21
    -1, -7, 0, -7, -7, -2, -7, -8, 1,
    -- filter=254 channel=22
    0, 1, -4, 2, 2, 5, -4, -7, -4,
    -- filter=254 channel=23
    1, 0, -3, 0, 0, -5, 5, 7, 6,
    -- filter=254 channel=24
    0, -3, -3, 7, 0, 0, 2, 4, 6,
    -- filter=254 channel=25
    -2, 0, -6, -4, -9, 4, 4, -8, 4,
    -- filter=254 channel=26
    6, 0, 2, -3, 6, 6, -1, 0, -3,
    -- filter=254 channel=27
    0, -2, -6, -10, -2, 5, -6, -5, -1,
    -- filter=254 channel=28
    0, -1, -6, -3, -7, 0, 1, 2, 3,
    -- filter=254 channel=29
    7, -1, -8, 0, 1, -5, 1, -5, -5,
    -- filter=254 channel=30
    -3, 5, 0, -1, -1, 7, 1, 7, 2,
    -- filter=254 channel=31
    0, -1, -1, -6, 0, -5, -2, -7, 3,
    -- filter=254 channel=32
    5, 6, -3, 3, -8, 4, 4, -4, 5,
    -- filter=254 channel=33
    0, 2, 0, 2, -1, 3, 0, 5, 5,
    -- filter=254 channel=34
    6, -1, 6, 0, -5, -3, 0, -6, 4,
    -- filter=254 channel=35
    5, -5, 4, 5, -2, 5, -6, -2, -4,
    -- filter=254 channel=36
    -6, 2, -5, -3, 3, 2, -5, 0, 1,
    -- filter=254 channel=37
    3, -4, 8, -7, -5, 8, 2, 0, 1,
    -- filter=254 channel=38
    5, 0, -3, -6, 2, 4, 0, 5, 4,
    -- filter=254 channel=39
    -2, 5, 6, -5, -6, -3, 8, -4, 7,
    -- filter=254 channel=40
    3, 7, 1, -5, 5, -5, 3, -4, -1,
    -- filter=254 channel=41
    12, -8, -6, 6, -1, -2, 11, 1, 2,
    -- filter=254 channel=42
    7, 4, 1, 0, 1, 1, 3, 1, 4,
    -- filter=254 channel=43
    5, -1, 4, 6, 2, 3, -2, -1, -1,
    -- filter=254 channel=44
    -2, 1, -3, 5, 1, -4, -5, -7, -6,
    -- filter=254 channel=45
    -5, -4, 0, 4, 6, 7, 3, 0, 5,
    -- filter=254 channel=46
    -5, -5, -6, -1, 2, 0, -2, 3, 5,
    -- filter=254 channel=47
    3, 4, 4, -6, -2, -1, 5, 5, 0,
    -- filter=254 channel=48
    -6, -4, -5, 1, -2, 5, -1, 2, -3,
    -- filter=254 channel=49
    -1, -7, -1, -1, 0, 2, 4, 2, -1,
    -- filter=254 channel=50
    -5, -2, 0, -8, 5, 2, -1, -2, 5,
    -- filter=254 channel=51
    4, -7, -2, 0, 7, -3, -1, 4, 3,
    -- filter=254 channel=52
    -4, -4, 5, -5, -6, -6, 0, 2, 4,
    -- filter=254 channel=53
    0, -5, 0, 6, -1, 6, 6, 7, 0,
    -- filter=254 channel=54
    -3, 3, 3, -7, 0, -7, 4, -2, 5,
    -- filter=254 channel=55
    -1, -4, -1, 4, -8, -1, 9, 5, 7,
    -- filter=254 channel=56
    -3, 2, -2, 0, 3, 0, 6, -2, -2,
    -- filter=254 channel=57
    3, 0, -1, -5, -3, 2, -3, 5, -6,
    -- filter=254 channel=58
    -3, 1, 3, 4, -3, -5, -3, 1, 0,
    -- filter=254 channel=59
    4, -4, 5, -4, 4, 3, -6, 3, 2,
    -- filter=254 channel=60
    -1, -6, -6, -1, 2, 1, 6, 0, 4,
    -- filter=254 channel=61
    -5, -7, -6, 2, -1, 2, 6, -2, 3,
    -- filter=254 channel=62
    -2, -5, 1, 0, 1, -6, -4, -1, -6,
    -- filter=254 channel=63
    2, -3, -5, 1, 6, 1, 7, -1, 6,
    -- filter=254 channel=64
    3, -5, 5, 3, 5, -4, -5, -6, -3,
    -- filter=254 channel=65
    -1, -1, 1, 5, 4, -3, -2, -1, 4,
    -- filter=254 channel=66
    8, -7, -6, 7, 1, 4, -4, 1, 4,
    -- filter=254 channel=67
    -4, -2, 5, 4, 3, 5, 1, 1, -3,
    -- filter=254 channel=68
    1, 0, 3, 4, 1, 1, 6, 7, 2,
    -- filter=254 channel=69
    7, -6, 3, 7, 1, -1, -5, 5, 0,
    -- filter=254 channel=70
    -3, -7, 3, 0, 0, -6, -6, -1, -5,
    -- filter=254 channel=71
    3, 1, -2, 6, 0, 2, 2, 3, -2,
    -- filter=254 channel=72
    7, 4, 1, -1, 0, 0, 0, -1, -4,
    -- filter=254 channel=73
    -3, 6, 3, 0, -5, -6, 7, 2, -1,
    -- filter=254 channel=74
    -3, 4, 1, 5, -2, -5, -7, -6, -7,
    -- filter=254 channel=75
    1, 0, 3, 3, 6, -1, 1, -6, 4,
    -- filter=254 channel=76
    4, -2, -7, 5, 0, -6, 1, 0, 2,
    -- filter=254 channel=77
    -3, -2, -2, 2, -2, -2, -1, 4, -2,
    -- filter=254 channel=78
    -2, -5, 6, 2, 3, 0, 6, 5, 0,
    -- filter=254 channel=79
    7, 3, -4, 2, 1, -1, 1, 0, -6,
    -- filter=254 channel=80
    -3, 3, -6, -6, 0, 1, -6, 4, -2,
    -- filter=254 channel=81
    0, 2, 5, 1, 1, -3, -3, -3, 5,
    -- filter=254 channel=82
    -7, 2, 2, -2, 3, 0, -2, 0, -5,
    -- filter=254 channel=83
    0, 0, 6, -6, -6, -7, -4, 7, 4,
    -- filter=254 channel=84
    1, -8, 6, 1, -4, 0, 3, 4, -2,
    -- filter=254 channel=85
    -2, 0, -3, 2, 3, 7, 5, -4, -7,
    -- filter=254 channel=86
    -4, 0, 2, -4, -5, 6, 1, -6, 3,
    -- filter=254 channel=87
    -2, 2, -7, 1, -1, -3, 1, -3, 3,
    -- filter=254 channel=88
    -7, 0, 2, -5, -3, 0, 0, -6, -1,
    -- filter=254 channel=89
    0, 4, 2, 2, -5, -8, 2, -4, -3,
    -- filter=254 channel=90
    -4, 0, 0, 0, 0, 1, -4, 0, 0,
    -- filter=254 channel=91
    2, 0, 2, 5, -8, -4, 4, -4, -7,
    -- filter=254 channel=92
    1, -1, -5, -1, -3, -5, 1, 0, -6,
    -- filter=254 channel=93
    -1, 3, 1, -4, 0, 7, -7, -3, -6,
    -- filter=254 channel=94
    1, -4, 0, 5, 6, 2, 5, -6, 4,
    -- filter=254 channel=95
    0, 5, 0, 5, 1, 0, 0, -5, 5,
    -- filter=254 channel=96
    -6, 3, 3, 0, 0, 0, -4, 6, 4,
    -- filter=254 channel=97
    -5, -5, 0, 4, 4, -6, 4, -5, 1,
    -- filter=254 channel=98
    5, -3, 0, 0, -8, 0, 3, 3, -2,
    -- filter=254 channel=99
    -7, 5, -4, -6, -6, 4, -6, 1, 3,
    -- filter=254 channel=100
    0, 4, 0, -1, 1, -4, 0, 1, 6,
    -- filter=254 channel=101
    4, 3, 2, -3, 6, 0, 7, 5, -4,
    -- filter=254 channel=102
    2, -6, 2, 7, -7, 5, -2, 2, -2,
    -- filter=254 channel=103
    4, 0, -3, -2, 3, -3, -3, -7, 1,
    -- filter=254 channel=104
    6, -4, -2, -2, -1, -6, 4, 5, -7,
    -- filter=254 channel=105
    -5, 6, 3, -1, -7, -4, 0, 3, -1,
    -- filter=254 channel=106
    6, -4, 2, 4, -7, -2, 2, 1, -4,
    -- filter=254 channel=107
    4, 6, -2, -3, 5, 0, 4, -3, -5,
    -- filter=254 channel=108
    -5, -5, -5, 5, 5, -4, 6, -1, 6,
    -- filter=254 channel=109
    4, 1, -7, 4, -1, 5, 2, 1, -7,
    -- filter=254 channel=110
    4, -6, -6, -2, 0, -1, -3, -4, -5,
    -- filter=254 channel=111
    2, -3, 6, 1, -7, -1, 4, -1, -5,
    -- filter=254 channel=112
    1, -3, -2, 2, 3, 7, 3, -4, 2,
    -- filter=254 channel=113
    1, -4, 3, 5, 2, 0, 2, -6, 5,
    -- filter=254 channel=114
    -4, 5, -6, 0, -8, 5, -5, 0, -7,
    -- filter=254 channel=115
    -1, 5, -7, 6, 4, 4, 3, 7, 0,
    -- filter=254 channel=116
    5, 0, -7, 6, -3, -2, -4, 3, 4,
    -- filter=254 channel=117
    6, -4, 6, -4, 5, 0, 1, 7, 1,
    -- filter=254 channel=118
    6, -5, 5, 1, 3, -1, -1, -3, -4,
    -- filter=254 channel=119
    1, 0, 1, -1, 4, 2, -4, -3, -7,
    -- filter=254 channel=120
    5, 2, -5, -5, 5, -2, 0, 4, -1,
    -- filter=254 channel=121
    -5, 0, -3, 6, -4, 6, 4, 0, 6,
    -- filter=254 channel=122
    -6, -6, 0, -5, 0, 0, 6, -1, 0,
    -- filter=254 channel=123
    4, 2, 4, 0, 6, -3, 0, 6, -2,
    -- filter=254 channel=124
    -1, -2, 2, 6, -5, 0, 0, 3, 0,
    -- filter=254 channel=125
    -1, 3, -7, 0, 0, 7, 2, -2, 1,
    -- filter=254 channel=126
    9, -1, -1, 6, -8, 0, -5, 0, 3,
    -- filter=254 channel=127
    4, 0, 3, 8, 3, -2, -3, -2, 5,
    -- filter=255 channel=0
    -1, 2, 7, -4, 5, 1, 0, 1, -2,
    -- filter=255 channel=1
    2, 0, -3, 5, -2, 6, 2, 0, 3,
    -- filter=255 channel=2
    0, 1, 6, 6, -3, 4, -6, 1, 1,
    -- filter=255 channel=3
    0, 8, 3, -1, -6, 5, -7, 5, 3,
    -- filter=255 channel=4
    -3, -6, -7, 6, 5, 0, 0, 9, 0,
    -- filter=255 channel=5
    -7, 2, -1, -2, 7, 11, 0, -6, 0,
    -- filter=255 channel=6
    0, 0, -6, -3, 0, 0, 6, 0, 0,
    -- filter=255 channel=7
    7, 4, -2, -3, 7, 7, 0, -2, 0,
    -- filter=255 channel=8
    -3, -5, -2, -6, 1, 6, -4, 2, -3,
    -- filter=255 channel=9
    -5, -3, -7, -1, 3, -3, -3, 0, 5,
    -- filter=255 channel=10
    0, -4, -8, 5, 1, -1, -5, 5, 5,
    -- filter=255 channel=11
    6, 7, 4, 0, -1, -1, 8, 3, 0,
    -- filter=255 channel=12
    3, 6, -2, 5, 0, -3, -2, -2, -1,
    -- filter=255 channel=13
    0, 2, -2, 5, -5, 1, 8, -4, 1,
    -- filter=255 channel=14
    6, 0, -6, 4, 1, -6, 1, -1, -2,
    -- filter=255 channel=15
    2, 7, -9, -1, 6, -3, -4, 4, -6,
    -- filter=255 channel=16
    6, -2, 3, 1, -3, 6, -2, 5, 3,
    -- filter=255 channel=17
    3, 1, -2, -3, 6, -2, -7, 3, -3,
    -- filter=255 channel=18
    0, 0, -5, 3, 4, -8, 3, -2, 2,
    -- filter=255 channel=19
    -5, 7, -5, -6, 5, 0, 5, 2, -2,
    -- filter=255 channel=20
    8, -1, -3, 7, -6, 0, 4, 6, -3,
    -- filter=255 channel=21
    3, 3, -1, -9, -1, -5, 5, 3, 7,
    -- filter=255 channel=22
    0, 5, 5, -5, -2, 0, 0, 0, -3,
    -- filter=255 channel=23
    -2, 0, -10, 5, 0, -3, -6, -5, 3,
    -- filter=255 channel=24
    4, -1, 4, 0, 0, 2, 2, -2, -6,
    -- filter=255 channel=25
    0, 3, -2, -6, 4, 0, 1, -3, 2,
    -- filter=255 channel=26
    0, 1, 0, 5, 0, 4, -2, 5, 2,
    -- filter=255 channel=27
    -6, 1, -1, -6, -1, -7, -5, 3, -7,
    -- filter=255 channel=28
    -4, -1, 1, 6, -3, -6, -5, -2, 7,
    -- filter=255 channel=29
    1, -3, -4, 5, -3, -7, -2, 8, 0,
    -- filter=255 channel=30
    3, 0, -5, -9, 4, 4, 3, -4, 0,
    -- filter=255 channel=31
    -4, -3, -2, -4, -11, 1, -4, -8, -8,
    -- filter=255 channel=32
    1, 7, 0, -8, -2, -7, -5, -2, 0,
    -- filter=255 channel=33
    -5, 1, -4, -7, 4, -3, -5, 1, -5,
    -- filter=255 channel=34
    -3, 2, -7, -2, 1, 0, -5, 3, -9,
    -- filter=255 channel=35
    2, 5, 0, 2, -7, -4, 3, -5, 0,
    -- filter=255 channel=36
    -4, 3, -1, 1, 1, 4, 2, 3, 4,
    -- filter=255 channel=37
    -1, -5, 5, -2, 5, 14, 2, -5, 9,
    -- filter=255 channel=38
    1, 0, -3, -4, 2, 3, 3, 7, 5,
    -- filter=255 channel=39
    -1, 2, 4, 4, -3, 1, -4, 5, 0,
    -- filter=255 channel=40
    0, -4, -5, -6, 1, 0, 7, 0, 0,
    -- filter=255 channel=41
    1, 0, 1, 2, -8, -8, 8, -3, -5,
    -- filter=255 channel=42
    -2, -6, -3, 1, 5, 7, -7, 2, 2,
    -- filter=255 channel=43
    -2, 0, 0, -4, 0, 4, -5, 1, -7,
    -- filter=255 channel=44
    2, -2, 7, -7, 2, 0, -9, -6, 4,
    -- filter=255 channel=45
    -2, 0, -1, -2, 0, 5, 5, -4, 4,
    -- filter=255 channel=46
    -4, -3, 3, 0, 5, 1, 2, 2, 4,
    -- filter=255 channel=47
    5, 3, 3, -5, -1, 2, 1, -4, 1,
    -- filter=255 channel=48
    3, -7, 0, 2, -1, 2, -7, 1, -5,
    -- filter=255 channel=49
    2, 3, 0, 1, 2, -2, 7, 0, -4,
    -- filter=255 channel=50
    1, 6, -6, -7, 0, -7, 1, 3, 1,
    -- filter=255 channel=51
    4, 5, 7, 0, -1, -5, -4, 2, -7,
    -- filter=255 channel=52
    -2, 6, -6, -1, 6, -4, 5, -3, 0,
    -- filter=255 channel=53
    1, 5, 0, 1, 3, 0, 5, 0, -6,
    -- filter=255 channel=54
    3, 3, -5, 6, 4, -4, 5, 0, 3,
    -- filter=255 channel=55
    0, -4, -2, 9, -8, -7, 9, 0, -6,
    -- filter=255 channel=56
    -3, -2, -2, 4, -3, -8, 6, -4, 2,
    -- filter=255 channel=57
    3, 1, -3, 6, 0, 1, 7, 2, 0,
    -- filter=255 channel=58
    5, 3, 10, -3, 8, 10, 2, 3, 8,
    -- filter=255 channel=59
    1, -7, -6, -6, -7, 0, 5, 4, -1,
    -- filter=255 channel=60
    4, 5, 1, 1, 3, -1, -1, -6, 5,
    -- filter=255 channel=61
    1, 5, -5, 7, -6, 4, 1, -6, 1,
    -- filter=255 channel=62
    1, 6, 5, 7, 2, 2, -3, -5, -4,
    -- filter=255 channel=63
    -4, -1, -2, -1, -5, -1, -3, -5, -2,
    -- filter=255 channel=64
    5, -6, -3, 1, -3, -6, 0, -5, 1,
    -- filter=255 channel=65
    -3, 0, -1, 6, -1, 0, 0, 1, 7,
    -- filter=255 channel=66
    -6, 3, -3, 5, 1, -4, 4, -7, -4,
    -- filter=255 channel=67
    3, -5, -2, 4, -3, 0, 7, 2, -2,
    -- filter=255 channel=68
    6, -7, 1, 4, 4, 3, -3, 0, 2,
    -- filter=255 channel=69
    5, -2, -1, -5, 6, -4, -1, -5, 4,
    -- filter=255 channel=70
    -2, -3, -4, 0, -4, -8, 3, 4, -5,
    -- filter=255 channel=71
    -3, 6, 3, -6, 2, -1, -2, 4, 3,
    -- filter=255 channel=72
    2, 5, -1, -7, -6, -7, 5, -4, -6,
    -- filter=255 channel=73
    0, 1, -3, 1, 0, 5, 0, 8, 2,
    -- filter=255 channel=74
    -4, -9, -5, 2, 4, 0, -7, -6, -7,
    -- filter=255 channel=75
    0, 9, -1, -1, 5, 6, 0, -1, 9,
    -- filter=255 channel=76
    8, -1, 1, -4, -1, -9, 3, 0, 4,
    -- filter=255 channel=77
    5, 0, 3, 4, 6, 4, -6, -2, 6,
    -- filter=255 channel=78
    5, 1, 3, -2, -3, 0, 2, -7, 2,
    -- filter=255 channel=79
    -3, 7, 1, 6, 5, -11, -5, -2, -3,
    -- filter=255 channel=80
    7, -5, 1, 3, -8, -8, -1, -5, 3,
    -- filter=255 channel=81
    1, -1, 7, 0, -1, 0, 3, 2, -2,
    -- filter=255 channel=82
    -4, 1, 0, 0, -1, 1, 1, -4, -6,
    -- filter=255 channel=83
    -5, 0, 2, 5, 1, -5, 3, 5, 5,
    -- filter=255 channel=84
    1, -5, -2, -4, -5, 4, 3, -1, -3,
    -- filter=255 channel=85
    1, 1, -3, 5, -5, -5, -3, 5, -4,
    -- filter=255 channel=86
    -4, 3, 0, 0, 1, -4, 0, 3, 0,
    -- filter=255 channel=87
    7, -1, 2, -2, 0, -3, 1, 4, -7,
    -- filter=255 channel=88
    4, -8, -4, 6, -6, -4, 0, -6, 2,
    -- filter=255 channel=89
    11, 5, -2, -2, 0, -9, 8, -1, -8,
    -- filter=255 channel=90
    0, 3, -6, -6, 0, 4, 7, 4, -2,
    -- filter=255 channel=91
    0, -8, -10, 1, 0, -1, -1, -5, 2,
    -- filter=255 channel=92
    -6, 5, 4, -3, -5, -8, -2, 5, -5,
    -- filter=255 channel=93
    2, 4, -6, 4, -1, 12, 0, 2, 2,
    -- filter=255 channel=94
    5, 0, -4, -3, 6, 6, -6, 1, -1,
    -- filter=255 channel=95
    2, -5, -3, 0, 6, -6, 5, 0, 0,
    -- filter=255 channel=96
    3, -3, 0, 0, 3, -2, 0, -5, 0,
    -- filter=255 channel=97
    6, 0, 7, 6, 7, 0, 4, 7, 3,
    -- filter=255 channel=98
    -6, 1, 0, 0, -4, 0, -7, 6, -3,
    -- filter=255 channel=99
    -1, 0, -7, -2, -1, -8, 0, 5, -5,
    -- filter=255 channel=100
    2, -1, 0, 3, -7, -3, 0, -3, -3,
    -- filter=255 channel=101
    1, 0, 4, 0, -3, 5, 0, 5, -4,
    -- filter=255 channel=102
    1, 7, 2, -5, -5, 4, 5, 3, 6,
    -- filter=255 channel=103
    -2, 5, -4, -7, -4, 7, -8, -6, 2,
    -- filter=255 channel=104
    -3, 4, -7, -8, -7, -1, 5, 1, 6,
    -- filter=255 channel=105
    2, 5, -4, 2, 0, 0, 6, -6, -4,
    -- filter=255 channel=106
    4, -5, 3, 0, 0, -5, -2, -7, 6,
    -- filter=255 channel=107
    -2, 5, -5, 7, -3, 0, 1, 1, -4,
    -- filter=255 channel=108
    3, 0, 8, 0, 7, 6, 0, 4, 6,
    -- filter=255 channel=109
    -4, -5, -9, 4, 0, -5, 2, 8, 0,
    -- filter=255 channel=110
    -5, -6, -7, 6, 3, -7, -3, -3, -2,
    -- filter=255 channel=111
    1, -1, 7, 4, -3, -3, 2, 0, 4,
    -- filter=255 channel=112
    -3, -9, 0, -5, 3, 3, 1, -4, 5,
    -- filter=255 channel=113
    0, -7, -7, -4, -8, -5, -3, 4, -6,
    -- filter=255 channel=114
    0, 1, 2, -2, -2, -3, -3, 3, -5,
    -- filter=255 channel=115
    0, 0, -4, 0, 5, -7, 4, 2, 3,
    -- filter=255 channel=116
    -4, -6, -6, 6, 1, 0, 4, 4, -3,
    -- filter=255 channel=117
    0, -2, 2, 4, -8, 1, -4, 1, -2,
    -- filter=255 channel=118
    0, 1, -6, 6, 4, 6, -2, -5, -1,
    -- filter=255 channel=119
    1, -9, 0, -7, -2, -6, -6, -6, -8,
    -- filter=255 channel=120
    4, -6, 0, -4, 0, -3, -1, 0, 0,
    -- filter=255 channel=121
    0, 2, -4, 5, -6, -7, 5, 6, -2,
    -- filter=255 channel=122
    -7, -2, 0, -1, -2, 4, -2, -2, 5,
    -- filter=255 channel=123
    -1, -6, -6, 6, -7, -5, 3, -1, -6,
    -- filter=255 channel=124
    4, 0, -4, 8, 0, 5, 2, 0, 0,
    -- filter=255 channel=125
    7, -2, -2, 5, 0, -1, -5, -3, 1,
    -- filter=255 channel=126
    3, 9, 6, -6, 6, 1, -2, -6, -2,
    -- filter=255 channel=127
    0, -5, 0, 4, 1, 1, 0, 1, -1,

    -- ifmap
    -- channel=0
    861, 879, 868, 823, 508, 353, 561, 
    433, 795, 649, 283, 217, 135, 174, 
    159, 741, 520, 262, 304, 149, 55, 
    51, 369, 450, 165, 292, 153, 124, 
    22, 107, 78, 114, 171, 58, 131, 
    0, 245, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=1
    945, 985, 1021, 837, 527, 380, 603, 
    610, 1003, 805, 421, 284, 336, 237, 
    440, 787, 794, 610, 445, 380, 236, 
    328, 591, 502, 453, 404, 345, 315, 
    257, 414, 289, 304, 213, 37, 190, 
    0, 358, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=2
    0, 12, 0, 0, 0, 0, 0, 
    121, 136, 156, 53, 12, 18, 0, 
    24, 0, 0, 157, 154, 0, 103, 
    129, 50, 0, 0, 0, 0, 40, 
    70, 273, 263, 209, 0, 0, 17, 
    0, 13, 0, 0, 30, 137, 97, 
    0, 0, 25, 121, 142, 112, 134, 
    
    -- channel=3
    175, 24, 73, 642, 35, 0, 302, 
    0, 0, 0, 0, 66, 0, 181, 
    0, 638, 168, 0, 0, 84, 0, 
    0, 0, 720, 431, 308, 351, 11, 
    0, 0, 0, 0, 449, 9, 0, 
    690, 160, 1222, 935, 32, 0, 0, 
    486, 1291, 241, 0, 0, 142, 47, 
    
    -- channel=4
    0, 15, 2, 0, 1, 0, 0, 
    348, 494, 584, 292, 0, 3, 0, 
    0, 0, 18, 603, 418, 0, 389, 
    247, 121, 0, 0, 0, 0, 34, 
    38, 843, 785, 638, 0, 146, 0, 
    0, 0, 0, 0, 138, 312, 124, 
    0, 0, 5, 205, 242, 51, 113, 
    
    -- channel=5
    1372, 1421, 1219, 1124, 543, 453, 976, 
    674, 1179, 606, 70, 86, 0, 328, 
    0, 931, 146, 0, 0, 0, 0, 
    0, 387, 266, 0, 73, 0, 200, 
    0, 0, 0, 0, 0, 0, 262, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=6
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 132, 19, 0, 
    60, 0, 0, 0, 0, 25, 0, 
    134, 127, 33, 35, 0, 103, 0, 
    242, 344, 421, 373, 520, 650, 584, 
    715, 374, 644, 649, 739, 777, 855, 
    
    -- channel=7
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=8
    7, 0, 7, 0, 105, 0, 0, 
    283, 136, 99, 8, 184, 0, 43, 
    71, 147, 81, 0, 464, 0, 26, 
    0, 108, 36, 0, 139, 0, 59, 
    0, 370, 220, 76, 0, 174, 90, 
    49, 252, 0, 0, 81, 98, 24, 
    77, 0, 106, 23, 60, 26, 62, 
    
    -- channel=9
    429, 451, 387, 255, 125, 98, 292, 
    185, 387, 132, 51, 144, 66, 96, 
    253, 242, 260, 23, 46, 64, 77, 
    87, 159, 192, 113, 131, 77, 234, 
    97, 24, 36, 50, 4, 0, 196, 
    171, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 0, 
    
    -- channel=10
    330, 322, 327, 404, 212, 222, 300, 
    148, 201, 111, 137, 183, 204, 207, 
    356, 354, 299, 157, 58, 294, 113, 
    304, 249, 473, 419, 345, 332, 207, 
    410, 97, 43, 165, 355, 119, 214, 
    531, 426, 584, 476, 180, 85, 212, 
    347, 770, 213, 109, 92, 178, 173, 
    
    -- channel=11
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 64, 46, 0, 
    0, 0, 0, 0, 23, 56, 138, 
    141, 0, 0, 0, 0, 98, 9, 
    294, 133, 125, 215, 127, 318, 92, 
    627, 316, 670, 811, 1032, 1202, 1182, 
    1217, 742, 1145, 1197, 1321, 1411, 1495, 
    
    -- channel=12
    0, 0, 267, 98, 96, 14, 0, 
    0, 0, 126, 0, 199, 52, 0, 
    315, 0, 55, 149, 338, 0, 84, 
    461, 53, 497, 54, 374, 0, 74, 
    519, 265, 0, 378, 178, 0, 138, 
    201, 961, 0, 138, 0, 62, 68, 
    0, 787, 32, 0, 59, 22, 174, 
    
    -- channel=13
    42, 19, 235, 239, 129, 93, 60, 
    0, 0, 93, 244, 209, 316, 50, 
    504, 49, 441, 477, 275, 404, 275, 
    605, 233, 508, 495, 383, 453, 186, 
    810, 359, 45, 447, 363, 167, 210, 
    717, 964, 577, 468, 379, 333, 391, 
    293, 1075, 411, 342, 353, 386, 486, 
    
    -- channel=14
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 283, 191, 22, 
    343, 0, 362, 147, 327, 266, 157, 
    490, 23, 296, 328, 264, 278, 133, 
    712, 533, 263, 285, 243, 340, 137, 
    1153, 805, 1123, 1068, 969, 1102, 1139, 
    1321, 1198, 1168, 1163, 1237, 1404, 1447, 
    
    -- channel=16
    871, 875, 835, 767, 418, 313, 672, 
    431, 755, 358, 142, 175, 13, 273, 
    132, 540, 208, 0, 85, 4, 95, 
    0, 360, 313, 110, 205, 69, 264, 
    0, 0, 0, 0, 103, 0, 286, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=17
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=18
    0, 0, 0, 0, 0, 12, 0, 
    0, 0, 0, 194, 121, 398, 17, 
    628, 0, 449, 590, 271, 537, 224, 
    998, 123, 284, 456, 313, 463, 84, 
    1157, 665, 408, 598, 358, 194, 55, 
    1026, 1212, 1292, 1045, 914, 1021, 1075, 
    1217, 1396, 1131, 1150, 1228, 1328, 1499, 
    
    -- channel=19
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 13, 0, 
    0, 0, 0, 0, 48, 58, 39, 
    0, 0, 12, 43, 45, 37, 24, 
    
    -- channel=20
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 161, 53, 0, 
    0, 0, 0, 0, 193, 54, 217, 
    259, 0, 0, 0, 0, 123, 24, 
    478, 324, 30, 212, 195, 541, 181, 
    1173, 669, 1247, 1509, 1771, 2135, 2100, 
    2254, 1525, 2062, 2157, 2365, 2576, 2687, 
    
    -- channel=21
    1204, 1317, 1178, 964, 655, 635, 932, 
    790, 1118, 831, 505, 432, 431, 554, 
    504, 788, 541, 448, 326, 379, 432, 
    214, 626, 542, 495, 496, 362, 634, 
    208, 110, 283, 298, 348, 123, 561, 
    0, 55, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=22
    0, 0, 0, 0, 0, 0, 10, 
    41, 0, 0, 0, 124, 0, 58, 
    109, 107, 101, 0, 196, 0, 0, 
    0, 60, 122, 62, 91, 48, 56, 
    14, 169, 0, 0, 11, 109, 14, 
    353, 180, 282, 240, 176, 164, 142, 
    382, 232, 248, 199, 202, 269, 258, 
    
    -- channel=23
    187, 0, 75, 228, 178, 31, 304, 
    69, 0, 0, 0, 798, 74, 248, 
    521, 889, 600, 0, 757, 178, 0, 
    202, 210, 1195, 454, 910, 364, 444, 
    532, 347, 0, 52, 372, 302, 467, 
    1507, 1264, 1225, 1139, 668, 869, 885, 
    1518, 1424, 1015, 841, 943, 1178, 1138, 
    
    -- channel=24
    134, 133, 111, 57, 18, 8, 64, 
    67, 119, 34, 0, 0, 0, 0, 
    0, 44, 0, 0, 0, 0, 0, 
    0, 26, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=25
    463, 492, 621, 311, 122, 197, 295, 
    323, 423, 358, 201, 257, 300, 33, 
    821, 173, 664, 542, 362, 294, 277, 
    779, 401, 515, 407, 429, 253, 390, 
    903, 485, 159, 578, 188, 0, 396, 
    470, 968, 0, 0, 0, 0, 0, 
    0, 493, 0, 0, 0, 0, 0, 
    
    -- channel=26
    655, 703, 563, 403, 287, 176, 429, 
    336, 650, 288, 60, 14, 0, 159, 
    0, 254, 0, 0, 0, 0, 61, 
    0, 133, 0, 0, 0, 0, 133, 
    0, 0, 0, 0, 0, 0, 149, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=27
    568, 483, 612, 182, 326, 228, 457, 
    555, 595, 348, 115, 823, 239, 189, 
    1100, 702, 1216, 265, 1064, 252, 313, 
    867, 580, 1087, 435, 840, 222, 698, 
    1037, 960, 511, 759, 209, 82, 774, 
    1314, 1520, 236, 269, 281, 477, 493, 
    609, 645, 293, 351, 367, 421, 439, 
    
    -- channel=28
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=29
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 24, 0, 82, 
    389, 0, 0, 0, 0, 0, 0, 
    494, 305, 83, 273, 135, 350, 11, 
    998, 660, 1164, 1348, 1640, 2002, 2017, 
    2038, 1431, 1863, 1985, 2192, 2372, 2529, 
    
    -- channel=30
    622, 617, 664, 414, 286, 209, 422, 
    365, 608, 373, 168, 265, 79, 100, 
    422, 371, 466, 173, 344, 75, 153, 
    255, 312, 373, 71, 226, 52, 294, 
    247, 245, 130, 324, 41, 0, 419, 
    202, 385, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=31
    854, 825, 799, 538, 577, 379, 746, 
    470, 773, 298, 75, 698, 136, 384, 
    500, 693, 629, 0, 464, 20, 302, 
    90, 450, 845, 310, 613, 118, 746, 
    124, 64, 24, 192, 175, 73, 746, 
    536, 240, 0, 0, 0, 0, 0, 
    0, 102, 0, 0, 0, 0, 0, 
    
    -- channel=32
    152, 112, 277, 52, 29, 14, 74, 
    134, 5, 0, 8, 258, 142, 0, 
    696, 51, 509, 245, 424, 193, 163, 
    711, 203, 540, 321, 433, 237, 247, 
    857, 451, 44, 488, 156, 57, 300, 
    937, 1196, 528, 563, 440, 555, 572, 
    633, 1115, 598, 570, 633, 677, 835, 
    
    -- channel=33
    379, 305, 351, 457, 276, 201, 346, 
    81, 195, 73, 0, 397, 182, 136, 
    539, 612, 772, 44, 219, 225, 37, 
    434, 251, 882, 586, 587, 307, 337, 
    669, 199, 0, 153, 372, 70, 243, 
    956, 876, 725, 748, 70, 14, 145, 
    357, 1154, 131, 42, 11, 125, 132, 
    
    -- channel=34
    100, 0, 0, 0, 51, 0, 268, 
    760, 164, 0, 0, 713, 0, 205, 
    431, 593, 0, 0, 1322, 0, 0, 
    0, 178, 493, 0, 724, 0, 136, 
    0, 781, 103, 0, 0, 114, 363, 
    433, 778, 0, 0, 0, 115, 8, 
    617, 0, 231, 0, 9, 112, 52, 
    
    -- channel=35
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=36
    47, 60, 101, 0, 137, 159, 68, 
    202, 100, 167, 242, 186, 175, 195, 
    140, 0, 0, 267, 255, 152, 313, 
    202, 167, 0, 48, 135, 132, 208, 
    177, 271, 219, 319, 135, 225, 301, 
    50, 188, 0, 39, 279, 361, 333, 
    227, 127, 270, 290, 327, 293, 345, 
    
    -- channel=37
    1111, 1177, 1158, 884, 627, 432, 697, 
    613, 1151, 942, 421, 323, 200, 286, 
    146, 967, 682, 401, 408, 134, 174, 
    0, 536, 521, 180, 401, 180, 313, 
    0, 47, 183, 178, 67, 0, 205, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=38
    303, 269, 287, 246, 119, 94, 270, 
    101, 99, 0, 0, 220, 36, 116, 
    386, 288, 318, 0, 130, 10, 22, 
    154, 97, 497, 209, 314, 80, 258, 
    254, 0, 0, 32, 114, 0, 245, 
    487, 428, 171, 288, 7, 39, 83, 
    204, 522, 58, 61, 64, 107, 125, 
    
    -- channel=39
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 61, 61, 59, 0, 
    0, 0, 0, 50, 53, 66, 140, 
    159, 0, 0, 0, 0, 63, 9, 
    243, 100, 78, 194, 92, 233, 108, 
    419, 265, 394, 552, 740, 903, 883, 
    807, 597, 798, 873, 972, 1010, 1094, 
    
    -- channel=40
    0, 0, 0, 0, 64, 101, 19, 
    0, 0, 0, 75, 187, 172, 198, 
    32, 26, 12, 26, 74, 162, 210, 
    96, 9, 123, 144, 173, 245, 189, 
    168, 26, 31, 112, 215, 327, 185, 
    417, 184, 499, 646, 584, 679, 663, 
    801, 642, 656, 716, 754, 820, 824, 
    
    -- channel=41
    58, 310, 201, 506, 99, 226, 0, 
    0, 108, 514, 970, 0, 829, 201, 
    6, 0, 463, 1578, 0, 1427, 566, 
    773, 460, 0, 951, 0, 1311, 0, 
    731, 32, 455, 576, 575, 423, 0, 
    0, 0, 1409, 256, 373, 0, 0, 
    0, 797, 140, 49, 0, 0, 0, 
    
    -- channel=42
    442, 504, 498, 372, 271, 181, 251, 
    127, 440, 407, 248, 136, 170, 57, 
    59, 413, 416, 234, 91, 158, 101, 
    76, 181, 278, 180, 161, 160, 146, 
    171, 0, 158, 192, 64, 0, 81, 
    0, 145, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=43
    0, 0, 0, 238, 0, 0, 81, 
    0, 0, 0, 0, 132, 0, 94, 
    59, 285, 29, 0, 20, 83, 0, 
    0, 0, 406, 235, 247, 206, 0, 
    71, 0, 0, 0, 306, 177, 0, 
    623, 322, 993, 884, 357, 337, 393, 
    813, 1052, 557, 412, 440, 594, 580, 
    
    -- channel=44
    978, 1019, 989, 683, 521, 422, 677, 
    682, 967, 736, 234, 394, 148, 306, 
    388, 911, 693, 170, 456, 65, 148, 
    69, 544, 630, 203, 454, 48, 460, 
    0, 107, 187, 214, 44, 0, 407, 
    0, 189, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=45
    229, 238, 189, 144, 164, 147, 215, 
    71, 228, 171, 52, 160, 92, 109, 
    54, 90, 169, 0, 30, 0, 139, 
    36, 52, 99, 45, 92, 27, 202, 
    73, 0, 67, 68, 37, 109, 174, 
    139, 0, 0, 161, 115, 180, 145, 
    140, 79, 151, 227, 233, 240, 213, 
    
    -- channel=46
    22, 20, 0, 62, 0, 53, 22, 
    57, 22, 69, 123, 0, 104, 101, 
    27, 96, 0, 151, 0, 185, 42, 
    45, 87, 0, 90, 8, 153, 0, 
    0, 62, 159, 7, 93, 92, 0, 
    0, 0, 220, 0, 24, 0, 0, 
    66, 0, 26, 0, 0, 0, 0, 
    
    -- channel=47
    1597, 1691, 1597, 1312, 834, 732, 1170, 
    923, 1503, 1053, 474, 447, 374, 530, 
    593, 1216, 838, 408, 312, 306, 322, 
    154, 788, 792, 499, 573, 299, 645, 
    96, 9, 205, 271, 332, 0, 613, 
    0, 131, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=48
    847, 953, 944, 425, 297, 380, 524, 
    747, 903, 847, 444, 301, 296, 219, 
    638, 479, 626, 596, 504, 259, 318, 
    463, 587, 413, 172, 339, 121, 471, 
    362, 392, 488, 561, 0, 0, 397, 
    0, 361, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=49
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 150, 116, 14, 20, 0, 
    14, 0, 61, 299, 270, 10, 179, 
    345, 0, 0, 0, 0, 0, 0, 
    326, 551, 443, 428, 0, 112, 0, 
    109, 241, 0, 0, 462, 612, 528, 
    232, 0, 481, 569, 626, 576, 637, 
    
    -- channel=50
    340, 278, 302, 161, 288, 188, 330, 
    238, 365, 131, 61, 435, 114, 165, 
    459, 358, 594, 0, 389, 73, 185, 
    304, 254, 507, 230, 371, 108, 419, 
    326, 336, 186, 289, 78, 73, 420, 
    608, 426, 85, 153, 119, 178, 213, 
    268, 165, 133, 151, 130, 178, 88, 
    
    -- channel=51
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 16, 0, 
    0, 0, 0, 0, 54, 77, 69, 
    85, 0, 70, 63, 71, 82, 69, 
    
    -- channel=52
    18, 0, 0, 0, 69, 0, 57, 
    308, 23, 0, 0, 305, 0, 110, 
    285, 123, 41, 0, 561, 0, 59, 
    100, 198, 236, 22, 316, 31, 170, 
    106, 442, 50, 83, 41, 231, 214, 
    440, 547, 135, 202, 272, 325, 288, 
    519, 355, 383, 268, 328, 372, 437, 
    
    -- channel=53
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 69, 36, 8, 
    76, 0, 0, 0, 126, 53, 82, 
    184, 0, 33, 39, 61, 52, 40, 
    289, 179, 82, 152, 46, 185, 85, 
    531, 402, 457, 538, 584, 743, 749, 
    819, 614, 680, 747, 828, 901, 967, 
    
    -- channel=54
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=55
    0, 0, 0, 0, 0, 54, 0, 
    52, 0, 0, 71, 330, 301, 95, 
    637, 0, 229, 302, 477, 397, 270, 
    874, 143, 384, 407, 377, 330, 216, 
    1070, 737, 395, 568, 428, 386, 357, 
    1352, 1266, 1296, 1301, 1215, 1432, 1522, 
    1680, 1599, 1418, 1471, 1596, 1765, 1925, 
    
    -- channel=56
    22, 0, 0, 0, 32, 0, 94, 
    276, 138, 0, 14, 111, 0, 156, 
    49, 220, 83, 0, 281, 105, 0, 
    0, 95, 0, 88, 33, 83, 14, 
    0, 311, 191, 0, 0, 223, 0, 
    88, 0, 268, 0, 120, 25, 0, 
    219, 0, 151, 17, 0, 34, 0, 
    
    -- channel=57
    0, 70, 66, 20, 0, 89, 0, 
    30, 22, 213, 216, 0, 121, 92, 
    0, 24, 0, 334, 0, 210, 103, 
    133, 100, 0, 0, 0, 157, 0, 
    42, 0, 202, 208, 37, 73, 0, 
    0, 0, 79, 0, 17, 5, 0, 
    0, 0, 0, 13, 22, 0, 48, 
    
    -- channel=58
    762, 809, 679, 639, 362, 143, 487, 
    226, 702, 325, 97, 9, 0, 89, 
    0, 521, 34, 0, 0, 0, 0, 
    0, 88, 16, 0, 4, 0, 41, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=59
    565, 640, 653, 450, 290, 376, 392, 
    414, 540, 547, 364, 155, 397, 203, 
    628, 308, 584, 612, 162, 415, 332, 
    658, 483, 384, 474, 270, 335, 349, 
    674, 339, 287, 505, 275, 0, 291, 
    183, 468, 0, 0, 0, 0, 0, 
    0, 160, 0, 0, 0, 0, 0, 
    
    -- channel=60
    28, 36, 21, 0, 7, 0, 15, 
    48, 20, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 0, 0, 18, 19, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=61
    66, 30, 100, 0, 83, 27, 79, 
    245, 93, 0, 0, 182, 0, 21, 
    263, 0, 0, 0, 367, 0, 77, 
    144, 110, 102, 5, 181, 0, 113, 
    156, 350, 0, 105, 58, 79, 227, 
    191, 419, 0, 72, 179, 206, 209, 
    182, 174, 199, 158, 189, 190, 268, 
    
    -- channel=62
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 
    0, 25, 0, 0, 0, 40, 0, 
    0, 0, 25, 22, 0, 44, 0, 
    7, 0, 0, 0, 64, 14, 0, 
    82, 0, 221, 174, 75, 93, 109, 
    173, 184, 118, 116, 120, 167, 150, 
    
    -- channel=63
    878, 965, 806, 721, 337, 214, 569, 
    352, 707, 348, 119, 0, 0, 194, 
    0, 394, 0, 0, 0, 0, 0, 
    0, 112, 0, 0, 0, 0, 96, 
    0, 0, 0, 0, 0, 0, 53, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=64
    9, 0, 0, 38, 98, 96, 74, 
    68, 9, 0, 102, 71, 82, 133, 
    4, 0, 0, 46, 34, 146, 166, 
    46, 91, 0, 69, 0, 136, 92, 
    1, 102, 107, 96, 128, 268, 150, 
    195, 0, 280, 235, 351, 372, 374, 
    365, 215, 330, 364, 375, 417, 398, 
    
    -- channel=65
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=66
    0, 8, 234, 87, 25, 0, 0, 
    0, 0, 63, 16, 0, 139, 0, 
    350, 0, 96, 382, 0, 75, 228, 
    613, 125, 288, 158, 150, 93, 65, 
    639, 87, 0, 472, 277, 0, 80, 
    151, 756, 0, 201, 0, 0, 20, 
    0, 1141, 0, 0, 6, 0, 132, 
    
    -- channel=67
    0, 0, 0, 0, 21, 27, 25, 
    50, 0, 0, 31, 0, 32, 59, 
    0, 0, 0, 11, 0, 74, 32, 
    0, 0, 0, 52, 0, 68, 30, 
    0, 39, 84, 0, 0, 131, 0, 
    44, 0, 159, 99, 143, 118, 128, 
    130, 0, 166, 154, 144, 181, 126, 
    
    -- channel=68
    0, 0, 0, 0, 0, 4, 0, 
    31, 0, 126, 145, 0, 93, 0, 
    8, 0, 0, 225, 72, 55, 136, 
    169, 0, 0, 0, 0, 0, 0, 
    91, 134, 183, 244, 0, 69, 47, 
    0, 59, 0, 0, 152, 229, 192, 
    57, 0, 161, 215, 248, 182, 247, 
    
    -- channel=69
    139, 195, 204, 189, 77, 66, 74, 
    0, 88, 128, 78, 0, 81, 0, 
    46, 0, 0, 122, 0, 44, 54, 
    85, 9, 0, 92, 0, 32, 0, 
    114, 0, 0, 37, 61, 0, 0, 
    0, 8, 0, 37, 0, 0, 0, 
    0, 195, 0, 0, 0, 0, 0, 
    
    -- channel=70
    86, 0, 53, 0, 249, 103, 138, 
    293, 236, 155, 114, 685, 209, 206, 
    459, 633, 800, 131, 847, 212, 197, 
    325, 308, 770, 404, 668, 273, 429, 
    515, 750, 419, 304, 199, 290, 280, 
    832, 906, 486, 361, 247, 318, 322, 
    549, 417, 346, 250, 249, 334, 271, 
    
    -- channel=71
    125, 62, 28, 276, 177, 161, 214, 
    0, 0, 0, 0, 112, 101, 222, 
    33, 291, 176, 0, 0, 95, 16, 
    0, 65, 304, 332, 212, 198, 122, 
    8, 0, 0, 0, 249, 217, 88, 
    356, 0, 452, 534, 74, 0, 17, 
    219, 534, 90, 0, 0, 35, 1, 
    
    -- channel=72
    342, 372, 408, 293, 296, 355, 326, 
    302, 303, 334, 273, 298, 349, 224, 
    540, 179, 421, 351, 218, 322, 341, 
    565, 345, 482, 413, 339, 260, 404, 
    612, 275, 252, 492, 299, 78, 433, 
    398, 510, 165, 263, 140, 153, 251, 
    83, 428, 84, 148, 146, 136, 173, 
    
    -- channel=73
    0, 0, 0, 0, 0, 51, 0, 
    198, 8, 165, 105, 165, 83, 23, 
    301, 0, 85, 240, 445, 60, 105, 
    423, 90, 83, 0, 141, 0, 40, 
    422, 511, 394, 437, 42, 26, 205, 
    245, 728, 129, 91, 366, 598, 548, 
    539, 113, 412, 503, 603, 577, 733, 
    
    -- channel=74
    365, 243, 275, 0, 399, 114, 349, 
    650, 584, 57, 0, 764, 0, 142, 
    488, 503, 449, 0, 1078, 0, 87, 
    100, 406, 605, 0, 552, 0, 450, 
    13, 782, 143, 162, 0, 187, 587, 
    627, 718, 0, 0, 30, 248, 186, 
    384, 0, 61, 48, 84, 153, 76, 
    
    -- channel=75
    1383, 1409, 1325, 1395, 702, 498, 967, 
    519, 1157, 758, 396, 290, 356, 367, 
    407, 1281, 963, 368, 103, 489, 94, 
    103, 615, 856, 736, 571, 569, 354, 
    174, 0, 0, 0, 445, 62, 205, 
    98, 188, 315, 0, 0, 0, 0, 
    0, 384, 0, 0, 0, 0, 0, 
    
    -- channel=76
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 37, 103, 175, 81, 
    125, 0, 0, 85, 82, 219, 254, 
    367, 0, 0, 104, 61, 285, 36, 
    493, 246, 0, 242, 310, 467, 128, 
    882, 570, 1227, 1312, 1440, 1659, 1641, 
    1740, 1390, 1693, 1705, 1857, 2010, 2148, 
    
    -- channel=77
    0, 0, 10, 13, 0, 0, 0, 
    0, 0, 0, 6, 0, 0, 8, 
    0, 0, 0, 13, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 12, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=78
    570, 617, 488, 414, 177, 93, 345, 
    210, 481, 189, 0, 53, 0, 122, 
    0, 465, 0, 0, 16, 0, 0, 
    0, 120, 93, 0, 33, 0, 83, 
    0, 0, 0, 0, 0, 0, 69, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=79
    0, 0, 7, 25, 64, 38, 0, 
    0, 0, 0, 147, 403, 327, 0, 
    772, 111, 788, 471, 536, 470, 248, 
    1017, 205, 781, 602, 560, 464, 216, 
    1284, 740, 176, 620, 448, 221, 224, 
    1336, 1567, 1209, 1070, 757, 813, 860, 
    918, 1716, 949, 854, 913, 1002, 1150, 
    
    -- channel=80
    1265, 1370, 1362, 1043, 685, 669, 928, 
    733, 1148, 881, 504, 455, 533, 396, 
    965, 695, 917, 652, 312, 463, 461, 
    753, 699, 837, 680, 605, 426, 693, 
    859, 330, 263, 657, 433, 0, 771, 
    362, 711, 0, 0, 0, 0, 0, 
    0, 315, 0, 0, 0, 0, 0, 
    
    -- channel=81
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=82
    69, 53, 43, 109, 42, 48, 74, 
    0, 0, 0, 0, 19, 0, 115, 
    0, 187, 0, 0, 0, 8, 0, 
    0, 5, 104, 39, 48, 92, 7, 
    0, 0, 0, 0, 69, 95, 21, 
    57, 0, 186, 169, 66, 40, 47, 
    220, 65, 113, 72, 71, 108, 102, 
    
    -- channel=83
    309, 385, 272, 78, 228, 241, 227, 
    414, 508, 445, 199, 133, 180, 133, 
    250, 111, 268, 260, 148, 130, 227, 
    234, 259, 0, 123, 47, 12, 222, 
    155, 357, 459, 273, 9, 128, 192, 
    0, 0, 0, 0, 69, 68, 75, 
    0, 0, 0, 26, 5, 0, 0, 
    
    -- channel=84
    0, 0, 18, 0, 49, 0, 0, 
    167, 144, 160, 79, 153, 78, 0, 
    288, 0, 201, 272, 439, 73, 197, 
    450, 108, 1, 0, 82, 3, 69, 
    444, 640, 330, 412, 0, 155, 148, 
    371, 576, 69, 160, 463, 589, 564, 
    443, 287, 460, 537, 602, 618, 702, 
    
    -- channel=85
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=86
    242, 210, 340, 157, 232, 0, 141, 
    244, 257, 100, 0, 307, 0, 0, 
    190, 144, 94, 0, 540, 0, 0, 
    41, 129, 383, 0, 326, 0, 105, 
    94, 294, 0, 71, 7, 0, 207, 
    166, 620, 0, 0, 0, 15, 0, 
    0, 281, 0, 0, 0, 0, 50, 
    
    -- channel=87
    0, 0, 0, 0, 0, 0, 0, 
    125, 0, 0, 0, 178, 0, 34, 
    217, 0, 0, 0, 393, 0, 39, 
    89, 4, 52, 2, 211, 56, 71, 
    161, 353, 0, 29, 1, 237, 92, 
    480, 538, 386, 434, 620, 709, 649, 
    803, 604, 818, 688, 801, 876, 961, 
    
    -- channel=88
    204, 195, 192, 124, 223, 232, 256, 
    390, 257, 156, 197, 352, 173, 335, 
    287, 122, 0, 105, 465, 107, 277, 
    136, 221, 132, 65, 296, 100, 323, 
    77, 349, 245, 222, 154, 236, 435, 
    141, 233, 0, 0, 227, 323, 298, 
    329, 0, 226, 245, 267, 276, 252, 
    
    -- channel=89
    1, 26, 199, 263, 0, 182, 43, 
    0, 0, 46, 268, 113, 464, 140, 
    673, 114, 502, 504, 0, 500, 209, 
    811, 135, 681, 642, 481, 561, 243, 
    1076, 81, 7, 496, 498, 0, 173, 
    744, 1109, 879, 750, 297, 245, 383, 
    415, 1316, 430, 362, 384, 400, 574, 
    
    -- channel=90
    232, 176, 135, 158, 275, 178, 329, 
    368, 274, 22, 69, 437, 103, 350, 
    119, 437, 6, 0, 478, 36, 196, 
    0, 249, 309, 155, 389, 160, 342, 
    0, 251, 117, 0, 180, 338, 311, 
    324, 167, 106, 169, 215, 251, 230, 
    444, 68, 279, 207, 220, 309, 229, 
    
    -- channel=91
    37, 29, 133, 0, 179, 36, 0, 
    272, 352, 356, 191, 420, 183, 0, 
    466, 0, 598, 382, 690, 138, 348, 
    603, 248, 216, 113, 241, 51, 304, 
    680, 900, 564, 671, 0, 173, 283, 
    580, 774, 0, 33, 425, 607, 556, 
    284, 149, 418, 511, 556, 539, 583, 
    
    -- channel=92
    16, 0, 0, 58, 0, 41, 107, 
    205, 0, 0, 0, 75, 0, 243, 
    24, 393, 0, 0, 145, 60, 0, 
    0, 94, 80, 11, 134, 50, 0, 
    0, 14, 140, 0, 80, 138, 47, 
    95, 0, 353, 129, 28, 35, 21, 
    429, 0, 98, 9, 20, 79, 37, 
    
    -- channel=93
    1316, 1446, 1436, 946, 612, 455, 802, 
    797, 1413, 1077, 488, 289, 214, 244, 
    373, 896, 695, 513, 467, 153, 218, 
    74, 605, 472, 160, 336, 103, 394, 
    0, 198, 276, 320, 0, 0, 349, 
    0, 41, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=94
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=95
    10, 6, 35, 150, 20, 66, 29, 
    0, 0, 45, 36, 0, 34, 25, 
    0, 88, 0, 6, 0, 63, 0, 
    40, 15, 130, 14, 6, 48, 0, 
    37, 0, 19, 26, 184, 18, 55, 
    74, 71, 178, 197, 37, 53, 107, 
    106, 307, 8, 34, 47, 72, 81, 
    
    -- channel=96
    74, 101, 94, 131, 110, 121, 61, 
    37, 93, 202, 188, 0, 206, 58, 
    85, 56, 225, 284, 0, 217, 119, 
    200, 62, 48, 244, 32, 191, 36, 
    266, 101, 173, 163, 142, 99, 5, 
    92, 93, 242, 167, 143, 46, 87, 
    0, 166, 84, 71, 60, 35, 77, 
    
    -- channel=97
    164, 100, 30, 352, 203, 136, 259, 
    0, 29, 0, 0, 83, 74, 173, 
    0, 374, 195, 0, 0, 72, 0, 
    0, 34, 302, 381, 181, 190, 97, 
    0, 0, 0, 0, 235, 165, 0, 
    294, 0, 617, 570, 6, 0, 0, 
    160, 500, 55, 0, 0, 0, 0, 
    
    -- channel=98
    535, 572, 716, 530, 170, 186, 352, 
    95, 290, 264, 38, 158, 122, 0, 
    643, 430, 684, 153, 77, 114, 0, 
    538, 224, 878, 363, 461, 122, 217, 
    776, 0, 0, 360, 190, 0, 339, 
    574, 1051, 29, 150, 0, 0, 0, 
    0, 763, 0, 0, 0, 0, 0, 
    
    -- channel=99
    289, 248, 287, 54, 234, 170, 322, 
    513, 300, 31, 0, 722, 135, 266, 
    770, 415, 350, 0, 897, 64, 227, 
    488, 350, 817, 230, 769, 79, 567, 
    601, 686, 234, 431, 206, 154, 695, 
    968, 1178, 260, 468, 440, 706, 751, 
    962, 718, 597, 597, 713, 814, 874, 
    
    -- channel=100
    0, 0, 0, 41, 0, 0, 0, 
    0, 0, 17, 176, 0, 90, 171, 
    0, 316, 0, 123, 0, 258, 0, 
    0, 11, 0, 98, 0, 268, 0, 
    0, 0, 221, 0, 0, 158, 0, 
    0, 0, 388, 0, 56, 0, 0, 
    169, 0, 90, 0, 0, 0, 0, 
    
    -- channel=101
    0, 0, 0, 0, 0, 0, 0, 
    253, 281, 370, 168, 0, 0, 0, 
    0, 0, 0, 344, 247, 0, 227, 
    152, 66, 0, 0, 0, 0, 1, 
    0, 490, 503, 432, 0, 78, 40, 
    0, 0, 0, 0, 73, 215, 113, 
    0, 0, 7, 131, 159, 30, 100, 
    
    -- channel=102
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=103
    1500, 1571, 1427, 1293, 769, 725, 1165, 
    854, 1274, 917, 276, 397, 262, 542, 
    529, 1221, 724, 111, 135, 127, 125, 
    37, 626, 869, 497, 598, 175, 581, 
    15, 0, 20, 8, 330, 0, 534, 
    0, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=104
    844, 913, 860, 563, 499, 494, 655, 
    630, 871, 666, 290, 367, 331, 339, 
    593, 447, 554, 358, 288, 215, 361, 
    407, 505, 454, 368, 404, 175, 541, 
    414, 248, 327, 447, 219, 43, 577, 
    112, 299, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=105
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 32, 57, 36, 
    144, 0, 0, 0, 0, 78, 0, 
    272, 117, 0, 70, 126, 244, 0, 
    542, 480, 988, 950, 1067, 1300, 1251, 
    1417, 967, 1317, 1328, 1487, 1595, 1734, 
    
    -- channel=106
    0, 0, 0, 16, 0, 76, 0, 
    0, 0, 0, 196, 0, 129, 123, 
    0, 0, 0, 155, 0, 241, 126, 
    85, 16, 0, 61, 0, 218, 0, 
    45, 51, 115, 80, 173, 224, 26, 
    142, 4, 565, 380, 554, 567, 556, 
    610, 305, 610, 584, 630, 657, 704, 
    
    -- channel=107
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 146, 0, 0, 
    0, 0, 0, 0, 265, 0, 33, 
    68, 0, 27, 0, 79, 52, 0, 
    249, 222, 49, 84, 109, 286, 0, 
    599, 554, 727, 837, 936, 1191, 1101, 
    1336, 828, 1197, 1210, 1355, 1460, 1553, 
    
    -- channel=108
    233, 274, 186, 298, 43, 95, 118, 
    29, 169, 145, 252, 0, 183, 82, 
    0, 94, 4, 340, 0, 318, 90, 
    49, 82, 0, 191, 0, 311, 0, 
    38, 0, 62, 4, 138, 55, 0, 
    0, 0, 418, 36, 94, 0, 0, 
    0, 104, 93, 54, 21, 45, 29, 
    
    -- channel=109
    358, 353, 411, 14, 154, 201, 237, 
    613, 542, 401, 119, 448, 202, 92, 
    970, 296, 700, 401, 796, 204, 228, 
    893, 478, 520, 225, 477, 63, 400, 
    904, 999, 569, 708, 66, 0, 486, 
    769, 1214, 85, 25, 183, 361, 380, 
    381, 327, 209, 281, 322, 341, 433, 
    
    -- channel=110
    199, 206, 233, 236, 229, 78, 157, 
    46, 121, 48, 78, 183, 107, 71, 
    124, 281, 195, 34, 132, 116, 78, 
    109, 108, 379, 274, 277, 202, 163, 
    250, 68, 0, 93, 175, 118, 111, 
    338, 383, 375, 354, 171, 134, 187, 
    196, 545, 251, 132, 162, 215, 241, 
    
    -- channel=111
    87, 70, 36, 135, 54, 130, 120, 
    211, 102, 89, 131, 0, 132, 118, 
    188, 0, 6, 201, 0, 184, 94, 
    140, 159, 0, 149, 0, 127, 18, 
    82, 172, 147, 45, 138, 93, 57, 
    52, 0, 212, 48, 94, 8, 32, 
    6, 78, 55, 40, 11, 14, 21, 
    
    -- channel=112
    395, 326, 283, 105, 282, 103, 342, 
    399, 481, 131, 0, 458, 0, 113, 
    327, 502, 514, 0, 523, 0, 14, 
    14, 244, 442, 84, 348, 0, 345, 
    37, 334, 98, 50, 0, 64, 332, 
    488, 321, 0, 0, 0, 0, 0, 
    115, 0, 0, 0, 0, 0, 0, 
    
    -- channel=113
    314, 233, 245, 430, 249, 227, 374, 
    159, 105, 13, 3, 335, 131, 247, 
    370, 612, 475, 0, 209, 188, 3, 
    179, 300, 722, 455, 519, 286, 255, 
    332, 56, 0, 2, 368, 114, 227, 
    670, 591, 623, 600, 43, 0, 31, 
    341, 797, 107, 0, 0, 34, 50, 
    
    -- channel=114
    9, 0, 148, 0, 0, 11, 0, 
    218, 36, 169, 93, 301, 132, 0, 
    609, 136, 467, 423, 756, 180, 108, 
    793, 200, 368, 66, 350, 77, 77, 
    886, 846, 339, 592, 103, 58, 206, 
    726, 1465, 605, 465, 656, 944, 815, 
    918, 757, 837, 902, 1024, 1033, 1241, 
    
    -- channel=115
    0, 0, 6, 0, 7, 0, 0, 
    0, 0, 0, 0, 26, 0, 0, 
    0, 0, 1, 0, 56, 0, 11, 
    0, 0, 22, 0, 1, 0, 15, 
    0, 11, 0, 28, 0, 0, 0, 
    7, 63, 0, 0, 0, 29, 29, 
    0, 24, 0, 2, 23, 17, 35, 
    
    -- channel=116
    229, 299, 384, 52, 145, 258, 112, 
    409, 375, 466, 382, 133, 304, 39, 
    671, 0, 390, 652, 372, 348, 373, 
    852, 347, 84, 172, 114, 168, 223, 
    806, 709, 564, 801, 126, 24, 419, 
    365, 742, 53, 0, 376, 492, 517, 
    147, 172, 280, 398, 424, 356, 495, 
    
    -- channel=117
    27, 49, 126, 29, 30, 55, 15, 
    22, 0, 53, 168, 62, 156, 78, 
    145, 18, 170, 242, 92, 180, 155, 
    167, 55, 109, 134, 92, 206, 114, 
    211, 66, 75, 203, 61, 36, 69, 
    40, 215, 35, 0, 82, 62, 55, 
    0, 86, 68, 66, 67, 27, 53, 
    
    -- channel=118
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 10, 0, 37, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 43, 32, 0, 4, 23, 0, 
    0, 0, 74, 0, 95, 79, 65, 
    13, 0, 80, 85, 77, 86, 61, 
    
    -- channel=119
    32, 0, 0, 0, 0, 0, 203, 
    631, 173, 0, 0, 219, 0, 452, 
    108, 629, 0, 0, 586, 184, 0, 
    0, 207, 0, 37, 133, 138, 21, 
    0, 567, 488, 0, 0, 336, 18, 
    156, 0, 498, 0, 147, 58, 0, 
    673, 0, 217, 34, 0, 108, 0, 
    
    -- channel=120
    185, 129, 145, 0, 218, 93, 159, 
    504, 492, 206, 0, 767, 0, 97, 
    471, 470, 476, 0, 1161, 0, 145, 
    298, 311, 556, 0, 487, 0, 407, 
    283, 851, 629, 622, 0, 213, 790, 
    873, 1065, 0, 107, 597, 1112, 977, 
    1109, 0, 623, 800, 963, 1009, 1044, 
    
    -- channel=121
    198, 173, 197, 326, 130, 163, 207, 
    176, 139, 104, 156, 73, 204, 161, 
    340, 167, 184, 258, 61, 335, 129, 
    343, 246, 230, 358, 220, 315, 109, 
    320, 205, 79, 120, 296, 117, 127, 
    310, 269, 417, 257, 28, 0, 13, 
    78, 602, 45, 0, 0, 0, 0, 
    
    -- channel=122
    2168, 2244, 2108, 1741, 1192, 1010, 1653, 
    1414, 2020, 1362, 705, 689, 517, 880, 
    796, 1494, 945, 525, 546, 426, 601, 
    89, 1166, 986, 692, 760, 463, 1028, 
    0, 67, 236, 304, 445, 46, 881, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=123
    59, 0, 0, 32, 36, 44, 194, 
    308, 97, 0, 0, 253, 0, 209, 
    185, 322, 0, 0, 332, 26, 0, 
    0, 123, 162, 57, 262, 13, 92, 
    0, 263, 204, 0, 72, 165, 146, 
    312, 39, 193, 140, 43, 63, 92, 
    378, 20, 88, 9, 0, 94, 0, 
    
    -- channel=124
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 
    0, 0, 0, 0, 14, 0, 0, 
    54, 0, 0, 0, 0, 0, 0, 
    176, 56, 0, 12, 48, 191, 0, 
    513, 305, 526, 708, 728, 890, 885, 
    962, 730, 858, 888, 990, 1080, 1157, 
    
    -- channel=125
    362, 427, 448, 87, 245, 224, 262, 
    382, 506, 382, 137, 374, 203, 49, 
    558, 49, 433, 303, 435, 90, 330, 
    548, 304, 359, 154, 330, 0, 426, 
    611, 526, 280, 562, 104, 0, 453, 
    348, 680, 0, 0, 83, 221, 264, 
    0, 220, 0, 113, 147, 116, 186, 
    
    -- channel=126
    201, 240, 252, 442, 13, 147, 152, 
    0, 0, 0, 195, 0, 309, 139, 
    355, 95, 274, 401, 0, 470, 61, 
    438, 106, 203, 585, 73, 541, 4, 
    565, 0, 0, 67, 338, 6, 0, 
    289, 243, 943, 562, 130, 0, 0, 
    102, 879, 226, 53, 16, 49, 162, 
    
    -- channel=127
    0, 31, 0, 100, 0, 35, 0, 
    0, 0, 32, 146, 0, 139, 52, 
    0, 43, 0, 220, 0, 246, 27, 
    56, 30, 0, 92, 0, 224, 0, 
    47, 0, 79, 40, 140, 3, 0, 
    0, 0, 217, 62, 49, 0, 23, 
    0, 186, 16, 21, 7, 24, 11, 
    
    
    others => 0);
end inmem_package;
