library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    64, 70, 71, 69, 68, 67, 72, 76, 68, 51, 44, 53, 59, 58, 56, 
    71, 74, 74, 69, 74, 85, 54, 55, 35, 40, 18, 15, 29, 52, 55, 
    28, 64, 72, 73, 72, 59, 34, 18, 21, 47, 14, 21, 2, 20, 58, 
    0, 56, 63, 76, 55, 58, 34, 12, 13, 46, 21, 17, 9, 0, 54, 
    6, 45, 47, 88, 68, 43, 22, 11, 3, 61, 34, 6, 21, 3, 17, 
    0, 41, 49, 45, 66, 48, 38, 22, 0, 86, 14, 4, 23, 12, 7, 
    13, 12, 43, 44, 58, 69, 36, 28, 1, 73, 11, 7, 19, 28, 12, 
    22, 29, 13, 38, 50, 59, 8, 23, 17, 62, 26, 4, 24, 23, 43, 
    20, 35, 0, 46, 23, 32, 27, 22, 38, 26, 24, 0, 19, 46, 56, 
    41, 36, 0, 46, 4, 22, 54, 31, 8, 20, 0, 5, 30, 62, 53, 
    53, 36, 0, 92, 25, 6, 30, 16, 0, 0, 0, 0, 0, 0, 0, 
    0, 37, 27, 82, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 60, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    
    -- channel=1
    24, 23, 24, 27, 25, 24, 25, 24, 25, 26, 19, 17, 18, 20, 19, 
    24, 25, 26, 27, 27, 36, 32, 24, 10, 13, 21, 16, 11, 16, 23, 
    23, 15, 23, 25, 24, 34, 7, 10, 9, 23, 33, 26, 19, 13, 17, 
    35, 19, 29, 26, 25, 20, 37, 20, 15, 26, 23, 16, 8, 6, 13, 
    40, 53, 32, 36, 73, 41, 34, 16, 11, 1, 40, 25, 20, 17, 3, 
    26, 45, 30, 0, 21, 15, 35, 32, 23, 23, 38, 15, 23, 21, 11, 
    25, 40, 21, 22, 24, 22, 57, 27, 34, 31, 32, 19, 12, 21, 25, 
    25, 49, 30, 37, 27, 62, 34, 17, 21, 28, 21, 19, 17, 22, 16, 
    38, 46, 18, 27, 18, 8, 18, 23, 30, 16, 24, 5, 1, 16, 26, 
    37, 42, 35, 22, 45, 8, 18, 50, 25, 21, 9, 4, 22, 28, 27, 
    38, 39, 34, 45, 59, 59, 42, 43, 31, 12, 18, 20, 22, 29, 23, 
    38, 28, 48, 63, 43, 0, 5, 5, 12, 18, 20, 19, 21, 24, 23, 
    26, 23, 21, 61, 20, 18, 19, 16, 18, 20, 24, 29, 29, 24, 33, 
    27, 19, 24, 47, 19, 22, 20, 19, 17, 22, 21, 24, 18, 30, 26, 
    26, 19, 7, 33, 15, 14, 20, 20, 23, 25, 25, 20, 32, 44, 26, 
    
    -- channel=2
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 25, 11, 0, 0, 0, 29, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 20, 0, 0, 
    53, 0, 0, 0, 1, 0, 20, 10, 2, 0, 18, 0, 5, 8, 0, 
    65, 10, 17, 0, 58, 29, 13, 18, 0, 0, 19, 32, 4, 31, 0, 
    9, 0, 25, 0, 0, 0, 34, 23, 40, 0, 8, 15, 0, 17, 35, 
    33, 0, 0, 8, 0, 0, 0, 24, 26, 0, 21, 23, 0, 1, 17, 
    24, 21, 31, 28, 0, 0, 0, 0, 7, 0, 4, 13, 0, 0, 1, 
    21, 0, 42, 0, 8, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 50, 0, 9, 0, 0, 34, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 31, 0, 127, 55, 0, 0, 23, 28, 24, 27, 5, 0, 3, 
    0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 9, 2, 0, 0, 0, 2, 5, 5, 0, 0, 12, 
    12, 2, 0, 0, 4, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 3, 12, 3, 0, 6, 16, 30, 
    
    -- channel=3
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 1, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 7, 5, 0, 0, 8, 9, 0, 
    0, 30, 0, 0, 0, 41, 0, 0, 0, 35, 5, 4, 0, 8, 18, 
    0, 20, 0, 0, 0, 2, 0, 0, 4, 50, 1, 12, 0, 0, 38, 
    0, 29, 0, 9, 3, 0, 2, 0, 4, 36, 6, 0, 5, 0, 5, 
    0, 44, 0, 0, 93, 22, 8, 0, 0, 62, 0, 0, 17, 0, 0, 
    0, 38, 12, 0, 61, 26, 36, 0, 0, 83, 0, 0, 8, 11, 0, 
    0, 28, 0, 0, 20, 61, 6, 28, 0, 61, 11, 0, 19, 22, 3, 
    4, 43, 0, 40, 0, 45, 9, 3, 17, 15, 24, 0, 21, 22, 2, 
    36, 39, 0, 54, 0, 0, 22, 13, 0, 15, 5, 3, 22, 18, 0, 
    76, 31, 0, 61, 0, 0, 42, 43, 0, 0, 0, 0, 11, 24, 5, 
    82, 66, 12, 83, 30, 16, 38, 34, 14, 15, 19, 24, 23, 23, 15, 
    12, 66, 53, 56, 0, 17, 18, 18, 15, 14, 19, 17, 25, 27, 22, 
    13, 23, 73, 53, 3, 21, 11, 15, 21, 20, 24, 30, 23, 22, 39, 
    11, 26, 32, 51, 14, 28, 29, 19, 20, 18, 14, 22, 29, 18, 5, 
    
    -- channel=4
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 10, 7, 0, 9, 6, 8, 0, 0, 
    15, 0, 0, 0, 0, 0, 0, 5, 6, 0, 4, 6, 14, 9, 0, 
    20, 0, 0, 0, 0, 0, 7, 11, 12, 0, 5, 10, 6, 9, 0, 
    30, 0, 0, 0, 0, 0, 0, 7, 13, 0, 8, 18, 6, 9, 9, 
    27, 10, 0, 0, 0, 0, 0, 2, 15, 0, 18, 18, 11, 8, 2, 
    23, 18, 10, 0, 0, 0, 6, 7, 5, 0, 6, 20, 9, 0, 0, 
    22, 20, 29, 0, 2, 9, 11, 8, 0, 0, 9, 15, 7, 0, 0, 
    10, 13, 28, 12, 22, 1, 1, 6, 10, 1, 13, 20, 0, 0, 0, 
    14, 15, 30, 0, 6, 18, 3, 21, 25, 30, 38, 33, 34, 39, 44, 
    50, 23, 14, 0, 47, 67, 60, 62, 57, 53, 54, 56, 59, 58, 62, 
    66, 46, 16, 15, 67, 52, 52, 52, 54, 55, 58, 59, 57, 61, 62, 
    73, 62, 36, 40, 50, 52, 54, 54, 53, 57, 62, 65, 67, 68, 67, 
    70, 65, 59, 64, 56, 55, 52, 49, 48, 55, 61, 60, 53, 65, 71, 
    
    -- channel=5
    2, 1, 2, 3, 6, 2, 3, 10, 13, 14, 11, 6, 1, 0, 1, 
    6, 3, 3, 5, 3, 0, 3, 16, 13, 0, 0, 0, 0, 3, 3, 
    15, 15, 8, 6, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 10, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=6
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 43, 1, 0, 0, 0, 16, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 16, 5, 8, 2, 0, 0, 
    19, 29, 0, 0, 0, 0, 27, 9, 0, 0, 0, 0, 0, 0, 0, 
    30, 66, 0, 11, 97, 55, 0, 0, 0, 0, 22, 15, 8, 14, 0, 
    0, 0, 0, 0, 0, 0, 15, 16, 16, 40, 0, 0, 0, 7, 27, 
    6, 0, 0, 0, 0, 7, 0, 2, 1, 5, 0, 0, 0, 11, 17, 
    4, 6, 16, 8, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 1, 43, 0, 0, 0, 0, 25, 16, 0, 
    0, 0, 0, 62, 104, 89, 14, 0, 0, 0, 28, 46, 16, 0, 0, 
    0, 0, 16, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 5, 11, 19, 0, 0, 25, 
    0, 0, 0, 0, 0, 2, 7, 0, 0, 2, 0, 0, 0, 16, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 16, 17, 2, 0, 38, 26, 0, 
    
    -- channel=7
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 7, 0, 0, 0, 15, 0, 0, 0, 7, 0, 
    0, 27, 0, 0, 0, 10, 0, 0, 1, 31, 0, 0, 0, 0, 13, 
    0, 26, 0, 0, 0, 22, 0, 0, 0, 34, 0, 0, 0, 0, 37, 
    0, 14, 0, 47, 12, 0, 0, 0, 0, 48, 0, 0, 0, 0, 0, 
    0, 5, 0, 0, 47, 0, 0, 0, 0, 71, 0, 0, 10, 0, 0, 
    0, 0, 0, 0, 43, 10, 0, 0, 0, 59, 0, 0, 0, 10, 0, 
    0, 2, 0, 0, 24, 24, 0, 0, 0, 26, 0, 0, 11, 0, 0, 
    0, 0, 0, 25, 0, 9, 0, 0, 26, 0, 1, 0, 7, 19, 0, 
    0, 0, 0, 37, 0, 0, 29, 0, 0, 0, 0, 9, 28, 7, 0, 
    43, 0, 0, 77, 0, 0, 0, 0, 0, 0, 8, 2, 0, 1, 0, 
    23, 20, 0, 29, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 8, 39, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 1, 11, 
    0, 0, 21, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 20, 0, 0, 0, 0, 2, 0, 0, 4, 25, 0, 0, 
    
    -- channel=8
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=9
    24, 27, 27, 26, 29, 27, 29, 35, 34, 27, 22, 22, 20, 23, 24, 
    29, 31, 30, 28, 24, 10, 26, 36, 24, 0, 0, 3, 18, 14, 19, 
    35, 14, 30, 31, 33, 30, 14, 11, 0, 0, 0, 0, 0, 6, 8, 
    0, 5, 21, 32, 36, 4, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 7, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=10
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 19, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 38, 0, 0, 0, 17, 10, 0, 
    28, 37, 0, 0, 0, 47, 14, 16, 0, 0, 0, 0, 0, 20, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 11, 0, 0, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 19, 70, 16, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 20, 0, 25, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 12, 16, 28, 0, 4, 0, 0, 4, 6, 0, 
    0, 0, 0, 0, 0, 50, 0, 0, 0, 0, 37, 31, 13, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 42, 30, 9, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 34, 6, 0, 0, 0, 0, 20, 19, 
    78, 27, 0, 0, 63, 60, 42, 39, 16, 5, 0, 0, 0, 0, 0, 
    0, 57, 4, 14, 39, 0, 0, 0, 0, 0, 0, 0, 1, 4, 0, 
    0, 0, 62, 46, 4, 0, 0, 0, 0, 0, 1, 11, 0, 0, 33, 
    0, 0, 11, 50, 15, 23, 22, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=11
    35, 39, 36, 38, 36, 36, 37, 42, 38, 31, 23, 23, 26, 32, 34, 
    36, 41, 39, 39, 36, 40, 25, 31, 19, 4, 1, 4, 11, 22, 32, 
    29, 24, 38, 40, 42, 47, 7, 3, 0, 8, 0, 0, 5, 8, 26, 
    11, 16, 35, 37, 32, 9, 15, 0, 1, 7, 0, 4, 0, 3, 22, 
    0, 20, 17, 8, 15, 0, 0, 0, 5, 0, 0, 0, 5, 3, 6, 
    0, 2, 7, 22, 16, 0, 4, 0, 10, 8, 0, 0, 4, 0, 0, 
    0, 13, 1, 31, 33, 0, 10, 0, 4, 17, 0, 0, 0, 0, 3, 
    0, 0, 0, 15, 13, 20, 0, 0, 0, 24, 0, 0, 0, 7, 7, 
    0, 0, 0, 2, 0, 0, 0, 10, 0, 14, 16, 0, 3, 14, 32, 
    0, 0, 0, 0, 0, 0, 0, 10, 0, 2, 0, 0, 12, 29, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=12
    64, 67, 67, 71, 69, 67, 67, 69, 69, 62, 55, 52, 59, 59, 56, 
    64, 66, 67, 72, 70, 98, 88, 66, 52, 56, 69, 54, 40, 44, 58, 
    58, 37, 68, 70, 67, 79, 75, 50, 39, 66, 99, 82, 65, 26, 44, 
    95, 31, 71, 69, 80, 70, 93, 71, 58, 52, 111, 64, 63, 30, 15, 
    140, 96, 97, 74, 157, 135, 125, 83, 52, 36, 116, 93, 61, 54, 14, 
    144, 123, 112, 67, 84, 122, 141, 100, 76, 38, 150, 95, 58, 69, 47, 
    150, 133, 73, 79, 50, 105, 145, 125, 94, 61, 142, 88, 59, 67, 73, 
    158, 156, 99, 93, 61, 111, 154, 89, 82, 69, 119, 89, 51, 70, 69, 
    176, 152, 136, 81, 96, 76, 89, 82, 67, 92, 59, 68, 30, 47, 60, 
    159, 153, 149, 83, 110, 72, 88, 132, 89, 68, 62, 23, 29, 61, 79, 
    116, 154, 148, 105, 213, 130, 107, 139, 112, 71, 48, 53, 62, 70, 75, 
    74, 125, 151, 158, 200, 103, 71, 70, 68, 64, 68, 73, 81, 87, 89, 
    91, 67, 116, 191, 149, 76, 73, 69, 70, 71, 78, 87, 89, 88, 103, 
    97, 72, 66, 171, 94, 80, 84, 70, 69, 77, 83, 82, 85, 89, 97, 
    105, 77, 69, 82, 68, 57, 68, 76, 80, 92, 88, 79, 96, 129, 96, 
    
    -- channel=13
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 17, 11, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 7, 11, 0, 2, 2, 0, 0, 
    19, 11, 0, 0, 0, 0, 0, 0, 6, 5, 5, 1, 5, 2, 0, 
    36, 20, 0, 0, 7, 0, 0, 0, 3, 15, 11, 4, 10, 9, 3, 
    31, 26, 0, 0, 0, 0, 8, 1, 5, 25, 12, 8, 11, 11, 1, 
    29, 27, 10, 0, 0, 15, 14, 7, 0, 5, 4, 8, 13, 4, 0, 
    40, 42, 24, 6, 0, 6, 0, 3, 6, 0, 0, 0, 5, 0, 0, 
    28, 38, 23, 35, 15, 3, 5, 12, 15, 0, 4, 9, 2, 0, 0, 
    38, 31, 25, 38, 26, 35, 43, 38, 28, 23, 40, 49, 61, 55, 50, 
    94, 53, 31, 40, 51, 59, 68, 68, 70, 74, 81, 86, 89, 90, 88, 
    104, 84, 45, 44, 58, 76, 77, 73, 76, 81, 91, 95, 94, 97, 103, 
    109, 96, 85, 53, 65, 81, 78, 77, 79, 87, 97, 101, 100, 111, 109, 
    104, 102, 90, 77, 76, 81, 81, 78, 81, 88, 91, 92, 98, 111, 100, 
    
    -- channel=14
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 28, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 19, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 10, 3, 0, 0, 15, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 23, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 2, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 2, 0, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 20, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 2, 6, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 8, 17, 0, 15, 8, 14, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 18, 0, 0, 0, 2, 1, 8, 
    27, 15, 0, 0, 31, 0, 0, 0, 3, 0, 12, 8, 10, 2, 0, 
    11, 30, 0, 0, 4, 0, 10, 0, 6, 13, 10, 8, 9, 4, 4, 
    15, 5, 1, 0, 0, 18, 16, 20, 3, 13, 9, 14, 15, 15, 0, 
    20, 22, 24, 1, 0, 18, 3, 6, 0, 0, 28, 16, 16, 0, 0, 
    20, 27, 17, 12, 19, 3, 0, 0, 23, 17, 12, 9, 0, 0, 0, 
    22, 18, 19, 0, 0, 6, 28, 32, 19, 4, 17, 19, 35, 29, 26, 
    86, 33, 5, 15, 69, 63, 63, 61, 56, 52, 57, 60, 60, 65, 64, 
    76, 79, 17, 48, 50, 52, 56, 54, 54, 57, 59, 62, 68, 66, 58, 
    78, 68, 77, 52, 48, 54, 52, 58, 57, 61, 71, 78, 70, 75, 97, 
    75, 74, 73, 69, 63, 70, 67, 53, 51, 55, 68, 63, 53, 73, 71, 
    
    -- channel=16
    58, 59, 59, 58, 55, 56, 59, 55, 51, 51, 49, 48, 47, 45, 38, 
    51, 50, 59, 59, 60, 76, 60, 54, 47, 43, 43, 35, 37, 41, 41, 
    54, 51, 56, 56, 59, 89, 64, 30, 28, 74, 90, 70, 44, 31, 43, 
    31, 37, 54, 56, 55, 50, 65, 55, 52, 89, 91, 68, 48, 22, 36, 
    88, 90, 71, 78, 113, 113, 102, 64, 45, 65, 92, 62, 48, 26, 24, 
    133, 137, 86, 89, 153, 144, 117, 70, 34, 95, 136, 74, 59, 50, 24, 
    132, 130, 76, 44, 82, 124, 144, 104, 58, 115, 118, 64, 53, 61, 56, 
    153, 130, 82, 49, 70, 155, 147, 105, 66, 113, 117, 66, 60, 78, 61, 
    170, 161, 111, 93, 87, 99, 77, 68, 67, 68, 77, 58, 43, 57, 63, 
    171, 168, 113, 100, 94, 78, 89, 95, 87, 87, 51, 13, 31, 60, 60, 
    144, 158, 114, 145, 148, 94, 142, 154, 94, 37, 22, 39, 61, 73, 64, 
    132, 161, 135, 201, 200, 109, 86, 84, 72, 65, 71, 77, 83, 90, 86, 
    88, 119, 158, 209, 122, 76, 73, 69, 65, 67, 75, 85, 95, 95, 99, 
    91, 79, 147, 167, 87, 81, 74, 69, 73, 80, 89, 94, 87, 99, 117, 
    97, 84, 90, 85, 68, 76, 85, 79, 81, 87, 84, 81, 100, 117, 78, 
    
    -- channel=17
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 9, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 17, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 16, 2, 0, 11, 11, 0, 0, 0, 0, 
    35, 31, 0, 11, 55, 37, 17, 3, 0, 21, 30, 8, 4, 0, 0, 
    28, 30, 0, 0, 21, 28, 37, 14, 0, 44, 21, 0, 2, 5, 0, 
    39, 30, 0, 0, 4, 41, 32, 24, 3, 41, 22, 7, 5, 18, 0, 
    49, 48, 8, 0, 14, 39, 6, 4, 0, 20, 22, 2, 6, 0, 0, 
    58, 55, 19, 25, 8, 1, 7, 14, 10, 0, 0, 0, 0, 0, 0, 
    49, 52, 29, 43, 14, 0, 26, 46, 1, 0, 0, 0, 0, 0, 0, 
    53, 51, 24, 77, 88, 47, 45, 31, 11, 5, 15, 29, 22, 13, 11, 
    21, 48, 48, 84, 33, 11, 17, 18, 20, 23, 28, 32, 39, 39, 37, 
    35, 22, 55, 56, 11, 32, 29, 26, 27, 32, 40, 43, 38, 42, 55, 
    40, 36, 33, 27, 26, 34, 34, 29, 31, 36, 37, 36, 40, 52, 30, 
    40, 41, 33, 11, 16, 20, 23, 31, 41, 45, 36, 37, 64, 59, 35, 
    
    -- channel=18
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 7, 0, 0, 1, 0, 0, 
    0, 11, 0, 0, 0, 0, 24, 35, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 18, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 
    0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 9, 0, 2, 8, 0, 0, 10, 
    0, 0, 0, 0, 0, 29, 18, 0, 0, 0, 0, 41, 8, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 34, 21, 0, 0, 0, 
    0, 0, 13, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 4, 14, 
    0, 0, 0, 0, 0, 83, 38, 38, 25, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 86, 0, 0, 2, 4, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 26, 19, 0, 0, 0, 0, 0, 0, 1, 15, 0, 0, 
    1, 0, 0, 48, 16, 4, 4, 2, 0, 0, 0, 7, 0, 0, 19, 
    
    -- channel=19
    42, 40, 44, 43, 45, 39, 42, 46, 45, 33, 28, 30, 35, 37, 38, 
    46, 39, 43, 43, 46, 47, 39, 33, 27, 33, 25, 19, 22, 32, 36, 
    20, 38, 43, 46, 45, 19, 38, 26, 20, 17, 7, 20, 15, 19, 33, 
    12, 36, 40, 44, 39, 42, 19, 16, 17, 9, 20, 9, 17, 15, 25, 
    23, 15, 40, 50, 26, 25, 14, 16, 8, 33, 18, 15, 15, 14, 16, 
    18, 16, 40, 30, 9, 25, 21, 16, 10, 22, 14, 18, 11, 16, 19, 
    28, 2, 32, 27, 10, 32, 4, 25, 7, 12, 18, 16, 18, 17, 14, 
    24, 12, 29, 28, 22, 0, 15, 13, 16, 13, 25, 13, 12, 8, 32, 
    19, 9, 17, 21, 23, 17, 22, 16, 24, 25, 1, 12, 14, 31, 36, 
    18, 13, 13, 19, 2, 20, 32, 10, 10, 8, 12, 10, 12, 23, 31, 
    7, 13, 11, 23, 34, 6, 0, 0, 7, 15, 8, 7, 6, 17, 20, 
    0, 10, 18, 11, 0, 9, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 30, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    
    -- channel=20
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 7, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 21, 10, 5, 0, 15, 18, 11, 0, 0, 
    21, 0, 0, 0, 0, 0, 16, 4, 6, 2, 38, 24, 20, 11, 0, 
    22, 0, 0, 0, 9, 0, 15, 27, 15, 14, 36, 24, 12, 12, 0, 
    47, 25, 30, 1, 36, 64, 50, 32, 15, 0, 32, 38, 9, 8, 15, 
    89, 47, 42, 22, 16, 62, 39, 28, 15, 0, 76, 42, 13, 16, 14, 
    89, 51, 34, 0, 0, 32, 53, 46, 26, 5, 61, 33, 14, 10, 25, 
    95, 46, 65, 12, 0, 44, 79, 37, 20, 7, 41, 31, 13, 26, 8, 
    90, 68, 83, 18, 52, 26, 22, 16, 16, 19, 16, 28, 2, 0, 3, 
    59, 67, 64, 17, 61, 48, 22, 25, 59, 34, 22, 0, 0, 1, 10, 
    28, 70, 60, 23, 74, 70, 65, 74, 65, 23, 12, 21, 38, 40, 41, 
    57, 59, 62, 53, 113, 62, 38, 40, 38, 33, 36, 37, 39, 44, 47, 
    58, 55, 58, 90, 81, 38, 39, 35, 31, 33, 35, 45, 51, 48, 48, 
    55, 47, 72, 67, 43, 39, 40, 38, 36, 41, 45, 46, 43, 51, 68, 
    61, 43, 50, 29, 35, 34, 39, 38, 36, 41, 46, 38, 37, 64, 53, 
    
    -- channel=21
    16, 16, 13, 13, 11, 12, 17, 18, 10, 9, 12, 15, 12, 11, 10, 
    10, 16, 14, 13, 12, 0, 2, 10, 15, 0, 0, 0, 10, 15, 10, 
    9, 27, 17, 15, 16, 32, 11, 9, 0, 0, 0, 0, 0, 6, 13, 
    0, 0, 13, 12, 4, 3, 0, 0, 0, 8, 0, 0, 0, 0, 13, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 16, 43, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 19, 11, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 7, 4, 6, 0, 0, 0, 3, 6, 
    0, 0, 0, 0, 0, 22, 7, 0, 0, 0, 23, 9, 9, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 6, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 2, 0, 0, 3, 13, 4, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=22
    31, 37, 32, 30, 28, 34, 32, 32, 27, 27, 31, 33, 33, 24, 21, 
    25, 33, 32, 32, 34, 39, 22, 31, 41, 35, 17, 10, 20, 31, 21, 
    21, 49, 32, 33, 30, 51, 48, 25, 16, 37, 31, 29, 7, 9, 33, 
    3, 2, 27, 33, 26, 39, 25, 14, 16, 42, 44, 29, 28, 0, 26, 
    44, 18, 27, 49, 52, 33, 47, 24, 14, 42, 41, 18, 17, 4, 0, 
    54, 63, 40, 41, 114, 94, 64, 28, 1, 42, 55, 39, 24, 18, 1, 
    59, 51, 50, 32, 47, 69, 72, 51, 22, 50, 61, 24, 19, 28, 12, 
    69, 70, 16, 30, 31, 70, 66, 56, 40, 44, 65, 27, 27, 31, 31, 
    80, 79, 39, 57, 25, 66, 48, 26, 32, 26, 43, 34, 23, 33, 21, 
    95, 79, 51, 52, 36, 26, 54, 41, 11, 48, 30, 12, 9, 21, 30, 
    88, 77, 55, 68, 60, 10, 52, 82, 45, 14, 0, 3, 9, 30, 30, 
    51, 98, 71, 78, 95, 74, 47, 47, 34, 21, 18, 22, 25, 20, 23, 
    10, 43, 93, 86, 72, 25, 20, 19, 15, 13, 16, 16, 23, 33, 28, 
    20, 18, 53, 96, 39, 22, 19, 16, 22, 20, 21, 28, 27, 22, 30, 
    20, 22, 26, 42, 16, 23, 30, 26, 22, 22, 16, 21, 28, 20, 16, 
    
    -- channel=23
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 11, 7, 12, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 
    9, 3, 10, 0, 29, 11, 11, 15, 9, 2, 6, 19, 18, 6, 0, 
    40, 20, 21, 14, 18, 9, 20, 19, 24, 32, 41, 45, 50, 51, 48, 
    62, 32, 6, 7, 13, 39, 43, 39, 40, 44, 52, 52, 55, 56, 60, 
    66, 55, 18, 27, 26, 44, 44, 41, 44, 48, 54, 56, 59, 55, 67, 
    66, 61, 46, 41, 35, 36, 42, 44, 47, 51, 53, 54, 60, 71, 70, 
    
    -- channel=24
    72, 76, 76, 77, 75, 76, 75, 76, 74, 63, 54, 57, 63, 63, 61, 
    75, 74, 76, 77, 79, 123, 72, 66, 40, 66, 68, 51, 47, 57, 64, 
    53, 56, 77, 77, 78, 74, 61, 37, 47, 88, 79, 68, 51, 38, 65, 
    51, 83, 75, 80, 77, 73, 86, 57, 57, 74, 78, 57, 48, 35, 52, 
    82, 117, 73, 89, 142, 99, 82, 61, 43, 78, 96, 61, 61, 43, 31, 
    81, 124, 80, 71, 115, 92, 114, 71, 52, 121, 94, 53, 60, 54, 44, 
    90, 110, 68, 57, 82, 126, 114, 90, 56, 119, 85, 64, 61, 75, 61, 
    111, 112, 72, 71, 77, 127, 77, 71, 62, 104, 93, 60, 61, 66, 64, 
    124, 125, 78, 100, 78, 60, 74, 81, 78, 66, 72, 29, 43, 73, 81, 
    130, 127, 88, 101, 74, 54, 88, 110, 69, 54, 27, 23, 59, 79, 67, 
    133, 122, 83, 160, 154, 99, 108, 92, 60, 39, 50, 60, 61, 66, 60, 
    76, 113, 106, 183, 101, 56, 56, 53, 56, 53, 60, 62, 72, 74, 68, 
    68, 74, 125, 150, 51, 63, 57, 57, 58, 62, 69, 76, 70, 68, 90, 
    67, 63, 92, 102, 64, 66, 65, 58, 59, 65, 67, 67, 66, 87, 65, 
    67, 66, 66, 53, 49, 55, 57, 61, 71, 78, 66, 66, 98, 95, 56, 
    
    -- channel=25
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=26
    57, 58, 60, 60, 61, 53, 63, 64, 61, 49, 38, 41, 47, 55, 56, 
    60, 61, 63, 62, 59, 60, 60, 53, 35, 23, 23, 25, 26, 39, 53, 
    42, 34, 61, 63, 63, 31, 36, 19, 21, 11, 13, 12, 23, 21, 41, 
    29, 33, 59, 59, 59, 29, 33, 20, 15, 2, 19, 15, 14, 22, 25, 
    8, 25, 57, 33, 37, 31, 20, 22, 15, 5, 18, 25, 17, 21, 23, 
    0, 5, 52, 47, 0, 8, 27, 21, 26, 9, 14, 11, 10, 14, 23, 
    0, 12, 28, 55, 12, 20, 11, 17, 18, 2, 9, 16, 12, 12, 23, 
    1, 3, 18, 37, 20, 9, 6, 7, 15, 16, 13, 14, 7, 13, 29, 
    0, 0, 11, 11, 29, 0, 15, 23, 10, 28, 11, 7, 10, 30, 56, 
    0, 0, 10, 0, 12, 13, 5, 21, 16, 13, 7, 6, 14, 42, 46, 
    0, 0, 4, 0, 26, 19, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=27
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=28
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 
    0, 0, 0, 0, 0, 0, 20, 0, 14, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 36, 8, 0, 0, 13, 12, 34, 0, 0, 
    78, 0, 0, 0, 3, 0, 3, 16, 3, 0, 42, 0, 30, 21, 0, 
    89, 0, 35, 0, 0, 0, 35, 29, 12, 0, 9, 49, 0, 38, 0, 
    49, 0, 50, 0, 0, 16, 39, 33, 48, 0, 44, 58, 0, 20, 21, 
    52, 17, 10, 42, 0, 0, 8, 31, 61, 0, 69, 35, 0, 0, 21, 
    34, 27, 27, 22, 0, 0, 55, 4, 35, 0, 42, 41, 0, 0, 17, 
    36, 0, 79, 0, 0, 0, 24, 0, 0, 10, 0, 47, 0, 0, 0, 
    0, 0, 94, 0, 42, 0, 0, 17, 0, 4, 45, 5, 0, 0, 7, 
    0, 0, 81, 0, 101, 22, 0, 8, 64, 26, 0, 0, 0, 0, 0, 
    0, 0, 36, 0, 89, 51, 0, 0, 11, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 106, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 0, 0, 56, 28, 0, 9, 0, 0, 0, 0, 0, 2, 0, 2, 
    24, 0, 0, 0, 3, 0, 0, 0, 0, 0, 5, 0, 0, 4, 52, 
    
    -- channel=29
    55, 58, 57, 57, 57, 53, 59, 64, 57, 46, 42, 47, 49, 48, 49, 
    56, 58, 60, 58, 59, 51, 44, 47, 42, 33, 11, 14, 31, 45, 48, 
    36, 61, 60, 61, 60, 68, 41, 30, 14, 23, 9, 13, 2, 21, 47, 
    5, 29, 52, 59, 48, 45, 21, 7, 8, 27, 20, 15, 15, 1, 40, 
    4, 14, 40, 51, 27, 11, 21, 11, 10, 26, 20, 3, 14, 2, 12, 
    2, 28, 40, 35, 62, 34, 26, 16, 3, 26, 15, 14, 17, 7, 0, 
    2, 14, 41, 44, 44, 33, 31, 20, 9, 31, 18, 8, 13, 13, 7, 
    2, 24, 1, 35, 27, 32, 25, 26, 23, 37, 24, 12, 15, 20, 36, 
    7, 20, 0, 27, 11, 39, 30, 15, 22, 29, 29, 20, 21, 33, 35, 
    32, 22, 3, 21, 5, 11, 30, 15, 3, 24, 15, 7, 13, 36, 46, 
    35, 21, 13, 29, 0, 0, 0, 17, 0, 1, 0, 0, 0, 3, 0, 
    5, 24, 15, 29, 13, 9, 4, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 26, 22, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=30
    30, 34, 28, 33, 28, 29, 29, 32, 29, 25, 23, 22, 24, 25, 27, 
    24, 29, 27, 32, 29, 35, 25, 25, 20, 17, 11, 8, 11, 18, 25, 
    30, 21, 31, 33, 28, 42, 46, 23, 10, 9, 38, 32, 13, 0, 20, 
    39, 0, 26, 27, 30, 21, 28, 20, 16, 3, 54, 22, 35, 9, 0, 
    55, 1, 35, 4, 42, 12, 52, 38, 25, 0, 37, 31, 20, 20, 0, 
    54, 48, 51, 24, 64, 59, 68, 38, 32, 0, 64, 53, 18, 24, 6, 
    56, 49, 35, 52, 7, 32, 61, 51, 46, 0, 69, 38, 14, 18, 27, 
    55, 67, 8, 34, 0, 34, 85, 45, 54, 12, 62, 45, 13, 28, 38, 
    71, 54, 60, 25, 27, 34, 46, 31, 14, 18, 38, 51, 15, 26, 18, 
    80, 57, 78, 3, 48, 18, 21, 42, 19, 46, 38, 5, 0, 3, 27, 
    41, 54, 76, 10, 69, 17, 12, 64, 52, 15, 1, 0, 0, 6, 14, 
    15, 54, 59, 17, 101, 74, 31, 34, 32, 17, 15, 16, 22, 17, 25, 
    18, 10, 32, 75, 107, 22, 18, 17, 16, 13, 13, 17, 20, 23, 25, 
    32, 10, 0, 115, 47, 18, 22, 16, 15, 17, 19, 26, 25, 19, 33, 
    35, 19, 8, 46, 24, 19, 26, 25, 15, 22, 23, 19, 13, 34, 33, 
    
    -- channel=31
    55, 53, 55, 53, 54, 51, 57, 59, 53, 46, 43, 48, 47, 47, 47, 
    55, 55, 57, 53, 56, 49, 38, 47, 35, 30, 11, 21, 39, 49, 48, 
    38, 64, 59, 55, 60, 57, 22, 22, 25, 35, 2, 5, 1, 38, 50, 
    0, 61, 50, 58, 42, 41, 16, 8, 13, 45, 0, 17, 4, 11, 59, 
    0, 29, 30, 58, 10, 12, 0, 1, 11, 50, 5, 0, 16, 0, 41, 
    0, 16, 22, 50, 45, 10, 0, 0, 0, 76, 0, 0, 21, 4, 6, 
    0, 0, 32, 27, 56, 36, 4, 0, 0, 67, 0, 0, 17, 16, 7, 
    0, 0, 1, 19, 42, 40, 0, 14, 5, 58, 0, 0, 22, 24, 25, 
    0, 0, 0, 21, 20, 24, 7, 12, 24, 22, 28, 1, 32, 34, 45, 
    1, 2, 0, 27, 0, 23, 27, 0, 13, 18, 1, 12, 31, 52, 41, 
    29, 3, 0, 53, 0, 0, 22, 0, 0, 0, 1, 0, 0, 10, 0, 
    22, 12, 0, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 20, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end ifmap_package;
