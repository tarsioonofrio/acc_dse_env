LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
	PACKAGE gold_package is
		type padroes is array(0 to 4000000) of integer;
		constant gold: padroes := ( 0, 
		
		240, 
		
		0, 
		
		0, 
		
		0, 
		
		0, 
		
		188, 
		
		140, 
		
		0, 
		
		0, 
		
		181, 
		
		0, 
		
		468, 
		
		0, 
		
		185, 
		
		0, 
		
		334, 
		
		13, 
		
		272, 
		
		0, 
		
		0, 
		
		311, 
		
		0, 
		
		164, 
		
		0, 
		
		0, 
		
		0, 
		
		234, 
		
		0, 
		
		0, 
		
		0, 
		
		0, 
		
		0, 
		
		0, 
		
		0, 
		
		0, 
		
		98, 
		
		0, 
		
		278, 
		
		0, 
		
		0, 
		
		218, 
		
		0, 
		
		608, 
		
		206, 
		
		0, 
		
		0, 
		
		0, 
		
		0, 
		
		0, 
		
		0, 
		
		0, 
		
		0, 
		
		0, 
		
		386, 
		
		0, 
		
		0, 
		
		0, 
		
		0, 
		
		10, 
		
		0, 
		
		224, 
		
		0, 
		
		0, 
		
		0, 
		
		0, 
		
		181, 
		
		0, 
		
		89, 
		
		362, 
		
		0, 
		
		53, 
		
		0, 
		
		39, 
		
		0, 
		
		118, 
		
		0, 
		
		3, 
		
		0, 
		
		0, 
		
		0, 
		
		179, 
		
		0, 
		
		248, 
		
		0, 
		
		0, 
		
		130, 
		
		0, 
		
		0, 
		
		0, 
		
		69, 
		
		0, 
		
		0, 
		
		0, 
		
		0, 
		
		353, 
		
		0, 
		
		105, 
		
		166, 
		
		0, 
		
		0, 
		
		0, 
		
		0, 
		
		0, 
		
		124, 
		
		340, 
		
		0, 
		
		0, 
		
		0, 
		
		0, 
		
		0, 
		
		0, 
		
		0, 
		
		0, 
		
		146, 
		
		145, 
		
		0, 
		
		0, 
		
		0, 
		
		0, 
		
		240, 
		
		0, 
		
		0, 
		
		0, 
		
		123, 
		
		0, 
		
		258, 
		
		256, 
		
		others=>0 );
END gold_package;
