library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 4000000) of integer;

  constant input_wght : mem := (
    -- bias
    -9328, -16224, 26112, -8563, -3485, -5337, 114, -587, -6114, 18302, -20091, 11361, -20330, -17242, -9964, -1451,

    -- weights
    -- filter=0 channel=0
    -32, -35, -38, 29, -49, 1, 35, -35, -12,
    -- filter=0 channel=1
    -9, 0, 35, -26, 15, -36, -8, 41, -21,
    -- filter=0 channel=2
    11, 40, 15, 14, -21, -38, -31, 46, 11,
    -- filter=1 channel=0
    -18, -18, -24, -10, -57, -44, -22, -24, 28,
    -- filter=1 channel=1
    7, 14, -6, -10, -11, 28, -36, 2, 16,
    -- filter=1 channel=2
    -11, 22, 28, 80, 65, -25, 72, 85, -7,
    -- filter=2 channel=0
    29, 0, 2, -45, 66, 71, -53, -27, 59,
    -- filter=2 channel=1
    56, 112, 60, -25, 100, 107, 22, 0, 68,
    -- filter=2 channel=2
    -89, -65, -4, -115, -48, 2, -111, -86, -36,
    -- filter=3 channel=0
    17, -38, -19, 47, 25, -36, -41, 34, 25,
    -- filter=3 channel=1
    0, -49, -47, -25, 0, -12, 37, 19, 20,
    -- filter=3 channel=2
    -24, -35, -37, -28, -4, -40, 0, -40, 41,
    -- filter=4 channel=0
    114, 38, -24, 148, 27, -43, 103, 73, 10,
    -- filter=4 channel=1
    -8, -92, -145, -17, -21, -131, 70, 35, -14,
    -- filter=4 channel=2
    26, 3, -94, -13, 25, -98, 60, -3, 16,
    -- filter=5 channel=0
    -26, 5, -14, 16, -10, 9, 5, 43, 33,
    -- filter=5 channel=1
    -53, -58, 25, 18, 37, 38, -40, 11, 45,
    -- filter=5 channel=2
    -47, -6, 0, 0, 3, 28, -50, 2, 45,
    -- filter=6 channel=0
    -12, -7, -22, 27, -39, 2, -47, 16, -5,
    -- filter=6 channel=1
    -38, -1, -43, 41, 41, -26, -40, -13, 3,
    -- filter=6 channel=2
    -10, 28, 44, -44, -3, -33, 33, -16, -23,
    -- filter=7 channel=0
    34, -29, 27, -1, -18, 12, 15, -3, -27,
    -- filter=7 channel=1
    -23, -41, -31, 35, 5, 18, 31, 30, 33,
    -- filter=7 channel=2
    26, 40, -40, -17, -45, -23, -43, -30, 13,
    -- filter=8 channel=0
    20, -44, -53, -15, -50, -42, 33, 32, -78,
    -- filter=8 channel=1
    15, -8, -26, 48, 69, 29, 49, 48, -31,
    -- filter=8 channel=2
    67, -12, 41, 32, 77, -3, 10, 56, 49,
    -- filter=9 channel=0
    -66, -100, -40, -17, -96, -90, -60, 13, -63,
    -- filter=9 channel=1
    -66, -60, -34, -12, -14, 2, 52, 23, 44,
    -- filter=9 channel=2
    -9, 49, 87, 9, 105, 31, 100, 128, 110,
    -- filter=10 channel=0
    -41, -21, -18, -5, -17, -41, -73, 7, -58,
    -- filter=10 channel=1
    -68, 30, -54, -3, -5, -29, -9, 41, -21,
    -- filter=10 channel=2
    75, 69, 80, 60, 95, 38, 28, 85, 68,
    -- filter=11 channel=0
    -28, -72, -77, -37, 12, -2, 36, 18, -37,
    -- filter=11 channel=1
    57, 25, 3, 90, 88, 60, 126, 111, 77,
    -- filter=11 channel=2
    -44, -39, -92, -17, -61, -45, 55, -8, -55,
    -- filter=12 channel=0
    -57, 44, -8, 10, 83, 37, -28, 56, 17,
    -- filter=12 channel=1
    10, -34, 26, 71, 66, 26, 28, 33, -8,
    -- filter=12 channel=2
    -25, 9, -52, 34, 77, 16, 26, 15, 46,
    -- filter=13 channel=0
    -17, 31, 28, -18, 77, 78, -25, 42, 87,
    -- filter=13 channel=1
    -56, -36, -14, 8, -25, 8, -62, 14, 36,
    -- filter=13 channel=2
    -41, 37, 34, 64, 75, 78, -1, 52, 28,
    -- filter=14 channel=0
    49, 70, 2, 14, 33, 62, 10, -30, 23,
    -- filter=14 channel=1
    -1, 15, 81, -5, 25, 75, -17, -4, 53,
    -- filter=14 channel=2
    -41, 18, -1, -35, 34, -34, -10, -62, -40,
    -- filter=15 channel=0
    56, 79, 85, 31, 51, 39, -2, 37, 13,
    -- filter=15 channel=1
    -61, 12, -43, -67, -56, 21, 10, -73, -3,
    -- filter=15 channel=2
    33, 35, -45, -36, 9, 39, -34, 36, -8,

    others => 0);
end iwght_package;
