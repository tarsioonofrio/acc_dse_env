library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    29, 34, 33, 34, 34, 29, 30, 27, 
    4, 19, 32, 6, 27, 0, 22, 19, 
    0, 52, 0, 0, 14, 0, 0, 28, 
    0, 17, 21, 0, 13, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=1
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 
    22, 0, 0, 0, 0, 0, 0, 0, 
    23, 0, 0, 0, 0, 0, 0, 0, 
    22, 1, 3, 0, 0, 0, 6, 0, 
    
    -- channel=2
    89, 110, 240, 245, 154, 270, 122, 0, 
    384, 307, 519, 472, 421, 615, 314, 0, 
    1060, 795, 1031, 1021, 676, 852, 410, 63, 
    1322, 978, 1009, 1146, 794, 957, 453, 243, 
    1575, 1390, 1052, 926, 808, 517, 383, 305, 
    1548, 1771, 1794, 1114, 909, 847, 1041, 971, 
    1368, 1752, 1682, 953, 993, 1140, 1332, 1260, 
    1141, 1140, 970, 857, 1029, 1126, 1356, 1220, 
    
    -- channel=3
    79, 54, 67, 60, 61, 57, 48, 59, 
    89, 45, 92, 22, 99, 44, 14, 54, 
    150, 59, 86, 48, 111, 64, 27, 51, 
    178, 49, 103, 54, 109, 19, 39, 31, 
    186, 59, 56, 51, 47, 21, 71, 55, 
    179, 136, 20, 37, 26, 62, 52, 41, 
    163, 111, 30, 69, 77, 84, 98, 100, 
    161, 83, 72, 57, 74, 75, 91, 54, 
    
    -- channel=4
    561, 575, 606, 559, 528, 399, 473, 484, 
    539, 612, 643, 573, 457, 415, 410, 483, 
    483, 676, 682, 515, 462, 422, 328, 360, 
    501, 660, 713, 631, 565, 541, 380, 419, 
    487, 462, 660, 662, 580, 537, 444, 504, 
    531, 598, 487, 402, 345, 208, 227, 302, 
    369, 644, 501, 202, 90, 0, 0, 31, 
    59, 345, 238, 87, 94, 90, 125, 82, 
    
    -- channel=5
    66, 0, 17, 0, 37, 21, 0, 0, 
    108, 11, 48, 0, 102, 59, 0, 0, 
    241, 0, 127, 0, 104, 81, 0, 0, 
    303, 0, 130, 29, 112, 44, 35, 0, 
    337, 0, 82, 24, 38, 6, 52, 0, 
    326, 191, 28, 87, 25, 115, 119, 70, 
    289, 253, 0, 96, 130, 137, 164, 128, 
    204, 206, 103, 122, 140, 150, 192, 67, 
    
    -- channel=6
    31, 27, 7, 97, 29, 74, 60, 154, 
    63, 55, 71, 160, 74, 177, 125, 152, 
    157, 253, 175, 248, 178, 249, 130, 157, 
    217, 290, 35, 263, 201, 260, 119, 207, 
    245, 319, 192, 156, 218, 166, 58, 227, 
    199, 270, 414, 193, 228, 119, 122, 380, 
    155, 184, 418, 212, 176, 198, 217, 453, 
    207, 186, 295, 159, 162, 209, 230, 429, 
    
    -- channel=7
    54, 54, 123, 139, 90, 157, 93, 21, 
    210, 145, 250, 244, 256, 404, 221, 19, 
    639, 445, 553, 545, 382, 515, 256, 116, 
    821, 573, 542, 625, 456, 570, 279, 182, 
    958, 809, 651, 566, 489, 331, 262, 233, 
    985, 1034, 1122, 778, 682, 693, 783, 782, 
    986, 1140, 1106, 778, 838, 936, 1078, 1089, 
    989, 936, 818, 755, 873, 930, 1121, 1078, 
    
    -- channel=8
    352, 397, 427, 427, 356, 319, 324, 312, 
    335, 452, 474, 423, 325, 312, 294, 300, 
    385, 487, 495, 456, 388, 359, 284, 255, 
    397, 498, 502, 513, 434, 374, 304, 310, 
    384, 471, 464, 456, 437, 362, 306, 365, 
    407, 535, 474, 397, 358, 210, 237, 279, 
    260, 521, 432, 204, 110, 56, 82, 88, 
    93, 239, 213, 72, 77, 94, 108, 109, 
    
    -- channel=9
    17, 2, 73, 61, 46, 90, 7, 0, 
    101, 72, 199, 173, 177, 311, 122, 0, 
    451, 299, 463, 424, 295, 399, 152, 0, 
    588, 392, 504, 510, 352, 465, 182, 84, 
    762, 596, 457, 424, 320, 257, 155, 101, 
    773, 782, 825, 519, 434, 393, 490, 447, 
    692, 840, 815, 493, 501, 571, 668, 631, 
    621, 614, 519, 450, 531, 571, 699, 622, 
    
    -- channel=10
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 40, 0, 145, 83, 0, 
    213, 167, 172, 174, 67, 169, 101, 33, 
    288, 228, 107, 238, 119, 207, 103, 66, 
    379, 258, 130, 181, 128, 133, 78, 43, 
    355, 254, 418, 315, 303, 163, 222, 230, 
    357, 344, 486, 325, 270, 308, 341, 395, 
    370, 346, 411, 280, 275, 313, 373, 429, 
    
    -- channel=11
    66, 67, 68, 57, 65, 46, 56, 41, 
    15, 13, 18, 7, 3, 0, 10, 0, 
    22, 29, 16, 0, 23, 0, 0, 1, 
    0, 5, 3, 0, 21, 0, 0, 0, 
    0, 13, 0, 0, 0, 7, 25, 3, 
    46, 19, 21, 23, 42, 32, 36, 23, 
    43, 14, 6, 8, 8, 15, 18, 8, 
    20, 8, 17, 18, 32, 40, 37, 44, 
    
    -- channel=12
    373, 395, 428, 436, 337, 316, 297, 317, 
    364, 446, 467, 429, 299, 344, 280, 288, 
    414, 479, 516, 495, 338, 387, 272, 219, 
    441, 467, 491, 516, 354, 411, 268, 309, 
    475, 454, 444, 456, 381, 360, 280, 342, 
    451, 478, 550, 353, 318, 184, 209, 249, 
    231, 493, 490, 136, 79, 45, 72, 146, 
    45, 224, 155, 50, 64, 69, 101, 127, 
    
    -- channel=13
    68, 54, 91, 82, 41, 106, 43, 25, 
    144, 104, 140, 156, 144, 222, 127, 2, 
    378, 254, 323, 350, 215, 290, 163, 80, 
    486, 360, 314, 367, 242, 325, 169, 136, 
    563, 495, 403, 358, 275, 152, 158, 140, 
    543, 607, 622, 418, 410, 418, 463, 491, 
    542, 602, 575, 448, 479, 534, 625, 620, 
    516, 468, 462, 418, 487, 519, 619, 590, 
    
    -- channel=14
    590, 603, 688, 630, 518, 488, 470, 514, 
    562, 675, 717, 602, 525, 502, 403, 494, 
    566, 725, 776, 627, 579, 559, 363, 363, 
    576, 656, 768, 705, 585, 560, 407, 454, 
    593, 540, 636, 597, 549, 520, 447, 528, 
    587, 750, 652, 533, 351, 240, 278, 357, 
    332, 715, 471, 144, 66, 28, 52, 103, 
    54, 253, 122, 35, 56, 46, 99, 69, 
    
    -- channel=15
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 
    25, 0, 0, 0, 0, 0, 0, 0, 
    18, 33, 11, 10, 12, 26, 22, 16, 
    
    -- channel=16
    223, 134, 195, 151, 165, 166, 109, 101, 
    322, 210, 291, 167, 265, 224, 105, 112, 
    452, 239, 337, 258, 333, 285, 104, 106, 
    528, 187, 367, 265, 342, 268, 155, 116, 
    571, 308, 323, 280, 228, 148, 204, 171, 
    558, 525, 365, 295, 170, 215, 243, 248, 
    454, 510, 280, 177, 208, 224, 276, 263, 
    355, 330, 107, 162, 227, 239, 294, 214, 
    
    -- channel=17
    236, 206, 228, 359, 199, 291, 236, 304, 
    383, 321, 387, 443, 180, 454, 353, 312, 
    631, 608, 563, 632, 411, 571, 359, 292, 
    771, 756, 388, 667, 419, 581, 329, 392, 
    827, 769, 569, 539, 567, 394, 243, 464, 
    745, 722, 963, 515, 617, 399, 460, 726, 
    538, 649, 1011, 514, 480, 504, 590, 880, 
    534, 569, 701, 436, 477, 528, 641, 821, 
    
    -- channel=18
    107, 97, 101, 115, 86, 76, 88, 88, 
    91, 92, 84, 68, 50, 74, 69, 82, 
    107, 124, 84, 79, 29, 90, 59, 85, 
    81, 106, 63, 84, 60, 89, 77, 106, 
    100, 63, 78, 31, 84, 65, 75, 104, 
    86, 55, 94, 44, 59, 1, 15, 69, 
    53, 45, 61, 10, 5, 11, 5, 95, 
    83, 25, 24, 27, 36, 37, 48, 64, 
    
    -- channel=19
    407, 229, 318, 113, 268, 143, 189, 229, 
    421, 344, 316, 112, 356, 149, 144, 267, 
    545, 377, 404, 69, 407, 176, 101, 172, 
    593, 169, 495, 68, 342, 114, 177, 140, 
    651, 161, 215, 241, 159, 126, 257, 198, 
    665, 277, 0, 54, 0, 123, 126, 70, 
    446, 350, 0, 12, 38, 48, 58, 48, 
    329, 104, 31, 37, 68, 58, 122, 0, 
    
    -- channel=20
    45, 16, 60, 56, 48, 99, 47, 0, 
    138, 79, 92, 91, 120, 212, 79, 22, 
    315, 200, 256, 225, 203, 275, 107, 69, 
    372, 233, 259, 289, 206, 284, 136, 92, 
    455, 332, 303, 272, 224, 135, 143, 115, 
    486, 482, 499, 350, 327, 372, 391, 392, 
    490, 522, 482, 373, 410, 441, 528, 509, 
    495, 443, 374, 381, 434, 439, 546, 486, 
    
    -- channel=21
    0, 0, 0, 0, 0, 0, 0, 0, 
    32, 0, 0, 18, 58, 160, 53, 0, 
    280, 127, 218, 238, 134, 231, 79, 0, 
    411, 229, 205, 274, 181, 258, 87, 50, 
    531, 426, 283, 267, 195, 57, 43, 11, 
    532, 564, 609, 385, 362, 437, 475, 487, 
    541, 577, 575, 493, 544, 604, 686, 702, 
    599, 510, 437, 477, 569, 595, 727, 680, 
    
    -- channel=22
    107, 115, 130, 151, 116, 109, 116, 126, 
    116, 123, 153, 177, 98, 133, 126, 127, 
    122, 184, 165, 151, 75, 149, 112, 131, 
    141, 201, 169, 192, 128, 166, 106, 126, 
    117, 133, 161, 173, 168, 182, 85, 153, 
    116, 110, 205, 115, 126, 58, 53, 138, 
    55, 158, 220, 43, 20, 0, 0, 121, 
    50, 121, 115, 49, 64, 56, 74, 105, 
    
    -- channel=23
    621, 678, 736, 677, 619, 493, 512, 508, 
    601, 716, 789, 693, 557, 552, 447, 486, 
    634, 898, 946, 784, 584, 568, 439, 294, 
    647, 830, 987, 924, 787, 730, 509, 483, 
    756, 727, 845, 882, 709, 704, 526, 569, 
    786, 968, 779, 630, 495, 233, 288, 339, 
    526, 985, 770, 308, 119, 29, 47, 30, 
    85, 443, 337, 141, 184, 201, 252, 147, 
    
    -- channel=24
    94, 81, 133, 131, 57, 132, 44, 6, 
    213, 148, 227, 244, 228, 368, 169, 0, 
    632, 445, 611, 583, 346, 510, 242, 30, 
    809, 577, 569, 659, 423, 549, 245, 156, 
    992, 830, 610, 551, 454, 260, 222, 166, 
    980, 1024, 1083, 658, 587, 587, 666, 648, 
    870, 1027, 1001, 650, 702, 798, 919, 890, 
    787, 740, 693, 612, 715, 770, 931, 855, 
    
    -- channel=25
    0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 2, 1, 
    0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=26
    24, 13, 26, 89, 22, 97, 64, 67, 
    149, 52, 142, 157, 119, 286, 193, 35, 
    478, 357, 340, 406, 255, 358, 224, 137, 
    611, 480, 284, 440, 303, 378, 231, 142, 
    668, 569, 417, 351, 391, 221, 160, 162, 
    652, 666, 766, 585, 498, 409, 486, 515, 
    660, 726, 850, 557, 532, 603, 689, 766, 
    709, 668, 607, 507, 565, 619, 743, 821, 
    
    -- channel=27
    48, 47, 54, 40, 48, 11, 35, 37, 
    60, 51, 50, 19, 19, 0, 31, 43, 
    0, 58, 51, 0, 17, 0, 0, 16, 
    0, 22, 66, 2, 8, 0, 12, 8, 
    0, 0, 26, 33, 0, 17, 32, 35, 
    23, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=28
    22, 12, 14, 61, 17, 55, 43, 81, 
    54, 18, 7, 64, 0, 71, 77, 86, 
    73, 115, 41, 111, 4, 99, 66, 74, 
    57, 126, 0, 100, 15, 105, 22, 108, 
    47, 99, 75, 63, 98, 45, 14, 131, 
    2, 0, 125, 29, 120, 42, 32, 181, 
    0, 0, 133, 7, 10, 0, 0, 177, 
    0, 0, 54, 0, 0, 6, 10, 158, 
    
    -- channel=29
    0, 0, 0, 0, 0, 0, 0, 22, 
    0, 0, 0, 0, 0, 0, 0, 21, 
    0, 0, 0, 0, 0, 0, 0, 22, 
    0, 0, 0, 0, 0, 0, 0, 24, 
    0, 0, 0, 0, 0, 0, 0, 17, 
    0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=30
    20, 26, 28, 48, 50, 52, 52, 49, 
    65, 56, 35, 80, 83, 48, 71, 53, 
    24, 83, 22, 60, 118, 67, 80, 84, 
    23, 100, 38, 59, 105, 84, 89, 57, 
    22, 99, 88, 81, 59, 98, 84, 52, 
    13, 88, 135, 97, 143, 126, 87, 118, 
    93, 34, 200, 133, 118, 98, 109, 112, 
    102, 66, 154, 95, 86, 114, 87, 127, 
    
    -- channel=31
    4, 0, 0, 2, 0, 0, 0, 0, 
    18, 25, 1, 12, 9, 6, 0, 0, 
    40, 26, 33, 9, 7, 20, 0, 0, 
    6, 0, 0, 0, 4, 0, 0, 10, 
    12, 0, 24, 12, 11, 0, 0, 0, 
    0, 0, 50, 0, 0, 5, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end gold_package;
