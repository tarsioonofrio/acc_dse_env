library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    118, 367, 0, 
    50, 0, 0, 
    158, 305, 176, 
    
    -- channel=1
    0, 412, 0, 
    14, 177, 193, 
    0, 74, 169, 
    
    -- channel=2
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=3
    0, 0, 297, 
    0, 0, 0, 
    0, 149, 0, 
    
    -- channel=4
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=5
    0, 0, 0, 
    0, 0, 0, 
    42, 0, 0, 
    
    -- channel=6
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=7
    0, 0, 0, 
    0, 5, 138, 
    67, 0, 20, 
    
    -- channel=8
    0, 276, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=9
    0, 27, 0, 
    0, 90, 0, 
    0, 0, 0, 
    
    -- channel=10
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=11
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=12
    0, 381, 239, 
    61, 326, 106, 
    0, 0, 0, 
    
    -- channel=13
    0, 0, 0, 
    0, 98, 238, 
    121, 133, 82, 
    
    -- channel=14
    0, 0, 0, 
    0, 0, 99, 
    0, 5, 144, 
    
    -- channel=15
    0, 57, 0, 
    0, 0, 0, 
    433, 0, 361, 
    
    -- channel=16
    198, 0, 344, 
    0, 0, 99, 
    0, 0, 0, 
    
    -- channel=17
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=18
    0, 0, 60, 
    0, 0, 0, 
    0, 83, 148, 
    
    -- channel=19
    0, 0, 0, 
    0, 0, 0, 
    499, 0, 23, 
    
    -- channel=20
    0, 0, 0, 
    0, 0, 0, 
    0, 296, 270, 
    
    -- channel=21
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=22
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=23
    0, 0, 0, 
    0, 0, 97, 
    0, 197, 0, 
    
    -- channel=24
    0, 0, 219, 
    183, 341, 0, 
    194, 0, 216, 
    
    -- channel=25
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 21, 
    
    -- channel=26
    30, 0, 0, 
    0, 0, 0, 
    0, 0, 80, 
    
    -- channel=27
    36, 0, 0, 
    0, 94, 0, 
    0, 435, 179, 
    
    -- channel=28
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=29
    187, 264, 262, 
    249, 0, 0, 
    0, 0, 0, 
    
    -- channel=30
    0, 50, 53, 
    520, 86, 5, 
    0, 0, 0, 
    
    -- channel=31
    0, 0, 0, 
    16, 0, 92, 
    0, 0, 0, 
    
    -- channel=32
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=33
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=34
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=35
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=36
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=37
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=38
    201, 354, 50, 
    252, 107, 0, 
    0, 0, 0, 
    
    -- channel=39
    24, 0, 0, 
    0, 0, 0, 
    352, 578, 539, 
    
    -- channel=40
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=41
    0, 39, 408, 
    0, 0, 0, 
    194, 421, 355, 
    
    -- channel=42
    0, 217, 0, 
    418, 130, 13, 
    265, 0, 0, 
    
    -- channel=43
    0, 0, 27, 
    142, 0, 33, 
    0, 0, 0, 
    
    -- channel=44
    0, 222, 0, 
    0, 0, 0, 
    559, 505, 0, 
    
    -- channel=45
    0, 0, 0, 
    0, 0, 0, 
    545, 0, 0, 
    
    -- channel=46
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=47
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=48
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=49
    0, 0, 0, 
    0, 0, 0, 
    0, 62, 0, 
    
    -- channel=50
    0, 98, 199, 
    271, 40, 0, 
    0, 0, 0, 
    
    -- channel=51
    0, 199, 0, 
    285, 215, 249, 
    0, 0, 0, 
    
    -- channel=52
    121, 16, 190, 
    0, 184, 47, 
    0, 0, 0, 
    
    -- channel=53
    22, 0, 0, 
    0, 0, 0, 
    0, 24, 0, 
    
    -- channel=54
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=55
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=56
    294, 0, 373, 
    272, 0, 131, 
    126, 0, 0, 
    
    -- channel=57
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=58
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=59
    0, 0, 0, 
    485, 166, 0, 
    190, 0, 0, 
    
    -- channel=60
    0, 0, 0, 
    0, 0, 0, 
    0, 41, 77, 
    
    -- channel=61
    0, 16, 0, 
    54, 388, 325, 
    50, 329, 411, 
    
    -- channel=62
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=63
    16, 258, 0, 
    0, 0, 247, 
    0, 0, 0, 
    
    -- channel=64
    0, 53, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=65
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=66
    0, 0, 0, 
    0, 0, 0, 
    0, 12, 60, 
    
    -- channel=67
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=68
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=69
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=70
    40, 0, 0, 
    325, 0, 94, 
    0, 0, 0, 
    
    -- channel=71
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=72
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=73
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=74
    0, 0, 21, 
    167, 341, 0, 
    149, 0, 0, 
    
    -- channel=75
    0, 0, 0, 
    5, 89, 0, 
    0, 0, 0, 
    
    -- channel=76
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=77
    0, 0, 0, 
    0, 0, 84, 
    0, 192, 31, 
    
    -- channel=78
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=79
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=80
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=81
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=82
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=83
    272, 0, 204, 
    523, 0, 116, 
    0, 0, 0, 
    
    -- channel=84
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=85
    0, 148, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=86
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=87
    93, 233, 0, 
    53, 410, 0, 
    0, 0, 0, 
    
    -- channel=88
    422, 603, 0, 
    20, 0, 0, 
    0, 0, 0, 
    
    -- channel=89
    0, 0, 0, 
    0, 3, 0, 
    0, 0, 81, 
    
    -- channel=90
    0, 0, 0, 
    0, 0, 0, 
    0, 281, 0, 
    
    -- channel=91
    72, 0, 0, 
    0, 0, 105, 
    0, 0, 0, 
    
    -- channel=92
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=93
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=94
    0, 0, 0, 
    0, 0, 0, 
    0, 293, 175, 
    
    -- channel=95
    0, 78, 0, 
    0, 0, 0, 
    0, 323, 388, 
    
    -- channel=96
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=97
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=98
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=99
    0, 118, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=100
    0, 499, 0, 
    509, 0, 79, 
    0, 0, 0, 
    
    -- channel=101
    77, 0, 24, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=102
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=103
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=104
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=105
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=106
    244, 0, 0, 
    207, 0, 0, 
    0, 0, 0, 
    
    -- channel=107
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=108
    0, 0, 150, 
    142, 147, 393, 
    0, 0, 0, 
    
    -- channel=109
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=110
    0, 0, 0, 
    0, 0, 0, 
    0, 123, 227, 
    
    -- channel=111
    3, 121, 105, 
    0, 59, 146, 
    0, 484, 212, 
    
    -- channel=112
    0, 102, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=113
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=114
    85, 0, 0, 
    237, 286, 0, 
    0, 149, 68, 
    
    -- channel=115
    0, 0, 0, 
    0, 75, 111, 
    493, 0, 0, 
    
    -- channel=116
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=117
    23, 0, 0, 
    0, 208, 204, 
    172, 0, 0, 
    
    -- channel=118
    191, 0, 235, 
    338, 0, 0, 
    0, 0, 0, 
    
    -- channel=119
    0, 187, 0, 
    0, 48, 0, 
    163, 564, 35, 
    
    -- channel=120
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=121
    26, 0, 292, 
    0, 57, 0, 
    0, 0, 0, 
    
    -- channel=122
    416, 0, 196, 
    0, 38, 188, 
    0, 0, 0, 
    
    -- channel=123
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=124
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=125
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=126
    0, 0, 213, 
    0, 18, 0, 
    0, 0, 0, 
    
    -- channel=127
    39, 96, 53, 
    17, 236, 162, 
    105, 0, 0, 
    
    -- channel=128
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=129
    69, 387, 0, 
    424, 341, 490, 
    0, 0, 0, 
    
    -- channel=130
    0, 0, 0, 
    0, 0, 0, 
    0, 10, 0, 
    
    -- channel=131
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=132
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=133
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=134
    0, 0, 0, 
    0, 72, 0, 
    483, 448, 582, 
    
    -- channel=135
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=136
    0, 0, 0, 
    0, 0, 462, 
    109, 0, 0, 
    
    -- channel=137
    0, 0, 239, 
    0, 62, 0, 
    0, 0, 32, 
    
    -- channel=138
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=139
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=140
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=141
    0, 53, 0, 
    0, 31, 0, 
    0, 0, 0, 
    
    -- channel=142
    0, 230, 0, 
    107, 0, 0, 
    0, 0, 0, 
    
    -- channel=143
    240, 322, 0, 
    304, 338, 23, 
    0, 0, 0, 
    
    -- channel=144
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=145
    101, 0, 31, 
    0, 0, 127, 
    0, 12, 0, 
    
    -- channel=146
    0, 0, 139, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=147
    198, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=148
    0, 141, 0, 
    0, 37, 152, 
    215, 148, 95, 
    
    -- channel=149
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=150
    208, 0, 24, 
    182, 0, 0, 
    0, 0, 0, 
    
    -- channel=151
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=152
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=153
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=154
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=155
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=156
    0, 0, 0, 
    0, 0, 0, 
    136, 0, 148, 
    
    -- channel=157
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=158
    0, 49, 0, 
    0, 0, 0, 
    0, 166, 0, 
    
    -- channel=159
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=160
    170, 311, 290, 
    220, 330, 414, 
    64, 0, 173, 
    
    -- channel=161
    0, 81, 0, 
    0, 0, 0, 
    139, 0, 0, 
    
    -- channel=162
    0, 21, 78, 
    300, 0, 454, 
    181, 235, 164, 
    
    -- channel=163
    0, 0, 0, 
    0, 36, 0, 
    0, 0, 0, 
    
    -- channel=164
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=165
    0, 0, 199, 
    0, 0, 139, 
    96, 0, 0, 
    
    -- channel=166
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=167
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=168
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=169
    0, 0, 0, 
    156, 0, 0, 
    0, 30, 0, 
    
    -- channel=170
    0, 0, 0, 
    0, 0, 15, 
    0, 537, 0, 
    
    -- channel=171
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=172
    506, 0, 361, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=173
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=174
    0, 276, 0, 
    196, 0, 0, 
    0, 0, 0, 
    
    -- channel=175
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=176
    0, 0, 0, 
    0, 0, 0, 
    15, 0, 18, 
    
    -- channel=177
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=178
    0, 0, 0, 
    0, 0, 0, 
    55, 0, 0, 
    
    -- channel=179
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=180
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=181
    0, 0, 291, 
    187, 0, 0, 
    0, 112, 0, 
    
    -- channel=182
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=183
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=184
    16, 263, 175, 
    146, 65, 0, 
    70, 108, 338, 
    
    -- channel=185
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=186
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=187
    0, 0, 0, 
    91, 264, 150, 
    440, 0, 0, 
    
    -- channel=188
    0, 0, 0, 
    0, 0, 0, 
    0, 486, 130, 
    
    -- channel=189
    688, 686, 454, 
    437, 0, 0, 
    0, 0, 0, 
    
    -- channel=190
    0, 0, 0, 
    0, 6, 45, 
    0, 0, 0, 
    
    -- channel=191
    0, 0, 0, 
    0, 198, 0, 
    0, 0, 0, 
    
    -- channel=192
    0, 313, 23, 
    0, 120, 33, 
    0, 0, 0, 
    
    -- channel=193
    0, 65, 0, 
    0, 0, 0, 
    0, 260, 512, 
    
    -- channel=194
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=195
    153, 0, 266, 
    97, 0, 363, 
    0, 236, 0, 
    
    -- channel=196
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=197
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=198
    179, 0, 204, 
    251, 371, 475, 
    352, 705, 218, 
    
    -- channel=199
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=200
    0, 0, 0, 
    62, 0, 0, 
    249, 0, 0, 
    
    -- channel=201
    7, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=202
    0, 0, 0, 
    90, 0, 0, 
    0, 0, 0, 
    
    -- channel=203
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=204
    39, 0, 57, 
    246, 275, 0, 
    0, 0, 0, 
    
    -- channel=205
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=206
    0, 0, 0, 
    260, 0, 0, 
    63, 0, 130, 
    
    -- channel=207
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=208
    107, 0, 0, 
    0, 0, 30, 
    0, 0, 0, 
    
    -- channel=209
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=210
    7, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=211
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=212
    167, 0, 58, 
    0, 34, 0, 
    0, 0, 0, 
    
    -- channel=213
    250, 0, 187, 
    90, 0, 151, 
    110, 0, 0, 
    
    -- channel=214
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=215
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 353, 
    
    -- channel=216
    0, 70, 0, 
    0, 285, 0, 
    0, 0, 0, 
    
    -- channel=217
    184, 0, 171, 
    65, 0, 151, 
    0, 6, 179, 
    
    -- channel=218
    42, 0, 210, 
    0, 334, 0, 
    0, 0, 0, 
    
    -- channel=219
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=220
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=221
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=222
    300, 0, 283, 
    140, 30, 181, 
    387, 131, 396, 
    
    -- channel=223
    0, 61, 198, 
    126, 164, 0, 
    6, 106, 0, 
    
    -- channel=224
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=225
    0, 0, 0, 
    261, 44, 30, 
    0, 0, 0, 
    
    -- channel=226
    0, 0, 35, 
    5, 0, 0, 
    0, 556, 109, 
    
    -- channel=227
    67, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=228
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=229
    0, 55, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=230
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=231
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=232
    0, 0, 0, 
    0, 0, 0, 
    0, 12, 222, 
    
    -- channel=233
    0, 226, 0, 
    0, 0, 0, 
    363, 0, 0, 
    
    -- channel=234
    265, 65, 16, 
    288, 166, 31, 
    0, 0, 0, 
    
    -- channel=235
    62, 317, 0, 
    279, 0, 329, 
    0, 0, 449, 
    
    -- channel=236
    116, 261, 0, 
    89, 0, 46, 
    0, 0, 0, 
    
    -- channel=237
    344, 649, 333, 
    366, 0, 129, 
    100, 573, 505, 
    
    -- channel=238
    0, 73, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=239
    0, 0, 38, 
    146, 2, 131, 
    0, 0, 0, 
    
    -- channel=240
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=241
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=242
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=243
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=244
    0, 53, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=245
    0, 0, 0, 
    11, 0, 0, 
    86, 290, 133, 
    
    -- channel=246
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=247
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=248
    78, 275, 0, 
    0, 0, 102, 
    0, 0, 0, 
    
    -- channel=249
    0, 0, 0, 
    0, 0, 0, 
    0, 299, 502, 
    
    -- channel=250
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=251
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=252
    0, 0, 126, 
    167, 124, 221, 
    0, 69, 0, 
    
    -- channel=253
    0, 0, 148, 
    503, 0, 151, 
    108, 0, 239, 
    
    -- channel=254
    0, 0, 0, 
    0, 0, 64, 
    0, 0, 0, 
    
    -- channel=255
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    
    others => 0);
end gold_package;
