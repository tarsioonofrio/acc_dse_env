library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    16, 16, 10, 9, 6, 8, 12, 13, 5, 11, 20, 15, 7, 2, 1, 
    0, 3, 9, 11, 10, 0, 3, 5, 41, 0, 0, 0, 0, 5, 0, 
    15, 31, 8, 10, 12, 76, 44, 19, 0, 0, 33, 18, 0, 0, 0, 
    0, 0, 1, 3, 0, 3, 0, 8, 1, 41, 45, 36, 28, 0, 0, 
    39, 0, 17, 14, 0, 10, 51, 19, 13, 0, 17, 11, 0, 0, 0, 
    105, 43, 39, 58, 127, 124, 37, 20, 0, 0, 83, 60, 14, 3, 0, 
    94, 42, 46, 19, 30, 26, 79, 44, 23, 0, 86, 19, 1, 0, 2, 
    88, 59, 7, 0, 11, 59, 128, 80, 44, 30, 77, 35, 15, 37, 32, 
    95, 79, 65, 14, 19, 105, 50, 0, 1, 18, 53, 72, 21, 3, 0, 
    113, 94, 64, 12, 46, 36, 27, 0, 23, 75, 53, 0, 0, 0, 15, 
    53, 84, 80, 0, 0, 0, 34, 114, 60, 0, 0, 0, 0, 0, 1, 
    86, 103, 76, 33, 196, 135, 71, 72, 39, 17, 12, 21, 20, 23, 30, 
    16, 68, 81, 109, 163, 21, 22, 19, 15, 7, 6, 7, 31, 42, 14, 
    35, 10, 77, 144, 57, 21, 15, 16, 22, 20, 31, 44, 36, 11, 74, 
    41, 24, 28, 80, 36, 38, 49, 28, 12, 11, 27, 26, 3, 27, 31, 
    
    -- channel=1
    122, 124, 128, 128, 128, 124, 129, 139, 135, 113, 97, 100, 105, 113, 112, 
    129, 131, 135, 130, 131, 123, 114, 116, 78, 60, 37, 45, 70, 93, 107, 
    96, 103, 130, 133, 135, 113, 62, 53, 49, 47, 23, 25, 23, 62, 89, 
    20, 92, 114, 136, 114, 89, 53, 37, 27, 59, 20, 35, 14, 31, 85, 
    0, 61, 89, 135, 67, 61, 26, 25, 22, 62, 36, 24, 34, 20, 66, 
    4, 34, 77, 95, 54, 40, 24, 32, 13, 92, 20, 12, 38, 22, 27, 
    9, 3, 68, 80, 85, 67, 32, 23, 11, 70, 1, 17, 30, 31, 32, 
    12, 0, 44, 53, 82, 69, 10, 26, 22, 75, 17, 13, 36, 36, 61, 
    1, 5, 0, 35, 49, 32, 28, 32, 51, 39, 49, 13, 36, 60, 102, 
    13, 13, 0, 25, 16, 51, 48, 15, 44, 40, 10, 20, 52, 98, 104, 
    15, 15, 0, 71, 0, 22, 31, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 2, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 25, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=2
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 0, 0, 13, 0, 8, 0, 0, 0, 7, 0, 0, 0, 0, 
    22, 23, 0, 0, 37, 11, 15, 0, 0, 0, 16, 0, 0, 0, 0, 
    18, 33, 0, 0, 0, 0, 42, 0, 0, 0, 23, 0, 0, 0, 0, 
    29, 50, 0, 0, 0, 35, 11, 0, 0, 0, 7, 0, 0, 0, 0, 
    50, 60, 7, 5, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    46, 47, 32, 11, 28, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 
    53, 44, 34, 23, 44, 22, 24, 54, 14, 0, 0, 0, 6, 27, 27, 
    65, 54, 40, 50, 98, 48, 37, 41, 32, 24, 27, 30, 37, 37, 41, 
    38, 41, 32, 87, 56, 26, 25, 20, 20, 22, 32, 39, 42, 45, 50, 
    53, 35, 42, 88, 27, 26, 26, 24, 25, 32, 38, 49, 44, 55, 57, 
    48, 42, 30, 60, 19, 25, 30, 23, 26, 35, 38, 32, 45, 66, 46, 
    
    -- channel=3
    17, 26, 21, 21, 16, 25, 15, 10, 10, 11, 17, 21, 24, 10, 6, 
    11, 14, 17, 19, 25, 80, 14, 16, 17, 56, 55, 28, 20, 15, 11, 
    17, 22, 15, 16, 13, 65, 53, 25, 28, 107, 112, 102, 48, 5, 29, 
    43, 29, 12, 17, 27, 51, 77, 61, 65, 94, 121, 70, 72, 15, 18, 
    132, 106, 34, 61, 158, 118, 126, 83, 56, 84, 121, 70, 70, 42, 0, 
    152, 176, 61, 44, 193, 161, 161, 91, 56, 120, 155, 93, 76, 73, 34, 
    163, 163, 54, 28, 89, 151, 172, 135, 81, 143, 149, 83, 71, 88, 64, 
    184, 201, 68, 54, 59, 175, 175, 120, 91, 127, 148, 85, 77, 88, 67, 
    220, 215, 130, 128, 75, 110, 97, 90, 85, 64, 77, 74, 54, 67, 33, 
    232, 216, 159, 143, 103, 78, 125, 144, 79, 90, 64, 26, 38, 41, 30, 
    208, 201, 159, 212, 225, 110, 165, 200, 125, 67, 56, 76, 90, 95, 83, 
    166, 226, 186, 247, 229, 162, 133, 132, 122, 114, 125, 137, 153, 154, 153, 
    148, 151, 215, 249, 187, 137, 127, 124, 123, 128, 144, 154, 157, 164, 186, 
    168, 138, 166, 250, 145, 142, 136, 123, 133, 145, 155, 162, 162, 178, 175, 
    172, 159, 137, 147, 115, 127, 141, 142, 145, 159, 146, 151, 186, 200, 150, 
    
    -- channel=4
    113, 109, 108, 111, 113, 98, 113, 124, 119, 110, 104, 98, 95, 98, 106, 
    109, 104, 108, 115, 108, 60, 97, 103, 117, 58, 29, 42, 70, 92, 98, 
    109, 118, 114, 118, 119, 143, 127, 88, 38, 13, 41, 40, 44, 58, 81, 
    56, 3, 104, 110, 103, 76, 38, 40, 44, 34, 79, 61, 72, 47, 55, 
    48, 0, 101, 57, 0, 3, 61, 54, 62, 12, 35, 47, 36, 40, 38, 
    67, 42, 106, 118, 101, 88, 62, 48, 47, 0, 81, 87, 40, 43, 18, 
    49, 58, 98, 123, 55, 37, 73, 64, 62, 0, 92, 54, 39, 27, 41, 
    43, 47, 28, 73, 37, 25, 120, 92, 77, 36, 93, 71, 35, 56, 82, 
    52, 34, 70, 32, 59, 102, 81, 48, 26, 85, 76, 112, 56, 53, 64, 
    82, 49, 76, 4, 45, 51, 36, 19, 36, 96, 101, 43, 2, 54, 109, 
    37, 48, 88, 0, 3, 0, 0, 75, 63, 43, 0, 0, 0, 28, 40, 
    30, 55, 40, 0, 157, 116, 56, 55, 31, 12, 2, 2, 0, 0, 4, 
    0, 22, 24, 78, 136, 4, 4, 7, 8, 0, 0, 0, 0, 5, 0, 
    4, 0, 0, 139, 50, 0, 3, 0, 0, 0, 2, 9, 7, 0, 28, 
    5, 0, 5, 67, 35, 20, 25, 9, 0, 0, 0, 0, 0, 0, 10, 
    
    -- channel=5
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 19, 15, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 44, 0, 0, 0, 5, 13, 0, 
    18, 50, 0, 0, 0, 62, 5, 10, 0, 0, 0, 0, 0, 10, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 84, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 13, 0, 28, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 17, 12, 22, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 48, 0, 0, 0, 0, 34, 38, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 42, 15, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 46, 7, 0, 0, 0, 0, 7, 4, 
    72, 29, 0, 0, 46, 49, 28, 25, 7, 0, 0, 0, 0, 0, 0, 
    0, 38, 0, 0, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 20, 79, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 20, 
    0, 0, 0, 73, 3, 12, 20, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=6
    1, 0, 6, 0, 0, 2, 0, 0, 0, 0, 0, 9, 3, 0, 0, 
    1, 1, 6, 0, 13, 29, 0, 0, 0, 27, 0, 0, 4, 18, 0, 
    0, 57, 3, 0, 9, 7, 0, 0, 11, 81, 0, 0, 0, 10, 31, 
    0, 101, 0, 12, 0, 32, 0, 0, 0, 104, 0, 0, 0, 0, 85, 
    0, 29, 0, 102, 0, 0, 0, 0, 0, 148, 0, 0, 0, 0, 30, 
    0, 8, 0, 30, 104, 0, 0, 0, 0, 257, 0, 0, 13, 0, 0, 
    0, 0, 0, 0, 97, 86, 0, 0, 0, 203, 0, 0, 4, 21, 0, 
    0, 0, 0, 0, 67, 95, 0, 0, 0, 128, 0, 0, 33, 0, 0, 
    0, 0, 0, 47, 0, 9, 0, 0, 31, 0, 14, 0, 31, 32, 14, 
    0, 0, 0, 85, 0, 8, 57, 0, 0, 0, 0, 0, 45, 46, 0, 
    94, 0, 0, 220, 0, 0, 75, 0, 0, 0, 0, 20, 13, 10, 0, 
    78, 65, 0, 150, 0, 0, 0, 0, 0, 0, 2, 6, 5, 0, 0, 
    0, 82, 133, 0, 0, 0, 0, 0, 0, 3, 8, 5, 0, 4, 14, 
    0, 0, 172, 0, 0, 4, 0, 0, 6, 4, 0, 0, 0, 35, 0, 
    0, 0, 11, 0, 0, 22, 8, 0, 12, 0, 0, 4, 58, 0, 0, 
    
    -- channel=7
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 34, 27, 40, 24, 0, 0, 
    27, 7, 0, 0, 0, 0, 5, 21, 23, 0, 6, 0, 13, 13, 0, 
    52, 41, 0, 0, 39, 21, 5, 22, 15, 17, 23, 21, 32, 38, 0, 
    26, 16, 0, 0, 0, 0, 10, 22, 42, 36, 1, 7, 20, 38, 46, 
    43, 14, 0, 0, 0, 0, 0, 15, 24, 21, 3, 28, 28, 33, 23, 
    33, 50, 23, 0, 0, 0, 0, 0, 1, 0, 0, 15, 21, 0, 0, 
    42, 42, 34, 14, 0, 0, 0, 18, 22, 0, 0, 0, 2, 0, 0, 
    9, 25, 40, 47, 16, 14, 25, 46, 17, 0, 0, 30, 28, 0, 0, 
    28, 22, 28, 78, 102, 89, 47, 23, 44, 65, 98, 114, 104, 66, 59, 
    62, 39, 45, 31, 0, 32, 59, 65, 91, 108, 121, 124, 135, 129, 131, 
    149, 64, 47, 0, 50, 118, 115, 113, 117, 129, 143, 150, 132, 133, 167, 
    157, 140, 57, 27, 88, 124, 126, 118, 121, 134, 136, 131, 142, 167, 116, 
    154, 149, 110, 72, 96, 101, 103, 120, 130, 142, 133, 137, 162, 166, 151, 
    
    -- channel=8
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=9
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 63, 5, 0, 0, 29, 54, 19, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 31, 72, 34, 34, 26, 0, 1, 
    20, 67, 1, 2, 0, 30, 55, 33, 28, 33, 11, 7, 3, 4, 8, 
    62, 104, 3, 61, 125, 87, 16, 14, 0, 71, 59, 31, 34, 25, 0, 
    28, 45, 0, 0, 0, 7, 46, 35, 19, 127, 13, 0, 25, 30, 41, 
    51, 28, 0, 0, 19, 76, 27, 37, 9, 96, 9, 23, 33, 56, 29, 
    61, 52, 48, 27, 62, 60, 0, 0, 1, 44, 15, 3, 29, 9, 0, 
    60, 65, 18, 54, 33, 0, 7, 39, 50, 13, 0, 0, 0, 24, 29, 
    36, 56, 20, 83, 21, 11, 56, 86, 21, 0, 0, 9, 52, 36, 0, 
    68, 57, 7, 155, 151, 119, 81, 4, 7, 29, 69, 96, 72, 48, 44, 
    14, 40, 67, 142, 0, 0, 1, 4, 30, 52, 60, 61, 74, 71, 64, 
    70, 24, 81, 36, 0, 58, 53, 52, 57, 70, 81, 86, 65, 66, 101, 
    65, 68, 51, 0, 36, 64, 66, 57, 59, 67, 64, 55, 64, 98, 29, 
    61, 68, 58, 0, 30, 35, 35, 55, 81, 84, 65, 69, 125, 96, 55, 
    
    -- channel=10
    125, 123, 128, 131, 131, 121, 137, 145, 133, 108, 87, 90, 100, 113, 108, 
    130, 136, 135, 136, 130, 117, 139, 114, 77, 35, 31, 41, 54, 81, 105, 
    86, 86, 134, 138, 139, 118, 73, 47, 20, 18, 29, 16, 24, 41, 76, 
    48, 51, 133, 134, 119, 74, 60, 25, 13, 24, 44, 31, 9, 9, 50, 
    30, 58, 130, 96, 87, 88, 61, 28, 12, 8, 55, 41, 17, 9, 33, 
    34, 41, 126, 99, 28, 56, 60, 47, 26, 7, 65, 28, 16, 12, 11, 
    34, 44, 85, 105, 47, 51, 65, 48, 32, 21, 50, 27, 14, 12, 33, 
    41, 36, 55, 86, 54, 51, 57, 33, 29, 46, 40, 30, 6, 33, 59, 
    38, 33, 32, 19, 67, 38, 43, 32, 26, 83, 33, 17, 8, 38, 97, 
    36, 37, 30, 11, 40, 31, 28, 46, 49, 25, 10, 0, 9, 91, 114, 
    9, 46, 37, 12, 48, 37, 11, 14, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 31, 63, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 68, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=11
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 0, 0, 27, 10, 0, 
    20, 47, 0, 0, 0, 86, 2, 22, 0, 0, 0, 0, 0, 40, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 0, 20, 0, 0, 42, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 39, 
    0, 0, 0, 26, 107, 13, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 6, 33, 0, 58, 0, 3, 0, 0, 26, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 18, 40, 0, 33, 0, 0, 8, 23, 0, 
    0, 0, 0, 0, 0, 92, 3, 0, 0, 19, 49, 36, 35, 0, 0, 
    0, 1, 0, 5, 0, 0, 0, 0, 6, 33, 31, 6, 0, 0, 0, 
    18, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 21, 3, 
    136, 37, 0, 0, 88, 74, 77, 65, 14, 1, 0, 6, 0, 0, 0, 
    0, 108, 8, 28, 31, 0, 0, 0, 0, 0, 0, 0, 6, 7, 0, 
    0, 7, 112, 46, 0, 0, 0, 0, 0, 0, 8, 22, 3, 0, 63, 
    0, 1, 31, 90, 28, 36, 29, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=12
    3, 0, 0, 3, 5, 0, 5, 2, 5, 11, 9, 0, 0, 10, 11, 
    0, 0, 0, 7, 0, 0, 46, 20, 25, 0, 10, 21, 0, 0, 6, 
    46, 0, 3, 3, 1, 0, 52, 5, 0, 0, 28, 0, 48, 0, 0, 
    92, 0, 11, 0, 31, 0, 9, 36, 14, 0, 57, 18, 33, 44, 0, 
    62, 0, 65, 0, 0, 38, 56, 58, 36, 0, 0, 77, 0, 39, 0, 
    91, 0, 80, 80, 0, 18, 42, 27, 70, 0, 92, 74, 0, 17, 30, 
    77, 45, 7, 66, 0, 0, 1, 48, 59, 0, 81, 56, 0, 0, 38, 
    77, 0, 48, 17, 0, 0, 103, 16, 30, 0, 44, 60, 0, 3, 4, 
    65, 0, 152, 0, 81, 0, 11, 15, 0, 43, 0, 68, 0, 0, 0, 
    0, 0, 117, 0, 56, 34, 0, 3, 55, 22, 56, 0, 0, 0, 17, 
    0, 2, 97, 0, 95, 51, 0, 15, 76, 36, 0, 0, 0, 0, 12, 
    0, 0, 3, 0, 163, 63, 0, 0, 6, 0, 0, 0, 0, 0, 5, 
    31, 0, 0, 48, 117, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 0, 0, 62, 31, 0, 13, 2, 0, 0, 0, 0, 0, 0, 40, 
    43, 0, 12, 0, 17, 0, 0, 0, 0, 0, 15, 0, 0, 18, 49, 
    
    -- channel=13
    101, 112, 111, 111, 107, 107, 116, 121, 107, 81, 70, 79, 93, 100, 95, 
    110, 119, 115, 113, 108, 123, 106, 94, 58, 42, 36, 40, 50, 71, 90, 
    68, 70, 111, 117, 110, 84, 65, 37, 30, 38, 37, 37, 32, 32, 80, 
    45, 56, 104, 110, 99, 62, 62, 32, 25, 25, 56, 34, 28, 24, 55, 
    35, 62, 100, 74, 102, 79, 65, 46, 27, 29, 58, 46, 35, 31, 31, 
    15, 51, 106, 72, 51, 65, 83, 54, 43, 33, 54, 35, 28, 28, 34, 
    28, 48, 70, 97, 53, 64, 57, 53, 43, 32, 45, 36, 26, 28, 43, 
    39, 53, 38, 74, 38, 49, 49, 38, 44, 52, 49, 36, 21, 39, 72, 
    40, 39, 28, 43, 47, 33, 48, 41, 35, 58, 28, 28, 25, 62, 94, 
    42, 37, 40, 26, 38, 35, 42, 58, 37, 31, 20, 8, 34, 83, 87, 
    21, 40, 38, 40, 72, 32, 15, 20, 15, 9, 0, 0, 0, 0, 0, 
    0, 4, 36, 55, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=14
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 9, 1, 0, 0, 0, 0, 
    0, 9, 0, 0, 0, 24, 3, 0, 0, 49, 37, 34, 3, 0, 0, 
    0, 3, 0, 0, 0, 6, 11, 10, 20, 59, 35, 26, 21, 0, 12, 
    33, 35, 0, 21, 34, 24, 32, 14, 14, 50, 37, 6, 20, 0, 0, 
    55, 75, 0, 5, 107, 68, 47, 21, 0, 75, 50, 24, 31, 19, 0, 
    56, 61, 14, 0, 49, 63, 71, 41, 14, 90, 49, 17, 25, 35, 11, 
    66, 77, 10, 0, 27, 88, 62, 56, 26, 71, 57, 20, 35, 36, 16, 
    83, 99, 30, 57, 13, 60, 33, 25, 34, 16, 34, 21, 24, 22, 0, 
    105, 101, 45, 74, 28, 23, 54, 45, 19, 38, 20, 7, 14, 9, 0, 
    111, 88, 51, 112, 60, 22, 81, 95, 39, 17, 16, 28, 34, 43, 29, 
    116, 122, 76, 130, 103, 80, 75, 74, 60, 60, 67, 74, 82, 83, 80, 
    77, 102, 118, 113, 76, 68, 65, 65, 64, 69, 78, 80, 85, 92, 96, 
    88, 75, 115, 117, 70, 75, 66, 63, 71, 77, 85, 93, 90, 97, 101, 
    86, 86, 79, 90, 63, 77, 83, 75, 76, 80, 76, 84, 102, 98, 73, 
    
    -- channel=15
    56, 56, 58, 57, 56, 53, 66, 73, 59, 38, 32, 39, 43, 49, 44, 
    58, 67, 61, 60, 56, 23, 49, 45, 30, 0, 0, 0, 8, 33, 40, 
    17, 50, 65, 66, 64, 35, 16, 0, 0, 0, 0, 0, 0, 0, 29, 
    0, 0, 59, 63, 36, 19, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 39, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 37, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 22, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 36, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end gold_package;
