LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
	PACKAGE gold_package is
		type padroes is array(0 to 4000000) of integer;
		constant gold: padroes := ( 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 150, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 238, 0, 0, 0, 132, 0, 0, 
		88, 193, 0, 0, 0, 78, 149, 58, 0, 0, 0, 0, 0, 238, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 220, 0, 182, 170, 0, 161, 
		0, 0, 0, 0, 0, 0, 0, 0, 123, 0, 0, 0, 0, 0, 247, 
		115, 0, 0, 220, 28, 170, 0, 0, 0, 0, 0, 130, 0, 0, 0, 
		0, 0, 40, 0, 217, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 212, 103, 0, 0, 134, 81, 0, 0, 0, 
		0, 0, 0, 0, 0, 229, 100, 0, 0, 141, 154, 180, 212, 0, 0, 
		0, 0, 0, 0, 0, 199, 0, 0, 0, 19, 248, 28, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51, 83, 
		100, 125, 0, 0, 67, 156, 46, 38, 160, 0, 0, 0, 0, 0, 0, 
		0, 21, 0, 0, 160, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 2, 12, 225, 0, 0, 0, 0, 0, 149, 36, 165, 0, 38, 
		0, 0, 54, 59, 23, 176, 242, 0, 0, 0, 0, 0, 0, 0, 0, 
		
		23, 170, 28, 61, 139, 40, 36, 58, 226, 117, 249, 47, 143, 149, 39, 
		59, 184, 26, 207, 253, 111, 110, 242, 240, 197, 81, 152, 40, 204, 41, 
		179, 80, 127, 101, 147, 69, 204, 189, 116, 201, 109, 7, 63, 41, 228, 
		239, 243, 39, 247, 187, 6, 21, 97, 134, 152, 155, 92, 192, 120, 12, 
		122, 251, 32, 107, 247, 104, 212, 221, 85, 93, 5, 150, 94, 223, 141, 
		0, 16, 92, 31, 255, 28, 72, 22, 0, 232, 14, 135, 41, 170, 189, 
		212, 101, 252, 130, 71, 220, 223, 254, 0, 240, 70, 206, 191, 255, 102, 
		148, 65, 154, 137, 156, 72, 0, 80, 108, 21, 156, 72, 164, 51, 185, 
		130, 200, 0, 177, 77, 171, 56, 115, 84, 22, 235, 0, 108, 24, 113, 
		58, 235, 0, 237, 187, 180, 82, 137, 35, 128, 159, 96, 26, 47, 172, 
		130, 87, 0, 193, 78, 11, 164, 47, 104, 45, 77, 201, 101, 107, 216, 
		148, 107, 46, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 9, 128, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 237, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		
		55, 233, 225, 76, 85, 113, 151, 183, 61, 192, 154, 120, 169, 216, 135, 
		213, 105, 82, 96, 161, 74, 180, 252, 152, 106, 36, 87, 144, 71, 64, 
		71, 245, 239, 248, 80, 208, 56, 78, 175, 212, 189, 40, 223, 21, 144, 
		93, 212, 145, 145, 211, 25, 85, 199, 15, 194, 243, 178, 230, 254, 151, 
		94, 145, 146, 205, 238, 76, 135, 51, 207, 100, 77, 214, 63, 244, 228, 
		216, 90, 127, 150, 108, 197, 63, 232, 52, 162, 168, 178, 10, 171, 13, 
		20, 193, 211, 178, 182, 144, 60, 73, 11, 103, 212, 110, 10, 135, 23, 
		118, 197, 173, 115, 21, 242, 31, 75, 85, 151, 176, 120, 2, 247, 46, 
		131, 147, 213, 118, 209, 60, 67, 70, 32, 231, 36, 177, 1, 117, 173, 
		4, 44, 65, 232, 86, 173, 180, 170, 206, 179, 28, 198, 85, 57, 166, 
		15, 187, 159, 107, 251, 162, 249, 45, 20, 178, 132, 182, 53, 36, 93, 
		137, 18, 215, 90, 207, 34, 192, 108, 22, 121, 16, 229, 66, 1, 8, 
		188, 124, 81, 53, 248, 136, 101, 210, 35, 52, 163, 50, 253, 33, 199, 
		153, 199, 226, 197, 105, 242, 73, 188, 117, 142, 30, 246, 248, 33, 103, 
		150, 81, 183, 74, 47, 164, 227, 158, 51, 92, 233, 151, 53, 188, 238, 
		
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 49, 0, 0, 0, 143, 118, 0, 0, 0, 
		166, 0, 0, 0, 0, 0, 0, 181, 132, 0, 76, 82, 17, 0, 0, 
		20, 0, 0, 0, 0, 0, 67, 209, 89, 0, 12, 174, 27, 240, 0, 
		179, 225, 86, 0, 165, 199, 75, 72, 217, 0, 101, 66, 10, 107, 0, 
		121, 194, 15, 0, 0, 204, 69, 161, 62, 0, 160, 238, 19, 61, 169, 
		160, 243, 153, 135, 0, 0, 220, 97, 105, 0, 69, 137, 149, 238, 69, 
		18, 87, 55, 9, 0, 0, 48, 72, 13, 0, 49, 163, 0, 208, 94, 
		109, 125, 48, 0, 67, 0, 45, 83, 135, 236, 0, 60, 0, 0, 124, 
		172, 120, 154, 0, 2, 0, 0, 159, 38, 0, 83, 135, 124, 0, 189, 
		0, 228, 24, 0, 49, 50, 99, 47, 105, 33, 97, 40, 31, 96, 174, 
		0, 0, 163, 0, 184, 28, 236, 126, 168, 13, 74, 250, 26, 213, 224, 
		243, 0, 0, 59, 67, 202, 124, 96, 200, 118, 140, 65, 243, 36, 158, 
		66, 156, 0, 38, 136, 170, 173, 187, 137, 89, 45, 54, 210, 74, 97, 
		43, 216, 26, 130, 241, 54, 202, 27, 239, 73, 96, 74, 153, 70, 14, 
		
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 220, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 209, 0, 0, 0, 0, 0, 0, 
		255, 49, 0, 0, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 110, 0, 0, 
		0, 118, 0, 0, 0, 0, 100, 68, 0, 0, 0, 194, 211, 0, 0, 
		152, 184, 105, 0, 0, 83, 0, 0, 0, 0, 96, 144, 76, 0, 0, 
		53, 108, 170, 117, 254, 0, 0, 0, 134, 0, 55, 221, 0, 0, 0, 
		53, 233, 225, 0, 0, 0, 0, 180, 72, 244, 189, 140, 198, 50, 147, 
		17, 16, 135, 0, 170, 206, 128, 168, 35, 71, 147, 103, 88, 7, 64, 
		183, 190, 58, 199, 176, 217, 58, 154, 175, 245, 18, 40, 48, 103, 203, 
		137, 3, 23, 32, 230, 68, 73, 75, 195, 197, 202, 112, 177, 108, 195, 
		229, 49, 206, 116, 128, 26, 110, 2, 221, 137, 166, 11, 86, 135, 10, 
		
		209, 142, 76, 137, 16, 60, 61, 255, 205, 78, 166, 241, 85, 165, 170, 
		2, 249, 114, 231, 50, 86, 230, 33, 185, 253, 0, 15, 139, 185, 211, 
		135, 111, 19, 178, 196, 159, 232, 196, 113, 116, 0, 0, 0, 98, 179, 
		0, 119, 74, 114, 173, 25, 0, 0, 0, 56, 0, 0, 0, 0, 171, 
		0, 122, 0, 12, 52, 0, 0, 0, 0, 40, 0, 0, 0, 0, 110, 
		0, 30, 0, 217, 96, 99, 0, 0, 0, 241, 0, 0, 0, 0, 0, 
		0, 0, 138, 78, 222, 75, 0, 0, 0, 82, 0, 0, 0, 166, 0, 
		0, 0, 0, 0, 7, 174, 0, 222, 0, 236, 0, 0, 184, 0, 0, 
		0, 0, 0, 190, 0, 226, 0, 0, 231, 0, 75, 0, 20, 7, 106, 
		15, 0, 0, 64, 0, 0, 44, 0, 0, 38, 0, 21, 149, 179, 43, 
		75, 0, 0, 209, 0, 0, 44, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 144, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 195, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 101, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 120, 0, 228, 0, 0, 0, 
		0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 95, 0, 0, 106, 215, 0, 0, 0, 233, 99, 0, 11, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 197, 0, 0, 0, 0, 74, 
		0, 0, 0, 0, 0, 55, 0, 0, 0, 132, 0, 0, 73, 22, 0, 
		0, 123, 0, 0, 219, 0, 0, 0, 0, 211, 0, 0, 216, 0, 0, 
		0, 97, 0, 0, 0, 0, 0, 0, 202, 0, 0, 0, 0, 0, 0, 
		0, 121, 0, 97, 0, 0, 205, 10, 0, 0, 0, 0, 105, 0, 0, 
		40, 0, 0, 10, 190, 154, 176, 0, 0, 0, 189, 131, 152, 48, 0, 
		112, 0, 150, 108, 0, 0, 0, 141, 17, 223, 107, 111, 222, 197, 89, 
		176, 80, 222, 0, 0, 67, 69, 227, 72, 106, 13, 99, 133, 106, 176, 
		237, 21, 12, 0, 197, 145, 30, 99, 27, 158, 77, 60, 189, 207, 34, 
		107, 157, 206, 2, 86, 127, 37, 95, 233, 226, 75, 192, 99, 237, 223, 
		
		9, 83, 219, 173, 97, 89, 55, 23, 117, 226, 114, 93, 87, 73, 84, 
		23, 59, 205, 40, 147, 17, 64, 122, 182, 58, 150, 246, 93, 155, 189, 
		134, 0, 45, 18, 249, 71, 218, 112, 247, 202, 203, 77, 34, 197, 112, 
		52, 206, 94, 84, 186, 37, 218, 168, 89, 221, 137, 201, 5, 225, 47, 
		229, 84, 190, 236, 131, 50, 48, 148, 169, 26, 90, 175, 64, 255, 196, 
		121, 5, 20, 22, 0, 155, 147, 251, 105, 77, 123, 118, 184, 233, 190, 
		191, 215, 72, 109, 77, 18, 142, 79, 172, 240, 2, 73, 10, 20, 201, 
		29, 131, 194, 149, 248, 81, 212, 197, 136, 139, 220, 224, 53, 185, 50, 
		54, 0, 228, 35, 182, 247, 31, 110, 242, 74, 210, 119, 182, 217, 6, 
		247, 12, 134, 229, 23, 220, 251, 245, 123, 103, 248, 142, 138, 99, 27, 
		196, 76, 81, 49, 86, 90, 251, 235, 141, 220, 197, 154, 232, 255, 100, 
		0, 102, 152, 45, 229, 9, 172, 30, 214, 96, 112, 103, 101, 190, 218, 
		97, 74, 242, 239, 62, 10, 152, 238, 55, 237, 85, 168, 253, 148, 34, 
		132, 71, 0, 255, 192, 118, 57, 125, 129, 50, 162, 169, 65, 132, 14, 
		187, 6, 164, 0, 125, 60, 214, 14, 40, 91, 63, 242, 189, 135, 153, 
		
		202, 248, 63, 5, 12, 198, 67, 34, 87, 21, 108, 32, 187, 92, 156, 
		249, 65, 216, 182, 60, 0, 138, 193, 71, 9, 74, 247, 39, 243, 70, 
		111, 0, 235, 131, 50, 27, 197, 51, 139, 171, 36, 1, 85, 130, 165, 
		249, 140, 73, 57, 135, 25, 90, 239, 180, 138, 100, 246, 113, 249, 202, 
		116, 212, 187, 223, 133, 89, 61, 142, 228, 153, 211, 239, 178, 1, 254, 
		150, 85, 215, 127, 143, 139, 0, 197, 58, 142, 221, 146, 235, 204, 55, 
		47, 192, 29, 59, 136, 85, 2, 203, 76, 220, 64, 121, 252, 203, 107, 
		31, 53, 99, 134, 1, 247, 36, 162, 245, 191, 122, 244, 238, 179, 66, 
		56, 183, 239, 253, 95, 23, 243, 91, 217, 192, 152, 145, 35, 88, 11, 
		123, 34, 137, 217, 188, 21, 135, 59, 179, 42, 224, 25, 133, 176, 5, 
		29, 81, 56, 148, 124, 148, 11, 10, 4, 146, 186, 102, 107, 132, 29, 
		24, 150, 10, 189, 156, 137, 28, 107, 130, 162, 93, 97, 7, 239, 211, 
		42, 185, 9, 23, 141, 37, 11, 238, 53, 53, 89, 57, 222, 183, 216, 
		184, 109, 206, 50, 169, 21, 184, 203, 209, 57, 61, 118, 249, 226, 245, 
		141, 121, 183, 3, 62, 41, 93, 234, 109, 239, 160, 152, 150, 4, 176, 
		
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 122, 108, 0, 0, 0, 94, 36, 218, 0, 0, 
		0, 0, 0, 0, 128, 0, 0, 0, 137, 74, 0, 0, 189, 70, 0, 
		0, 177, 0, 0, 193, 0, 60, 0, 0, 0, 0, 0, 0, 210, 0, 
		0, 39, 116, 133, 0, 140, 0, 0, 0, 180, 25, 110, 0, 0, 170, 
		210, 0, 0, 116, 0, 0, 0, 0, 0, 186, 0, 0, 0, 0, 118, 
		40, 0, 0, 0, 0, 167, 0, 0, 0, 249, 0, 70, 1, 196, 8, 
		72, 0, 21, 0, 102, 0, 0, 0, 0, 186, 0, 0, 0, 0, 0, 
		0, 0, 38, 0, 153, 0, 0, 90, 0, 215, 0, 0, 0, 0, 171, 
		0, 0, 0, 207, 0, 64, 0, 0, 246, 0, 0, 0, 0, 164, 0, 
		0, 0, 0, 209, 0, 204, 0, 0, 0, 18, 194, 75, 92, 0, 0, 
		0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 113, 0, 
		237, 0, 0, 0, 0, 0, 0, 0, 0, 0, 94, 138, 0, 0, 206, 
		0, 26, 219, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 42, 0, 
		0, 0, 8, 0, 0, 0, 0, 0, 0, 211, 0, 0, 39, 139, 0, 
		
		218, 4, 27, 146, 193, 96, 253, 44, 2, 210, 184, 170, 85, 74, 20, 
		231, 239, 175, 3, 78, 112, 122, 153, 50, 61, 180, 4, 234, 16, 38, 
		38, 156, 59, 122, 50, 116, 36, 109, 227, 72, 30, 222, 154, 253, 161, 
		90, 247, 127, 118, 252, 164, 238, 229, 120, 222, 40, 244, 68, 49, 113, 
		220, 230, 90, 225, 193, 132, 130, 187, 41, 0, 218, 142, 117, 128, 164, 
		230, 123, 73, 65, 60, 13, 36, 218, 82, 0, 37, 202, 253, 162, 93, 
		212, 99, 67, 54, 197, 236, 47, 12, 141, 0, 210, 59, 50, 108, 138, 
		115, 188, 57, 70, 223, 63, 25, 206, 148, 17, 190, 96, 243, 57, 142, 
		214, 116, 68, 113, 114, 115, 36, 178, 26, 158, 173, 105, 125, 94, 243, 
		165, 69, 90, 0, 200, 4, 35, 156, 26, 24, 28, 57, 155, 220, 241, 
		0, 76, 64, 0, 47, 134, 0, 135, 153, 33, 0, 0, 0, 0, 0, 
		0, 0, 95, 0, 146, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 81, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 130, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		
		243, 158, 196, 254, 105, 92, 225, 97, 76, 95, 150, 7, 123, 132, 221, 
		186, 188, 146, 237, 226, 241, 244, 15, 246, 3, 213, 148, 0, 207, 140, 
		140, 0, 163, 186, 62, 130, 150, 27, 0, 0, 25, 138, 121, 0, 71, 
		107, 0, 255, 226, 25, 86, 44, 118, 2, 0, 162, 226, 248, 70, 0, 
		252, 0, 44, 0, 25, 238, 25, 149, 242, 0, 98, 41, 227, 1, 0, 
		157, 27, 177, 0, 242, 18, 142, 123, 219, 0, 106, 33, 185, 73, 67, 
		163, 186, 140, 96, 0, 0, 196, 114, 231, 0, 99, 218, 98, 185, 247, 
		202, 248, 215, 148, 0, 0, 184, 22, 96, 0, 205, 175, 0, 197, 245, 
		212, 23, 116, 105, 63, 77, 122, 74, 93, 27, 14, 231, 0, 248, 237, 
		107, 230, 41, 0, 68, 0, 48, 66, 111, 3, 2, 67, 0, 0, 140, 
		0, 142, 131, 0, 222, 0, 0, 73, 119, 133, 42, 0, 0, 0, 120, 
		0, 200, 186, 0, 80, 154, 24, 232, 242, 120, 61, 197, 183, 237, 200, 
		232, 0, 0, 235, 185, 27, 27, 214, 207, 229, 162, 31, 80, 22, 158, 
		167, 255, 0, 209, 33, 28, 110, 32, 79, 67, 202, 211, 164, 0, 133, 
		217, 116, 70, 59, 154, 0, 146, 99, 29, 19, 83, 73, 0, 69, 182, 
		
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 236, 0, 156, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 177, 0, 235, 115, 200, 252, 0, 0, 
		95, 0, 0, 0, 0, 0, 16, 191, 208, 51, 7, 222, 223, 0, 0, 
		174, 0, 0, 0, 118, 182, 20, 16, 224, 0, 74, 49, 199, 252, 0, 
		18, 36, 0, 0, 153, 94, 93, 248, 25, 0, 109, 204, 80, 122, 220, 
		195, 139, 0, 0, 230, 0, 6, 144, 190, 0, 237, 94, 216, 117, 95, 
		40, 127, 106, 0, 72, 244, 159, 63, 201, 0, 86, 5, 237, 236, 0, 
		39, 147, 115, 0, 41, 22, 189, 0, 0, 133, 0, 143, 163, 0, 0, 
		244, 5, 248, 69, 138, 179, 121, 231, 38, 192, 6, 37, 0, 0, 0, 
		147, 106, 189, 0, 66, 22, 202, 178, 87, 214, 166, 222, 27, 224, 132, 
		235, 125, 183, 5, 33, 189, 133, 190, 100, 182, 30, 248, 123, 173, 217, 
		231, 136, 202, 81, 140, 108, 6, 187, 194, 244, 248, 173, 254, 100, 66, 
		2, 129, 73, 171, 121, 56, 29, 233, 153, 125, 200, 8, 168, 71, 44, 
		116, 222, 178, 59, 158, 99, 207, 37, 52, 34, 109, 149, 185, 54, 182, 
		
		209, 173, 209, 253, 146, 89, 176, 221, 165, 214, 189, 60, 59, 85, 122, 
		168, 186, 123, 184, 171, 0, 131, 247, 151, 168, 99, 182, 150, 72, 166, 
		144, 54, 157, 39, 100, 181, 31, 99, 0, 0, 193, 66, 2, 185, 46, 
		105, 0, 58, 23, 208, 245, 99, 125, 159, 0, 86, 189, 16, 39, 0, 
		248, 0, 184, 0, 0, 84, 134, 69, 161, 0, 67, 88, 0, 250, 0, 
		83, 0, 66, 238, 0, 170, 191, 142, 78, 0, 56, 47, 0, 37, 153, 
		128, 160, 132, 119, 0, 0, 74, 189, 46, 0, 152, 230, 0, 0, 164, 
		130, 242, 246, 88, 0, 0, 216, 44, 51, 0, 206, 254, 0, 0, 203, 
		215, 0, 174, 0, 251, 40, 244, 189, 0, 155, 0, 91, 0, 0, 0, 
		30, 0, 13, 0, 2, 0, 0, 84, 112, 241, 106, 22, 0, 0, 166, 
		0, 0, 225, 0, 57, 0, 0, 33, 215, 169, 0, 0, 0, 0, 200, 
		0, 0, 197, 0, 98, 150, 93, 117, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 128, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 242, 147, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 253, 
		
		126, 122, 204, 231, 149, 1, 35, 58, 177, 204, 62, 252, 58, 116, 28, 
		236, 62, 225, 12, 24, 165, 102, 130, 75, 0, 0, 226, 66, 89, 142, 
		14, 108, 190, 119, 164, 77, 239, 37, 0, 0, 0, 0, 208, 184, 8, 
		113, 229, 39, 181, 47, 6, 182, 0, 0, 0, 0, 74, 0, 93, 134, 
		0, 0, 95, 184, 0, 136, 68, 0, 0, 0, 0, 33, 0, 0, 254, 
		0, 0, 251, 223, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 26, 88, 254, 0, 0, 0, 0, 0, 0, 0, 0, 0, 170, 
		0, 0, 229, 1, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 98, 
		0, 0, 0, 0, 15, 26, 0, 0, 0, 3, 0, 171, 0, 83, 172, 
		0, 0, 0, 0, 0, 180, 0, 0, 70, 0, 145, 0, 0, 205, 2, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
		
		others=>0 );
END gold_package;
