library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=1
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=2
    0, 0, 0, 
    0, 221, 0, 
    0, 0, 0, 
    
    -- channel=3
    399, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=4
    0, 0, 0, 
    0, 0, 123, 
    0, 0, 0, 
    
    -- channel=5
    0, 133, 249, 
    0, 0, 252, 
    0, 0, 0, 
    
    -- channel=6
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=7
    0, 0, 0, 
    0, 0, 0, 
    0, 506, 383, 
    
    -- channel=8
    4, 0, 0, 
    0, 0, 134, 
    0, 0, 0, 
    
    -- channel=9
    0, 0, 0, 
    0, 0, 39, 
    0, 0, 0, 
    
    -- channel=10
    0, 0, 0, 
    273, 0, 0, 
    0, 0, 0, 
    
    -- channel=11
    0, 372, 0, 
    129, 766, 0, 
    0, 0, 0, 
    
    -- channel=12
    251, 0, 0, 
    0, 0, 861, 
    0, 0, 0, 
    
    -- channel=13
    698, 518, 294, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=14
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=15
    0, 498, 0, 
    0, 0, 0, 
    0, 823, 157, 
    
    -- channel=16
    0, 0, 0, 
    0, 0, 0, 
    0, 25, 0, 
    
    -- channel=17
    0, 0, 501, 
    0, 0, 162, 
    0, 0, 0, 
    
    -- channel=18
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=19
    468, 0, 0, 
    0, 121, 0, 
    781, 0, 123, 
    
    -- channel=20
    0, 0, 0, 
    0, 0, 264, 
    0, 270, 983, 
    
    -- channel=21
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=22
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=23
    0, 0, 0, 
    0, 54, 0, 
    0, 0, 0, 
    
    -- channel=24
    267, 0, 207, 
    193, 0, 701, 
    193, 0, 0, 
    
    -- channel=25
    0, 0, 0, 
    0, 571, 368, 
    453, 0, 504, 
    
    -- channel=26
    0, 142, 0, 
    0, 0, 9, 
    0, 0, 0, 
    
    -- channel=27
    184, 141, 346, 
    575, 898, 1005, 
    867, 765, 0, 
    
    -- channel=28
    0, 449, 0, 
    318, 657, 694, 
    0, 0, 0, 
    
    -- channel=29
    517, 1139, 0, 
    0, 0, 751, 
    793, 0, 97, 
    
    -- channel=30
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=31
    0, 193, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=32
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=33
    0, 0, 0, 
    0, 0, 0, 
    235, 968, 489, 
    
    -- channel=34
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=35
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=36
    153, 0, 0, 
    206, 757, 547, 
    0, 0, 0, 
    
    -- channel=37
    0, 652, 0, 
    0, 0, 0, 
    0, 821, 1487, 
    
    -- channel=38
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=39
    490, 531, 827, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=40
    235, 0, 415, 
    144, 459, 0, 
    0, 0, 0, 
    
    -- channel=41
    0, 767, 0, 
    103, 147, 0, 
    0, 0, 414, 
    
    -- channel=42
    512, 0, 350, 
    0, 0, 0, 
    0, 0, 209, 
    
    -- channel=43
    0, 0, 0, 
    0, 505, 0, 
    0, 0, 0, 
    
    -- channel=44
    300, 732, 0, 
    0, 0, 8, 
    0, 0, 437, 
    
    -- channel=45
    286, 0, 0, 
    839, 376, 540, 
    0, 0, 0, 
    
    -- channel=46
    171, 68, 987, 
    0, 0, 0, 
    0, 0, 187, 
    
    -- channel=47
    0, 0, 49, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=48
    382, 0, 219, 
    0, 154, 0, 
    847, 0, 0, 
    
    -- channel=49
    0, 0, 0, 
    0, 38, 655, 
    325, 65, 362, 
    
    -- channel=50
    179, 0, 0, 
    0, 435, 873, 
    622, 0, 0, 
    
    -- channel=51
    169, 0, 0, 
    0, 141, 0, 
    0, 372, 0, 
    
    -- channel=52
    635, 0, 0, 
    0, 39, 505, 
    0, 0, 0, 
    
    -- channel=53
    0, 0, 0, 
    829, 0, 0, 
    0, 0, 0, 
    
    -- channel=54
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=55
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 270, 
    
    -- channel=56
    0, 30, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=57
    0, 0, 1073, 
    343, 0, 0, 
    644, 216, 996, 
    
    -- channel=58
    0, 0, 0, 
    0, 0, 0, 
    899, 1369, 1442, 
    
    -- channel=59
    0, 0, 0, 
    0, 0, 0, 
    0, 341, 285, 
    
    -- channel=60
    0, 0, 359, 
    0, 121, 0, 
    0, 0, 0, 
    
    -- channel=61
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=62
    879, 0, 427, 
    196, 407, 462, 
    507, 0, 0, 
    
    -- channel=63
    460, 651, 837, 
    250, 782, 1087, 
    0, 1738, 755, 
    
    
    others => 0);
end gold_package;
