-- https://docs.xilinx.com/r/en-US/ug953-vivado-7series-libraries/BRAM_SINGLE_MACRO

library UNISIM;
use UNISIM.vcomponents.all;
library UNIMACRO;
use unimacro.Vcomponents.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use IEEE.std_logic_arith.all;

-- BRAM_SINGLE_MACRO: Single Port RAM
--                    7 Series
-- Xilinx HDL Language Template, version 2021.2

-- Note -  This Unimacro model assumes the port directions to be "downto".
--         Simulation of this model with "to" in the port directions could lead to erroneous results.

---------------------------------------------------------------------
--  READ_WIDTH | BRAM_SIZE | READ Depth  | ADDR Width |            --
-- WRITE_WIDTH |           | WRITE Depth |            |  WE Width  --
-- ============|===========|=============|============|============--
--    37-72    |  "36Kb"   |      512    |    9-bit   |    8-bit   --
--    19-36    |  "36Kb"   |     1024    |   10-bit   |    4-bit   --
--    19-36    |  "18Kb"   |      512    |    9-bit   |    4-bit   --
--    10-18    |  "36Kb"   |     2048    |   11-bit   |    2-bit   --
--    10-18    |  "18Kb"   |     1024    |   10-bit   |    2-bit   --
--     5-9     |  "36Kb"   |     4096    |   12-bit   |    1-bit   --
--     5-9     |  "18Kb"   |     2048    |   11-bit   |    1-bit   --
--     3-4     |  "36Kb"   |     8192    |   13-bit   |    1-bit   --
--     3-4     |  "18Kb"   |     4096    |   12-bit   |    1-bit   --
--       2     |  "36Kb"   |    16384    |   14-bit   |    1-bit   --
--       2     |  "18Kb"   |     8192    |   13-bit   |    1-bit   --
--       1     |  "36Kb"   |    32768    |   15-bit   |    1-bit   --
--       1     |  "18Kb"   |    16384    |   14-bit   |    1-bit   --
---------------------------------------------------------------------

entity bram_single is
    generic (
        INPUT_SIZE : integer := 8;
        ADDRESS_SIZE    : integer := 12;
        DEVICE     : string := "7SERIES";
        BRAM_NAME  : string := "default"
        );

    port (
        RST  : in std_logic;
        CLK  : in std_logic;
        EN   : in std_logic;
        WE   : in std_logic;
        DI   : in std_logic_vector(INPUT_SIZE-1 downto 0);
        ADDR : in std_logic_vector(ADDRESS_SIZE-1 downto 0);
        DO   : out std_logic_vector(INPUT_SIZE-1 downto 0)
    );
 end bram_single;

  architecture a1 of bram_single is
    signal bram_wr_en    : std_logic_vector(2-1 downto 0);
    signal bram_addr     : std_logic_vector(10-1 downto 0);

    begin
    bram_wr_en <= (others => '1') when WE = '1' else (others => '0');
    bram_addr <= ADDR(10-1 downto 0);
          

    MEM_IWGHT_LAYER0_ENTITY0 : if BRAM_NAME = "iwght_layer0_entity0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"f05b04fefa570894001d08a4112a1869fcf0deecfeba13d2188d0a4bcfa01da3",
            INIT_01 => X"001f0022000afff7ffcaffe5000000040003002c002effd30038ffffffdd0018",
            INIT_02 => X"0035002100200018ffc9ffccffc3ffedffc6ffda000bffe6001b001fffd3ffc0",
            INIT_03 => X"ffc6ffe20010fff5001700180025000fffd8ffd8fff6ffd3000700070032fff3",
            INIT_04 => X"0026001d0033ffd80006000cffcf0013fff3002000050024fffffffb000bffeb",
            INIT_05 => X"ffdffffaffc1ffdcfff4ffec000effdb003200090027ffe100060037002d0018",
            INIT_06 => X"002400120002ffe60021002dffee0016ffe7ffc6fff8fffbffc20037fffcffd2",
            INIT_07 => X"ffe6001effc20040001f000000340010fff50052001effccffe5ffc6ffe6fff6",
            INIT_08 => X"002bffeb004d002bfffaffbeffaffffcffcdfffd002b002200440039ffe1ffc2",
            INIT_09 => X"ffe100010039000b0033fffafff9002c00280026001f002f003b0045002ffffa",
            INIT_0A => X"001bffeffff0ffe60018ffe40021fff8ffd5ffd6ffd20004ffe5ffcaffc6fff4",
            INIT_0B => X"ffe9ffd600190000001c000400300033ffd6000d0044ffbefffc0005ffb3ffc1",
            INIT_0C => X"0022fff0ffd0fff50009ffe4001cffbc00100025000f0000000e002600400011",
            INIT_0D => X"0033002dffea001f00340000fff0ffcdfff6fff50009ffc9ffc4ffbbffd30021",
            INIT_0E => X"001c000affc7ffba0000fff2ffc600280015002dffff0034003c0033fff7ffcb",
            INIT_0F => X"ffc7002f0003ffdefff8fff70017ffd1ffc9ffc5fff8000afffc000b0039001c",
            INIT_10 => X"fff7ffd5fff900030002fffbfffafff80016ffc1ffc5fff0002b001effdf001d",
            INIT_11 => X"001b00170031002dfff30020003b0028ffe900290006fff7002c00270014003d",
            INIT_12 => X"00250025fff5ffd2fff1ffd8ffc8001d00100031001effe400120021ffbfffae",
            INIT_13 => X"ffe6001d0045fff3ffdcffda00350010ffcbffedffdd001cffd0fff7ffe6ffd5",
            INIT_14 => X"ffecffe0ffd9fffd0026ffe3ffe2fff900150001001f002f00160033ffea002c",
            INIT_15 => X"0033ffe5fffb0033ffc5ffdb003effe0fff9001bffd70028fff8ffd700050026",
            INIT_16 => X"0003000a004bfff3003a0030ffd8fffefff9ffc70029ffffffd7ffebfffaffdd",
            INIT_17 => X"ffc9ffd9ffdfffe40034fff9004dfffeffd6ffffffbfffec00190013003d0003",
            INIT_18 => X"001bffdbfff2ffbcffe90007ffff0036ffe8003efffb0038000f00240012000a",
            INIT_19 => X"0023002d000affe40010fffa00150029ffd1fff7fffdffd1ffdfffe000090019",
            INIT_1A => X"ffda0010fff7001affebfff5000dffdd0018ffe1ffef0013ffe4ffd200020031",
            INIT_1B => X"001400460026fff00042002bfff5ffdbffcffff8fff7ffe4ffda0023fff2ffcc",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER0_ENTITY0;


    MEM_IFMAP_LAYER0_ENTITY0 : if BRAM_NAME = "ifmap_layer0_entity0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"009e009f00a500a600a0009c00a2009f009e009f00a100a000a100a600a900aa",
            INIT_01 => X"00a700a200a000a0009c0095009600940095008f008c008d008f0089007e0074",
            INIT_02 => X"00980097009f00a600a200a000a400a200a3009c009b009f00a300aa00ab00ab",
            INIT_03 => X"00a900a0009a00970091008b008c008d009500930091008e008f0088007d0077",
            INIT_04 => X"00970097009e00a700a000a300a500a500a300a2009e009d00a100a600a700a9",
            INIT_05 => X"00aa009f00910079006e00620065007200780086008f008c008e008b00820078",
            INIT_06 => X"009b009b00a000ae00a700a700a900a900a500a500a700bf00b1009d00a200a4",
            INIT_07 => X"009e0095006800670062005c0050004a0056005300710084008c008c0088007f",
            INIT_08 => X"009b009c00a100aa00a900a300a900a600a400a400ad00f600c300970092008e",
            INIT_09 => X"006f004e005500710070006a0061005d004a0054005500690080008a00850081",
            INIT_0A => X"009400850082009300a100a500a700a700a300a500a300b4009d008000610042",
            INIT_0B => X"0045004200590076007a00770072005e0063005b003a0043006c008c008a0086",
            INIT_0C => X"007f006d002f0058009900aa00a800aa00a900a600a400930081007f00640044",
            INIT_0D => X"004e0048005300840092007c0069006b00730055003f002e004f0084008d0086",
            INIT_0E => X"00830063002a0046008f00a700a500a800ab00a1008c00780082009000740058",
            INIT_0F => X"005b0055004d007c00a300880066006a00640055003600310039006b008a0088",
            INIT_10 => X"00aa00670036007c009900a100a300a600a500ae0071007d009d009c00790056",
            INIT_11 => X"0052005400500051008a00920071005700530056004700380028004a00850089",
            INIT_12 => X"00b40086005e009a00ae009e009c009900cf00ed00cf009c00ae0094007d005d",
            INIT_13 => X"0056004a003b004c0089008f0085006a005600570054004b00320028005f0084",
            INIT_14 => X"00b7006c008e00a500b1009b009f007a00d500ed00dc00a400b7009c007d0078",
            INIT_15 => X"004e0050002d005b00af009d009b006b005700670058004e003b0029003b0068",
            INIT_16 => X"00bc0064008700aa00bb00a600ad0086007500c200c700aa00b900bd00860075",
            INIT_17 => X"006600540026007d00d200a00092005d0053005e0068005500490037003e004c",
            INIT_18 => X"00bd005a007f00af00ae00a600b2009f006100a800a8008900ba00d800a0007b",
            INIT_19 => X"007800730032009600c2009b007b005b00540054005f005600540049004f0049",
            INIT_1A => X"00bd005d009800b90077008800ad00a700670093009100a700bd00e200b4008d",
            INIT_1B => X"007e00750047009a00ba00950072005700500048005000630064005a0061005e",
            INIT_1C => X"00c2006c00a800ba00690063009c00a700640073008a00c600be00ac0091009a",
            INIT_1D => X"009200670047009800b300890082006e0055005b005f006d0073006400610075",
            INIT_1E => X"00c5008400ac00b80082004e008c009b00730082008f00e600f2009100870083",
            INIT_1F => X"0079006c005f009000a800980070005700470057006900700078006700790088",
            INIT_20 => X"00cb009200a800bf00a8004e007e008a008a0060009a00ad00a2008c00710071",
            INIT_21 => X"00650069007000ab009c00940087006d004e004f005e0065006b007d00970090",
            INIT_22 => X"00d600a300a400b700b0005e0060009c0094006a008100760072007400660073",
            INIT_23 => X"0056006500900076004400800085004b003c003a004700660074008f0096008c",
            INIT_24 => X"00d400b200a700ad00b0007c0056008d009900870068004d0086007c00810093",
            INIT_25 => X"0055005c009600840075006b004b0040002c004100560085009b00a0009a0097",
            INIT_26 => X"00c700bb00ab00ae00b1009000560077007a0089009000460081006c009100b8",
            INIT_27 => X"00740049008300890086005900330034002f005a007900a300ab00a4009e0095",
            INIT_28 => X"00a500c300b300b100b500980063008300ab0067005d0050005d007a00b200bf",
            INIT_29 => X"0096006400590057003c002e00260018002e003c006c009000900080007f0078",
            INIT_2A => X"007500c300b100b200b5008a0053009600f500db00850086009500b000be00c2",
            INIT_2B => X"00a8007d006e003d002300220031003a003d003a00450048004e0045003b0037",
            INIT_2C => X"004f00af00ae00b000b1008c006d00d300fd00fc00d0007c0072007c0074007a",
            INIT_2D => X"006800440044003c003400320033003800380033002b0033003b0030002b002a",
            INIT_2E => X"00290060009000a800b200a500a500f600fd00e3006e003c0035003100310030",
            INIT_2F => X"002d002a002e002a0026002e002e002b002a002e002e0032003700350033002d",
            INIT_30 => X"001d001d003b008300a6008400c200fe00f1008d003d00320032003300310032",
            INIT_31 => X"002f002a00270022002300270026002a002d0038003e003b00380032002e0033",
            INIT_32 => X"0030001e002200490080008000d7010000bb00420036003200340034002e002d",
            INIT_33 => X"002b00290024002700280028002b002e003b003e0040003b0036003200460053",
            INIT_34 => X"00340023001f00290042008000e000f0007c003a003100380036002c002c002f",
            INIT_35 => X"002e002b002b002c002c002d0036003a0036002e002b0024003300490055004c",
            INIT_36 => X"00320023001d0023002c004e00ca00d30061004100360030003a00300028002d",
            INIT_37 => X"002f0030002f002e0033002700270030002f0027001c002800430043002e0033",
            INIT_38 => X"00320023002000210029002e006800aa0040003600340035003d003a0036002d",
            INIT_39 => X"002a0029002e0031002e002a0028002700250028002c003f002f001f000f0033",
            INIT_3A => X"0044002a001f00260025002b002a00470031001f001b002600310038003a0035",
            INIT_3B => X"0038003c003900350032002d00270021002a003e004f004900380026000d0028",
            INIT_3C => X"003d00310023002b0027002a002c0028002a001b0017001e001b001d0024002f",
            INIT_3D => X"0038003e0042004b00450031002b002b003c0055006d005d003c001a001d0014",
            INIT_3E => X"00360038002d002b00280028002800260024001a0016001d0019001d00130012",
            INIT_3F => X"0020002f003d004a004200350034002d00430059006900590030001800220015",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY0;


    MEM_IFMAP_LAYER0_ENTITY1 : if BRAM_NAME = "ifmap_layer0_entity1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0070006f007400760070006d00730071006f00710074006f006f007500750077",
            INIT_01 => X"00750071006f0070006d006b006b006a006b0065006200610061005f005b0055",
            INIT_02 => X"0070006e0072007400700071007500720074006e006f006e0071007700750073",
            INIT_03 => X"0073006f00700073006e00680066006400690066006600610062005f005b0058",
            INIT_04 => X"006e006d006f006f006a007300750075007300730072006d006f007300720071",
            INIT_05 => X"00740072006f0060005a004e004d0055005600600067006300630062005f0059",
            INIT_06 => X"006b006e006d0070006e00750078007700730075007b00920082006f00730072",
            INIT_07 => X"0070006f00500057005a005a004b003f0046003e00550062006600650063005e",
            INIT_08 => X"006b007200730072007200710078007400710074008000d6009c0072006f006c",
            INIT_09 => X"0050003500450067006e00720066005e0048004e0049005300600065005e005d",
            INIT_0A => X"006d0068006400700073007100740073006f00740076008a007a0066004b0032",
            INIT_0B => X"003a0038005300710079007a007400600064005b003a003a005400690062005f",
            INIT_0C => X"0064005f0025004a0075007600730076007500740078006b0062006c00570043",
            INIT_0D => X"0053004b00540082008e007600630066006f00530047002f003d00620063005d",
            INIT_0E => X"00730060002b0040006f00750072007400770071006d005e006e0083006a0057",
            INIT_0F => X"005f0058004d00760099007c005d0062005d0051003c0035002f005300670061",
            INIT_10 => X"00a10069003a0079007c00710075007a0079008700590069008d008f006f0050",
            INIT_11 => X"00510055004e0047007d00870067004f004d0052004900390023003b006a0067",
            INIT_12 => X"00b0008b0064009a009500740074007600b400d600b4008300990083006e0055",
            INIT_13 => X"0054004a00390044007d0085007c0062005100550055004c0031001e004b0067",
            INIT_14 => X"00b70074009700a9009c00700076005900c500e000bf0087009f0089006c006f",
            INIT_15 => X"004c0050002c005500a5009300930064005300660058004f003b0024002e0051",
            INIT_16 => X"00bf006c009000af00a70078007b005d005f00b600ab008e00a100ab0077006b",
            INIT_17 => X"006200540026007900c90098008b00590050005d00680057004b003500370038",
            INIT_18 => X"00c20060008600b4009c007b007b006d0044009a0090007200a600ca00950071",
            INIT_19 => X"007200720032009300bb00950076005800530054005f005700570049004a0037",
            INIT_1A => X"00c0005f009a00bc006e006a007c007400480084007d009500ae00d800ac0083",
            INIT_1B => X"007500720047009800b50090006e005500500049005000640065005800590049",
            INIT_1C => X"00c4006b00a700ba006d00590077007a004a006a007b00b900b400a5008c008f",
            INIT_1D => X"008800640047009800af00850080006d0056005d0060006e007400600055005f",
            INIT_1E => X"00c5008100a700b2008900530078007d005e0078008300dd00ec008a00820079",
            INIT_1F => X"0070006800580086009f0093006c0055004800580068006d006e005600600068",
            INIT_20 => X"00cb009200a400b600aa0056007d007e00790050008f00a300980084006a006a",
            INIT_21 => X"00650065005a008f008a008d00820069004c004f005d005b00530058006c0068",
            INIT_22 => X"00d700a600a700b800b60066006000950089005d0074006900660069005b006e",
            INIT_23 => X"005b00670080006000380078007e0045003800380046005d005e00700074006e",
            INIT_24 => X"00d300b800af00b500b800830058008b00940080005a00400079006f0075008f",
            INIT_25 => X"005c0060008b0075006d00630044003b0029003e00450069007700780073006f",
            INIT_26 => X"00c000bd00b000b300b60095005a0079007c00880086003b00760061008600b0",
            INIT_27 => X"0076004b0077007c00810056003100330031005a005b007600790071006f006b",
            INIT_28 => X"009c00c100b200ad00b5009d0067008700af0069005a004d005a007600ad00b6",
            INIT_29 => X"00940064004e004d003d0034002e0021003900470064007d007b006d00710069",
            INIT_2A => X"007800c800b200a900b300900057009900f700de008c008d009c00b600c400c0",
            INIT_2B => X"00ac0085006d003e0031003600460051005500540063006500680060005c005a",
            INIT_2C => X"006900c500b700ac00b10092007000d300fc00fd00e0008f0084008d00850085",
            INIT_2D => X"007c005d00570052005400540055005d005e005b00600068006c00610061005f",
            INIT_2E => X"0059008900a800ae00b600aa00a600f500fb00e7008800580050004c004b0048",
            INIT_2F => X"004f0051005100520056005a005900570059005d005e00600060005e005f005a",
            INIT_30 => X"005b00570066009900b3008800bd00fa00f5009f005e00540054005500530054",
            INIT_31 => X"005600540052004f0053005600550059005c00670067006500660063005e0067",
            INIT_32 => X"006f005e0055006a0094008800d500fd00c6005d005b0058005a005a00530052",
            INIT_33 => X"005200510050005300560059005c005f006c006e006d006c006c0069007b0089",
            INIT_34 => X"0072006300560053005f009100e500f5008f005c0057005e005c005200520053",
            INIT_35 => X"0054005300560058005a0061006a006e00690061005f005b006c0082008a007d",
            INIT_36 => X"006e0062005900560053006a00db00e4007e0068005e00570061005700500052",
            INIT_37 => X"00540057005900590061005c005d00660065005d005500650081007e00620060",
            INIT_38 => X"006c0061005c005800580054008500c500640061005e005f0067006400600053",
            INIT_39 => X"004f00500058005c005c005f005d005c005a005d0066007d006e005a003c005d",
            INIT_3A => X"007c00640058005b00570059004f006b0059004d00470052005d00640066005c",
            INIT_3B => X"005e006300630061005f005e00580053005b0070008400830074006100400055",
            INIT_3C => X"007400660055005b005a005c00580051005500480043004a0047004900500056",
            INIT_3D => X"005f0065006d00770071005f0058005800690082009c00910073005200520040",
            INIT_3E => X"006b0069005900560059005c00570051004f00450042004900450049003f003a",
            INIT_3F => X"0046005700680077006f0060005f0057006d0083009200870063004d00540043",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY1;


    MEM_IFMAP_LAYER0_ENTITY2 : if BRAM_NAME = "ifmap_layer0_entity2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0031002f00330035002e0029002f002d002c00290029003400310029002d002c",
            INIT_01 => X"002800260027002b002c002d002d002b002c0027002b00290026002400240021",
            INIT_02 => X"00330028002d00380031002b002f002d002e0026002900360034002900280021",
            INIT_03 => X"001e00210029003200350037003400300032002e002d00260022001f00200022",
            INIT_04 => X"002f002100240030002a002c002d002d002b002b003000390033002600250023",
            INIT_05 => X"0027002f0036003100340032002f003200300037003300270023002200220021",
            INIT_06 => X"00280020001f002c002b002e00300030002c002d0039005f004b0029002f0036",
            INIT_07 => X"003a0043002f0041004c00540042003200340027002d002e002b002700270024",
            INIT_08 => X"002900300031002f002b0028002f002c0029002a003b00a4006b0038003c0047",
            INIT_09 => X"0032001f00380062006f00760069005d00430046002f002d0030002e00240024",
            INIT_0A => X"0036004000390035002c00270029002900250027002a0055004e003a002b001f",
            INIT_0B => X"002b002d004c006e0078007a0074006000610056002f00250031003a002c0028",
            INIT_0C => X"003900500011001c0030002b0028002b002a002500270034003b004b00460039",
            INIT_0D => X"00480040004a00790084006c005a005e0067004d004500270024003a00300027",
            INIT_0E => X"005a005c002600290038002a002400270031003300330031004d006b005d004f",
            INIT_0F => X"005800520045006b008c0070005100580054004a003a00310020003200330027",
            INIT_10 => X"00900069003b00710052002b002900320042005f003b004e007900800065004a",
            INIT_11 => X"004d00520049003d0070007b005d00460045004c00430035001b0023003b002d",
            INIT_12 => X"00a3008f0069009500700033002f003c009200c600a600770091007d006b004f",
            INIT_13 => X"004f00470035003a0070007a00720059004a004e004e0047002b000f002c0039",
            INIT_14 => X"00af007a009e00a8007a00320033002f00b300e200bc0083009b008400680068",
            INIT_15 => X"0045004d0028004d009a0089008a005c004d0060004f0049003b0021001f002e",
            INIT_16 => X"00bd0074009900b20088003b0037002c005000bc00a400850097009f006a005f",
            INIT_17 => X"0059004f0022007100c0008e00820052004b0058005e0051004e00370030001a",
            INIT_18 => X"00c20069009000b9008500440035002f002c0098007e005e009400b700810062",
            INIT_19 => X"0069006d002f008c00b2008c006f0053004f0050005500510059004900400018",
            INIT_1A => X"00c1006700a300c000620042003a0032002700780067007f009b00c8009d0075",
            INIT_1B => X"006b006d0044009300ae008800680050004c00460048005e0063005100450022",
            INIT_1C => X"00c4007000ac00bc006d0043003e003700220058006700a900a9009f008c0086",
            INIT_1D => X"007d005f0046009500aa007f007a00690053005b005a0068006f00500035002f",
            INIT_1E => X"00c5008800ae00b5008e004d0058004d0034005d007400d300e6008900820070",
            INIT_1F => X"0065005f004b00760092008a006500500044005700630063005d003600300030",
            INIT_20 => X"00cc00a000b200bc00ac005a007e0071005200250085009b008d00750058005a",
            INIT_21 => X"005c0057003a0068006d007e007600610048004d005e00520037002d0037002e",
            INIT_22 => X"00d700b400b800c200ba006900660091006f003d0069005f0059005900490062",
            INIT_23 => X"0058005f00660040002000690073003d003300350041004e0040004400400036",
            INIT_24 => X"00cd00c000bd00c100bc00850060008f008d006f00500037006c006000640085",
            INIT_25 => X"005d005d0078005d005c0056003a00340027003c0028003b003e0036002d002e",
            INIT_26 => X"00b400bb00b500b900b800980063008400820087007e0033006c0056007b00a8",
            INIT_27 => X"00760049006700690076004e002c00320034005d003c0044004000340032002e",
            INIT_28 => X"009200bb00af00ac00b400a0006f009200b9006f005700490056007400ad00b1",
            INIT_29 => X"009400650042003f003900360033002900450053004b0052004c003d0045003f",
            INIT_2A => X"007c00c800b000a800b30093005b009f00fa00e10090009300a400c000d000c5",
            INIT_2B => X"00b5008f006d003e003a004400570066006e006f007a00770078007000700073",
            INIT_2C => X"008500d500c000b100b60096007100d100f700fc00e8009d009500a2009c0098",
            INIT_2D => X"0094007700680065006f006e0073007d008300820087008d008e008400890084",
            INIT_2E => X"008700a800bc00bc00c000ae00a400ed00f100e40099006f00690069006b0065",
            INIT_2F => X"0073007800710074007d007d007e00800084008b0089008900870086008b0085",
            INIT_30 => X"008d0082008600b000bf008900b500f200f500af007f00760077007900780074",
            INIT_31 => X"00750075007300710078007d007d008200860091008e008e00920090008c0095",
            INIT_32 => X"00a2008c007c008800a7008f00d100f900cd00760080007d007f007f00790073",
            INIT_33 => X"0071007000710075007b00830086008a0096009800930095009a009800a700b6",
            INIT_34 => X"00a500930082007a007e00a400ea00f700990072007b00830081007700770077",
            INIT_35 => X"00770077007b007f0083008d0096009a0096008d008c008a009e00b200b600a9",
            INIT_36 => X"00a20095008a0085007e008a00e900ea008c007e0081007c0085007b00740077",
            INIT_37 => X"007a007e00820084008c008a008b00940093008b0085009900b600b0008e008b",
            INIT_38 => X"00a10093008f008d008a007d009f00d30077007900800082008b008700830078",
            INIT_39 => X"00760078008200870088008b008a00880087008a009700b200a4008c00670088",
            INIT_3A => X"00b1009400890092008b00840071008500720069006900750080008700890080",
            INIT_3B => X"00830089008b008a008900880083007d0085009a00b300b500a80092006c007f",
            INIT_3C => X"00a800940084008f008b0086007d0070007300680066006d006a006c00730078",
            INIT_3D => X"008000870090009c00980086007f007f009000aa00c500be00a40082007e006b",
            INIT_3E => X"00a000950084008600860084007b0073007200690065006c0068006c00620059",
            INIT_3F => X"0064007600890098009100830082007b009100a700b600af0091007c0081006e",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY2;


    MEM_GOLD_LAYER0_ENTITY0 : if BRAM_NAME = "gold_layer0_entity0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00120012000f00140017000d000f001d001d000a000000010006000c00150016",
            INIT_01 => X"0012000f00130013000400080003000000040000000000000005000b0000000b",
            INIT_02 => X"0013001b0012001b0020001e000000000000000000000000000100010000000c",
            INIT_03 => X"0019000b00110000000000000000000000000000000000000000000000030003",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_05 => X"0000000000000000000000000001000000000000000000000004001c00000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000002000000000000",
            INIT_07 => X"0000000000000000000000000000000b000000000000000000000000000b0000",
            INIT_08 => X"000000000000000b000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000b00000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000200000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"000b000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"00000000000000000000000000000000000000000000000000000000000d0000",
            INIT_16 => X"0000000000000000000400070000000000000000000000060000000000000000",
            INIT_17 => X"0000000000010000000000000000000000000000000000000000000000000000",
            INIT_18 => X"000000000000000f001a000f003f000a0000000000000032003a003800250020",
            INIT_19 => X"00220029002500270020002c003a00000000001e001d001d00200020001f0024",
            INIT_1A => X"001e0022002800210030002f002f000e000f00210019001d00220023002f0033",
            INIT_1B => X"00340028003a0029003300310041002a0030002a001f0017001c0021002d001a",
            INIT_1C => X"001c002900000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000030018000e00060000000000000000",
            INIT_1F => X"000b0000000000000000000200010000001b000000060000000000000000001e",
            INIT_20 => X"0000000000110014000500030000001d00100000000800000003000f00170000",
            INIT_21 => X"0000001a000a000600040000004400030000000b000000020017000b00000000",
            INIT_22 => X"000c001e000b00000000003700000004000a0011000200200014000600000006",
            INIT_23 => X"002d000000000000002000000000001100080000001d00280004001100080000",
            INIT_24 => X"0000000b000b0000001000000006000000000018002400000027000e00090012",
            INIT_25 => X"00120015000000000000000c00000000002b002300000058000d0028002d0011",
            INIT_26 => X"00000000001b0022001f000b0000003600230012004500000007001f0021001a",
            INIT_27 => X"001e00220028002e002f002f002a00380033002500000027002500240024002a",
            INIT_28 => X"002f0036002f002e003a002c002e005200000013002b0026002a002a002f002e",
            INIT_29 => X"002f002a00450028002b0033002c00190019002800230024002e0031002d002e",
            INIT_2A => X"0043003a001f0000000000000000000000000000000000000002000a00000000",
            INIT_2B => X"000000000000000000000000000000000010000800170000001f001c00030000",
            INIT_2C => X"0000002a00000000000000000000002b0011000000000042002d003f00000000",
            INIT_2D => X"0071000000000000000e00000028002c00250000005a0026003b002a0000006c",
            INIT_2E => X"00050023000000340024005d0048003c0000002f0052001e003e000000590031",
            INIT_2F => X"003700000000002c0061003e006000000073005c001200310025004800730015",
            INIT_30 => X"003800000000005a004a006a0000007500470012000c0037004d006500280031",
            INIT_31 => X"00000006008b003800460000004f0050000600250013006800420084000b002a",
            INIT_32 => X"0013002e002c000000290016005b000400000000004a003a009f000000640018",
            INIT_33 => X"0000004d0030003b005a001700000000000c000f003c009400000093004c0020",
            INIT_34 => X"007100830041001a001d002300200031001d002b004e000000d80073003a003c",
            INIT_35 => X"00470038003d003c003e0040004f005f00120000008200af00420049003f003e",
            INIT_36 => X"00390038004000500048003d006a0045000000cb005a0039004d0042003c0041",
            INIT_37 => X"0048004d004e0038007b0076004b003e00540048003500430044003800440055",
            INIT_38 => X"003a001a006f0080000000000008000800060003000500000004000000000000",
            INIT_39 => X"0000000600050007000a000c0007000a0049001a000000000000002400060000",
            INIT_3A => X"0000000400000000000400040007000000000000000d001a0015000700170000",
            INIT_3B => X"00000028002500090005000d00000037001b0005000000000000000000010000",
            INIT_3C => X"0026005a0013000b008000560006000e0000000000250025000f001800000000",
            INIT_3D => X"00000008000000000000002a001a001f003a0000000000000009002700060007",
            INIT_3E => X"00000004000000210000000a000900110000000b00000017001d00150007001c",
            INIT_3F => X"00100019001600000000000000000000000000000000000000100004000b0004",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY0;


    MEM_GOLD_LAYER0_ENTITY1 : if BRAM_NAME = "gold_layer0_entity1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"001c00000000001a000400000000000000000003002f00000000000900040011",
            INIT_01 => X"00000000004a000c000000000000001b001f00000000000000000046009c0085",
            INIT_02 => X"002800000000000000200041001b0000000000000000000f0046000000000000",
            INIT_03 => X"0000000000000000000000000000000000020000000000000000000000000000",
            INIT_04 => X"0000000400070012000000000011000000000000000000000000000800000000",
            INIT_05 => X"0000000000000000001300000000000000000000000000000000000000140013",
            INIT_06 => X"00040000002800220000009d00a300a200a500a4009d00ac00b700ad0094007c",
            INIT_07 => X"007c00840092009200a200ad00a800ac00a0008c00a900a0007a003a002e003e",
            INIT_08 => X"004e006e008b0089006a00ac00b000af008e00730048002d0007001e000a0027",
            INIT_09 => X"003a0067004d002b00a400aa00a20059004d00270015000c0033002d001b0025",
            INIT_0A => X"003a0017001f00940060004e00470043002f001f0000003100390017001c002f",
            INIT_0B => X"00160012008e00990025003b00450031002d0000003e002a001000120017000e",
            INIT_0C => X"002a0062009f002f0032003e002d002f0000003200280010000e0026001c000a",
            INIT_0D => X"002c006200370026002e00270029001e002f002d00090022004100140000002b",
            INIT_0E => X"000e0055002200360030000d005400420026000f002d00790010000500240000",
            INIT_0F => X"0035002000080028002d0034001d000600090062008a00000015002300000017",
            INIT_10 => X"001a0000000000060000000000000000000000000000000000000006003a0000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000034000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000022002300250020001e002700260024001d0017",
            INIT_15 => X"001a00260024001e00180023002c002a001f00280020000f001d000e001d0000",
            INIT_16 => X"00090020002b001c00060039002800210027001a000000060021002e00000000",
            INIT_17 => X"00000025002c0000004c00210029000f00240004000000000048000000090000",
            INIT_18 => X"0000004a00000026000200560009000b00000000000000590000000000060000",
            INIT_19 => X"002b0000000a0000001a003e0013000000000000008e00000000001400000000",
            INIT_1A => X"0000000000200000003f0036000000000000006600000000000a001500000000",
            INIT_1B => X"00000000000000380042000000000000004200000000001d000f000800000002",
            INIT_1C => X"0000002100040011000000000024000000250000001e00210023000000000000",
            INIT_1D => X"002c0000000f00270000000200050000000c003000340014002a000400000078",
            INIT_1E => X"0000000000220000000000000008000900010000000000200014000000400000",
            INIT_1F => X"0000000000000000000000000000000000000000000000210043000000000000",
            INIT_20 => X"00000000000000000000000000000000000000000000005d0000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000400000000002b0030002d002c002f00290030003a0037",
            INIT_23 => X"002a002500260027002a0031002c00350030002e002d0000001f0029003b000c",
            INIT_24 => X"00000000000e001f0025001c0029002e00350032003b002d0023000000000000",
            INIT_25 => X"000000000004001a000000000023003200250019000000000000000000000000",
            INIT_26 => X"0006000000110000000000120018000000000000000000000000000000000000",
            INIT_27 => X"0000000500000000000b00380003000300000000000000000000000000000000",
            INIT_28 => X"0000000000000007003a00070000000000000000000000000000000000000000",
            INIT_29 => X"00000000000000000002000000000000000000000000000000000000000d0000",
            INIT_2A => X"0000000000000000001a000500000000000f0003001800040000000800000000",
            INIT_2B => X"000000000000000000000000000000080011000a00000000001f000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"00000000000000000000000000000000000a0011000800080004000c000c000b",
            INIT_31 => X"000b0021002d00230011000800060000000a000a000c00080000000500230042",
            INIT_32 => X"000000000000000a0017000a0035003300050008000500370016000900000000",
            INIT_33 => X"000000000000000e000c000000000005000800080000000000020000001a0004",
            INIT_34 => X"001000060000000e000100000002000e00000000000900000007000000000000",
            INIT_35 => X"000000000000000f000000060003003e00280000000000000000001400150007",
            INIT_36 => X"0000000000000000001c00180012000000310000001100000011000000000000",
            INIT_37 => X"000000000000000000000002003500350021000e0000000900000005000e0000",
            INIT_38 => X"000000010000000000000026000000000000000000260030000000000000000c",
            INIT_39 => X"00000004000000230009000000000000004e0036001100000000001800030000",
            INIT_3A => X"0007000000000000001e0051003700000000000000000005000a00350021000c",
            INIT_3B => X"0000005600280004000500030000000000000000000000000000001600000018",
            INIT_3C => X"003f0000000000000000000000000000000000000000000000000018004f000b",
            INIT_3D => X"0000000000000000000000000000000000000014000000000000002200000003",
            INIT_3E => X"001200000000000000000000000000000000000d0013000a000e000900150008",
            INIT_3F => X"0006000c001c0022001b0013000600020008000b0009000d000f0036000f001a",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY1;


    MEM_GOLD_LAYER0_ENTITY2 : if BRAM_NAME = "gold_layer0_entity2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"001f0034003500240021001a000a00260024000b000a00080051003300280020",
            INIT_01 => X"0053005e004b002b0019001a00330014000e00120019002e0045002f0036005b",
            INIT_02 => X"005d0042003b0015001b0071005e00150035007e00440064003b0033003b0067",
            INIT_03 => X"0038003900250001007f009e0028001300bd007e007d004b002e005b007f0050",
            INIT_04 => X"0047003c0015007a009400430017005a007500a80065004e007800810046003b",
            INIT_05 => X"004c0033008e00a500400039003900a50085006a0050005f0078004c0048004b",
            INIT_06 => X"002600b000b800660073003800660059004e0051003300650041002c002b000e",
            INIT_07 => X"00c000b300860075006f0033005f00790042005a00400025002f0027002700c7",
            INIT_08 => X"00ab008b00a2009e0065009100b90079003c00400047005a0071006800c100cb",
            INIT_09 => X"009d00c900e700a5008a0085007c006f007800800088008a008e008c00a100b1",
            INIT_0A => X"00e500af007a00750070007100760084008c0095009a00a3009d008500a600ef",
            INIT_0B => X"008800800079007300770082008c009b009300a300ab0097008f007f00a70074",
            INIT_0C => X"007f0089007e007c008800860085009a00af008d000000000000000000000000",
            INIT_0D => X"0000000000000013001c000b000000000000000000000000000000000000000b",
            INIT_0E => X"00140033000000000014001e00000000003f0000000000000000003e001c0028",
            INIT_0F => X"00000000000000000007001e00000019000000000000000c0000000000000000",
            INIT_10 => X"00000000001a0006000e0000000000000009000000000000000f0004001d0000",
            INIT_11 => X"00000008000000000025002f00000002004f0003000000000000000600000026",
            INIT_12 => X"001c00000000000000000018000d000d00000000000500000009000000180008",
            INIT_13 => X"000000000000000200000007000000000000003d001e000000000000001c0000",
            INIT_14 => X"0010000000000000002e00000022003200030000000000360026003a000d0000",
            INIT_15 => X"000000000000000a00000012001500000000002e001f00310001000000000008",
            INIT_16 => X"00000000002200000000000000000019000f000d000000000000001600210041",
            INIT_17 => X"00000000000000a20052003f0037000c000600000002000000000000000d0036",
            INIT_18 => X"0000004100560000000200000000000000000000000300000000000200000025",
            INIT_19 => X"003e0006000000000001000000000007000a000000000042000c000000180036",
            INIT_1A => X"0024001300090000000000000005000000000000000400000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"00000004001f000000000000000000000000000b000000000000000000000000",
            INIT_1E => X"0005002d00000007000000020001000000020000000000000000000000000002",
            INIT_1F => X"003b000000000003000000100001000600000000002c0000000000000000005d",
            INIT_20 => X"00000000000e000000000000000000000000001c000f00000000000000520000",
            INIT_21 => X"00000012001300000004000000000000000c0017000000050000002d00000000",
            INIT_22 => X"001d00030000000000160000001100000012000000000008000000110000001b",
            INIT_23 => X"00000000000900190000003b0000000300100000000500000000001200120000",
            INIT_24 => X"00000033000d0000005800000000002d00040000000200280033003e002c001d",
            INIT_25 => X"007000360000003b0000002e004e004e00440049004f00560058005a0053005a",
            INIT_26 => X"006f00480008000000490048004a004c0054005b005b0057005d005e005a0060",
            INIT_27 => X"008a0000003100500045004d005300570061006400610074005e005000670067",
            INIT_28 => X"00410049005f00550049005200520052005e006b00530045002f002e0033002e",
            INIT_29 => X"002f002f0031002f002b0023001c0027002600270024003200320035002d0034",
            INIT_2A => X"00550013002500040021001300150024002d0028001a003b0034002e0038002c",
            INIT_2B => X"00000000001a004f000a000b00040027003900000079002c003600250023001a",
            INIT_2C => X"000800180053000000120000000e005300000063000a0049002c001a00000000",
            INIT_2D => X"0008005f000b0000001e00000039000000380000002e00490000000000000000",
            INIT_2E => X"00bf0000000000230004000d00000015000c000000610050000a0000000000a4",
            INIT_2F => X"00000000001e0027000d000000000001000000450068000000080000007c0000",
            INIT_30 => X"0000002a00220012000000170000003c001100030000001c0031000600220000",
            INIT_31 => X"0026003a0044000a00180000004a00000019002a000e0017000a000000050048",
            INIT_32 => X"0056001c00510011000000a30000000b005600000000000000140028002d001e",
            INIT_33 => X"0000004000280000009800000000000000000000000900100010000e00110000",
            INIT_34 => X"000300410048001f000000090005000a00080010001400170010000800170000",
            INIT_35 => X"0010007400000000001100000009000d0010000d00090000002600000000000d",
            INIT_36 => X"0019000000000016000c0009001800100000000b003100030000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000400000000000000000001000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000400120000000000000000",
            INIT_3A => X"0005000000000000000000000000000000000001002700000000003800080000",
            INIT_3B => X"0000000000000000000000000004000000000000000000000000000000000000",
            INIT_3C => X"000000140000000000000000000f000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000120000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY2;


    MEM_GOLD_LAYER0_ENTITY3 : if BRAM_NAME = "gold_layer0_entity3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"001100000000000000000000001e0030003e0000000000000000001c00240001",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000002",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"00000000000000000000000000000000000000000000001300000000002f0036",
            INIT_05 => X"00330035003500300039003b0036002b00200020002500280027003000380036",
            INIT_06 => X"003900330042003b003900230002000200060006001100270030001300360039",
            INIT_07 => X"0037003d001e0000000000000004000000010000001700150000003200370040",
            INIT_08 => X"0012001e00000000000000170000000000000000000000120034001000440033",
            INIT_09 => X"0025000600000000001000090000000000000000000f00310038000b000d002b",
            INIT_0A => X"0008000b0000002a00000000000000000000002c0007003d000e0011002e0017",
            INIT_0B => X"0008000300130000000000000000000400190000002500000022002e000a0000",
            INIT_0C => X"0013000f00000000000200000015001100090000001c00000000000c0000002c",
            INIT_0D => X"000000000000000000210016000e00140000000300000000001f000600050000",
            INIT_0E => X"00000000001e00280005001400150000002c0006001100170000000000000000",
            INIT_0F => X"0000000000000000000000000032003c00000000000000000000000000000000",
            INIT_10 => X"00000000000000000000004f0000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000002800000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000027",
            INIT_13 => X"002200230029002c00200028002b002f00320029001d001e0029002e00280024",
            INIT_14 => X"0024002c0021000e00430030002e00050021002900190015002c003f00020028",
            INIT_15 => X"0029002a00200028002400100000001c000c0032001a000b005c0000002e0024",
            INIT_16 => X"0038000c002700250019000000230018001a00260000002c0005004100000013",
            INIT_17 => X"0027002a002400250000001400380012002b001a002400000037002f00000000",
            INIT_18 => X"00160025004300000034002a0007001d002000110024000e0046000000000015",
            INIT_19 => X"001c00390000002b0028000d00000025000b000600290034000200000035000b",
            INIT_1A => X"001800000011002c00000011000d000d0000003f000000340000000e001b0000",
            INIT_1B => X"003f0005002b00000000001a0000000000390000002a00140000001d002c000f",
            INIT_1C => X"002f000f00000010002f000000000038000000290032000000050027002b000f",
            INIT_1D => X"0008000800110021000000000000000000520005000000000000000700030000",
            INIT_1E => X"0000000000030014000000000022002e00000006000200050001000000000002",
            INIT_1F => X"000000000009000000000022000d000000090006000000000001000000000000",
            INIT_20 => X"00150013000000000004001400000000000000000000000c000000000012001a",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY3;

    MEM_EMPTY_18Kb : if BRAM_NAME = "default" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST"      -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate;


end a1;