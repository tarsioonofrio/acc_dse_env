library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 4000000) of integer;

  constant input_wght : mem := (
    -- bias
    -2120, -710, -196, 2784, 2029, -2302, 679, -74, 893, -1124,

    -- weights
    -- filter=0 channel=0
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 2, 0, 0, 0, 0, 1, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 2, 0, 0, 1, 1, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 2, 1, 1, 1, 1, 1, 2, 1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -2, -2, 0, -1, -1, 0, 0, 1, 2, 0, 0, 0, 1, 0, 0, 1, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, -2, -1, 0, -1, -1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -1, -1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -2, 0, -2, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 0, 1, 0, 0, -1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -2, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, -1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -2, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -2, 0, -1, -2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 1, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 2, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, -1, 0, 0, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, -1, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, -1, 0, -1, -1, -1, -2, -1, -1, 0, -1, -2, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -2, -2, -2, -1, -1, -1, -1, 0, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, 0, -1, -1, -1, -3, -1, 0, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, -2, -3, -2, -1, -1, -2, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -3, -2, -2, -1, -2, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, -2, -1, -1, -2, 0, 0, -2, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -2, -1, -1, -2, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -2, -2, -2, 0, 0, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, -3, -2, -1, -1, 0, -2, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -2, -1, -1, -1, -3, -2, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -3, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -2, -1, -2, -1, -1, -1, 0, -2, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -3, -3, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -1, -2, -2, 0, -1, -2, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, -2, -2, -2, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -2, -1, -1, -1, -1, -2, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -2, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, -1, -1, 0, -1, -1, -2, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -2, -1, -1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 2, 1, 1, 2, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 3, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 3, 1, 3, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 1, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 2, 3, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 2, 2, 2, 1, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, 1, 0, 1, 1, 0, 0, 1, 1, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 1, 1, 1, 1, 1, 2, 0, 2, 2, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 2, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 2, 1, 2, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 3, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 1, 2, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 2, 2, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 2, 1, 2, 2, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 1, 0, 1, 1, 1, 1, 1, 1, 0, 1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 2, 0, 1, 1, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 2, 1, 0, 3, 1, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 2, 0, 2, 2, 1, 0, 0, 1, 1, 0, 0, -1, -2, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, -1, -1, -1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 1, 2, 2, 1, 1, 2, 1, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, -2, -1, -2, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 2, 2, 2, 2, 1, 2, 0, 0, -1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, -1, 0, 0, 1, 0, 0, 1, 0, 1, 2, 1, 2, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 2, 2, 2, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 2, 2, 1, 0, 0, 3, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 2, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 2, 1, -1, -1, 0, 0, 0, 1, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 1, 0, 0, 1, 0, -1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 1, 1, 1, 0, 2, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 1, 0, 0, 0, -1, -2, -2, -2, -1, 0, 0, 0, 0, 1, 1, 2, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -2, -2, -2, -2, -1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -2, -3, -3, -2, -2, -1, 0, 0, 0, 1, 0, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, -1, -2, -3, -1, -1, -1, -1, 0, 1, 2, 1, 2, 1, 2, 1, 0, 0, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -2, -1, -1, -1, -1, 0, 0, 1, 1, 2, 1, 2, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -2, 0, 0, 1, 1, 0, 0, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, -1, -2, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 1, 2, 1, 2, 2, 2, 1, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 2, 2, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 2, 2, 2, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, -2, -1, -1, 0, 0, 0, 1, 2, 2, 1, 1, 0, 1, 1, 0, 1, 0, 2, 1, 1, 2, 2, 1, 2, 0, 0, -1, -1, -1, -2, -3, -3, -1, 0, -1, 0, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 3, 2, 3, 3, 2, 3, 1, 0, -1, -1, -2, -2, -2, -2, 0, -1, 0, 1, 1, 1, 1, 0, -1, -2, -2, -2, -3, -3, -1, -1, 0, 1, 3, 4, 3, 5, 6, 4, 1, 0, 0, -1, -2, -1, -2, -1, -1, 0, 1, 0, 0, 1, 0, 0, -2, -2, -3, -3, -4, -4, -2, -2, 0, 0, 2, 3, 4, 6, 5, 5, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, -1, -3, -4, -3, -2, -2, -2, -1, 0, 1, 4, 5, 5, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, -2, 0, 0, 0, 1, 2, 5, 4, 4, 3, 0, 0, 1, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 3, 4, 3, 2, 1, 1, 1, 3, 2, 0, 0, 0, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 1, 0, 2, 1, 3, 2, 2, 1, 1, 1, 1, 2, 3, 1, 1, 1, 0, 0, 1, 1, 1, 0, 1, 1, 1, 1, 1, 0, 1, 1, 0, 0, 1, 2, 2, 1, 2, 1, 2, 1, 2, 3, 3, 4, 2, 2, 1, 1, -1, -1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 2, 2, 1, 1, 1, 0, 1, 2, 1, 3, 3, 3, 3, 1, 1, -1, -1, 0, 1, 2, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 2, 2, 1, 1, 0, 1, 1, 1, 1, 2, 3, 3, 4, 3, 3, 2, -1, 0, 0, 1, 1, 1, 0, 1, 1, 1, 1, 1, 2, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 3, 4, 3, 5, 3, 2, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 3, 3, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 2, 1, 3, 3, 4, 4, 5, 4, 2, 0, 0, 0, 1, 1, 1, 1, 0, 1, 3, 4, 3, 3, 2, 2, 1, 0, -2, -2, -1, -1, 0, 0, 1, 2, 3, 4, 4, 4, 5, 3, 2, -2, 0, 1, 1, 1, 0, 0, 1, 1, 3, 4, 3, 2, 2, 2, 1, 0, -3, -2, -3, -2, -1, -1, 0, 2, 4, 3, 5, 4, 4, 3, 1, -2, 0, 0, 1, 2, 1, 1, 1, 1, 3, 3, 3, 1, 2, 0, 0, 0, -2, -3, -4, -2, -1, 0, 0, 2, 3, 4, 4, 4, 4, 4, 3, 0, 0, 1, 2, 2, 1, 1, 1, 2, 2, 3, 3, 1, 0, 0, 0, 0, -2, -4, -2, -2, -2, 0, 0, 2, 3, 4, 4, 4, 6, 4, 3, -1, 0, 0, 2, 2, 1, 1, 1, 0, 1, 2, 1, 0, -1, 0, 0, 0, -1, 0, -2, -1, 0, 0, 2, 2, 4, 5, 5, 5, 5, 3, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 2, 1, 0, -1, 0, 1, 1, 0, 0, 0, 1, 0, 1, 1, 3, 2, 4, 3, 3, 4, 3, 2, -1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 3, 2, 2, 1, 1, 4, 2, 3, 1, 1, 0, -1, 0, 2, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 3, 1, 1, 2, 1, 2, 2, 2, 2, 1, 1, 3, 3, 2, 1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 3, 2, 2, 1, 2, 0, 1, 3, 1, 2, 1, 2, 1, 1, 2, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 2, 2, 0, 0, 2, 2, 3, 3, 3, 2, 2, 1, 0, 0, 1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 2, 4, 2, 2, 2, 1, 2, 2, 2, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 1, 1, 1, 0, 3, 3, 3, 3, 2, 1, 2, 2, 1, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, -2, -1, 0, 1, 2, 0, 1, 3, 3, 3, 4, 2, 1, 2, 1, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -2, -2, -3, -1, -1, 1, 1, 2, 3, 3, 4, 4, 3, 1, 1, 1, 1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -2, -2, -2, -2, -3, -1, -1, 0, 0, 2, 1, 3, 4, 4, 2, 2, 1, 1, 0, 0, 0, -2, -2, -2, -1, -2, -2, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 1, 1, 3, 3, 2, 1, 1, 0, 0, 0, -1, -3, -3, -2, -1, -1, -2, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, -1, 0, -1, -4, -4, -2, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, -2, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 2, 0, 1, 1, 1, 2, 0, 0, 0, 0, 0, -2, -2, -1, -1, -2, -2, -3, 1, 1, 1, 1, 1, 1, 2, 2, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 2, 1, 0, 0, 0, 1, 0, 0, -1, -2, -2, -3, -4, -2, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 1, 0, 0, 1, 0, 0, -1, -2, 0, -1, -3, -1, 1, 0, 2, 0, 0, 0, 1, 1, 1, 0, -1, -1, -1, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, 2, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 1, 2, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, -2, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 0, 1, 0, 0, 0, -1, 0, 0, -1, -2, 0, 2, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 2, 2, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 2, 1, 0, 1, 2, 1, 1, 2, 0, 0, 0, 0, -2, -1, 0, 0, 1, -1, -2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 1, 2, 0, 2, 1, 3, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 2, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 2, 1, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 1, 1, -1, 0, 0, 0, 1, 2, 1, 1, 2, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 1, 2, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 3, 2, 2, 1, 1, 2, 1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, -1, 1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 2, 1, 2, 2, 1, 1, 0, 1, 0, 0, 0, 0, -1, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 1, 1, 2, 2, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, 1, 2, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 2, 0, 2, 0, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 2, 1, 2, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 2, 0, 0, 0, 1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 1, 2, 2, 1, 3, 2, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 1, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, -1, -3, -3, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, -1, -1, -1, -1, -2, -3, -2, 1, 1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, -1, -1, 0, -2, -2, -3, -3, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, -2, -1, -2, 1, 1, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 1, 2, 2, 2, 2, 2, 3, 2, 2, 2, 1, 1, 1, 0, 0, 0, -1, -1, -2, -2, 1, 2, 2, 3, 1, 1, 3, 2, 1, 0, 0, 1, 1, 1, 3, 3, 4, 5, 6, 4, 3, 2, 2, 3, 0, 0, -2, -2, -2, -4, -6, -5, 2, 2, 2, 2, 2, 3, 3, 2, 0, 0, 0, 0, -1, 0, 0, 1, 2, 4, 5, 6, 4, 4, 3, 4, 1, 0, -1, -2, -3, -4, -5, -5, 1, 3, 2, 1, 1, 0, 2, 1, 0, -1, -3, -3, -4, -2, -1, 0, 1, 4, 4, 5, 4, 5, 6, 5, 4, 0, 0, 0, 0, -1, -3, -4, 1, 2, 1, 2, 0, 0, 0, 1, 0, -3, -3, -5, -4, -4, -2, -1, -1, 2, 2, 3, 5, 6, 6, 6, 4, 1, 1, 0, 2, 0, -1, -2, 3, 2, 1, 1, 0, 0, 0, 0, -1, -2, -3, -3, -3, -3, -2, -1, -1, 0, 2, 3, 5, 6, 6, 6, 4, 1, 1, 2, 2, 0, -1, -2, 1, 4, 1, 2, 1, 0, 1, 0, 0, 0, -2, -2, -1, -1, -1, -1, -1, -1, 1, 3, 5, 6, 5, 5, 4, 1, 1, 4, 3, 3, 1, -1, 2, 2, 2, 3, 2, 1, 2, 0, 1, 0, 0, 0, 2, 1, 0, -2, -1, 0, 2, 4, 3, 5, 4, 4, 2, 3, 2, 5, 5, 3, 1, 0, 2, 2, 1, 3, 2, 1, 2, 1, 0, 0, 1, 1, 3, 2, 1, -1, -1, 0, 2, 3, 4, 3, 2, 2, 2, 3, 4, 5, 5, 4, 2, 0, 2, 2, 1, 2, 2, 2, 2, 1, 0, 0, 0, 3, 4, 4, 0, -1, -1, 1, 0, 1, 1, 1, 1, 1, 3, 3, 5, 4, 6, 5, 3, 0, 1, 0, 1, 1, 1, 3, 3, 3, 1, 2, 3, 2, 2, 2, 1, -1, -2, 0, 0, 0, 1, 0, 2, 2, 3, 3, 3, 5, 5, 4, 2, 0, 0, 0, 0, 1, 0, 1, 3, 2, 1, 2, 3, 3, 2, 1, 0, -3, -2, -1, -1, 0, 0, 0, 0, 3, 2, 3, 4, 4, 6, 4, 4, 0, 0, 0, 0, 0, 1, 0, 2, 4, 3, 3, 4, 5, 3, 0, -1, -2, -4, -3, -4, -3, -1, 0, 1, 3, 3, 3, 5, 5, 6, 5, 3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 6, 6, 5, 3, 0, -1, -3, -5, -5, -5, -5, -3, -2, 1, 3, 4, 4, 4, 5, 6, 5, 2, 0, 1, 1, 0, 2, 1, 1, 1, 1, 4, 6, 7, 6, 4, 1, -1, -3, -5, -7, -7, -7, -6, -4, 0, 3, 4, 5, 6, 6, 4, 5, 2, 1, 1, 1, 0, 2, 0, 0, 2, 2, 4, 5, 7, 5, 3, 1, -1, -3, -6, -8, -7, -7, -7, -4, -1, 1, 5, 7, 7, 6, 4, 4, 4, 0, 2, 1, 1, 2, 1, 0, 1, 1, 3, 5, 6, 4, 2, 0, -1, -4, -6, -7, -7, -9, -6, -5, -1, 2, 5, 7, 7, 7, 5, 5, 2, 1, 2, 1, 0, 1, 1, 1, 1, 2, 3, 4, 5, 4, 1, -2, -4, -4, -6, -6, -8, -7, -5, -2, -1, 2, 5, 6, 7, 6, 5, 4, 4, 0, 1, 1, 0, 1, 0, 0, 0, 1, 3, 4, 4, 2, -1, -3, -4, -3, -3, -4, -5, -5, -3, -1, 0, 2, 5, 6, 5, 6, 4, 4, 2, 1, 2, 2, 1, 0, 0, 0, 0, 1, 3, 4, 3, 2, 0, -3, -2, -3, -1, -3, -2, -3, -1, 0, 1, 4, 5, 5, 5, 5, 5, 4, 1, 0, 1, 2, 0, 0, 0, 0, 0, 1, 3, 3, 2, 1, 0, -1, 0, -1, -1, -2, -1, -1, 0, 0, 2, 4, 5, 4, 5, 5, 4, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 2, 4, 4, 4, 5, 4, 3, 3, 0, 0, 2, 2, 1, 1, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 1, 3, 3, 4, 5, 4, 5, 4, 3, 2, 0, -1, 0, 1, 1, 0, 0, -2, -1, 0, 0, 0, 0, 1, 0, -1, 0, 1, 1, 1, 0, 0, 1, 2, 3, 4, 4, 4, 5, 5, 4, 2, 0, -1, 0, 1, 1, 0, 0, -1, 0, 0, 1, 0, 1, 0, -1, -1, 0, 0, 1, 1, 2, 1, 3, 4, 5, 5, 3, 3, 4, 6, 4, 3, 1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 0, -3, -2, -1, 1, 1, 3, 1, 2, 4, 6, 6, 4, 3, 4, 4, 5, 5, 2, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -3, -3, -3, -1, 0, 0, 1, 2, 5, 5, 6, 6, 4, 3, 2, 2, 4, 2, 2, 0, -1, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, -2, -3, -3, -4, -3, -1, 0, 1, 3, 5, 7, 7, 6, 5, 2, 2, 2, 1, 1, 0, -2, -3, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -2, -3, -3, -3, -3, -1, -1, 0, 2, 4, 5, 5, 6, 4, 1, 0, 0, 0, 0, -3, -5, -4, 0, -1, -2, -1, 0, 0, 1, 0, 0, 1, 0, -2, -1, -1, 0, 0, 0, 1, 1, 3, 3, 3, 3, 2, 0, 0, 0, -1, -3, -4, -5, -5, 0, -1, -2, 0, 0, 0, 2, 2, 2, 4, 3, 2, 1, 0, 2, 1, 1, 1, 1, 1, 3, 2, 2, 0, 0, -1, -3, -2, -4, -6, -5, -5, 0, 0, 0, -2, 0, 0, 1, 1, 1, 1, 3, 1, 2, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -4, -4, -4, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 2, 1, 0, 0, 0, 1, 1, 2, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 2, 3, 1, 1, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 2, 3, 3, 4, 3, 3, 2, 1, 1, 0, 0, 0, 0, -2, 0, 0, 0, -1, -1, -1, 0, 0, -1, -2, -1, -1, 0, 0, -1, 0, 0, 1, 1, 2, 2, 4, 4, 2, 3, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -2, -1, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, 1, 2, 3, 4, 2, 2, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, -1, -2, -1, -1, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 2, 3, 4, 5, 3, 2, 0, 0, 0, 1, 1, 0, 0, 0, -1, -2, -1, 0, -1, 0, -2, -1, 0, 0, -1, -2, -2, -2, -1, -1, 0, 0, 0, 3, 4, 5, 2, 1, 2, 1, 2, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, -2, -1, -1, -2, -1, 0, 0, 1, 1, 2, 2, 2, 3, 2, 2, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, -1, 0, -2, -1, -2, -1, -1, 0, 1, 2, 2, 2, 2, 3, 3, 3, 1, 0, 0, 0, -2, 0, 0, -1, 0, 0, 1, 1, 3, 2, 0, 0, 0, -1, -1, -3, -1, -1, -1, 0, 0, 1, 2, 1, 3, 2, 2, 3, 0, 0, 0, 0, -2, 0, 0, 0, 1, 1, 0, 2, 2, 1, 1, 0, -2, -1, -1, -2, -1, -1, -1, 0, 1, 1, 1, 1, 3, 3, 2, 2, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 2, 2, 2, 1, 0, -1, 0, -1, -1, -1, -2, 0, -2, 0, 0, 0, 0, 0, 1, 2, 3, 2, 2, 0, 0, 0, 0, 1, 2, 2, 1, 2, 1, 2, 2, 2, 0, 0, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 1, 0, 1, 2, 2, 2, 2, 0, 0, 0, 0, 2, 1, 1, 2, 1, 1, 2, 1, 0, 0, 0, -1, -1, -1, 0, -2, -3, -3, -1, 0, 0, 0, 0, 0, 1, 2, 4, 2, 1, 1, 0, 0, 2, 2, 2, 2, 2, 1, 0, 0, 1, 0, 1, 0, 0, 0, -2, -3, -3, -3, -3, -1, 0, 0, 0, 0, 1, 2, 2, 3, 2, 1, -1, -1, 1, 1, 1, 1, 1, 1, 2, 1, 1, 0, 0, -1, 0, 0, -3, -5, -4, -5, -2, -1, 0, -1, -1, 0, 1, 1, 2, 3, 2, 1, -1, 0, 0, 1, 0, 0, 1, 1, 2, 1, 1, 1, 0, 0, 0, 0, -2, -5, -5, -5, -4, -2, 0, 0, 0, 0, 1, 1, 2, 2, 0, 1, 0, 0, 0, 2, 1, 1, 0, 1, 1, 2, 1, 0, 0, 0, 0, -1, -1, -4, -3, -4, -2, 0, 0, 0, -1, 0, 0, 1, 3, 3, 1, 1, 0, 0, 1, 0, 2, 1, 0, 1, 1, 3, 1, 0, 0, 0, 0, 0, -1, -3, -1, -3, -1, 0, 1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, 2, 1, 1, 1, 0, 1, 2, 1, 2, 2, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 2, 1, 2, 0, 0, 0, 1, 2, 1, 2, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 2, 1, 1, 0, -2, -1, -2, -2, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -3, -2, -1, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 1, 0, 0, -2, -1, 0, 0, -2, 0, 0, 0, 2, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, 1, 0, 1, 2, 1, 0, 1, 0, 0, 1, 0, -1, -1, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 3, 2, 1, 1, 2, 0, 0, 0, 0, 0, -2, -2, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, -1, -1, -2, -1, -1, 1, 0, 2, 2, 4, 4, 2, 2, 1, 0, 0, -1, 0, -1, -1, -1, -1, 0, -1, 0, -1, -2, 0, 0, 0, 0, -1, 0, -2, -2, -2, 0, 0, 2, 2, 3, 4, 5, 3, 2, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 2, 3, 4, 4, 5, 2, 1, 0, 0, -1, 0, -1, -1, -2, -2, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 3, 2, 2, 2, 0, 0, -1, -1, -2, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, -2, -2, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, -1, -2, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -3, -1, -2, 0, -1, -2, -1, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -2, -1, -2, -2, 0, 0, -1, -1, 0, 1, 2, 1, 1, 2, 0, 1, 0, 0, -1, -1, -1, -2, -1, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, -1, -2, 0, -1, 0, -1, -2, -1, 0, 1, 1, 1, 2, 1, 0, 1, 0, 0, -2, -1, -2, -2, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, -2, -1, -2, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -2, -3, -2, -2, -2, -2, -2, -2, -1, 0, 0, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -3, -2, -2, -2, -2, -2, -2, 0, 0, 0, 0, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, -2, -2, -1, -1, -1, -2, -1, -1, 0, 0, 0, -2, -2, -1, -2, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, -1, -1, 0, -1, -1, -2, -2, -2, 0, 0, 0, -1, -2, -1, -2, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -2, -1, -1, -2, -1, -1, -2, -2, -2, -1, -2, -3, -1, 0, 0, -1, -2, -1, -2, -1, -2, -2, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -2, -2, -2, -2, -1, -1, -3, -1, 0, 0, 0, -1, -3, -2, 0, -1, -1, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -2, -1, -1, -1, -2, -1, 0, 0, 0, -1, -2, -1, -1, 0, -1, 0, -1, -2, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, -1, -2, -1, -1, 0, -1, 0, 0, 0, 0, -2, -2, -2, -1, -2, 0, -2, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, -2, 0, -1, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, -1, 0, -2, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -2, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, -1, -2, -2, -1, 0, 1, 0, 0, 0, -1, -2, -1, -1, -2, -1, -3, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, -2, -2, -2, 0, -1, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, -2, -2, -2, 0, -2, -2, -2, -2, -2, -2, 0, 0, -1, 0, 0, 0, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, -2, -3, -2, -1, -1, -2, -3, -3, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, -1, 0, -1, -1, 1, 0, -1, -3, -2, -2, -2, -2, -2, -3, -3, -2, 0, -2, 0, 0, 0, 0, 0, -2, -2, -2, -1, -2, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -1, -1, -2, -3, -2, -3, -1, -1, -1, 0, 0, 0, 0, -1, -1, -3, -2, -3, -3, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, -3, -3, -2, -2, -1, -1, -2, -2, -2, -1, -2, -1, -1, 0, 0, 0, -1, -1, -1, -1, -1, -3, -3, -2, -1, -1, 0, 0, 1, 0, 0, 0, -1, -2, -1, -2, -2, -2, -2, -3, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -2, -3, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -2, -2, -1, -2, -2, -2, -1, -1, -1, 0, 0, 0, -1, 0, 0, -2, -2, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -2, -3, -2, -2, -2, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -2, -2, -2, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, -1, -2, -2, -2, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -2, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -2, -2, -1, -2, -2, -2, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, -1, -2, -1, -1, -1, 0, -2, -2, -3, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -2, -2, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, -1, -3, -2, 0, -1, -3, -3, -3, -1, -3, -1, -1, -1, -1, -1, -1, -2, 0, -1, 0, 0, 0, 0, 1, 1, 1, 2, 0, 1, 0, 0, 0, -1, -3, -3, -2, -1, -3, -3, -3, -2, -3, -2, -2, -2, -3, 0, -2, -2, 0, -1, 0, 0, 0, 0, 1, 1, 2, 3, 2, 1, 2, 1, -1, 0, -2, -1, -2, -2, -2, -2, -2, -3, -2, -2, -2, -1, 0, -2, -1, 0, -1, 0, 0, 0, 1, 2, 0, 2, 1, 3, 3, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 1, 2, 1, 0, 0, 1, 2, 1, 1, 1, 2, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 2, 2, 2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 2, 1, 0, 0, 0, 1, 1, 1, 2, 2, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 1, 0, 1, 0, 1, 1, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 1, 2, 0, 1, 0, 1, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 2, 1, 2, 1, 1, 1, 2, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 1, 1, 1, 2, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -2, 0, -1, -2, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -2, -2, -2, 0, -1, -1, 0, -1, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, -1, -1, -2, -2, -1, -2, -1, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, -3, -3, -3, -2, 0, -1, -1, -1, -1, 0, 0, 2, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -3, -3, -2, -3, -1, -1, 0, 0, -1, -1, 0, 1, 1, 1, 1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, -1, -1, -1, -2, -3, -2, -3, -2, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, -2, -3, -3, -2, -1, -1, -2, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -2, -2, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -2, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 2, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 2, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, -1, -1, -2, -1, -2, -2, -2, -1, -2, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 2, 3, 4, 2, 1, 0, 0, -1, -3, -4, -5, -5, -5, -6, -6, -5, -4, -4, -4, -4, -5, -3, -1, 0, -1, -3, -2, 0, 0, 0, 0, 0, 1, 2, 2, 3, 4, 0, 0, -1, -4, -3, -4, -4, -5, -4, -3, -3, -3, -3, -2, -2, -2, -3, -1, 0, -1, -1, -2, 0, 0, -1, -1, 0, 1, 0, 2, 3, 1, 1, -1, 0, -2, -4, -3, -3, -3, -3, -2, -3, -2, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, -1, -2, -1, -1, -2, -3, -2, -2, -3, -3, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 2, 0, 0, -1, 0, -1, -2, -1, -2, -3, -4, -3, -4, -2, 0, 0, 1, 0, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -3, 0, 0, 0, 0, 0, 0, -2, -3, -3, -3, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -2, -2, -1, 0, -1, 1, 1, 3, 0, 1, 0, -1, -3, -3, -3, -1, -2, -1, -1, 0, -1, -1, -1, -1, -1, -2, 0, 0, -1, -1, -2, -1, -2, 0, 0, -1, 0, 1, 2, 2, 1, 0, 0, 0, -2, -3, -3, -4, -2, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, -1, -2, -1, -1, -1, -2, -2, -2, -2, -1, -1, 0, 1, 0, 0, 1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, -2, -2, -1, -1, -1, -1, -1, 0, 0, -2, -1, -3, -3, -2, -2, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, -2, -1, -2, -2, -1, 0, 0, 0, -1, -1, -1, -2, -3, -2, -2, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, -2, -2, -2, -1, -1, -2, -1, -3, -3, -3, -2, 0, 1, 0, 0, 2, 2, 3, 2, 1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -1, -3, -2, -1, -1, -1, -3, -3, -2, 0, 1, 1, 0, 1, 2, 1, 3, 1, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -2, -3, -3, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, -1, -2, -1, -2, -1, 0, 0, 0, 0, -2, -1, -1, -1, -1, -2, -2, -4, -3, -3, 0, 0, 0, -1, -1, -2, 0, 0, -1, -2, -3, -1, 0, -1, 0, -2, -2, -1, 0, 0, 0, -1, 0, -1, -1, -1, -2, -2, -2, -2, -2, -2, -2, 0, -1, -1, -3, -2, -2, -2, -2, -2, -2, -2, -1, -1, -1, 0, -2, 0, 0, 0, 0, 0, -1, -2, -2, -1, -1, -2, -1, -2, -3, -1, -2, -2, -1, -1, -2, -3, -2, -2, -1, -3, -3, -2, 0, 0, 0, 0, 0, 1, 0, 1, 1, -1, -2, -2, 0, 0, 0, -1, -2, -2, -1, -2, -3, -3, -2, -1, 0, 0, -2, -2, -3, -2, -3, -2, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, -2, -2, -2, -1, -1, -2, -2, -1, -3, -2, -2, -2, -2, -3, 0, -1, -3, -3, -4, -4, -4, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, 0, -1, 0, -1, -1, -1, 0, 0, 0, -1, -2, 0, -1, -2, -2, -3, -3, -5, -3, -3, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -3, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -2, -2, -2, -3, -4, -5, -6, -4, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, -3, -4, -4, -4, -4, -5, -5, -5, -3, -2, -2, -1, -1, -1, 0, 0, 0, 0, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -4, -4, -4, -2, -3, -4, -3, -3, -4, -3, -2, -1, 0, 0, 0, 0, 0, -2, -2, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -2, -4, -4, -5, -4, -3, -3, -3, -2, -2, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -3, -3, -4, -5, -5, -4, -4, -3, -2, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -2, -1, -1, -1, 0, 0, -1, -1, -2, -2, -3, -4, -3, -5, -4, -3, -3, -1, -1, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, -2, -2, -2, -2, 0, -1, -1, -2, -1, -1, -2, -2, -3, -2, -3, -1, 0, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, -2, -1, -1, -2, 0, 0, 0, 0, 0, 2, 3, 3, 4, 2, 2, 3, 4, 3, 4, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 3, 3, 3, 3, 1, 2, 2, 2, 1, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, -2, -2, -1, -2, -2, -1, -2, -1, -1, -1, -1, -2, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, -2, 0, 0, -2, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, -2, -2, -1, 0, -1, -1, -1, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, -1, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, 0, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, 0, 0, 0, -1, 1, 0, 0, 0, -2, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 2, 0, 2, 2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 2, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 2, 1, 1, 1, 2, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -2, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, -1, -1, -2, -1, -2, 0, -1, 0, 0, -1, 0, -1, 0, -1, -2, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -2, -2, -2, 0, 0, -2, -1, -1, -1, 0, -1, 0, -2, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, 0, 0, -1, 0, -1, 0, 0, 0, 0, -2, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -2, -3, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -3, -2, -2, -2, 0, -1, 0, -1, -1, -1, 0, -1, 0, -2, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -2, -2, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, -2, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 0, -1, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 2, 1, 1, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -2, 0, -2, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, -2, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, -1, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, -1, -2, -1, -2, -2, -2, -2, -1, 0, -2, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -3, -2, -3, -1, -1, -2, -2, 0, -2, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -3, -3, -3, -1, -1, -1, -2, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 1, 1, 0, -1, 0, 0, 0, 0, -1, -2, -1, -2, -1, -1, -2, -2, -1, -2, -2, -2, -2, -1, -1, -1, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -2, -1, -1, -2, -2, -2, -2, -3, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, -1, -1, -2, 0, -1, -3, -2, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -2, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, -2, -3, -1, -2, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, -2, -1, 0, 0, 0, -1, 0, 0, -1, -2, -1, -1, -1, -1, 0, -1, -1, -1, -1, -3, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, -1, -1, -2, -1, -1, -2, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, -1, -1, -2, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, -2, -1, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 2, 0, 1, 1, 0, 1, 1, 2, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 1, 0, 0, 1, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, -2, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 0, 0, 0, 0, 2, 1, 1, 1, 0, -1, -1, -1, 0, -1, 0, 0, -2, -1, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 2, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -2, -1, -1, -1, 0, 0, 0, 1, 0, 0, 1, 2, 2, 2, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 1, 1, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 2, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, -1, -1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 2, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 2, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 2, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 2, 0, 0, 0, 2, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 2, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 2, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 1, 0, 0, 2, 1, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 1, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 2, 1, 1, 1, 1, 3, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -2, -1, 0, 0, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, -1, -1, -1, -1, -1, -1, -2, -2, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, -1, 0, -2, -2, -1, -1, 0, -2, 0, -2, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, -1, -1, -2, 0, -1, -1, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, -1, -2, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, 0, -2, -1, -1, -1, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -2, -2, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, -1, -2, -2, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -2, -2, -2, -1, -1, -1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, -1, -2, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 2, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 2, 0, 1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -2, -1, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, -2, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -2, 0, -2, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, -2, -1, -2, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -2, -1, 0, -1, -1, 0, -1, -1, -1, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -2, -1, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -2, -2, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -1, -1, -2, -2, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, -1, 0, -2, -2, -2, -2, 0, -2, 0, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -2, 0, 0, 0, -2, -1, 0, -1, -1, -1, -2, -2, -1, -1, -1, -1, -2, 0, -1, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, -2, -1, -1, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -2, -1, 0, 0, 0, 0, -1, -2, 1, 1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 2, 3, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 2, 0, 0, -2, -1, 1, 0, 0, 2, 2, 1, 2, 0, 1, 2, 0, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, -1, -1, 0, 1, 1, 2, 2, 2, 2, 1, 2, 2, 0, 1, 4, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 1, 1, 1, 3, 2, 3, 2, 2, 1, 0, 2, 3, 2, 0, 0, -1, 0, -1, 2, 0, 0, 0, 0, -1, 0, 0, 3, 2, 1, 0, 0, 0, 2, 2, 2, 3, 4, 5, 2, 1, 3, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -2, -1, 0, -1, 1, 1, 0, 0, 0, 0, 2, 2, 2, 4, 3, 4, 3, 3, 3, 1, 1, 1, 0, -1, 0, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 1, 0, 0, 0, 1, 2, 3, 2, 4, 5, 4, 5, 2, 3, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 1, 3, 3, 2, 3, 6, 6, 4, 2, 3, 0, -1, 1, -1, -1, 0, -1, 0, -1, -1, -1, 0, -1, -2, 0, -1, -1, 0, 0, -1, -1, 0, 1, 2, 2, 3, 3, 5, 6, 4, 3, 1, 0, -1, 1, -1, -2, 0, 0, -2, 0, -1, -1, 0, -2, 0, 0, -1, -1, 1, 0, -1, 0, 0, 1, 1, 2, 3, 3, 4, 5, 4, 3, 3, 0, 0, 1, 0, -1, 0, 0, 0, -1, -2, -1, 0, -2, -1, -1, -3, -1, 0, 0, 0, 1, 1, 0, 1, 1, 2, 1, 3, 4, 4, 5, 4, 0, 2, 1, -1, -1, -1, 0, -1, -2, 0, -1, 0, -3, -1, -1, -2, -1, 0, 0, -1, 0, 1, 0, 0, 1, 2, 2, 4, 4, 3, 3, 3, 0, 1, 1, 0, -2, -1, -2, -1, -1, 0, 0, 0, -2, -1, -1, -1, 0, 0, 0, -2, 0, 1, 1, 0, 0, 2, 3, 3, 5, 4, 4, 2, 0, 2, 2, -1, -1, -1, -2, -2, -2, 1, 0, 0, -2, 0, 0, -2, 0, 0, -1, -1, -1, 0, 1, 1, 1, 3, 5, 3, 4, 5, 2, 1, 0, 2, 0, 0, -2, -2, -3, -3, -1, 1, 1, 0, -4, -2, -2, 0, 0, 1, -1, 0, 0, 0, 0, 2, 1, 2, 4, 3, 3, 5, 1, 2, 0, 1, 0, 0, -1, -1, -3, -2, -1, 0, 1, 0, -3, -2, -1, -2, 0, 0, 0, 0, -2, -1, 0, 2, 2, 3, 3, 3, 3, 5, 2, 2, 2, 1, 0, 0, -1, -1, -2, -2, 0, 0, 1, 0, -3, -1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 1, 3, 3, 4, 2, 5, 4, 1, 3, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 1, 0, -4, -3, -2, -1, 0, 0, 1, -1, -2, 0, 0, 1, 3, 3, 4, 4, 3, 5, 1, 1, 1, 0, 0, 0, -1, -2, -1, 0, -1, 0, 1, 0, -3, -1, -1, 0, 0, 0, 1, 0, -1, 0, 0, 1, 3, 3, 3, 3, 4, 4, 2, 2, 0, 0, 1, 1, 0, -1, 0, -1, 0, 0, 0, 0, -2, -1, -2, 0, 0, 0, 1, 0, -1, -1, 1, 2, 1, 4, 3, 4, 2, 5, 3, 2, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, 0, -3, -1, -2, 0, -1, 0, 2, 0, -2, 0, 0, 2, 1, 2, 5, 3, 3, 4, 2, 1, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 1, -1, -3, 0, 0, 1, 3, 3, 4, 3, 1, 5, 3, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, 0, -2, 0, 0, 0, 0, 0, -2, 0, 0, 1, 2, 1, 4, 2, 3, 3, 2, 1, 0, 1, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 1, 2, 2, 4, 2, 0, 2, 2, 2, 0, 0, -1, 0, 0, 0, 1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 2, 2, 3, 2, 2, 3, 3, 0, 0, 0, 1, 0, 0, 1, 0, 0, -2, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 2, 1, 1, 1, 1, 2, 1, 1, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 1, 0, 0, 0, -1, -1, 0, 0, 1, 2, 0, 0, 1, 2, 1, 0, 1, 3, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 1, 1, 0, 3, 3, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 3, 0, 0, 2, 2, 1, 1, 0, 2, 2, 1, 0, 0, 2, 1, 1, 1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 3, 2, 3, 3, 2, 2, 2, 2, 2, 2, 1, 1, 0, 1, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 2, 1, 2, 2, 2, 1, 1, 0, 1, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 1, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 1, 0, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 2, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 2, 1, 2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, -1, -1, 0, -1, 0, 1, 1, 0, 1, 1, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, -1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 2, 1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -2, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -2, -1, -1, -1, -1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, -1, -1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 1, 1, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 1, 1, 0, 0, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, -1, -2, -2, -2, -2, -1, -2, -2, -1, -2, -1, -2, -2, -1, -2, -2, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, -1, -1, -2, -1, 0, -1, -1, -2, -1, -2, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, -2, -1, -2, -1, -2, -1, -1, -2, 0, 0, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, 0, -2, -1, 0, -1, -1, -1, -1, 0, -2, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, -2, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, -1, 0, -1, -1, 0, -1, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -2, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, -1, 0, -1, -2, -1, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 3, 2, 1, 0, 0, 1, 1, 1, 2, 1, 2, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 2, 1, 1, 2, 3, 1, 2, 1, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 1, 2, 3, 4, 2, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 2, 4, 2, 3, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 2, 2, 3, 2, 3, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 4, 5, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 0, 1, 2, 2, 2, 1, 0, 0, 1, 2, 1, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 1, 2, 1, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 1, 1, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 1, 1, 2, 1, 1, 2, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 1, 2, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, -1, 0, 1, 1, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 2, 1, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 1, 1, 2, 3, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, -1, -2, -2, -2, -1, -2, 0, 0, 0, 0, 1, 2, 2, 2, 1, 2, -1, -1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -3, -3, -3, -3, -3, -1, 0, 0, 0, 0, 1, 2, 2, 2, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -2, -4, -4, -3, -4, -2, -1, 0, 0, 0, 0, 1, 2, 2, 3, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -2, -3, -3, -3, -3, -2, -1, -1, 0, 0, 2, 3, 2, 2, 2, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -3, -2, -1, -1, -1, -1, 0, 1, 2, 3, 2, 2, 2, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -2, -2, -1, 0, -1, 0, 0, -1, 0, 1, 1, 1, 2, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 1, 0, 1, 1, 1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, -1, -1, -1, -2, -1, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 1, 1, 2, 0, 1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 2, 2, 0, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, -1, 0, -1, 0, -2, -1, -1, -1, 0, -1, -1, 0, 0, 2, 1, 2, 2, 1, 1, 1, 1, 0, 0, 1, 0, -1, -1, 0, -1, -2, -1, -1, -2, 0, 0, -1, -1, -1, -2, -2, -1, 0, 0, 1, 1, 1, 1, 3, 3, 1, 2, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, -2, 0, -2, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 3, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 1, 1, 1, 2, 2, 2, 1, 1, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -1, -2, -3, -2, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 2, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -2, -3, -2, 2, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 1, 1, 0, 1, 0, 1, 1, -1, 0, 0, 0, -2, -3, -1, 1, 0, 0, 1, 0, 0, 1, 2, 0, 0, 0, -1, 0, -1, 0, 0, 0, 2, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -2, -2, 1, 1, 0, 0, 0, 0, 2, 0, 1, 0, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, 1, 2, 2, 0, 0, 0, 0, 0, -1, -1, 2, 2, 1, 1, 0, 0, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, -2, -1, 2, 1, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, -1, 2, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 2, 2, 2, 0, 1, 0, 2, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 2, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 2, 2, 1, 0, 0, 1, 2, 1, 1, 0, 0, 0, -1, -2, 0, 1, 0, 0, 0, -2, 1, 0, 1, 1, 0, 1, 1, 2, 0, 0, 0, 1, 1, 2, 0, 0, 0, 2, 2, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 2, 0, 0, 0, 0, 0, 2, 1, 1, 1, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, -1, 0, 0, 0, 2, 2, 0, 1, 3, 2, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 1, 0, 1, 1, 2, 2, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 1, 0, 1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 1, 2, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 2, 0, -1, 0, 0, 1, 2, 1, 2, 1, 1, 1, 1, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 1, 0, 0, 0, 0, 2, 2, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 2, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 2, 2, 2, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 1, 1, 3, 2, 1, 3, 1, 0, 0, 0, 1, 0, 0, 0, -2, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 1, 0, 1, 2, 3, 2, 0, 0, 0, 1, 0, -1, -2, -2, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -2, 0, -2, -2, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, -1, -1, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 2, 0, 1, 2, 0, 0, 0, 0, 0, 0, -2, -3, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 3, 2, 2, 2, 3, 2, 0, -1, -1, 0, -2, -3, -2, -2, 0, 0, 0, 0, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 2, 3, 2, 2, 1, 1, 0, 0, 0, 0, -3, -3, -2, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 2, 3, 3, 4, 4, 2, 2, 1, 0, 0, 0, -2, -3, -1, 0, 0, 0, 0, 1, 2, 2, 1, 0, -1, 0, -1, -1, -1, 0, -1, 1, 0, 2, 3, 2, 4, 3, 4, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, 1, 2, 3, 4, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 2, 3, 3, 2, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 1, 2, 1, 2, 2, 3, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 2, 3, 2, 0, 0, 2, 1, 1, 1, 1, 1, 1, 0, 0, 1, 2, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 2, 2, 2, 1, 0, 2, 1, 2, 2, 0, 1, 0, 0, 1, 0, 2, 3, 3, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 2, 1, 2, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 1, 1, 1, 2, 3, 3, 2, 2, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 3, 2, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 2, 2, 3, 3, 3, 3, 1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 3, 3, 2, 1, 0, 0, 1, 0, 0, 0, -1, -2, 0, 1, 2, 1, 2, 3, 2, 2, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 3, 4, 2, 1, 2, 1, 0, -1, -2, -2, -2, 0, 1, 1, 3, 3, 3, 3, 2, 2, 3, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 2, 4, 3, 2, 1, 1, 0, 0, -1, -1, -2, -2, -2, -1, 2, 3, 2, 2, 2, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 3, 1, 1, 1, 0, 0, -2, -2, -3, -3, -3, 0, 0, 2, 3, 3, 3, 3, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 1, 0, 0, -1, -1, -3, -3, 0, -1, 1, 1, 3, 2, 4, 3, 3, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 1, 0, 0, -1, 0, -2, 0, 0, 0, 2, 1, 3, 2, 3, 2, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 3, 2, 2, 2, 3, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 2, 1, 3, 2, 2, 3, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 2, 1, 2, 1, 2, 2, 1, 1, 2, 2, 2, 2, 3, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 1, 1, 1, 2, 3, 1, 0, 0, 1, 2, 2, 1, 2, 2, 3, 2, 2, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 3, 2, 1, 1, 1, 2, 3, 3, 1, 3, 2, 2, 3, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 2, 2, 2, 1, 2, 1, 3, 3, 2, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 2, 2, 1, 1, 2, 4, 4, 3, 1, 1, 1, 2, 3, 2, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, -2, -1, 0, 0, 2, 2, 3, 3, 3, 4, 3, 3, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -2, -1, 0, 0, 1, 3, 3, 3, 3, 3, 2, 2, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 1, 2, 3, 3, 3, 3, 2, 1, 0, 1, 0, -1, 0, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, -2, -2, -1, -1, -2, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 0, -1, 0, -1, -1, -2, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 2, 2, 1, 0, 0, -1, -2, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 2, 1, 0, 2, 1, 1, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, -2, -1, 1, 1, 0, 2, 1, 2, 2, 1, 0, 1, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 2, 2, 0, 1, 0, 0, 0, -1, 0, -2, -2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, -2, 0, 0, 0, 1, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, -2, 0, -1, -1, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, -2, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -2, -1, 1, 0, 1, 0, 0, 0, 1, 2, 1, 1, 0, 1, 0, 0, -1, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, -1, -1, 0, 1, 1, 0, 1, 1, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -2, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 1, 1, 0, 2, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -2, -2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 2, 2, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 2, 1, 2, 2, 2, 1, 0, 0, 0, 1, 1, 0, 1, 0, -2, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, 0, 2, 0, -1, -2, -2, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 3, 2, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 0, 2, 0, 0, 1, 0, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 2, 2, 0, -1, 0, 0, 0, 1, 0, 1, 3, 2, 1, 2, 1, 0, 3, 3, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 3, 0, 0, -1, 0, 0, 0, 1, 2, 3, 4, 4, 2, 1, 1, 2, 2, 2, -1, 0, 0, -1, 0, 0, 0, 0, 0, -2, -2, 0, -1, 0, 0, 2, 0, 0, 0, 0, 0, 1, 1, 4, 3, 4, 3, 3, 2, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, 0, 1, -1, -1, -1, 0, 2, 2, 1, 2, 4, 4, 3, 2, 1, 1, 1, 0, -2, 0, 0, -1, 0, 0, -1, 0, 0, -2, -1, 0, -2, -1, 0, 1, 0, 0, 0, 0, 1, 2, 2, 3, 6, 5, 3, 2, 1, 1, 0, 0, -2, -2, -1, 0, 0, 0, -1, 0, 0, -1, -1, -2, -2, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 4, 5, 6, 3, 2, 1, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, -1, -2, 0, 0, 0, 1, 2, 2, 4, 6, 6, 5, 3, 2, 0, 0, 0, 0, -2, 0, 0, -1, 0, -1, 0, 0, -3, -2, -2, -3, 0, 0, -1, -2, 1, 1, 0, 0, 2, 1, 3, 7, 4, 5, 3, 3, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, -3, -1, -3, -2, 0, 0, -1, -2, 1, 1, 0, 0, 2, 3, 4, 6, 4, 5, 4, 3, 0, 1, 0, -1, -3, -2, -2, -1, 0, 0, 0, -1, -3, -2, -2, -2, -1, 0, -1, -1, 0, 0, 1, 0, 2, 3, 4, 5, 5, 5, 3, 2, 0, 1, 1, -2, -2, -2, -3, -2, 0, 2, 0, 0, -3, -1, -2, -1, -1, -1, -1, -2, 0, 1, 1, 0, 1, 4, 6, 5, 4, 4, 3, 1, 0, 2, 1, -1, -2, -3, -3, 0, -1, 2, 0, 0, -3, -1, -2, -2, 0, 0, 0, 0, -2, 0, 1, 2, 2, 6, 5, 4, 5, 3, 3, 2, 0, 0, 0, -1, -1, -2, -3, 0, 0, 3, 0, 0, -3, -2, -2, 0, 0, 0, 0, -1, -1, -1, 1, 3, 3, 6, 4, 4, 5, 5, 2, 1, 0, 0, 0, -1, -1, -3, -1, -1, 0, 2, 0, 0, -3, -2, -1, 0, 0, 1, -1, -1, 0, 0, 2, 3, 4, 5, 4, 4, 4, 4, 2, 2, 0, 0, 0, -1, -1, -2, -1, -1, 0, 3, 0, -1, -4, -1, -1, -1, -1, 0, 0, -1, -1, 0, 1, 2, 3, 4, 3, 3, 4, 4, 2, 1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 2, 0, 0, -3, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 2, 3, 3, 5, 4, 5, 3, 3, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 1, 0, 0, -3, -1, 0, -1, 0, 0, 1, 0, -1, 2, 1, 2, 2, 4, 6, 3, 4, 3, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -3, -2, -1, 0, 0, 0, 0, -2, 0, 0, 2, 1, 2, 5, 6, 4, 3, 6, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, -2, -2, -1, -1, 0, 0, 0, -1, 0, 1, 3, 1, 2, 3, 4, 5, 5, 4, 3, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -3, -1, 0, 0, 0, 0, 1, -1, 0, 2, 2, 2, 1, 2, 4, 3, 5, 6, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 1, 3, 2, 2, 3, 3, 1, 0, 2, 1, 0, -1, -1, 0, -1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 2, 0, 3, 4, 1, 0, 3, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 2, 3, 3, 2, 2, 3, 3, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, 2, 3, 2, 0, 3, 1, 0, 0, 0, 0, 1, 1, 1, -1, 0, -1, -1, -2, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 1, 0, 0, 1, 2, 1, 1, 1, 3, 1, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, -2, -1, 0, 0, 0, -1, -2, -1, 0, -1, -1, 0, 0, -1, 0, 2, 2, 0, 1, 1, 2, 2, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, -1, 0, -1, -1, 1, 1, -1, 0, 1, 0, 0, 1, 1, 1, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -2, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, -2, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -2, -1, -1, -2, -1, -2, -1, -3, -1, -2, -1, -1, -1, 0, -1, 0, -2, 0, 0, -1, -1, 0, 1, 2, 2, 3, 3, 1, 1, 0, -1, -1, -2, -2, -1, -3, -1, -1, -2, -2, -1, 0, -1, 0, -2, -1, -2, -2, -2, -2, 0, 0, 0, -1, 0, 2, 2, 3, 4, 3, 2, 1, 0, 0, -1, -2, -3, -2, -3, -3, -1, 0, -1, 0, 0, -1, -1, 0, -1, -2, -2, -2, 0, -1, -1, -1, -1, 0, 0, 3, 4, 3, 1, 0, 0, 0, 0, -2, -3, -2, -2, -2, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 0, 0, 0, 0, -1, -2, -2, -1, -2, -3, -1, -1, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, -1, -1, -3, -1, -1, -1, -2, -1, 0, 1, 0, -1, -1, -3, -2, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, -3, -2, -3, -1, 0, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -3, -2, -2, -2, -1, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, -1, -1, -3, -2, -1, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, -1, -1, -1, -1, -2, 0, -2, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, -1, -2, -2, 0, -1, -1, -2, -2, -2, -2, -2, 0, 0, -1, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, -2, -2, -2, 0, 0, 0, 0, -1, -3, -2, -1, -1, -1, 0, 0, 0, 1, 1, 2, 0, 0, -1, -1, 0, 0, 1, 1, 1, 0, -1, -1, -1, -1, -3, -2, -2, -1, -1, -1, -1, -2, -4, -2, -1, 0, 1, 0, 1, 1, 2, 1, 2, 0, 1, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, -2, -2, -2, -2, -2, -2, -2, -1, -1, -3, -2, -1, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 0, 0, -1, 0, 1, 1, 0, 0, -1, -2, 0, -1, -2, -1, -2, -2, -3, -3, -2, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -2, -1, -1, -2, -1, -2, -2, -4, -2, -2, -1, 0, 0, -2, -3, -1, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -2, -1, -1, -2, -2, -2, -2, -1, -1, 0, -1, -2, -4, -3, -1, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -3, -1, -1, -3, -2, -2, -2, -2, -3, -3, -1, 0, 0, -2, -2, -2, -2, 0, -1, -1, -1, 0, 0, 0, 1, 1, 0, 1, 1, -1, -1, -1, -2, -1, -2, -2, -1, -2, -2, -2, -2, -2, -2, -2, -1, -1, -1, -2, -3, -2, -3, -2, -1, -1, 0, 0, 1, 2, 2, 0, 0, 0, -1, -1, -2, -2, -1, -1, -1, -3, -2, -2, -3, -3, -2, -3, -2, -1, -2, -1, -1, -1, -3, -2, -1, 0, 0, 1, 0, 1, 0, 2, 0, 0, -1, -2, -2, -2, -3, -1, 0, -1, -2, -1, 0, -2, -3, -2, -2, -2, -1, -1, 0, -1, -2, -3, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -2, -1, -1, -2, -1, -1, -2, -2, -2, -2, -2, -1, -3, -2, -1, 0, 0, -1, -2, -2, -3, -1, -1, 0, 1, 0, 0, 0, 0, 0, -1, -2, -1, -3, -2, -1, -1, -1, -2, -2, -2, -2, -1, -1, -2, -3, -2, -2, -2, -1, -1, -2, -3, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, -2, -1, -2, -3, -3, -1, -2, -2, -1, -2, -2, -2, -1, -1, -1, -1, -1, -2, -2, -2, -2, -2, -2, -1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, -2, -2, -1, -2, -3, -3, -1, -1, 0, -1, -1, -1, -2, -1, -1, -1, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, -2, -1, -2, -1, -1, -1, -1, -1, -2, -1, -1, -2, -1, -1, -2, -1, -3, -1, -1, 0, 0, 0, 1, 0, 1, 0, 1, 0, -1, -1, -1, 0, -2, -1, -3, -3, -3, -1, -1, -2, -2, -1, -2, -2, -1, -2, -3, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -2, -2, -1, -1, -1, -3, -3, -3, -3, -2, -3, -1, -2, -1, -2, -2, -3, -2, -2, -1, -1, 0, 0, 0, 1, 0, 2, 2, 0, 0, -1, -2, -1, -1, -1, 0, 0, -2, -1, -2, -2, -3, -2, -1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 3, 3, 1, 2, 3, 2, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 2, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 2, 2, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 2, 3, 2, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 1, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 3, 2, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 1, 1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -2, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -2, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 1, 0, 1, 0, 1, 1, 1, 2, 2, 1, 1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 1, 1, 2, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 1, 2, 1, 2, 1, 1, 2, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, -1, 0, -1, -1, 0, -2, -1, -2, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 1, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, -1, -2, -1, -1, 0, -2, -2, -2, -1, -1, -1, 0, 0, 0, 1, 0, 1, 3, 2, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, -2, -1, -2, 0, -2, 0, -2, -1, 0, -1, -1, -1, -1, -2, 0, 0, -1, 0, 1, 1, 3, 3, 3, 3, 2, 1, 1, 0, 0, 0, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, -1, 0, 0, 0, 1, 3, 2, 2, 3, 2, 1, 1, 1, 1, 0, 0, -2, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, 0, 1, 1, 3, 2, 2, 1, 2, 2, 2, 1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, -2, 0, -2, -2, -1, -1, 0, 1, 1, 3, 3, 2, 1, 2, 1, 2, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 2, 2, 3, 2, 1, 1, 3, 1, 1, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, -1, -1, -2, -1, -1, 0, 0, 1, 2, 3, 1, 1, 1, 1, 2, 0, 1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 1, 2, 2, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 1, 1, 2, 1, 2, 1, 2, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 1, 1, -1, -1, 0, -1, -1, 0, 0, 0, 1, 2, 2, 0, 0, 2, 3, 1, 1, 1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 3, 2, 1, 2, 0, -1, -1, 0, 1, 1, 0, 1, 2, 1, 1, 2, 1, 0, 1, 0, 0, 0, -2, -2, 0, 0, 1, 1, 0, 0, 1, 0, 3, 2, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -2, 0, -2, 0, 1, 0, 0, 0, 0, 2, 2, 1, 1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 2, 1, 1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 1, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 1, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 2, 1, 2, 1, 0, -1, 0, 0, 1, 0, 0, 1, 1, 2, 1, 1, 2, 1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 2, 1, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 1, 1, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 2, 1, 2, 1, 1, 1, 0, 0, -1, -1, 0, 1, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, -1, 0, -2, -1, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, -1, -1, -1, 0, 0, 0, 1, 1, 2, 1, 0, 1, 1, 1, 1, 1, 0, -1, -1, -1, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, -1, -1, -1, 0, -1, 0, 1, 1, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, 2, 3, 2, 1, 1, 2, 0, 1, 2, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 2, 2, 2, 2, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 1, 2, 1, 2, 2, 2, 2, 0, 0, 1, 1, 0, 0, -1, 0, -2, 0, -1, 0, -1, 0, -1, 0, 0, -1, -2, -1, 0, -1, -1, 0, 0, 2, 3, 3, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, -2, -2, -1, -1, -1, 0, 0, 0, 1, 1, 3, 2, 2, 1, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, 0, 1, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, -1, 0, 0, -2, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -2, -2, -2, -2, -1, -1, 0, 0, 0, -1, 0, 1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, -1, -1, -1, -2, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 1, 2, 0, -1, 0, 0, 0, 1, 0, 1, 1, 2, 1, 0, 0, -1, 0, 1, 0, -1, -2, -2, 0, -1, -2, 0, 0, 0, 0, 0, -1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, -1, -1, 1, 1, 0, 0, 0, 1, 2, 3, 0, 0, 1, 1, 0, 1, 1, 2, 0, 0, 0, -1, -1, 0, 0, 2, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 1, 1, 1, 1, 0, 2, 0, 1, 0, 0, 0, 0, 0, 1, 1, -1, -1, -1, -1, 0, 0, -1, 0, 1, 0, 1, 1, 0, 0, 2, 2, 1, 1, 0, 1, 2, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, -3, -2, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 2, 0, 0, 1, 1, 3, 2, 0, 2, 1, 1, 1, 0, 0, -1, -1, 0, -2, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 4, 3, 0, 0, 3, 2, 0, 1, 0, 0, 0, 0, -2, -3, -2, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 2, 2, 2, 0, 2, 3, 2, 2, 0, -1, -1, -1, -2, -4, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 2, 2, 2, 2, 2, 0, 0, 2, 3, 1, 2, 0, -1, -1, -1, -2, -3, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 2, 2, 0, 2, 4, 2, 2, 1, 1, 0, 1, 1, 0, 1, 0, -2, 0, 0, -1, -4, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, 0, 3, 3, 3, 3, 2, 2, 1, 2, 1, 0, 1, 0, 0, 0, 0, -1, -2, -2, -2, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 2, 0, 0, 3, 4, 3, 3, 2, 1, 2, 1, 0, 1, 0, -1, -2, 0, 1, -1, -3, -2, -2, -2, -2, 0, 0, 0, -1, 0, 0, -1, 1, 1, 2, 2, 2, 3, 2, 3, 2, 1, 2, 1, 0, 0, 0, -1, -1, 0, 0, -1, -2, -1, -4, -2, -1, 0, 0, 0, -2, 0, 0, 0, 0, 1, 1, 2, 1, 2, 2, 2, 2, 3, 2, 0, 2, 1, 0, 0, -2, -1, 0, 0, 0, -2, -2, -2, 0, 1, 0, 0, 0, 0, 0, 1, 0, 2, 1, 3, 1, 2, 2, 3, 2, 3, 1, 0, 2, 2, 0, 0, -1, 0, 0, 0, 0, -1, -2, -2, -2, 0, 0, 0, -2, 0, 0, 0, 0, 2, 1, 2, 1, 3, 2, 2, 3, 3, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, -3, -2, -2, -1, 1, 0, 0, -2, 0, 0, 0, 0, 0, 2, 1, 2, 3, 2, 2, 2, 1, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, -1, -2, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 2, 1, 3, 3, 2, 0, 2, 1, 0, 0, 1, 0, -1, -1, -1, 0, -1, -1, -1, -2, -2, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 2, 1, 1, 4, 2, 2, 0, 1, 2, 0, 0, 1, 0, -1, -1, 0, 0, 0, -2, -1, -2, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 2, 1, 1, 3, 2, 2, 0, 0, 2, 1, 1, 0, 0, 0, -2, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 1, 0, 2, 2, 2, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 1, 2, 0, 0, 1, 2, 2, 0, 1, 0, 1, 1, 2, 0, 0, 0, 0, -1, 0, -1, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 2, 1, 0, -1, 0, 0, 0, -2, -1, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -2, -2, 0, -2, 0, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 1, 1, 0, 0, 2, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 1, 0, -1, 2, 1, 0, -1, -3, -1, -2, -1, -1, -1, 0, 0, -1, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, -1, -2, 0, 1, 0, 0, 0, 0, 1, 0, -3, -1, -2, -1, -1, -2, -3, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, -1, -3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, -1, 0, 1, 0, 2, 1, 0, 0, 0, -1, -1, -2, -1, -1, -1, -1, -2, -1, -1, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -2, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 1, 0, 1, 3, 1, 3, 1, 1, 1, 1, 1, 0, -1, -2, -1, -2, -3, -5, -3, -1, 1, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, -1, -1, -1, 1, 1, 1, 2, 2, 2, 1, 2, 3, 2, 0, 0, -2, -3, -3, -5, -4, -2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, -4, -2, -2, -1, 0, 0, 0, 2, 2, 2, 3, 3, 4, 0, -1, -1, 0, -1, -2, -3, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -3, -5, -4, -3, -2, -1, -1, 0, 1, 1, 3, 3, 4, 3, 0, 0, -1, 0, 0, -2, -2, -1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, -4, -3, -3, -3, -2, -1, -2, 0, 1, 2, 2, 4, 3, 4, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, 0, 0, -1, 0, 0, 2, 4, 4, 3, 0, 0, 0, 1, 1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 3, 3, 2, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 2, 1, -1, 0, 0, 0, 1, 1, 2, 2, 0, 0, 1, 0, 0, 2, 3, 1, 0, -1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 2, 1, 0, 0, 1, 2, 1, 1, 1, 0, 1, 0, 0, 0, 1, 3, 2, 2, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 2, 2, 0, 0, 1, 1, 2, 0, 0, 1, 0, 1, 1, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 2, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 3, 2, 3, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, 1, 1, 3, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 3, 4, 3, 2, 0, 0, 0, 0, -1, -2, -2, -1, 0, 1, 2, 1, 1, 2, 2, 1, 1, 2, 1, 0, 0, 1, 0, 1, 0, 0, 0, 2, 4, 5, 4, 1, 1, 0, 0, -1, -3, -3, -3, -3, -1, 0, 1, 2, 1, 1, 2, 2, 1, 1, 1, 1, 0, 1, 0, 0, 1, 1, 0, 3, 4, 5, 4, 2, 2, 0, -1, -1, -1, -3, -3, -3, -1, -1, 0, 2, 3, 3, 2, 3, 2, 1, 0, 0, 1, 1, 0, 1, 2, 1, 2, 3, 4, 4, 2, 0, 0, 0, 0, -2, -2, -4, -4, -4, -2, 0, 0, 1, 2, 2, 2, 3, 2, 2, 0, 0, 1, 1, 1, 1, 1, 1, 1, 3, 3, 4, 2, 0, 0, 0, 0, -2, -2, -3, -4, -2, -1, -1, 1, 2, 1, 2, 2, 2, 2, 2, 1, 0, 0, 0, 1, 1, 0, 1, 2, 3, 3, 2, 1, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 2, 2, 3, 1, 2, 2, 1, 1, 0, 1, 0, 0, 1, 1, 1, 2, 3, 2, 3, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 2, 1, 2, 1, 3, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 1, 1, 2, 2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 2, 2, 1, 2, 2, 1, 2, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 1, 1, 1, 0, 0, 0, 1, 2, 2, 2, 2, 2, 2, 1, 2, 2, 1, 0, 1, 2, 1, 0, 0, -1, 1, 1, 1, 0, 1, 0, 1, 0, 1, 2, 1, 0, 0, 0, 1, 1, 2, 1, 1, 1, 0, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 2, 2, 1, 1, 0, 0, 2, 1, 2, 1, 1, 1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 2, 3, 2, 2, 2, 3, 2, 2, 1, 1, 0, -1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 2, 1, 2, 2, 2, 2, 2, 3, 2, 1, 0, 2, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, -2, -2, -2, -1, 0, 1, 2, 2, 2, 4, 3, 2, 1, 0, 0, 1, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -1, -2, -2, -2, 0, 2, 1, 2, 3, 4, 3, 1, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -2, -1, -1, -2, -2, 0, 0, 1, 1, 3, 2, 3, 3, 1, 0, 0, 0, -1, -2, -2, -3, -2, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 2, 0, 1, 2, 0, -1, 0, 0, -1, -4, -4, -4, -3, 0, -1, -1, -1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -2, -2, -2, -4, -4, -4, -2, 0, -1, -2, 0, 0, 0, 1, 2, 1, 1, 1, 2, 2, 2, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, -2, -2, -2, -2, -2, -2, -2, -2, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 2, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 2, 2, 2, 1, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, 2, 2, 2, 1, 0, 0, 0, 1, 0, 2, 1, 0, 1, 1, 1, 2, 2, 2, 3, 1, 1, -1, -2, 0, 0, 0, 0, 0, 0, -2, -1, 0, 2, 1, 1, 0, 1, 0, 0, 0, 0, 2, 1, 1, 1, 2, 1, 0, 1, 3, 3, 0, 1, -1, 0, -1, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 2, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 2, 1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 2, 1, 2, 1, 1, 0, 2, 0, 0, -1, -1, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 2, 1, 1, 1, 1, 0, 1, 0, 1, 2, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -1, 0, -1, -1, 0, 0, 1, 1, 0, 2, 1, 0, 0, 1, 1, 0, 1, 0, -2, -2, -1, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, -2, -1, -3, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -1, 0, 0, 0, -1, -1, -1, -2, -1, -1, -1, 0, -1, -2, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -1, 0, 0, 0, -1, -1, -2, -1, -1, -2, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -2, 0, 0, -1, 0, 0, -1, -1, -2, -3, -4, -3, -2, -2, -2, -1, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, -1, -2, -3, -3, -2, -2, -3, -1, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 1, 3, 2, 0, 1, -1, -1, -1, 0, -1, -1, 0, 0, -1, -1, -2, -3, -4, -2, -2, -1, -1, 0, -2, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 0, 1, -1, -1, 0, -1, 0, -1, -2, -1, -2, -2, -2, -2, -3, -2, -2, -1, 0, -1, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, -1, 0, -1, -1, -1, -2, -1, -1, -3, -2, -2, -2, -3, -3, -2, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 1, 0, 0, -2, -1, 0, -1, 0, -2, -2, -2, -2, -1, -3, -1, -1, -3, -2, -3, -3, -2, -2, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, 0, -1, 0, -1, -2, -1, -3, -2, -3, -2, -2, -1, -1, -2, -2, -2, -2, -2, -2, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -2, -1, -1, -2, -1, -1, -3, -2, -2, -1, -2, -2, -1, -2, -1, -1, -2, 0, 0, 0, 0, 1, 1, 1, 2, 0, 1, -1, 0, 0, 0, -2, 0, 0, -2, -1, -2, -1, -2, -1, -2, -1, -1, 0, -2, -1, -2, -1, 0, -1, 0, 0, 0, 1, 1, 2, 1, 1, 0, -1, -1, -2, 0, -1, -1, 0, -1, -2, 0, -2, -2, -2, -2, -1, -1, -1, -2, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 2, 2, 0, 1, -1, -1, -1, 0, 0, -2, -1, -1, -1, -2, -1, -1, -2, -2, -1, -1, -2, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 2, 1, 1, 1, 1, 0, 0, -2, -1, -2, -1, -1, -1, -1, -1, 0, -1, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 1, 0, 0, 0, -1, -2, 0, 0, -2, 0, 0, -2, -2, -2, -2, 0, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 1, 2, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, -1, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 2, 1, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 1, 0, 1, 1, 2, 3, 2, 2, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 3, 2, 2, 2, 2, 1, 0, -1, 0, -1, -1, -1, -1, -2, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 2, 2, 1, 2, 1, 2, 3, 3, 3, 2, 1, 0, -1, -1, -1, -2, -1, -1, 0, -3, -1, -3, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 3, 2, 2, 2, 3, 4, 3, 1, 1, 0, -1, -1, -1, -1, -2, -1, -2, -2, -3, -2, -1, -1, -1, -1, 0, 0, 0, 1, 0, 1, 1, 1, 2, 2, 1, 2, 3, 3, 2, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 1, 3, 1, 2, 0, 1, -3, -2, -2, 0, -1, 0, 0, -1, -1, -1, -1, -2, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, 0, 0, 0, -1, 0, 0, 0, -1, -2, -2, -1, -2, 0, -1, 0, 1, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -2, -1, -2, -3, -2, -1, 0, -1, 0, 0, 0, -2, -3, -2, 0, -1, 0, -1, -1, 1, 2, 3, 2, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -2, -2, -1, -1, -1, -2, -2, 0, 0, -1, -2, -1, 0, 0, 0, -1, 0, 1, 1, 3, 1, 1, 1, 2, 0, 1, 0, -1, -1, -1, -2, -2, -4, -3, 0, 0, -1, -2, -1, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 2, 2, 1, 0, 1, 0, -1, -2, -1, -4, -2, -3, -3, -1, -1, -1, -3, -2, -1, -1, -2, -2, -2, -1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 3, 0, 0, 0, 0, -1, -3, -4, -4, -4, -4, -3, -2, -2, -4, -3, -1, -1, 0, -3, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -3, -5, -5, -3, -3, -2, -4, -4, -3, -2, 0, -1, -3, -2, 0, -2, 0, -1, 0, 0, 0, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, -3, -2, -2, -1, -3, -4, -4, -1, 0, 0, -1, -1, 0, -2, 0, -1, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, -1, -2, -3, -3, -3, -3, -1, -3, -4, -3, -2, 0, 0, -1, -1, -1, -1, -2, -1, 0, -1, 0, 0, 0, 2, 2, 1, 0, 0, 0, 0, -2, -1, -2, -2, -2, -1, -2, -1, -3, -4, -4, -1, -1, 0, -2, -2, -2, 0, -1, -1, 0, 0, 0, 1, 0, 1, 2, 1, 0, 1, 1, 0, -2, -2, -1, -1, -1, -3, -1, -1, -2, -2, -2, -2, -1, 0, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 0, -1, 0, 0, -2, -3, -2, -2, -1, 0, -3, -2, -1, -1, 0, -3, -2, -1, 0, -1, 0, 0, 0, -1, 0, 0, 2, 2, 2, 0, 1, 1, 0, 0, 0, 1, 0, -2, -1, -1, 0, 0, -2, 0, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 2, 1, 1, 1, 0, 1, 1, 0, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 3, 2, 1, 0, 1, 2, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -2, -2, -1, -1, -1, -1, -1, 0, 0, 0, 2, 1, 1, 0, 0, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, -1, -2, -1, -1, -1, -1, 0, 0, -2, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, -2, -2, 0, 0, 0, 0, -3, -3, -2, 0, -1, -1, -1, -1, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -2, -2, -2, -4, -2, -1, 0, 0, -2, -2, -2, -1, -1, 0, -2, -2, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 2, 2, 0, 0, 0, -1, -1, -3, -3, -5, -3, -1, 0, -1, -1, -3, -3, 0, -1, 0, -3, -1, -1, -1, -1, 0, -1, 0, -2, -1, 0, 0, 1, 0, 2, 0, -1, -3, -3, -3, -3, -5, -5, -3, -2, -2, 0, -2, -1, -1, 0, 0, -3, -2, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, -1, -3, -4, -4, -4, -4, -5, -4, -2, -1, -1, -2, -1, -1, -1, 0, -3, -2, -2, -2, 0, -1, -2, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, -1, -3, -4, -4, -5, -4, -4, -2, -1, -1, -2, -2, -1, -1, 0, -3, -2, -1, -1, 0, 0, 0, -2, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -2, -4, -4, -4, -5, -3, -3, -1, -2, -2, -2, 0, 0, -1, -2, -2, -2, -2, 0, 0, -1, -1, -2, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, -3, -5, -6, -5, -5, -1, -2, -1, -2, -1, 0, 0, 0, -2, -1, -1, -1, -1, 0, -1, -1, -2, 0, -1, 0, 0, 0, 1, 0, 0, -1, -2, -3, -4, -5, -5, -3, -1, -1, -1, -1, 0, 0, 0, 0, -3, -2, -2, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -3, -2, -3, -3, -3, -1, -1, -1, -2, -1, 0, 0, 0, -2, -1, 0, -1, -1, -1, -2, -3, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -3, -1, -2, -3, -3, 0, -2, -1, -1, -1, 0, -1, -1, -2, -3, -1, 0, 0, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -1, -1, -1, -1, -1, -1, 0, -1, 0, 0, -1, -1, -1, -3, -2, 0, -1, -1, -1, -2, -2, -2, -2, -1, -1, -1, -1, -1, -2, -1, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -4, -2, -3, -3, -3, -1, -2, -2, -3, -3, -2, -3, -2, -2, -1, -3, -3, -2, -2, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, -1, 0, -2, -2, -1, -3, -2, -3, -3, -3, -1, -2, -1, -2, -2, -2, -1, -2, 0, -1, 0, 0, 0, 1, 1, 2, 3, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, -2, -1, -2, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, -1, -2, 0, -1, 0, 0, 0, -1, -1, -1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 2, 0, -1, -1, -1, 0, 0, 2, 2, 2, 2, 2, 1, 0, 0, 1, 3, 2, 1, 0, 0, 1, 0, 0, -2, 0, 0, 0, -1, -1, 0, 3, 3, 2, 0, -1, 0, 1, 1, 2, 1, 2, 3, 3, 1, 2, 0, 0, 4, 4, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 3, 4, 3, 1, 0, 2, 2, 1, 2, 2, 3, 2, 2, 0, 1, 1, 0, 2, 3, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 6, 3, 2, 2, 3, 2, 2, 2, 3, 4, 4, 4, 1, 1, 1, 0, 2, 3, -1, 0, 0, -2, 0, 0, 0, 0, 0, -2, 0, 0, -1, 1, 5, 4, 3, 2, 3, 2, 3, 4, 4, 7, 6, 5, 2, 3, 0, 0, 1, 0, -1, 0, -1, -2, 0, 0, 0, 0, 0, -3, 0, 0, -1, 0, 2, 4, 0, 1, 1, 2, 5, 4, 3, 7, 7, 5, 4, 1, 0, 1, 1, 0, -3, -3, -1, -2, -1, 0, 0, 0, 0, -3, -2, -1, 0, 0, 1, 3, 0, 0, 1, 3, 5, 5, 4, 6, 9, 6, 4, 2, 0, 0, -1, 0, -3, -2, -2, -2, 0, 0, -1, 0, -1, -3, -2, 0, -1, 0, 2, 1, 0, -1, 0, 1, 6, 7, 5, 6, 10, 9, 6, 1, 1, 0, -1, -1, -4, -3, -1, -2, -1, 1, -2, 0, 0, -3, -2, -1, -3, 0, 1, 0, 0, 0, 0, 1, 3, 6, 4, 5, 9, 9, 6, 4, 1, -1, 0, -1, -3, -3, -1, -3, 0, 0, -1, 0, 0, -5, -1, -2, -3, -1, 3, 0, -1, 2, 1, 0, 3, 4, 3, 3, 7, 7, 6, 5, 0, 0, 0, 0, -4, -4, -3, -3, -2, 0, -1, 0, -1, -4, -3, -3, -2, 0, 0, 0, 0, 3, 4, 1, 2, 2, 2, 2, 6, 6, 4, 4, 2, 0, 0, 0, -4, -3, -2, -2, -1, 0, 0, 0, -1, -4, -2, -2, -3, 0, 0, -1, -1, 3, 3, 1, 1, 3, 4, 4, 7, 5, 5, 5, 1, 0, 2, 1, -3, -4, -4, -4, -3, 0, 3, 0, 0, -4, -2, -3, -1, 0, 0, -2, -3, 0, 1, 2, 0, 2, 4, 7, 6, 6, 6, 4, 1, 0, 2, 0, -2, -3, -4, -5, -2, 0, 2, 0, 0, -5, -2, -2, -2, 0, -1, -3, -3, -2, 0, 2, 1, 4, 7, 7, 4, 5, 6, 2, 1, 0, 0, 0, 0, -2, -4, -5, -3, 0, 4, 0, -1, -4, -2, -1, -1, 0, 0, -2, -1, -3, 0, 2, 1, 3, 7, 6, 4, 6, 5, 2, 2, -2, -1, -1, 0, -2, -4, -4, -2, -1, 3, 0, -1, -4, -2, -2, -3, -1, 0, 0, -1, -2, -2, 0, 3, 5, 7, 5, 3, 6, 4, 3, 1, 0, 0, -1, -2, -2, -3, -4, -3, 0, 3, 0, 0, -4, -2, -1, -3, 0, 1, -1, -2, -2, -1, 1, 2, 3, 5, 4, 4, 5, 4, 3, 2, 1, 0, -1, -1, -2, -3, -3, -2, 0, 4, 0, 0, -5, -3, -1, -2, -2, 0, 0, -2, -1, 0, 1, 3, 3, 3, 4, 4, 6, 4, 2, 2, 0, 0, 0, 0, -1, -3, -2, -2, 0, 2, 0, 0, -4, -3, -3, -2, -1, 0, 0, 0, 0, 1, 2, 1, 3, 4, 6, 4, 5, 5, 1, 1, -1, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, -3, -3, -1, -1, -1, 0, 1, -1, -1, 1, 2, 2, 2, 5, 6, 4, 5, 6, 2, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, -3, -2, -2, -1, 0, 0, 0, -3, -2, 2, 2, 1, 2, 5, 5, 5, 5, 7, 2, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -3, -2, -1, 0, -1, 1, 1, -3, -2, 0, 2, 2, 1, 4, 4, 5, 5, 6, 2, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, -4, -3, 0, -1, -1, 0, 0, -1, -2, 2, 2, 2, 2, 3, 3, 3, 6, 6, 1, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -4, -2, 0, 0, -2, 0, -1, 0, 0, 2, 2, 1, 0, 2, 3, 3, 5, 6, 1, 1, 2, 2, 0, -1, -2, 0, -1, 0, 2, 1, 0, 0, -2, -2, 0, 0, -1, 0, 0, 0, 1, 2, 1, 1, 1, 0, 2, 2, 3, 4, 2, 1, 4, 3, 2, 0, -2, 0, 0, 1, 2, 0, 0, -1, -3, -2, 0, 1, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, 1, 1, 3, 2, 2, 1, 4, 3, 1, 0, 0, 2, 0, 0, 1, 0, 0, 0, -3, -2, -1, 1, 1, 1, 0, 0, 0, 0, 0, 4, 3, 0, -1, 2, 3, 2, 1, 1, 5, 4, 1, 0, 0, 2, 1, 1, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 5, 3, 0, 0, 3, 2, 1, 0, 0, 3, 2, 0, -1, 0, 3, 1, 0, 0, -1, 0, 0, -2, -2, -2, 0, 0, -1, -2, 0, 0, 0, 0, 3, 4, 0, 1, 2, 2, 1, 1, 0, 2, 1, 0, 0, 0, 3, 0, 0, 0, -2, 0, 0, -1, -1, -2, -1, 0, -2, -2, -2, -1, -1, -1, 3, 2, 0, 1, 2, 0, 2, 2, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, -2, -1, 0, 0, -1, 0, 1, 0, 1, 2, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 2, 0, 1, 1, 0, 1, 1, 1, 1, 1, 0, 1, 2, 0, 1, 0, 1, 0, 0, -1, -1, 0, -1, -1, -2, -2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 2, 0, 1, 0, 0, -1, 0, -1, -2, -2, -1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 2, 2, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 1, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 1, 2, 3, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 2, 2, 1, 2, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 0, 0, 0, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 3, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 2, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 2, 1, 1, 2, 2, 2, 2, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, -1, 0, -2, -2, -1, -1, 0, 0, 2, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 2, 2, 1, 1, 1, 0, -1, -2, -1, -1, -3, -2, 0, 0, 0, 1, 1, 3, 2, 2, 2, 2, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 2, 1, 0, 0, -1, -1, -2, -1, -3, -2, -2, -1, 0, 0, 0, 3, 1, 3, 2, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 0, 0, -1, -2, -1, -1, -3, -2, -2, 0, 0, 0, 1, 1, 2, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, 1, 2, 2, 2, 1, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 1, 1, 2, 2, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 2, 1, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 1, 2, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 1, 1, 2, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 2, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 1, 0, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, -2, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -1, -1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 1, 2, 2, 0, 0, 0, 0, -1, 0, -2, -2, -3, -2, -3, -4, -1, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 2, 1, 0, 0, 0, 0, 0, -1, -2, -1, -3, -4, -1, 0, 1, 0, 0, 1, 0, 2, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 3, 2, 2, 1, 0, 0, 2, 0, 0, 0, -1, -1, -1, -1, -2, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, -1, -1, -1, -1, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -2, -2, 0, 1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 1, 2, 2, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 2, 2, 0, 1, 1, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 1, 0, 0, 2, 2, 0, 1, 0, 0, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 1, 1, 1, 2, 0, 1, 0, 0, 0, 0, 0, 1, 3, 2, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 2, 1, 2, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 1, 0, 0, -1, 0, 1, 0, 1, 0, 1, 1, 1, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 2, 2, 1, 2, 2, 1, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 3, 2, 3, 2, 1, 1, 0, 0, -1, 0, -2, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 1, 2, 2, 3, 4, 1, 0, 1, 0, 0, -1, -1, -1, -1, -2, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 3, 0, 0, -1, -1, -1, -1, 0, -1, -1, 0, 1, 2, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 3, 1, 0, 0, 0, -2, -2, -1, -2, -3, -2, -2, 0, 0, 2, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 1, 0, 0, -2, -2, -1, -1, -1, -2, -1, -1, 1, 3, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, -1, -1, -2, 0, 0, -1, 0, 0, 2, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 1, 1, 0, 0, -1, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 2, 0, 0, 0, 0, 0, 1, 1, 1, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, -1, 1, 0, -1, -1, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 2, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 2, 2, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, -1, -1, -1, 0, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, -1, 0, 0, 1, 0, 1, 0, 0, -1, -1, 0, -1, -1, -3, -2, 0, -1, -1, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, -2, -1, 0, -1, -2, -2, -2, 0, 0, -1, 0, 0, 0, 0, 1, 2, 1, 3, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -2, -3, -3, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, -1, -1, -1, -1, -2, -2, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, -3, -2, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -2, 0, -1, -2, -2, -3, -2, 0, -1, 0, 0, -1, -1, -2, -1, -2, -3, -3, -3, -4, -2, -1, -1, -1, -1, -2, -1, -1, -1, 0, 0, -1, -2, -2, -1, -2, -3, -2, -1, -1, 0, -1, 0, -2, -1, -1, 0, -2, -2, -4, -4, -3, -4, -3, -3, -2, -2, -1, -1, -1, 0, 0, 0, -2, -3, -1, -2, -1, -2, -1, -1, 0, -1, -1, -2, -2, -2, -2, -1, -2, -3, -2, -3, -4, -2, -2, -1, -1, -2, -1, -2, -1, 0, -1, 0, -1, -2, -2, -1, 0, -1, -1, 0, 0, -1, -1, -1, -2, -1, 0, -2, 0, 0, -1, -1, -2, -2, -2, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, 0, -1, -2, -2, -1, -2, -2, 0, 0, -1, 0, 0, 0, -1, -2, -3, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -2, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -2, -2, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 2, 1, 1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 1, 2, 1, 2, 3, 3, 2, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 1, 2, 2, 3, 4, 3, 1, 2, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 2, 0, 0, 0, 0, -2, 0, 0, 0, 0, 2, 2, 3, 2, 3, 4, 2, 1, 1, 1, 0, 0, -2, -2, -2, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, -1, -2, 0, 1, 1, 1, 2, 2, 1, 2, 2, 3, 1, 1, 1, 0, -1, -1, -2, -2, -3, -2, 0, 0, 0, 1, 1, 1, 2, 0, 0, 1, 0, -2, 0, 0, 1, 1, 1, 1, 1, 3, 3, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 2, 1, 1, 1, 0, 0, 0, 1, 1, 0, 2, 2, 3, 2, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, -1, -1, 0, 0, 0, 1, 1, 3, 3, 4, 4, 3, 1, 1, 1, 0, 1, 1, 1, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 1, 1, 3, 4, 3, 3, 1, 0, 0, 0, 2, 0, 1, 1, 0, 1, 2, 1, 1, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 1, 2, 1, 0, 1, 1, 2, 3, 3, 1, 0, 0, 1, 1, 1, 0, 2, 1, 1, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 1, 0, 1, 1, 2, 2, 1, 1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, -1, 0, 0, 1, 1, 1, 1, 1, 1, 1, 2, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, -2, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -2, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -2, -1, 0, -2, 0, 0, 1, 0, 0, 0, 0, -2, -2, -2, -2, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -2, 0, -1, -2, -1, -1, -1, -1, -1, -1, -1, -1, 0, 0, -2, -2, -2, -2, -4, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -2, -2, -3, -2, 0, 0, -2, 0, -1, 0, 0, 0, -1, 0, -1, -2, -2, -3, -3, -1, 0, -1, -1, -1, 0, 0, 0, -1, -1, -1, -3, -2, -1, -3, -3, -2, -1, 0, -2, -1, -1, 0, 0, 0, 0, 0, -1, 0, -2, -2, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -2, -2, -4, -4, -3, -5, -3, -3, -2, 0, 0, -2, -2, -2, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, -1, -1, -2, -2, -2, -1, -3, -4, -2, -3, -4, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 1, 2, 1, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, -2, -1, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 2, 2, 3, 2, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 2, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 2, 3, 3, 2, 2, 2, 3, 3, 2, 0, 1, 0, -1, -1, -1, -1, 0, 0, -2, -1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 4, 2, 2, 3, 2, 1, 1, 0, 0, 0, -1, -2, 0, -1, 0, -1, 0, 0, 2, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 3, 4, 2, 2, 3, 3, 2, 0, 0, 0, -1, -2, -2, 0, 0, -2, -2, -1, 0, 1, 1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 3, 3, 3, 2, 2, 3, 2, 1, 0, -1, -2, -1, 0, -1, -1, -2, -1, -2, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 1, 2, 2, 3, 3, 3, 2, 1, 1, 1, 0, 0, -1, -1, -1, 0, 0, -1, -3, -2, 0, 0, 1, -1, 0, -2, -1, -1, 0, 0, 0, 0, 0, 3, 2, 1, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 1, 0, 0, -1, -1, -1, 0, -1, 0, 1, 1, 3, 3, 2, 2, 2, 3, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, -2, -2, 0, 0, 1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 2, 3, 2, 3, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -2, -2, -1, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, -1, 1, 2, 3, 3, 2, 3, 0, 1, 0, 0, -1, -2, 0, 0, 0, 0, -1, -1, -2, 0, 0, 1, -1, -2, -2, -1, -1, 0, -1, 0, 0, 0, 0, 2, 2, 2, 3, 3, 1, 1, 0, 1, 0, 0, -1, -1, -1, -1, -1, -1, -1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 2, 2, 3, 2, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 0, 0, 1, 1, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, -2, -1, 0, 0, 0, 2, 2, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, 0, 0, 0, 1, 0, -2, -1, -1, -2, -1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, 0, -1, -1, 0, 1, 0, 0, 0, -1, -2, -2, -1, 0, 0, 1, 0, -2, 0, -2, -1, 0, -1, -2, -1, 0, 1, 2, 3, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, -1, -1, 0, 1, 1, 0, 0, -1, -2, -1, 0, 0, 0, -1, -2, 0, 1, 3, 3, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -2, -1, 1, 0, 1, 0, 0, -1, -1, -1, -1, 0, -1, -1, 0, 0, 2, 2, 2, 2, 2, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -2, 0, 0, 1, 1, 0, -2, 0, 0, 0, -1, -1, 0, -1, -1, 0, 1, 1, 3, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, 0, -1, -1, 0, 0, 0, 1, 2, 2, 3, 1, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 2, 0, -1, -1, -2, 0, 0, -1, 0, 0, 0, 0, 2, 1, 1, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, -2, -1, -2, -1, 0, -1, 0, 0, 1, 2, 2, 2, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 0, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, -1, 0, -1, 1, 0, 1, 1, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, -1, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, -1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 2, 1, 2, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 2, 0, 1, 1, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 2, 1, 2, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 2, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 2, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 1, 1, 2, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 2, 2, 2, 2, 3, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 3, 3, 3, 3, 4, 2, 2, 2, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 2, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 3, 3, 2, 3, 3, 3, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 1, 0, 0, -1, 0, -2, -1, -1, 0, 0, -1, 1, 0, 0, -1, -1, 0, -1, -1, -1, 0, 1, 0, 0, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, -2, -2, -2, -2, -1, -1, -1, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -2, -3, -3, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -4, -2, -2, -1, -2, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -2, -3, -3, -2, -3, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, -2, -2, -3, -1, -1, -3, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, -1, -3, -3, -3, 0, 0, -2, -2, -1, -1, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, 0, -1, -2, -2, -2, -4, -3, -1, -1, -1, -1, -3, -1, -2, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, -1, 0, -1, -3, -4, -3, -5, -2, -1, -2, -1, -1, -2, -2, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -2, 0, -1, 0, 0, -1, -2, -2, -4, -4, -4, -4, -3, -1, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, -1, -2, -2, -3, -3, -4, -3, -2, -1, 0, -1, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, -3, -2, -3, -2, -4, -3, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -2, -2, -1, -1, -1, 0, 0, 0, -2, -3, -2, -2, -4, -3, -2, -2, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, -3, -3, -3, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -2, -3, -2, -1, -1, -1, 0, 0, 1, 0, 1, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, -3, -3, 0, 0, 0, 0, 0, 0, 2, 0, 0, -2, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 0, -1, 0, 0, -1, -2, -2, -3, -1, -2, 0, 0, 1, 1, 1, 2, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, -1, 0, 0, 0, 0, -2, -2, -1, -1, 0, 1, 1, 2, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 2, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 2, 2, 2, 1, 1, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 1, 2, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -2, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -2, 0, -1, 0, 0, 0, -1, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, -2, -1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, 0, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -3, -3, -4, -2, -2, -3, -2, -2, -3, -2, -3, -2, -3, -3, -3, -2, -3, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 2, 2, 1, 0, 0, -3, -6, -5, -5, -5, -3, -3, -3, -5, -3, -4, -2, -4, -5, -4, -4, -4, -2, -2, 0, 0, 1, 1, 0, 0, 0, 0, 3, 3, 3, 2, 1, -5, -5, -4, -4, -4, -3, -5, -4, -5, -2, -1, -2, -3, -3, -4, -4, -3, -1, -1, 1, 2, 3, 3, 3, 0, 0, 3, 3, 4, 2, 3, 0, -4, -6, -6, -4, -3, -5, -5, -5, -5, -4, 0, 0, -1, -2, -4, -4, -3, 0, -1, 0, 2, 1, 2, 3, 1, 0, 2, 3, 3, 2, 3, 0, -4, -7, -5, -6, -5, -5, -3, -5, -4, -3, -1, 0, 0, -2, -3, -2, -2, -1, 0, 0, 1, 2, 0, 3, 0, 0, 1, 2, 3, 2, 1, 1, -3, -7, -6, -4, -4, -4, -4, -5, -5, -3, -3, -1, 0, -1, -1, -1, -3, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 2, 0, -3, -6, -6, -5, -3, -4, -3, -3, -4, -4, -4, -3, -2, -1, -2, -1, -3, -1, 0, 2, 2, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -3, -6, -4, -4, -4, -3, -3, -2, -4, -3, -2, -4, -3, -3, -3, -3, -3, -1, 0, 1, 2, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, -4, -4, -5, -5, -4, -4, -4, -3, -3, -3, -3, -2, -4, -4, -3, -3, -2, -2, 0, 1, 1, 1, 1, 1, 2, 0, 0, -1, -2, 0, 1, 0, -3, -6, -5, -4, -4, -5, -4, -5, -5, -4, -4, -2, -4, -3, -3, -1, -1, -1, -2, 0, 0, 1, 0, 1, 1, -1, 0, -1, -3, 0, 0, 0, -4, -6, -5, -4, -4, -4, -3, -3, -3, -5, -4, -4, -4, -2, -2, -1, 0, -1, -1, -1, 1, 1, -1, 0, 0, 0, 0, -2, -1, 0, 0, 0, -2, -5, -5, -4, -5, -4, -2, -3, -4, -4, -4, -4, -3, -1, -1, -2, 0, 0, -1, 0, 2, 1, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, -4, -5, -6, -4, -3, -5, -4, -3, -3, -4, -3, -4, -4, -2, -2, -2, 0, 1, 0, 0, 4, 2, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -3, -6, -5, -3, -4, -3, -3, -4, -4, -3, -4, -5, -3, -1, -2, -1, 0, 1, 1, 1, 5, 3, 1, 0, -1, 0, 0, 2, 1, 1, 1, 0, -3, -4, -4, -4, -5, -4, -3, -3, -4, -2, -3, -4, -4, -3, -1, 0, 0, 0, 1, 2, 5, 4, 1, 0, 0, -1, 0, 1, 4, 3, 1, 0, -2, -5, -4, -5, -5, -5, -3, -4, -3, -2, -3, -4, -4, -1, 0, 0, 1, 0, 0, 3, 4, 4, 2, 0, 0, 0, 0, 1, 3, 3, 1, 0, -4, -5, -5, -4, -4, -5, -3, -4, -4, -2, -3, -2, -5, -3, -1, 0, 0, 1, 0, 0, 2, 3, 1, 0, 1, 0, 0, 0, 2, 3, 3, 0, -3, -5, -4, -5, -4, -4, -4, -4, -4, -3, -3, -2, -3, -3, -1, -1, 0, 0, 0, -1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, -4, -6, -4, -4, -5, -3, -4, -5, -5, -4, -3, -3, -3, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 0, -5, -6, -5, -4, -5, -4, -5, -5, -6, -5, -5, -3, -3, -1, -1, 0, -1, -1, -1, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 2, 2, 0, -5, -6, -5, -5, -5, -5, -5, -5, -5, -5, -4, -3, -4, -2, -1, 0, 0, -1, -2, -1, -2, -1, 0, 0, -2, -1, 0, 2, 1, 2, 2, 0, -3, -6, -5, -4, -4, -4, -4, -5, -4, -4, -4, -4, -3, -2, 0, -1, 0, -1, -1, -2, -2, 0, 0, -1, -2, 0, 0, 1, 2, 3, 2, 0, -4, -5, -5, -6, -4, -4, -5, -4, -4, -5, -4, -5, -4, -4, -1, -2, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 2, 1, 2, 1, 0, -3, -5, -5, -5, -5, -5, -4, -4, -4, -5, -4, -4, -3, -4, -3, -3, -1, 0, 1, 0, -1, 0, 0, -1, 0, 0, 2, 1, 2, 2, 1, 0, -3, -6, -6, -5, -5, -5, -4, -5, -6, -5, -3, -5, -3, -4, -2, -2, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 2, 3, 1, 4, 3, 0, -2, -5, -5, -5, -5, -4, -5, -5, -5, -3, -3, -3, -3, -2, -3, -2, -1, 0, 0, 1, 0, 1, 0, 0, 0, 3, 2, 2, 2, 4, 3, 0, -4, -4, -5, -5, -4, -4, -6, -6, -5, -4, -3, -3, -1, -2, -3, -2, -1, -1, 0, 0, 0, 1, 0, 0, 1, 2, 3, 2, 3, 3, 4, 1, -2, -5, -5, -4, -5, -4, -6, -7, -7, -4, -3, -4, -2, -2, -3, -3, -2, -1, -1, 0, 1, 1, 1, 0, 1, 2, 3, 4, 2, 4, 4, 0, -2, -4, -5, -5, -3, -3, -6, -6, -7, -5, -4, -5, -4, -5, -4, -3, -2, -3, -1, 0, 0, 1, 1, 1, 1, 2, 5, 5, 3, 4, 3, 1, -4, -5, -5, -4, -6, -4, -7, -8, -6, -6, -6, -7, -5, -6, -6, -5, -3, -4, -4, 0, 0, 1, 3, 2, 3, 3, 6, 6, 4, 3, 3, 1, -4, -6, -6, -6, -7, -7, -8, -8, -8, -8, -7, -8, -8, -8, -6, -5, -4, -4, -3, 0, 0, 1, 3, 3, 4, 4, 6, 7, 6, 5, 5, 2, -2, -3, -4, -4, -4, -5, -5, -3, -6, -4, -4, -5, -4, -4, -4, -4, -2, -1, -1, 0, 0, 0, 2, 3, 2, 1, 4, 4, 5, 2, 3, 2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, -1, -1, -1, -2, -2, -2, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 2, 1, 3, 2, 1, 1, 0, 0, -1, -2, -1, -2, -1, 0, 0, -1, 0, 0, 2, 2, 0, 0, 1, 0, 1, 2, 3, 2, 2, 1, 4, 3, 3, 4, 4, 3, 4, 1, 0, -1, -2, -1, -2, -2, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, -2, -1, -1, 0, 1, 0, 0, 2, 3, 3, 3, 4, 4, 5, 1, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, -1, -2, -2, -2, -2, 0, 0, 0, 1, 2, 4, 4, 6, 5, 4, 2, 0, 0, 0, 0, 0, 0, 1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -1, -1, 0, 0, 2, 3, 4, 6, 5, 4, 2, 1, 0, 0, 0, 0, 1, 1, 1, -2, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 2, 4, 5, 4, 1, 0, 1, 0, 0, 0, 1, 1, 0, -1, -2, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 2, 0, 2, 2, 2, 1, 1, 1, 1, 0, -1, -2, -1, 0, 0, -1, 0, 0, 1, 2, 2, 3, 2, 1, 0, 0, 2, 1, 0, 0, 0, 1, 1, 1, 1, 1, 3, 3, 3, 3, 1, 0, -2, -2, -1, 0, 0, 0, 1, 1, 1, 2, 2, 2, 2, 1, 1, 1, 2, 2, 1, 1, 0, 0, 0, 2, 2, 2, 2, 3, 2, 3, 2, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 2, 2, 1, 0, 1, 2, 3, 1, 0, 0, 0, 0, 0, 2, 3, 4, 4, 2, 3, 1, 0, 0, -2, 0, 1, 1, 0, 2, 2, 2, 2, 2, 1, 0, 1, 1, 1, 3, 2, 1, 1, 0, 0, 0, 1, 0, 1, 3, 4, 4, 3, 3, 1, 0, -1, 0, 0, 1, 2, 1, 2, 2, 2, 1, 1, 1, 0, 1, 1, 1, 1, 0, -1, 0, 1, 2, 1, 1, 1, 2, 4, 3, 5, 4, 2, 0, 0, 0, 1, 1, 0, 0, 1, 2, 3, 3, 3, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 2, 1, 2, 3, 3, 4, 5, 4, 3, -1, -1, 0, 1, 0, 1, 0, 1, 0, 2, 4, 4, 2, 1, 1, 2, 0, -2, -1, -2, -2, 0, 0, 0, 2, 2, 2, 3, 3, 3, 5, 3, -1, -1, 0, 1, 2, 1, 1, 0, 1, 3, 3, 4, 2, 1, 1, 1, 0, -2, -4, -4, -2, -2, 0, 1, 1, 2, 3, 3, 4, 5, 4, 4, -1, -1, 0, 0, 1, 0, 0, 0, 0, 2, 3, 4, 3, 1, 1, 0, -1, -2, -4, -3, -3, -1, 0, 0, 1, 3, 5, 4, 5, 4, 4, 3, -1, -2, -1, 0, 1, 1, 0, 0, 2, 2, 2, 2, 2, 1, 0, 1, 0, -2, -4, -4, -2, -2, 0, 1, 2, 3, 4, 5, 5, 4, 5, 2, -1, -2, 0, 1, 0, 1, 0, 0, 0, 2, 2, 0, 0, 1, 0, 2, 0, -1, -2, -2, 0, 0, 0, 1, 0, 2, 2, 4, 5, 4, 3, 3, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 1, 2, 2, 0, -1, 0, 0, 1, 0, 0, 2, 1, 1, 4, 4, 3, 2, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 1, 1, 2, 1, 0, 1, 0, 0, 0, 1, 2, 2, 1, 3, 3, 3, 2, 1, 0, -1, 1, 0, 1, 0, 0, 0, -1, 0, 2, 2, 1, 1, 3, 1, 1, 0, 1, 1, 0, 1, 1, 1, 0, 2, 1, 2, 2, 0, 1, 0, -1, 0, 0, 0, 0, 0, -2, -1, -2, -1, 0, 2, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 2, 0, 1, 1, 0, 0, -1, 0, 1, 0, 0, 0, -1, -1, -1, 0, 1, 1, 1, 1, 2, 0, 0, 0, -1, -1, 2, 0, 0, 1, 1, 2, 2, 1, 0, 1, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 1, 0, 0, 1, 1, 0, -1, -1, 0, 0, 1, 3, 2, 2, 1, 1, 2, 3, 2, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 2, 3, 3, 3, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, 0, -2, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 1, 2, 3, 3, 2, 2, 2, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -3, -2, -2, -3, -1, -1, 0, 0, 1, 2, 2, 3, 3, 3, 2, 3, 1, 2, 1, 0, -1, 0, 0, -2, -1, 0, -1, -1, -1, -1, -1, -2, -2, -3, -2, -3, -2, -1, -1, 0, 0, 2, 3, 4, 2, 2, 1, 1, 0, 1, 1, -1, 0, -2, 0, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 2, 3, 1, 2, 1, 0, 1, 1, 0, -2, -1, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 1, 1, 1, 1, 1, 0, 1, 1, 1, 0, 0, 0, -1, -1, -2, 0, 0, -1, -1, -1, -2, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 2, 2, 1, 1, 1, 1, 1, 0, 1, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 2, 2, 3, 2, 1, 0, 0, 0, -1, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 3, 2, 3, 3, 4, 4, 2, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, -1, -1, -1, -2, -3, -1, 0, 0, 0, 1, 3, 3, 3, 3, 5, 3, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, -1, -2, -2, -2, -3, -2, -1, -1, 0, 2, 2, 3, 4, 4, 5, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, -1, 0, -2, -2, -2, 0, 0, 0, 2, 2, 4, 5, 4, 1, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 2, 3, 4, 2, 2, 1, 0, 0, 2, 1, 1, 0, 0, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 0, 1, 1, 0, 2, 2, 2, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 3, 2, 2, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 2, 2, 3, 3, 1, 1, 0, -1, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 2, 1, 1, 0, 0, 0, 0, 0, 1, 2, 3, 2, 3, 3, 2, 0, -1, 0, 0, 0, 1, 2, 1, 2, 0, 1, 1, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 1, 1, 1, 1, 3, 3, 3, 3, 2, 0, -1, -1, 0, 0, 0, 1, 1, 0, 2, 2, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 2, 1, 2, 2, 1, 3, 3, 4, 4, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 3, 3, 1, 0, 1, 1, 0, -1, -1, 0, 0, -1, 0, 1, 1, 2, 1, 1, 3, 4, 3, 3, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 2, 3, 2, 1, 1, 0, 0, -1, 0, -1, -2, 0, -1, 0, 0, 3, 3, 4, 2, 3, 3, 3, 1, -1, -1, 0, 0, 0, 1, 1, 1, 2, 2, 2, 3, 1, 0, 2, 0, 0, -1, -3, -2, -2, -2, 0, 0, 2, 3, 3, 2, 4, 2, 3, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 2, 3, 2, 1, 1, 0, 0, -1, -1, -2, -2, -2, -1, 0, 0, 1, 2, 3, 4, 5, 3, 3, 1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 2, 3, 1, 0, 0, 1, 1, -1, -2, -2, -2, -2, -1, 0, 0, 1, 2, 3, 4, 4, 4, 3, 1, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 1, 0, 0, 1, 0, 1, -1, -1, 0, -1, -1, 0, 1, 2, 2, 2, 3, 3, 3, 2, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 1, 2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 2, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 1, 1, 1, 2, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 2, 2, 3, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 1, 2, 1, 2, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, -1, -2, -1, -1, 0, 0, 0, 2, 2, 2, 2, 2, 2, 1, 2, 2, 0, 0, -1, 0, 0, -2, 0, 0, 0, -1, -1, -1, -2, -2, -2, -3, -2, -2, -2, 0, 0, 0, 1, 2, 1, 2, 1, 2, 1, 2, 0, 0, 0, 0, -1, -1, -1, -2, -2, 0, -2, -1, -1, -2, -1, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, 2, 2, 2, 1, 0, 1, 0, 1, 0, -1, -1, 0, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -2, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -2, 0, -1, 0, -2, -1, -2, 0, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, -2, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -2, -1, 0, -1, -2, 0, 0, 0, -2, 0, -1, 0, -1, 0, 0, 0, 1, 2, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -2, -1, -2, -1, 0, 0, -3, -2, 0, -1, 0, -1, 0, -1, 2, 0, 1, 1, 2, 0, 0, 0, 1, 0, -2, -2, -1, -2, -1, -2, -2, -2, -1, -2, -2, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, -1, -2, -2, -1, -2, 0, -2, -3, -1, -2, -1, 0, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -3, -3, -3, -3, -2, -2, -4, -3, -3, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -2, -1, -3, -2, -3, -3, -1, -3, -2, -3, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, -2, -2, -2, -2, -2, -3, -2, -2, -2, -1, 0, -1, -1, -1, -2, 0, 0, -1, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, -2, 0, -2, -1, -1, -1, -1, -2, -2, -2, -3, -2, -2, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 2, 0, 1, 0, 0, -1, 0, -1, -2, 0, -2, -3, -2, -1, -2, -2, -2, -2, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -2, -2, -2, -2, -2, -2, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 0, 2, 1, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, -2, -2, -2, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -2, -1, -1, 0, -1, -1, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 1, 0, -1, -2, -2, 0, -1, -1, -2, -2, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -2, -2, -2, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 2, 0, 0, 2, 2, 0, 0, 0, 0, 1, 0, 1, 0, 0, -2, 0, -1, -2, -1, 0, -2, -2, 0, -1, -1, 0, 0, -1, 0, 1, 1, 1, 1, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -2, 0, 0, -1, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, -2, -1, 0, -1, -1, -1, 0, 0, -1, 1, 1, 0, 1, 0, 1, 1, 0, -1, 0, 0, -2, -3, -2, -1, -1, -1, -2, -3, -2, -2, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, -1, -1, -1, -2, -1, -3, -3, -2, -1, 0, -2, -2, -1, -3, -1, -1, -1, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -2, -1, -2, -1, -2, -2, -2, -1, -1, -2, -2, -3, 0, -2, 0, -2, 0, -2, -1, 0, -1, -1, -1, -1, 0, 1, 0, 1, 1, 1, 0, -1, -2, -2, -2, -3, -2, -3, -2, -2, -2, -2, -3, -1, -2, -1, 0, -2, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, -1, 0, -2, -2, -2, -3, -3, -3, -1, -2, -2, -2, -2, 0, 0, -1, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, -2, -1, -2, -3, -3, -3, -1, -1, -2, -1, -3, -2, -1, 0, -1, 0, -1, 0, 0, -1, -2, -1, 0, 0, -1, 0, 1, 0, 1, 0, -2, -2, -3, -1, -2, -3, -4, -2, -1, -1, -1, -3, -2, 0, 0, 0, -2, -1, 0, -1, 0, -1, -2, 0, 0, 0, 0, 0, 1, 1, 0, -1, -2, -2, -2, -3, -2, -3, -3, 0, -2, -2, -1, -1, -1, 0, -1, -1, -3, -2, 0, -1, -1, -2, -1, -1, -1, 0, 1, 0, 0, 1, 0, 1, -1, -2, -1, -2, -2, -3, -1, -1, 0, -2, -2, -1, -1, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, -2, 0, -2, -1, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -2, -2, -2, -1, 0, -2, -1, -2, -1, -1, -1, -1, -2, -1, 0, 0, -2, -1, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -2, -1, -1, -2, -1, -1, -1, -1, -2, -1, -2, -2, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 2, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 2, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 1, 2, 1, 1, 2, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 2, 2, 2, 2, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 3, 3, 2, 1, 2, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 3, 2, 1, 2, 1, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 2, 2, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 3, 2, 1, 1, 0, 0, 0, 0, -1, 1, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 3, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 2, 2, 2, 1, 1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 2, 2, 2, 1, 1, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 1, 3, 2, 1, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 1, 3, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 2, 2, 2, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 1, 1, 1, 3, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 1, 1, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 1, 1, 0, 1, 2, 2, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 2, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 1, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 1, 2, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, 1, 1, 1, 2, 2, 1, 1, 1, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 3, 4, 1, 0, 1, 2, 0, 2, 2, 1, 2, 1, 2, 1, 0, 0, 0, 2, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 3, 2, 2, 0, 1, 3, 1, 1, 1, 2, 0, 1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 2, 3, 2, 2, 0, 0, 2, 2, 2, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 1, 1, 1, 1, 2, 4, 4, 3, 2, 1, 1, 0, 0, 0, -1, 0, 0, -1, -1, -2, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 2, 1, 0, 1, 1, 2, 3, 2, 1, 2, 3, 0, 0, -1, 0, 0, 0, -1, -2, -2, -1, 0, 1, 0, 0, 1, 0, 0, 1, 1, 2, 2, 1, 1, 0, 0, 0, 3, 5, 3, 0, 2, 2, 1, 0, 0, -1, -2, 0, -2, -3, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 3, 2, 1, 2, 2, 0, 0, 0, 0, 0, -1, -2, -3, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 0, 1, 2, 0, 1, 2, 1, 0, 2, 1, 2, 2, 0, -1, -1, -1, -1, -2, -1, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -2, -2, -2, -2, 0, 0, 1, 0, 0, -1, 0, 0, -1, 1, 1, 1, 0, 2, 4, 3, 2, 1, 1, 0, 0, 0, 1, 0, -1, -1, 0, 1, -1, -1, -1, -2, 0, 0, 1, 0, 1, -2, 0, 0, 0, 0, 1, 0, 1, 1, 3, 4, 3, 0, 0, 1, 0, 1, 0, 0, -1, -1, 0, 1, 0, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 3, 2, 1, 1, 1, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, -2, -1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 1, 1, 0, 0, 0, 1, 0, 0, 0, -2, 0, 0, 0, -2, 0, 0, 0, 1, 0, 0, -2, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, 1, 0, 1, -1, -1, -1, 0, -1, 0, 0, 0, 1, 1, 2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, -1, 0, 1, 0, 1, 1, 1, 1, 0, 1, 0, 1, 0, 1, 0, -1, -1, 0, 1, -1, 0, 0, 0, 1, 0, -1, 0, -1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 2, 0, 0, 1, 0, 2, 2, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 0, 1, 2, 2, 2, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 1, 0, 0, 1, 0, -1, -1, 0, 0, -1, 0, 2, 1, 0, 0, 0, -1, -1, -2, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 1, 0, -1, 0, 1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 2, 1, 2, 0, 0, 2, 0, 0, -1, 0, 0, 0, 2, 0, 0, 0, -2, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 1, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 3, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 1, 2, 2, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 2, 2, 2, 2, 1, 1, 1, 2, 2, 4, 3, 2, 0, 0, -1, -1, 0, -1, -1, 0, 0, -2, -1, -2, 0, 0, -1, -2, -1, -1, -1, 0, 1, 2, 1, 2, 3, 2, 0, 1, 3, 3, 1, 3, 1, -1, -1, -2, -1, 0, 0, -1, -2, -2, -1, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, 1, 2, 2, 2, 1, 1, 1, 2, 3, 3, 1, 1, -1, 0, -2, -1, -1, 0, -2, -1, -1, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 2, 1, 2, 2, 2, 2, 2, 3, 1, 2, 0, -1, -1, -1, -1, -2, -2, 0, -1, 0, -2, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 2, 2, 1, 2, 2, 2, 1, 2, 3, 1, 1, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 2, 2, 1, 2, 1, 1, 2, 3, 2, 2, 2, 1, 0, -2, -2, -1, -1, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 2, 1, 1, 0, 2, 1, 2, 1, 0, 0, 1, -1, 0, -1, 0, -1, -1, 0, -1, 0, -1, -1, 0, -1, -1, -2, -1, -2, -1, -1, 0, 1, 1, 1, 0, 2, 1, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -2, -1, -2, -1, 0, 0, 1, 1, 2, 2, 2, 0, 1, 1, 1, 0, 0, -1, -1, -1, -1, 0, -1, 0, -1, 0, -1, -1, -2, -3, -2, -1, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -2, -2, -1, 0, 0, -1, -1, -1, -1, -2, -2, -1, -1, -2, -3, -2, -1, -2, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, -2, -1, -1, 0, -1, 0, 0, 0, -2, 0, -2, -2, -1, -3, -2, -3, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, -1, -1, -1, -1, -1, 0, 0, 0, -2, -1, -1, -2, -3, -2, -2, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -2, -1, -2, -2, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, -1, -2, -2, -3, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, -2, 0, -2, -2, -2, -2, -1, -2, -2, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, -2, 0, -1, 0, -1, -1, -1, -2, 0, -1, -1, -1, -3, -2, -2, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, -1, -1, -1, -1, -1, 0, -1, -1, -1, -1, -2, -1, -2, -2, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, -2, 0, -1, 0, -1, -1, 0, -2, -2, -2, -1, -2, -2, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -2, -1, -1, -2, -1, 0, 0, -1, -1, -1, -1, -1, -1, 0, -1, -1, -2, -1, -1, 0, 0, 1, 0, 1, 1, 1, 1, 2, 0, 1, 1, 0, -1, 0, 0, -1, 0, -1, -1, -2, 0, 0, -2, 0, 0, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 2, 0, 0, -1, -1, 0, -1, -1, 0, -1, -2, -2, 0, -2, -1, 0, -1, 0, -1, -1, 0, 0, -1, 0, 1, 1, 1, 1, 1, 2, 1, 2, 2, 1, 0, -1, -1, -1, 0, 0, 0, -1, 0, -2, -1, -2, -1, -2, -1, -1, -1, -2, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, -1, -2, -1, 0, 0, 0, -2, -1, 0, -1, 0, -1, -1, -1, -1, -1, -2, -1, 0, 1, 1, 0, 1, 1, 0, 0, 1, 1, 3, 2, 1, 0, 0, 0, -2, -1, -1, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 1, 0, 2, 2, 2, 1, 2, 0, 0, 0, -1, 0, 0, 0, -1, -2, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 2, 2, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 3, 1, 1, 1, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 2, 1, 1, 2, 3, 1, 2, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 1, 1, 3, 2, 2, 1, 0, 0, 0, -2, 0, 0, 0, -1, -1, -1, -2, 0, -1, -2, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 2, 2, 2, 3, 3, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -2, -2, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 2, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 2, 2, 2, 0, 0, 0, 3, 2, 1, 0, 0, 0, -2, 0, 0, -1, -1, -2, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, 0, 1, 1, 2, 2, 2, 1, 0, -1, -1, -1, 0, -1, -2, -1, -2, -1, -2, -2, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 3, 1, 1, 0, 1, 0, 2, 1, 1, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, -2, -2, 0, -1, -2, 0, -1, -1, 0, 0, 0, 1, 2, 3, 1, 1, 2, 1, 2, 1, 1, 0, 1, 0, -2, -2, -1, -1, 0, 0, 0, -1, -2, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 1, 2, 1, 1, 1, 1, 2, 3, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 2, 2, 2, 3, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 1, 0, 0, 2, 2, 3, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, -1, -2, -2, -1, -1, -1, -1, 0, 0, 1, 0, 0, 2, 2, 1, 0, 1, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -2, -2, 0, -2, -1, -1, -1, 0, 0, 1, 2, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, -1, 1, 1, 0, 0, 0, 0, 1, 2, 2, 1, 0, -1, 0, 1, 0, 0, 1, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -2, -2, -2, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -3, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 2, 2, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 2, 1, 2, 2, 2, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4, -4, -4, -3, -3, -2, -2, -4, -3, -3, -4, -3, -3, -4, -4, -5, -4, -2, -2, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 2, 2, 0, -5, -7, -4, -3, -5, -4, -4, -4, -5, -4, -3, -4, -4, -5, -5, -4, -5, -3, -1, 0, 0, 1, 2, 1, 0, 0, 1, 2, 3, 3, 3, 0, -6, -5, -5, -4, -4, -3, -4, -5, -5, -4, -3, -3, -3, -4, -4, -5, -4, -2, 0, -1, 0, 0, 2, 2, 1, 1, 1, 3, 3, 3, 2, 2, -5, -6, -5, -5, -4, -3, -4, -5, -5, -4, -3, -3, -2, -3, -4, -4, -3, -2, -1, 0, 0, 1, 1, 3, 1, 1, 3, 2, 4, 2, 3, 0, -5, -6, -5, -4, -3, -2, -3, -3, -5, -4, -2, -2, -3, -4, -4, -3, -3, -3, -1, 0, 0, 2, 1, 3, 1, 1, 1, 1, 1, 2, 1, 1, -6, -6, -5, -5, -4, -4, -4, -3, -4, -4, -2, -3, -3, -3, -3, -3, -2, -2, 0, 1, 2, 2, 1, 2, 1, 0, 0, 0, 1, 1, 2, 0, -5, -5, -3, -3, -3, -2, -2, -3, -3, -4, -3, -3, -3, -2, -3, -1, -1, -2, -1, 1, 1, 2, 2, 0, 1, 0, 1, 0, 1, 0, 0, 0, -5, -5, -4, -4, -2, -3, -2, -3, -2, -3, -3, -2, -2, -3, -3, -3, -3, -3, -1, 0, 1, 2, 0, 2, 1, 0, 1, 0, 1, 0, 1, 0, -5, -3, -3, -3, -3, -3, -2, -3, -2, -2, -2, -2, -2, -3, -3, -3, -2, -2, -1, 1, 1, 1, 1, 1, 1, 1, 0, 1, -1, 1, 2, 0, -4, -3, -4, -3, -2, -2, -2, -2, -3, -3, -2, -3, -2, -4, -3, -2, 0, -1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -3, -3, -3, -3, -2, -3, -2, -2, -2, -2, -3, -3, -4, -2, -2, -2, 0, 0, -1, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 1, -3, -4, -3, -3, -3, -1, -2, -1, -3, -2, -2, -3, -3, -3, -3, -2, 0, 0, 1, 0, 1, 2, 1, 1, 0, 1, 0, 0, 1, 2, 0, 0, -4, -5, -3, -4, -2, -3, -3, -2, -2, -3, -2, -3, -1, -2, -2, -1, 0, 0, 0, 1, 2, 2, 1, 1, 0, 0, 2, 1, 0, 2, 2, 0, -5, -4, -4, -2, -3, -3, -3, -3, -2, -2, -1, -2, -2, -1, -1, 0, 0, 1, 0, 1, 2, 2, 2, 1, 1, 1, 1, 1, 2, 1, 1, 0, -3, -4, -3, -2, -3, -1, -1, -2, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 2, 3, 3, 2, 2, 1, 0, 0, 2, 2, 3, 1, 0, -4, -4, -3, -3, -4, -2, -2, -1, -1, 0, 0, -2, -2, -2, 0, 0, 1, 1, 1, 1, 4, 3, 3, 1, 0, 0, 0, 1, 2, 3, 1, 0, -4, -3, -2, -2, -2, -3, -1, -2, -1, 0, -1, -1, -1, -1, -1, 0, 1, 1, 0, 2, 3, 3, 1, 1, 0, 0, 1, 1, 1, 3, 2, 0, -5, -3, -2, -3, -3, -3, -3, -2, -1, -1, 0, -1, -2, -1, 0, 0, 1, 2, 1, 0, 2, 1, 1, 0, 0, 0, 1, 1, 1, 2, 1, 0, -4, -4, -4, -3, -2, -3, -1, -3, -3, -1, -1, -1, -1, -2, 0, 1, 2, 0, 0, 0, 0, 2, 1, 0, 0, 0, 1, 0, 1, 2, 2, 1, -5, -5, -3, -4, -2, -3, -2, -2, -2, -2, -2, -1, -1, -2, -1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 2, 1, -3, -3, -4, -4, -4, -3, -2, -1, -3, -3, -2, -3, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, -4, -5, -3, -4, -2, -2, -2, -3, -3, -2, -1, -2, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 1, 0, -3, -4, -4, -4, -2, -2, -3, -3, -2, -4, -2, -1, -1, -1, -2, -1, -1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 1, 1, 2, 2, 1, 0, -3, -4, -4, -4, -2, -3, -3, -3, -4, -3, -3, -3, -2, -3, -2, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 1, 1, -4, -4, -3, -4, -3, -2, -3, -4, -3, -3, -2, -2, -1, -3, -1, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 2, 1, 2, 2, 1, -4, -4, -4, -2, -3, -4, -4, -3, -3, -3, -3, -1, -2, -3, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 1, 1, 1, 2, 2, 0, -3, -4, -4, -3, -3, -3, -4, -3, -3, -3, -3, -2, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 2, 2, 2, 1, -4, -3, -4, -2, -2, -4, -3, -5, -3, -3, -2, -3, -2, -3, -3, -1, -1, -1, -1, -1, 0, 0, 0, 0, 1, 2, 1, 1, 1, 2, 4, 2, -4, -4, -3, -3, -3, -4, -3, -4, -4, -4, -4, -3, -4, -4, -3, -3, -1, -2, -2, 0, 0, 0, 0, 1, 0, 1, 3, 3, 1, 3, 3, 2, -4, -5, -5, -5, -3, -5, -5, -4, -4, -5, -4, -5, -5, -4, -5, -3, -3, -3, -3, -1, -1, 0, 0, 1, 0, 2, 3, 2, 1, 2, 3, 1, -4, -4, -5, -5, -4, -5, -4, -6, -4, -5, -5, -5, -6, -6, -5, -6, -5, -5, -4, -2, -2, 0, 0, 0, 0, 1, 1, 1, 2, 1, 3, 2, -3, -3, -4, -4, -2, -3, -4, -4, -4, -4, -4, -4, -4, -4, -4, -3, -3, -3, -3, -2, 0, 0, 0, 0, 0, 1, 2, 1, 1, 2, 1, 0,
    -- filter=0 channel=1
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 2, 1, 1, 0, 2, 2, 2, 2, 1, 1, 2, 1, 2, 1, 0, 1, 2, 2, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 2, 1, 1, 2, 1, 2, 1, 1, 0, 1, 1, 0, 1, 1, 1, 0, 0, 2, 1, 0, 1, 0, 1, 0, 0, 1, 0, 1, 2, 0, 1, 2, 1, 2, 2, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 1, 0, 1, 0, 1, 0, 0, -1, -1, -1, -2, -3, -1, -1, -1, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 2, 0, 2, 0, 1, 1, 1, 1, 0, -1, -1, -3, -3, -2, -3, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, -2, -1, -2, -2, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -2, -2, -1, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -2, -1, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 1, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 2, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 1, 1, 0, 1, 1, 1, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, -2, -1, 0, 1, 1, 1, 0, 1, 0, 0, 0, -1, 0, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, -2, -2, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -3, -2, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -3, -2, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -3, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -3, -3, -3, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, -1, -1, -1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, -1, -2, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -2, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, -2, 0, 0, 0, 1, 1, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -1, 0, 1, 1, 2, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, -1, 0, -1, -1, -1, 0, 0, 0, 1, 2, 2, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 1, 1, 1, 1, 2, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -1, 0, -1, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -1, -1, 0, 0, 1, 1, 1, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, -2, -2, -1, 0, 1, 1, 2, 2, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, -2, -3, -1, 0, -1, 0, 1, 0, 1, 1, 1, 2, 1, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -2, -3, -2, -1, -1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 0, 2, 0, 1, 1, 0, 1, -1, -2, -1, -1, 0, 0, 1, 1, 1, 2, 1, 1, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 1, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 2, 2, 1, 1, 0, 1, 0, 0, -1, 0, 2, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 2, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 1, 0, 1, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 2, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, 0, 0, 0, 0, 1, 1, 2, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -2, -1, -1, 0, 0, 0, -1, -1, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 0, 0, 1, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, -1, -1, -1, -1, 0, -1, -1, 0, -1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, -2, -1, -2, -1, -1, -1, 0, -1, -1, -1, 0, -2, -1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, -2, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, -1, -2, -2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -2, -1, 0, -1, -2, -1, -1, 0, 0, 1, 1, 2, 1, 0, 1, 1, 1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -2, -2, -3, -1, -2, 0, -1, -1, 0, -1, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, -3, -2, -2, -1, -1, -1, 0, 1, 2, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, -2, -1, -2, -2, -2, -1, -1, 0, 0, -1, 0, 0, 0, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, -1, -2, -3, -1, 0, -2, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, 0, -1, -1, -1, -2, -1, 0, -1, 0, 0, 0, 0, 2, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, -1, -2, -1, 0, 0, -2, -1, -1, -2, -1, -1, -1, 1, 1, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, -1, -2, -2, -2, 0, -2, -1, -1, -2, -2, 0, -1, 0, 0, 0, 1, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, -3, -2, -1, -2, -1, -2, -2, 0, 0, 1, 0, 1, 1, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, -2, -2, -1, 0, 0, -1, -1, -1, 1, 2, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -2, -2, 0, 0, -1, -1, 0, 0, 0, 2, 1, 0, 1, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -2, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -2, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, -1, -2, -1, -3, -2, -2, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -2, -1, -3, -3, -3, -3, -3, -3, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -3, -3, -2, -2, -2, -2, -2, -2, -2, -2, -2, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, -2, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 2, 2, 2, 2, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 3, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 2, 2, 1, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 1, 1, 1, 0, 2, 2, 2, 2, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 2, 1, 0, 2, 2, 1, 0, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 1, 2, 1, 2, 3, 2, 1, 1, 2, 2, 1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 1, 1, 0, 1, 2, 1, 3, 1, 3, 2, 3, 3, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 2, 4, 3, 2, 3, 3, 3, 3, 2, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 2, 1, 2, 3, 1, 4, 3, 1, 2, 2, 2, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 5, 3, 2, 3, 2, 1, 2, 1, 1, 0, 0, 1, -1, -2, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 3, 3, 3, 3, 2, 2, 3, 2, 3, 2, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 2, 3, 4, 3, 1, 1, 3, 3, 2, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 2, 3, 3, 2, 1, 1, 1, 3, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 1, 1, 1, 2, 2, 4, 3, 0, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 3, 2, 1, 0, 1, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 3, 2, 2, 0, 1, 2, 1, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 2, 2, 2, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 1, 1, 2, 0, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 3, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 2, 1, 2, 2, 0, 1, 0, -2, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, -2, -1, -2, -1, -1, -1, 0, 0, 0, 0, 3, 3, 4, 3, 3, 2, 1, 1, 0, 0, 0, -1, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, -2, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 1, -1, -2, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 4, 2, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 0, 1, 3, 2, 0, 0, -1, 0, -1, -1, -1, 0, 1, 3, 4, 3, 4, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 4, 2, 2, 0, 0, -1, -1, -2, -2, -1, 1, 1, 4, 3, 3, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 2, 2, 3, 2, 0, -1, 0, -2, -2, -3, -2, 0, 1, 3, 4, 2, 2, 0, -1, -2, -2, -2, -2, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 3, 2, 1, 0, -1, -1, -2, -3, -2, -2, 0, 2, 2, 4, 2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, -2, -1, -2, -2, 0, 2, 3, 3, 3, 2, 0, 0, 0, -2, 0, -1, -1, 0, 0, 0, -2, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, -1, -2, -2, -1, 0, 0, 2, 2, 4, 4, 2, 2, 1, 0, -1, -1, -1, -1, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -2, -3, -1, 0, 1, 2, 3, 5, 5, 3, 3, 0, 0, -2, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, -2, -2, -2, 0, 0, 3, 3, 4, 4, 3, 1, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -2, -3, -2, -1, 0, 0, 1, 3, 4, 3, 3, 1, 0, 0, -3, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, -1, 0, -2, -3, -4, -2, -1, 0, 0, 0, 4, 3, 4, 1, 1, 1, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -4, -2, -2, -1, 0, 0, 3, 4, 3, 2, 1, 1, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -3, -2, -2, -1, -1, 0, 0, 3, 2, 3, 2, 1, 1, 1, 1, 0, 0, -1, -1, -1, 0, -1, 0, 1, 0, 0, -1, 0, 0, 1, -1, -2, -3, -1, -2, -1, -1, 0, 1, 2, 2, 3, 1, 1, 2, 0, 0, 1, 0, -1, -2, -1, -1, 0, 0, 0, 2, 0, 0, 0, 1, 0, 1, -1, -3, -3, -3, -2, -1, 0, 0, 1, 2, 2, 1, 1, 1, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, -2, -2, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 0, 0, -2, -3, -3, -2, -2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 2, 0, 0, -1, -2, -2, -3, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, -1, -1, -2, -2, -1, -1, 1, 0, 2, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, -1, 0, -1, -1, -1, 1, 1, 1, 2, 1, 0, 1, 0, 0, -1, 0, -1, -2, -1, -1, -1, -1, -2, 0, 1, 1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, -2, -1, -1, -2, -1, -2, -3, -2, -1, 0, 0, 2, 1, 0, 0, 1, 2, 0, 1, 0, 0, 1, 0, 2, 1, 1, 1, 0, -1, 0, -2, -2, -1, -1, -1, -2, -1, -2, -1, -2, 0, 0, 1, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -2, -3, -3, -2, -1, -1, 0, 0, -1, -2, -2, -1, 0, 2, 2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 1, 0, 0, -1, -1, 0, -2, 0, -2, -1, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -2, -1, -2, 0, 0, 0, 1, 1, 0, 0, 2, 1, -2, -3, -3, -5, -4, -5, -4, -2, -1, -1, 0, 2, 1, 1, 0, 0, 1, 0, -1, -2, -3, -3, -2, -1, 0, 1, 1, 1, 1, 2, 1, 0, -2, -6, -4, -5, -6, -4, -5, -4, -3, -2, 0, 1, 1, 2, 0, 1, 0, 1, 0, -1, -3, -1, -1, -2, 0, 0, 2, 0, 2, 2, 0, 0, -1, -4, -2, -3, -3, -3, -3, -1, -2, -1, 0, 0, 0, 0, -1, 1, 1, 1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -2, 0, 0, 0, 0, 1, 3, 3, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 2, 1, 0, 1, 2, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 3, 4, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 1, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 3, 3, 3, 5, 3, 2, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 2, 3, 1, 1, 3, 2, 1, 0, 0, 0, -2, -3, -2, 0, 0, 1, 2, 3, 4, 4, 3, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 2, 2, 1, 2, 4, 4, 3, 0, 0, 0, -2, -3, -3, -2, 0, 1, 3, 3, 3, 4, 3, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 2, 1, 2, 3, 4, 2, 0, 0, 0, -1, -1, -1, 0, 0, 1, 3, 4, 2, 2, 2, 1, 0, 0, 1, 0, -1, -1, 0, 0, -1, 0, 1, 1, 1, 2, 3, 3, 2, 0, 0, 0, 0, 0, 0, 0, 2, 2, 3, 4, 3, 3, 2, 2, 1, 1, 1, 1, 0, -1, 0, -1, 0, -1, 0, 1, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 4, 4, 5, 3, 4, 3, 3, 1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 1, 1, 1, 0, 0, -1, -2, 0, 0, 1, 1, 2, 4, 5, 5, 6, 4, 4, 5, 4, 2, 0, 0, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, 1, 0, -1, -3, -1, -2, -1, 1, 2, 2, 1, 2, 4, 6, 7, 6, 5, 4, 4, 2, 0, -1, 0, 0, -1, -1, -1, -1, -2, -2, 0, 0, 0, -1, -2, -3, -3, -3, 0, 1, 1, 1, 3, 4, 4, 6, 6, 5, 5, 3, 2, 1, 0, -1, -1, 0, 0, -1, -1, -1, -2, -2, 1, 0, 0, -1, -3, -3, -2, -1, 0, 0, 1, 0, 2, 4, 3, 4, 5, 3, 5, 2, 3, 1, 1, 0, 0, 0, -1, 0, -1, -3, -2, -1, 1, 1, 0, 0, -3, -3, -1, 0, -1, 0, 0, 0, 2, 1, 2, 4, 4, 3, 3, 3, 3, 2, 2, 0, 0, 0, 0, 0, -1, -2, -2, 0, 2, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, 1, 1, 2, 3, 3, 5, 4, 4, 2, 3, 2, 1, 1, 1, 1, 0, -2, -2, -2, -1, 1, 2, 0, -1, -2, -2, 0, 0, 0, -1, -1, 0, 0, 0, 1, 2, 3, 5, 4, 3, 3, 2, 1, 1, 1, 0, 0, -1, -2, -1, -2, 0, 2, 1, 0, 0, -1, -1, 1, 1, 0, 0, -1, -1, -1, 0, 0, 1, 1, 3, 2, 2, 2, 2, 2, 0, 0, 0, -1, -2, -1, -2, 0, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -2, 0, 1, 1, 1, 1, 0, 2, 3, 2, 1, 1, 0, 0, -1, -1, -1, 0, 0, 2, 3, 0, 0, 0, 0, 2, 1, 0, 0, -2, -3, -4, -2, 0, 1, 1, 0, 1, 1, 2, 2, 2, 1, 0, 0, -1, 0, 0, 0, 2, 2, 2, 1, 0, 1, 1, 2, 0, 0, 0, 0, -2, -3, -3, -2, 0, 1, 1, 0, 0, 1, 3, 3, 1, 0, 0, 0, 0, 0, 1, 2, 0, 2, 3, 3, 1, 1, 2, 1, 0, 0, -1, -1, -1, -3, -3, -2, 0, 1, 0, 1, 1, 3, 3, 2, 0, 0, 0, 0, 0, -1, 1, 0, 1, 2, 3, 2, 0, 0, 1, 0, 0, -2, -2, -1, -1, -1, -1, 0, 1, 2, 1, 1, 1, 1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 1, 0, 2, 3, 2, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 1, 2, 2, 1, 1, 0, 1, 2, 0, 0, -3, -2, -3, -3, -1, -1, 0, 0, 0, 0, 3, 1, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 1, 2, 2, 2, 0, 1, 0, 1, -1, -1, -4, -3, -3, -1, -2, -3, -3, -3, -1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 2, 1, -1, -1, -1, -1, -1, -3, -4, -3, -3, -2, 0, -1, -2, -2, -1, 1, 3, 1, 0, -1, -2, -1, 0, 0, 0, -1, -1, 0, 1, 2, 1, -1, -2, -2, -2, -3, -3, -3, -1, -1, -1, 0, 0, 0, -2, -1, 0, 2, 3, 1, 0, -1, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, -1, -1, -1, -2, -3, -2, -3, -1, 0, 0, 1, 2, 1, 0, 0, 1, 3, 2, 3, 1, -1, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 1, 1, 1, 2, 2, 1, 2, 1, 2, 0, 0, 0, -1, -1, -2, -2, -2, -1, -1, 0, -2, -2, -2, -1, -1, -2, -1, -1, -2, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, 0, -1, -1, -1, -1, -2, -1, -1, -3, -4, -4, -4, -3, -1, -2, -3, -1, -2, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, -1, -2, 0, -1, -3, -2, -1, -3, -2, -1, -2, -1, -2, -3, -4, -4, -2, -2, -1, -1, -1, -1, -3, -1, -2, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, -1, -3, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, 0, -1, -1, 0, 0, -1, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 0, 1, -1, -1, -1, -1, -1, 0, -1, -1, -2, -1, 0, 0, -1, 0, -1, -1, 0, 0, 1, 2, 2, 1, 0, 0, 0, 1, 1, 0, 2, 1, 3, 1, 0, 0, -1, -1, -1, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, -1, -1, 1, 0, 1, 2, 2, 1, 0, 0, 2, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 1, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 2, 2, 2, 1, 1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 1, 0, 0, -2, 0, 0, -1, -2, 0, 0, 0, 0, 0, 1, 0, 1, 1, 3, 2, 2, 3, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 4, 4, 3, 3, 1, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 4, 4, 5, 3, 4, 1, 0, 0, -1, -1, -2, 0, 0, 0, 0, 1, 0, 1, 0, -1, -2, -1, 0, 0, -1, 0, 0, 0, 1, 0, 2, 2, 4, 4, 4, 3, 3, 2, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, -1, -2, -1, -1, 0, 1, 0, -1, -1, 1, 1, 2, 1, 3, 4, 4, 2, 3, 3, 1, 0, -1, -1, -1, -2, -2, 0, 0, 0, 1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 1, 1, 3, 3, 3, 3, 4, 3, 3, 3, 3, 0, 0, 0, -1, -2, -3, 0, 0, 1, 0, 2, 0, 0, -2, -1, 0, 0, 1, 0, -1, 1, 0, 1, 2, 5, 4, 3, 4, 4, 3, 4, 1, 1, 0, -1, 0, -2, -2, -1, 0, 0, 0, 2, 0, -1, -2, -2, 0, 0, 1, 0, 0, 1, 3, 3, 4, 4, 3, 4, 3, 4, 2, 2, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 2, 2, 3, 3, 4, 3, 3, 2, 3, 2, 2, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, -1, -2, -1, 0, 0, 0, -1, 0, 1, 2, 2, 2, 3, 3, 2, 2, 2, 2, 3, 1, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 2, 3, 2, 2, 2, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 1, 1, 1, 2, 3, 3, 1, 2, 2, 2, 2, 1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 2, 3, 2, 1, 2, 3, 1, 1, 0, 1, 0, -2, 0, 0, 0, -1, -1, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 1, 2, 1, 1, 1, 2, 2, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 2, 2, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -2, -2, -2, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 2, 1, 2, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, -2, -2, -3, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 1, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, -2, -3, -3, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -2, -2, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -3, -3, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -2, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -1, -1, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, -2, -2, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -2, 0, -1, -1, -3, -2, -2, -1, -1, -3, -2, -2, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -2, -2, -1, -1, -2, -1, -1, -2, -2, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 1, 0, -1, -1, -1, 0, 0, -2, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, -3, -3, -3, -3, -3, -1, 0, -1, -1, -1, 0, 1, 0, 0, 0, 1, -1, -1, -2, -2, -4, -4, -3, -1, -1, -1, 0, 0, 0, 0, -4, -6, -7, -8, -7, -6, -4, -3, -3, -1, -1, 0, 1, 1, 0, 2, 2, 3, -2, -3, -4, -4, -4, -3, -3, -2, -3, -2, 0, 1, 1, -1, -4, -6, -8, -9, -8, -6, -5, -2, -2, -1, 0, 0, 0, 0, 0, 1, 3, 3, -2, -2, -3, -2, -3, -2, -1, -1, 0, 0, 1, 2, 2, 2, 0, -3, -5, -5, -6, -5, -2, -1, 0, 0, 0, 0, -2, -1, -2, 1, 3, 3, -2, -2, -1, -2, -1, -1, -1, 0, 0, 1, 2, 4, 5, 3, 0, 0, 0, 0, -1, -2, 0, 1, 1, 1, 0, -2, -2, -4, -2, 0, 3, 2, -1, -2, -2, 0, 0, -1, 0, 0, 0, 0, 1, 4, 4, 4, 3, 2, 2, 1, 0, -1, 0, 0, 2, 2, 0, 0, -2, -2, -2, 0, 2, 3, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 3, 3, 5, 5, 3, 4, 4, 1, 0, 0, 0, 1, 1, 0, 0, -2, -1, -1, 0, 3, 3, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 2, 4, 6, 6, 6, 6, 4, 3, 2, 0, 0, 0, 1, 0, -2, -1, -2, 0, 0, 3, 2, -1, 0, 1, 2, 1, 0, 1, 1, 0, -1, -2, 0, 3, 5, 5, 5, 6, 4, 4, 0, 0, 0, 0, 1, 0, -2, -2, 0, -1, 0, 1, 1, -2, 0, 1, 2, 2, 2, 0, 0, 0, -1, -2, 1, 2, 5, 5, 4, 6, 4, 3, 1, 0, 0, 0, 0, -1, -2, -3, 0, 0, 0, 2, 2, -2, 0, 3, 3, 2, 0, 0, -1, -1, -1, 0, 1, 4, 6, 6, 7, 4, 3, 1, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, -1, 0, 1, 1, 2, 0, 0, -1, 0, 0, 2, 2, 5, 7, 7, 7, 6, 2, 1, 1, -1, -1, 0, 0, -1, -2, -2, -1, -1, -1, 0, 0, -1, 1, 2, 0, 0, -1, 0, 0, 1, 2, 2, 4, 6, 7, 7, 6, 6, 4, 3, 2, -1, -1, -1, 0, -2, -3, -2, -3, -3, -2, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 3, 4, 3, 4, 7, 8, 8, 7, 6, 3, 2, 2, 0, -2, -1, -1, -1, -3, -2, -3, -3, -1, 0, 0, -2, 0, -1, -1, -1, -1, 0, 1, 4, 4, 4, 5, 6, 7, 8, 8, 8, 3, 1, 0, -1, -3, -2, -1, -2, -2, -2, -2, -2, -2, 0, 0, -1, 0, -1, -3, -2, -1, 0, 2, 3, 5, 4, 6, 6, 8, 7, 8, 8, 4, 1, 0, -2, -3, -2, -2, -1, -1, -3, -3, -2, 0, 0, 0, -1, -1, -2, -4, -3, 0, 1, 3, 4, 3, 5, 5, 6, 8, 7, 8, 8, 4, 1, 0, -1, -2, -1, -1, -1, -1, -3, -3, -3, -1, 1, 1, -1, -2, -2, -3, -3, 0, 2, 2, 4, 3, 5, 6, 5, 5, 7, 8, 7, 5, 2, 0, 0, -1, 0, 1, 0, -2, -3, -4, -3, 0, 1, 1, -1, -1, -2, -4, -2, 1, 2, 3, 2, 2, 4, 4, 3, 4, 5, 7, 7, 5, 3, 0, 0, 0, 0, 0, 0, -2, -4, -4, -3, 0, 2, 2, 0, -1, -2, -3, -2, 0, 2, 1, 1, 2, 2, 3, 2, 3, 4, 7, 7, 4, 3, 1, 2, 0, 0, 0, 0, -4, -4, -5, -3, 0, 1, 3, -1, 0, -1, -2, -2, 1, 2, 2, 1, 1, 2, 2, 1, 2, 4, 6, 7, 4, 1, 2, 2, 2, 0, 0, -2, -3, -5, -4, -2, 0, 2, 2, -1, 0, -2, -1, 0, 2, 3, 1, 0, 0, -1, 1, 1, 3, 3, 4, 2, 2, 0, 2, 3, 1, 0, -2, -2, -4, -4, -3, -1, 1, 3, 2, -1, 0, 0, 0, 0, 1, 3, 2, 0, -1, 0, 1, 1, 3, 3, 1, 1, 0, 0, 1, 1, 1, 0, -2, -3, -4, -3, -3, 0, 2, 3, 3, 0, 0, 0, 0, 0, 2, 2, 2, 0, -1, 0, 1, 2, 4, 4, 2, 2, 1, 0, 0, 1, 0, 0, 0, -2, -4, -4, -3, -1, 0, 3, 4, 0, 1, 1, 1, 0, 1, 0, 1, 0, -1, 0, 2, 2, 5, 4, 4, 3, 2, 1, 1, 0, -1, 0, -1, -1, -4, -3, -3, 0, 0, 4, 4, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, 2, 3, 5, 5, 4, 5, 5, 2, 0, 0, -1, -1, -1, -2, -3, -5, -3, -1, 0, 3, 2, -1, 0, 0, -1, 0, -1, -1, -1, -2, 0, 0, 3, 4, 3, 4, 4, 4, 3, 2, 0, 0, -1, -2, -2, -4, -4, -6, -5, -3, -1, 3, 3, 0, 0, 0, -1, 0, 0, -1, -2, -3, -2, 0, 2, 2, 1, 2, 2, 2, 1, 0, 0, -1, -1, -1, -3, -3, -4, -5, -5, -2, 0, 4, 2, 0, -1, 0, 0, -2, -2, -2, -2, -2, -1, 0, 1, 0, -1, 0, -1, -2, -1, -1, -2, -1, -2, -2, -2, -2, -4, -2, -2, -1, 1, 5, 3, 0, -1, -1, -1, -1, -2, -3, -2, -3, -3, -1, -1, -1, -2, -4, -4, -4, -4, -3, -3, -1, -2, 0, -1, -1, 0, 0, 0, 1, 4, 6, 5, 0, 0, 0, -1, -1, -1, -1, -2, -2, -4, -3, -3, -4, -3, -4, -6, -5, -4, -5, -3, -1, 0, 0, 0, 0, 1, 2, 1, 2, 5, 6, 4, 0, -1, -1, 0, -1, -1, -1, 0, -1, -1, -2, -1, -1, -3, -2, -3, -3, -2, -2, 0, 0, 1, 1, 1, 1, 0, 0, 3, 2, 2, 4, 2, 0, 0, -1, 0, 0, 0, 1, 1, 2, 1, 2, 3, 3, 2, 1, 1, 2, 0, 2, 1, 2, 3, 2, 3, 3, 5, 4, 5, 5, 3, 3, 0, 0, 0, -2, 0, 0, 1, 2, 2, 3, 3, 5, 4, 3, 3, 2, 1, 2, 2, 3, 3, 3, 5, 4, 4, 3, 3, 5, 5, 6, 8, 6, 3, 0, 0, 0, 0, 0, 1, 2, 4, 3, 3, 5, 4, 2, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 2, 2, 3, 6, 7, 6, 2, 0, 1, 0, 1, 0, 1, 2, 5, 5, 4, 2, 1, 0, 1, 0, 0, -2, -3, -3, -6, -4, -4, -2, -2, -2, -1, 0, 2, 3, 6, 4, 2, 0, 0, 0, 0, 0, 2, 2, 3, 4, 3, 0, 1, 0, 0, 0, -1, -2, -2, -5, -6, -6, -5, -5, -2, -2, -1, 0, 0, 3, 6, 5, 3, 1, 0, 0, 1, 0, 1, 0, 2, 1, 1, 0, 0, 1, 2, 1, 1, 0, 0, -4, -6, -6, -5, -4, -3, -2, -1, 0, 1, 3, 5, 3, 3, 1, 2, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 3, 1, 0, 0, -2, -5, -4, -4, -3, -2, 0, 0, 1, 2, 2, 4, 4, 2, 1, 2, 0, 2, 0, 0, 0, -1, -2, -3, -2, -1, 0, 3, 3, 2, 2, 2, 0, -3, -3, -3, -3, -3, 0, 0, 0, 1, 0, 3, 4, 2, 1, 2, 2, 1, 0, 0, 0, -1, -3, -5, -4, -2, 0, 1, 3, 3, 4, 2, 0, -3, -3, -3, -3, -3, -1, 0, 1, 0, 1, 3, 2, 2, 0, 3, 2, 3, 2, 2, 0, -2, -3, -5, -6, -3, -1, 1, 1, 3, 4, 1, 0, -2, -3, -3, -4, -3, -3, -1, 0, 0, 0, 1, 2, 1, 0, 2, 2, 3, 1, 1, 0, -2, -3, -4, -4, -3, -2, 0, 2, 3, 3, 2, 0, 0, -1, -3, -2, -3, -3, 0, 0, 0, 1, 1, 3, 2, 0, 2, 1, 1, 2, 1, 0, -1, -4, -5, -6, -4, -2, 0, 2, 3, 3, 3, 1, 1, 1, 0, -2, -3, -2, -3, 0, -1, 0, 2, 3, 1, 1, 1, 1, 1, 0, 0, 0, -2, -4, -5, -5, -5, 0, 2, 2, 2, 3, 4, 3, 4, 1, 0, 0, -2, -3, -3, -1, -3, 0, 2, 1, 1, 1, 1, 0, 0, -1, -1, 0, -3, -5, -5, -6, -4, -1, 1, 3, 3, 4, 4, 4, 4, 2, 1, 0, -2, -3, -3, -2, -3, -2, 0, 2, 1, 0, 0, 0, 0, -1, -2, -2, -3, -6, -8, -6, -5, -1, 1, 4, 4, 3, 4, 2, 1, 2, 0, -1, -3, -4, -3, -2, -1, -1, 0, 1, 2, 0, 0, -2, 0, 0, -1, -1, -5, -7, -8, -7, -6, -2, 0, 1, 2, 2, 3, 2, 2, 0, 0, -1, -3, -5, -3, -2, -3, -2, 1, 1, 1, 0, 0, 0, -1, 0, -1, -1, -4, -8, -8, -7, -5, -1, 0, 3, 3, 2, 1, 2, 0, 2, 0, -2, -3, -4, -5, -4, -3, -2, 0, 2, 1, 1, 1, 0, 0, 0, 0, -2, -4, -8, -8, -6, -5, -1, 0, 2, 4, 3, 2, 1, 1, 2, 0, 0, -3, -4, -5, -4, -2, -2, 2, 2, 1, 0, 1, -1, 0, 0, -1, -3, -4, -5, -7, -5, -6, -2, 0, 2, 3, 4, 4, 1, 0, 1, 0, -1, -4, -5, -5, -5, -2, -1, 1, 2, 2, 0, 1, -1, 0, 0, 0, 0, -3, -5, -7, -6, -5, -1, 1, 3, 3, 4, 3, 1, 0, 0, -2, -2, -4, -5, -5, -4, -1, 1, 4, 3, 3, 0, 0, 0, 0, 0, 0, -1, -3, -5, -5, -5, -4, -3, 0, 3, 4, 3, 1, 1, 0, -2, -2, -4, -4, -5, -4, -2, 0, 2, 4, 4, 2, 0, 1, 1, 3, 2, 1, -1, -4, -5, -6, -7, -4, -1, 0, 1, 3, 4, 3, 0, 0, -2, -2, -4, -4, -4, -3, 0, 2, 3, 4, 4, 4, 1, 2, 3, 2, 2, 0, -1, -3, -5, -7, -6, -3, -3, 0, 1, 1, 3, 2, 1, 0, -2, -3, -5, -4, -2, -2, 0, 3, 5, 5, 4, 3, 0, 3, 3, 3, 1, 0, -2, -3, -5, -5, -4, -2, -1, 0, 2, 2, 2, 0, -1, -1, -1, -4, -4, -3, -3, -1, 1, 3, 4, 5, 4, 2, 2, 2, 0, 1, 1, -1, -3, -3, -3, -5, -4, -1, -1, 1, 2, 1, 0, -1, -3, -3, -3, -5, -5, -3, -2, 0, 1, 4, 5, 6, 5, 3, 0, 0, 0, 1, -1, -2, -2, -2, -3, -3, -3, -1, 0, 1, 3, 2, 0, -2, -5, -6, -5, -5, -5, -4, -2, 0, 1, 3, 4, 7, 5, 2, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -2, 0, 1, 0, 1, 1, 0, -4, -6, -8, -8, -6, -4, -2, 0, 0, 0, 3, 5, 6, 6, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -3, -5, -7, -8, -7, -6, -4, -3, 0, 0, 1, 2, 3, 7, 6, 3, 0, 0, -2, 0, 1, 1, 1, 2, 2, 2, 0, 1, 0, 0, 0, -1, -2, -4, -6, -6, -4, -2, -1, 0, 0, 2, 3, 2, 4, 8, 6, 3, 0, 0, -2, -1, 0, 1, 2, 1, 2, 1, 2, 2, 0, 0, -1, -1, -2, -3, -4, -3, -2, 1, 2, 3, 3, 4, 4, 5, 6, 8, 6, 3, 0, -1, -3, 0, 0, 0, 1, 0, 2, 3, 3, 3, 1, 0, 0, 0, 0, 0, 0, 0, 2, 4, 4, 6, 5, 5, 7, 7, 7, 7, 5, 1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 2, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 3, 3, 3, 3, 3, 3, 3, 2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 1, 1, 2, 1, 2, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 2, 2, 1, 0, -1, -1, 0, 0, -1, 0, 1, 1, 2, 2, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, -1, -1, -1, 0, 0, 1, 2, 1, 2, 0, 0, 0, 0, 0, 1, 2, 2, 1, 2, 1, 0, 0, 0, 1, 2, 2, 0, 0, 0, 1, 1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, 0, -1, 0, 2, 1, 1, 1, 1, 0, 1, 1, 1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 1, 2, 1, 2, 3, 1, 0, 0, -1, 0, 2, 2, 2, 2, 2, 0, 0, 1, 0, 1, 1, 0, 1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 0, 2, 2, 0, 1, 2, 2, 3, 3, 1, 2, 1, 0, 1, 1, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 1, 1, 1, 0, 1, 0, 0, 1, 1, 2, 3, 3, 2, 1, 0, 0, 0, 1, 1, 1, 4, 5, 3, 1, 0, 1, 0, 0, 0, 0, 1, 1, 2, 2, 1, 1, 0, 0, 0, 0, 1, 1, 3, 2, 2, 0, 0, 0, 2, 3, 1, 3, 4, 5, 4, 1, 1, 1, 0, 0, 0, 1, 1, 2, 3, 1, 2, 0, 0, -1, 0, 0, 1, 1, 2, 1, 2, 1, 1, 1, 1, 0, 1, 2, 3, 4, 3, 1, 0, 0, 2, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, 0, -1, 0, 2, 3, 3, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 0, -1, 0, 0, 0, -1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 2, 3, 3, 0, 0, 0, 1, 1, 1, 0, 0, 0, 2, 2, 2, 0, -1, -2, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 2, 3, 3, 0, 0, 0, 1, 2, 1, 1, -1, 0, 0, 1, 2, -1, -1, -2, -2, -1, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 1, 1, 2, 2, 1, 0, -1, 0, 0, 2, 0, -1, 0, 1, 1, 1, 0, -2, -1, -2, 0, -1, 0, 0, 0, 2, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -2, -3, -1, 0, -1, 0, -1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 2, 0, -1, 0, 0, 1, 1, 0, -2, -2, -1, -1, -2, 0, 0, 1, 3, 2, 0, 0, -1, 0, 1, 1, 2, 2, 0, 1, 1, 0, 0, 0, 0, 1, -1, 1, 0, 0, 0, 0, 0, -2, -2, -2, -1, -2, -2, 0, 1, 2, 0, 1, 0, 0, 1, 2, 2, 2, 1, 0, 0, 2, 0, 0, 1, 1, 0, 2, 2, 1, 1, 0, 0, 0, 0, -1, 0, -2, -2, -1, 0, 1, 0, 1, 0, 0, 1, 3, 3, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, 0, 0, -1, -1, -2, -2, -1, 0, 0, 2, 1, 0, 1, 0, 3, 4, 5, 2, 2, 1, 0, 0, 1, 0, 0, 0, -1, 1, 2, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 2, 2, 1, 2, 1, 4, 6, 5, 2, 2, 0, -1, 0, 0, 0, 0, 0, -1, 0, 2, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 2, 2, 2, 4, 3, 3, 3, 2, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 1, 2, 1, 2, 2, 3, 3, 2, 4, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 3, 2, 2, 3, 1, 2, 2, 1, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 3, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 0, 1, 1, 0, 0, 0, 2, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 2, 2, 1, 1, 2, 0, 0, 0, 2, 3, 1, 0, 0, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 2, 2, 3, 2, 2, 2, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, -1, -1, 0, -1, 0, 1, 3, 3, 3, 3, 2, 0, 0, 0, 0, 1, 0, 0, 0, -2, -2, -1, 0, 0, -2, -2, -1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 3, 4, 5, 2, 2, 0, 1, -1, -1, -1, -1, -3, -3, -3, -4, -3, -3, -3, -2, -1, 0, 0, 3, 2, 2, 1, 1, 1, 2, 2, 2, 2, 3, 2, 3, 3, 1, 0, 1, 0, -1, -3, -4, -5, -6, -5, -5, -4, -3, -3, -3, -2, -1, 0, 0, 0, 2, 0, 1, 2, 2, 2, 1, 2, 2, 1, 0, 1, 0, 0, 1, 0, 0, -1, -2, -2, -4, -3, -3, -3, -3, -3, -2, -2, -1, 0, 0, -1, 0, -1, 1, 1, 1, 1, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 2, 1, 1, 2, 1, 2, 1, 1, 0, 0, -1, -1, -2, 0, 0, 0, 1, 1, 1, 2, 2, 3, 1, 1, 0, 0, 1, 0, 1, 2, 0, 0, 1, 1, 0, 2, 1, 2, 3, 2, 1, 0, 0, 0, 0, -1, 1, 0, 1, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -2, -4, -3, -3, -1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, -3, -2, -2, -2, -2, -2, -3, -2, 0, 0, 1, 1, 0, 1, 2, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, -3, -1, -2, -1, -1, 0, 2, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, -1, -2, -1, -1, -2, -1, 0, 0, 0, 0, 1, 2, 1, 0, 2, 2, 1, -1, 0, -1, -1, -2, -2, -1, -1, 0, 1, 0, 2, 2, 0, 0, -1, -1, -1, -2, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, 3, 2, 1, 1, 0, 0, -1, -2, -4, -3, -2, 0, 0, 0, 2, 2, 0, 0, -2, -3, -2, -2, -3, -3, -1, 0, 0, 0, 0, 1, 0, 1, 3, 3, 2, 1, 0, -1, -2, -2, -4, -5, -2, -1, 0, 1, 2, 1, 0, -1, -2, -2, -3, -2, -3, -3, -1, 0, 0, -1, -1, 0, 0, 1, 1, 2, 0, 0, 0, -1, -2, -2, -3, -4, -2, -1, -1, 0, 1, 0, 1, 0, -2, -1, -2, -3, -4, -3, -1, 0, -1, -1, 0, 0, 0, 0, 2, 0, 1, 0, 0, -1, -1, -2, -5, -4, -4, -2, -1, 0, 1, 1, 0, 0, 0, 0, -1, -3, -4, -2, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -3, -5, -6, -5, -3, -2, -1, 0, 1, 1, 2, 2, 0, 0, -1, -1, -3, -3, -2, -2, -2, -2, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -4, -4, -5, -4, -3, -2, 0, 0, 2, 1, 1, 2, 0, -1, -1, -1, -2, -3, -1, -1, -2, -2, 0, 0, 0, 1, 0, -1, -2, -3, -2, -1, -3, -5, -6, -6, -4, -3, 0, 0, 2, 2, 1, 2, 0, -1, -2, -1, -3, -2, -1, -1, -2, 0, -2, -1, 0, 1, 0, -1, -1, -2, -1, -1, -4, -6, -7, -6, -4, -3, -1, 1, 2, 1, 0, 1, 0, -1, -1, -2, -2, -2, -1, -2, -3, -1, -1, -1, 0, 0, 0, 0, 0, -2, -2, -2, -4, -5, -7, -6, -3, -3, 0, 1, 2, 2, 0, 1, 0, 0, 0, -2, -2, -2, -4, -3, -2, -1, -2, 0, 0, 0, 0, -1, -1, -1, -2, -3, -3, -4, -4, -4, -3, -2, -1, 0, 2, 1, 0, 1, 0, 0, -1, -1, -2, -4, -3, -3, -2, -1, -2, 0, 0, 0, 0, -1, 0, 0, -1, -3, -4, -5, -4, -4, -3, -2, -1, 0, 2, 0, 0, 0, 0, 0, -1, -2, -2, -5, -3, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -4, -4, -4, -4, -2, -1, 0, 2, 0, 0, 0, 0, -2, -2, -2, -2, -5, -5, -3, -2, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -3, -3, -4, -3, -4, -4, -3, 0, 0, 0, 0, 0, 0, 0, -3, -2, -3, -4, -3, -4, -2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -3, -2, -5, -3, -3, -3, -1, -1, 1, 0, 0, 0, -1, -2, -3, -2, -2, -3, -4, -3, -1, -1, 0, 1, 1, 0, 0, 2, 2, 2, 1, -1, -1, -2, -3, -4, -3, -2, -2, -1, 1, 1, 0, -1, 0, -1, -3, -2, -4, -4, -2, -1, -1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, -1, -1, -2, -2, -3, -1, 0, 0, 1, 0, 0, 0, 0, -2, -2, -3, -4, -4, -3, -2, -1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, -2, -1, -1, -3, -1, 0, 0, 0, 0, 0, -1, 0, -2, -2, -2, -4, -4, -3, -2, -1, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -2, -3, -1, -1, 0, 1, 1, 0, 0, -1, -2, -3, -5, -4, -3, -2, -3, -2, -3, -2, 0, 0, 2, 0, 1, 0, 0, 0, 1, 0, -1, 0, -2, -1, 0, 0, 0, 1, 1, 0, 0, -1, -3, -3, -4, -3, -4, -2, -2, -3, -1, -2, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 0, 1, 2, 2, 0, -1, -2, -4, -4, -4, -3, -2, -3, -4, -3, -1, 0, 0, 2, 2, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 3, 2, 0, 2, 1, 0, 0, 0, -1, -2, -3, -4, -4, -2, -3, -1, -2, -1, 0, 1, 4, 2, 0, -1, 0, 0, 1, 1, 1, 0, 0, 2, 2, 1, 2, 0, 1, 0, 0, -1, -1, -2, -2, -2, -1, -2, -1, -1, -1, 0, 1, 1, 3, 2, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 2, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 2, 1, 3, 1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 1, 0, 0, 0, 1, 1, 2, 1, 2, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 2, 1, 1, 0, 1, 0, 1, 3, 4, 5, 5, 4, 1, 1, 0, 0, 0, 1, 0, -1, -2, -2, -1, -1, -2, -1, -1, 0, 0, 1, 1, 1, 3, 2, 1, 0, -1, 0, 1, 2, 4, 5, 5, 5, 5, 3, 1, 0, 0, 1, 2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 2, 3, 2, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 1, 0, -1, -1, -3, -3, -3, -3, -4, -3, -2, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, -4, -3, -4, -2, -1, -2, -3, -1, -1, -3, -2, -3, -3, -2, -3, -3, -2, -2, 0, 2, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, -5, -5, -4, -5, -5, -4, -3, -1, -2, -2, -3, -3, -2, -2, -3, -2, -2, -1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -3, -3, -5, -5, -5, -4, -5, -2, -2, -1, 1, 0, 0, 0, -2, -1, -1, -1, -1, 0, 1, 1, 1, 1, 0, 0, -1, -1, -1, -2, -2, -3, -5, -6, -5, -5, -6, -6, -4, 0, 1, 0, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 3, 1, 0, 0, 0, -1, -1, -2, -4, -3, -4, -5, -6, -5, -3, -4, -5, -4, -1, -1, 0, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 1, 4, 4, 2, 2, 1, 0, 0, -3, -5, -4, -5, -5, -4, -4, -4, -4, -4, -5, -4, -2, -3, -1, -1, -2, 0, 0, -1, -1, -3, -1, 0, 0, 3, 2, 3, 1, 0, 0, -2, -4, -4, -7, -8, -8, -8, -6, -4, -4, -5, -4, -5, -4, -1, -1, -1, -1, 0, 0, -1, -2, -3, -2, 0, 0, 2, 1, 2, 0, 0, 0, -2, -4, -4, -5, -8, -7, -6, -7, -7, -7, -5, -4, -4, -2, 0, 1, 0, 1, 1, 1, -1, -3, -2, -2, -1, 0, 2, 2, 2, 1, -1, -1, -4, -5, -7, -8, -7, -6, -8, -7, -6, -6, -6, -3, -2, 0, 0, 1, 2, 1, 1, 1, -1, -2, -2, -1, 0, 0, 0, 1, 0, 0, -1, -1, -2, -4, -5, -6, -6, -4, -3, -4, -3, -3, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, -2, -3, -2, 0, 0, 2, 0, -1, 0, -1, -1, -3, -5, -6, -7, -7, -7, -3, -2, 0, -1, -4, -3, -1, -2, 0, 0, 0, 1, 0, 2, 0, -1, -2, -3, 0, 1, 1, 0, -1, 0, -1, -2, -3, -5, -7, -8, -8, -8, -7, -4, -2, -2, -2, -2, -1, 0, 0, 0, 0, 1, 1, 2, 1, 0, -1, -2, -1, 1, 2, 1, 0, -1, 0, -2, -3, -5, -6, -7, -6, -7, -7, -6, -5, -3, -4, -4, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, -2, -4, -1, 0, 1, 0, 0, 0, -1, -3, -4, -5, -5, -5, -5, -5, -5, -6, -6, -4, -2, -1, 0, 0, 2, 3, 2, 0, 0, 0, 0, -1, -4, -4, -2, 0, 1, 1, 0, -1, -1, -2, -3, -5, -6, -5, -7, -6, -7, -6, -5, -4, -1, 0, 2, 3, 2, 2, 2, 0, 0, -1, -2, -2, -4, -3, -2, 0, 1, 1, 0, 0, 0, 0, -1, -2, -2, -4, -5, -6, -6, -6, -3, -2, -2, 0, 2, 3, 1, 2, 0, -1, -3, -2, -1, -3, -3, -4, -1, 0, 1, 0, 0, 0, -1, 0, -2, -1, 0, -1, -3, -4, -5, -5, -5, -4, -3, -1, 0, 1, 1, 2, 0, -1, -3, -1, -2, -2, -4, -2, -1, 0, 2, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, -2, -4, -3, -2, -3, -2, -2, -2, -2, 0, 0, 0, -1, -2, -2, -3, -2, -3, -2, 0, 0, 4, 2, 0, 0, 0, 0, 0, -2, -1, -1, -2, -3, -2, -1, -2, -1, -2, -2, -1, -1, -2, -2, -2, -3, -2, -2, -2, -3, -2, -1, 0, 1, 3, 3, 2, 3, 1, 1, 1, 0, -1, -1, -2, -4, -4, -4, -4, -3, -1, 0, 1, 0, -1, -2, -2, -1, -3, -3, -2, -4, -4, -1, -1, 1, 4, 2, 2, 1, 0, 0, -1, 0, 0, 0, -2, -3, -2, -1, -2, -2, -2, 0, 1, 1, 0, -1, 0, 0, 0, -1, -3, -3, -4, -2, -1, 1, 4, 2, 0, 0, -1, 0, -1, -2, 0, -2, -1, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 3, 3, 1, -1, -2, -1, -2, -2, -1, -2, 0, 1, 1, 1, 1, 2, 1, 1, 3, 2, 1, 1, 0, -1, 0, 0, 0, -1, -2, -1, -1, 0, 2, 2, 0, 1, 0, -2, -2, -1, 0, 0, 0, 1, 3, 4, 4, 5, 4, 3, 1, 2, 1, 0, 0, -2, -2, -1, -2, -3, -2, -2, 0, 1, 4, 4, 2, 1, 0, 0, 0, 0, 0, 0, 0, 2, 3, 4, 4, 5, 4, 3, 0, -1, -1, -2, -3, -3, -3, -2, -2, -3, -3, -1, 0, 2, 1, 3, 3, 2, 1, 1, 1, 1, 0, 1, 1, 0, 0, 1, 0, -1, -1, -2, -4, -5, -4, -5, -4, -4, -6, -5, -4, -3, 0, 2, 1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, -2, -2, -2, -2, -2, 0, -1, -1, 0, -1, -1, -1, -2, -1, 0, 2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 1, 1, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, -1, 0, 0, 0, 0, -1, 0, -1, 0, -2, -1, -1, -1, 0, 0, 0, 1, 2, 1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, -1, -1, -2, 0, -1, -2, -1, -1, 0, -1, -1, -2, -2, -3, -2, -2, 0, 0, 0, 1, 0, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -1, -1, -1, 0, -1, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, -2, -2, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -2, -1, -2, -1, 0, -1, 0, 0, 2, 2, 1, 1, 1, 0, 0, 0, 0, -2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -2, -1, -2, -2, -2, -1, -1, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, -2, -2, -1, 0, -1, 0, 0, 2, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -2, -1, -1, -1, -1, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -1, -1, -1, -2, -2, -2, -2, 0, -1, 0, 0, 1, 2, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, -3, -2, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, 0, -2, -1, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, -2, -3, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -3, -2, 0, 0, -1, -1, 0, 1, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, -2, -2, -2, -1, -1, -1, 0, 1, 0, 1, 2, 2, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -2, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, -1, -2, -1, -2, -3, -3, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, -2, -2, -1, -1, -3, -2, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -2, -1, -1, -2, -2, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, -1, -2, -2, -2, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -2, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -2, -1, -2, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 0, -1, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, -1, 0, -1, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -2, -2, -2, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, -1, -2, -2, -1, -1, -1, -1, -3, -3, -2, -2, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -2, -2, -1, -1, -1, -3, -2, -2, -2, -1, -2, 1, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -2, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 2, 1, 1, 0, 1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, -2, -1, -1, -2, 0, -3, -3, -1, -2, -2, -1, 0, 0, -1, 0, 1, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -2, -2, -2, -1, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, -1, -1, -2, -2, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, -2, -3, -3, -2, -2, -1, -1, 0, 0, 1, 0, 1, 0, 0, -1, -1, -1, -1, -2, -1, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -3, -4, -4, -3, -2, 0, -1, 0, 0, 0, 0, 0, 0, -2, 0, -1, -3, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -3, -4, -4, -3, -5, -3, -2, 0, -1, 0, 0, 0, 0, 0, -1, 0, -2, 0, -1, -2, 0, -1, -2, 0, 0, -1, 0, 2, 0, 0, -1, 0, -3, -4, -4, -5, -5, -2, -3, -2, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -2, -2, -4, -6, -5, -5, -3, -1, -1, -1, 0, 1, 0, 1, 1, 1, 0, -1, -2, -1, -1, -2, -2, -2, 0, 0, 0, 1, 0, -1, 0, -1, -2, -3, -4, -6, -6, -5, -3, -2, 0, 0, 2, 0, 0, 1, 0, 0, 0, -1, -2, -3, -2, -2, -1, 0, -1, 0, -1, 0, 1, 0, 0, -2, -1, -3, -4, -6, -5, -5, -4, -3, -1, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, -3, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, -5, -6, -6, -5, -4, -2, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, -2, -3, -1, -2, -2, 0, 0, 0, 0, 0, 1, 0, 1, -1, -1, -3, -3, -4, -5, -4, -4, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -2, -2, -2, -1, -1, -2, 0, 0, 0, 0, 1, 1, 1, 0, -1, -3, -4, -4, -4, -3, -3, -2, 0, 0, 1, 0, 0, 1, 0, 0, 1, -1, -2, -3, -2, -2, -2, -1, -1, 0, 0, 1, 1, 1, 1, 0, -1, -2, -2, -2, -4, -3, -2, -2, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, -1, -1, -2, -2, -2, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, -1, -1, -1, -2, -2, -1, 0, 1, 1, 0, -1, 0, 0, -1, -1, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -1, -2, -1, -1, -1, 0, 0, 1, 2, 0, 0, -1, 0, -2, -2, -1, -1, 0, -1, 0, -1, 0, -1, 0, 0, 1, 0, 2, 1, 1, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -2, -2, -1, -2, -3, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, -2, -2, -3, -2, -3, -1, 0, -1, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, -2, 0, -2, -2, -2, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -3, -1, 0, -2, 0, -2, 0, -1, 0, 1, 0, 0, 1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, -1, -2, -2, -1, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 2, 2, 1, 1, 0, -1, -2, -1, -1, -2, 0, -1, -2, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 2, 2, 1, 2, 2, 2, 1, 2, 2, 1, 1, 0, -1, -1, -1, -1, 0, -2, -2, -2, -1, -2, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 2, 3, 3, 2, 2, 2, 1, 1, 1, 1, 1, 0, 0, -1, -1, -2, -1, -1, -2, -2, -1, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 1, 1, 2, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 2, 0, 2, 2, 1, 0, 0, 0, 0, 1, 0, 0, 1, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0, -3, -2, 0, -2, 0, 1, 0, 0, 0, 1, 3, 3, 1, 0, 1, 1, 1, 1, 1, 2, 2, 1, 3, 3, 3, 3, 2, 1, 3, 2, 0, 0, -1, 0, 0, 0, 0, 2, 2, 2, 3, 2, 3, 2, 1, 1, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 0, 0, -1, -1, 0, -1, 0, 2, 3, 2, 0, 2, 1, 2, 1, 0, 1, 1, 0, -1, 0, -1, -2, -1, 0, -1, -1, 0, 0, 1, 2, 2, 1, 0, -1, 0, 0, 0, 0, 0, 2, 1, 1, 2, 2, 0, 1, 1, 2, 0, -1, -3, -2, -2, -1, -2, -2, 0, 0, 0, 0, 0, 1, 3, 1, 0, -1, 0, 0, -1, 0, 1, 1, 1, 1, 1, 0, 1, 2, 2, 2, 0, -1, -3, -2, -3, -2, -1, 0, 0, 0, 0, 0, 1, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 3, 2, 2, 2, 0, -3, -3, -2, -1, 0, 0, 1, 2, 1, 0, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 3, 2, 3, 2, 0, -1, -3, -2, -2, 0, 0, 1, 2, 1, 0, 1, 2, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 1, 2, 2, 3, 3, 3, 1, -1, -2, -2, -2, -1, -1, 0, 2, 1, 1, 1, 0, 3, 2, 0, 0, 2, 1, 0, 0, 0, -1, 0, -2, -1, 0, 1, 2, 3, 4, 3, 0, -1, -3, -3, -1, -1, 0, 0, 0, 3, 1, 0, 0, 2, 1, 0, 0, 2, 1, 0, 0, 1, 0, 0, -2, -1, 0, 0, 0, 3, 3, 3, 0, 0, 0, -1, -2, 0, 0, 0, 1, 1, 1, 0, 0, 2, 0, 0, 0, 1, 0, 1, 2, 1, 0, 0, -2, -2, 0, 0, 2, 2, 2, 2, 2, 1, 0, -1, -1, 0, -2, -1, 1, 1, 0, 0, 0, 1, 2, 0, 0, 1, 0, 1, 1, 2, 1, -1, -2, -1, 0, 0, 2, 2, 3, 2, 2, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, -2, -2, 0, 0, 2, 2, 4, 3, 2, 1, 1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -2, -1, 0, 0, 0, 1, -1, -2, -3, 0, 0, 2, 3, 4, 3, 1, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, -1, 0, 2, 0, 0, -1, -1, 1, 0, 0, 0, 0, -2, -3, -3, -2, 0, 1, 2, 2, 3, 1, 0, 0, -1, -2, 0, -1, 0, 0, 0, -1, 0, 0, 2, 1, 0, -2, -1, 0, 0, 0, 0, 0, -3, -2, -2, -1, 0, 1, 3, 2, 3, 0, 1, 0, -1, -1, -1, -1, -2, -1, -1, -1, 0, 1, 1, 2, 0, -1, -2, 0, 1, 0, 0, -1, -3, -3, -1, -2, 0, 0, 2, 2, 3, 2, 0, 0, -1, 0, 0, 0, -2, -1, -1, 0, 0, 0, 1, 1, 0, -1, -1, 0, 0, 0, 0, -2, -2, -2, -1, -2, 0, 0, 3, 3, 4, 1, 0, 0, 0, 0, 0, 0, -2, -2, -2, -1, 1, 2, 3, 1, 0, -1, -1, 0, 0, 0, 0, -1, -1, -2, -2, -3, 0, 0, 3, 5, 4, 1, 0, 1, -1, -1, 0, -2, -2, 0, 0, 0, 0, 2, 3, 2, 0, -2, 0, 0, 0, 0, -1, -2, -2, -1, -3, -3, -2, 0, 2, 4, 4, 1, 1, 0, -1, -1, -2, -1, -2, 0, 0, 1, 1, 2, 3, 2, 0, -1, 0, 0, 1, 0, 0, -1, -1, -2, -2, -2, 0, 2, 3, 3, 3, 0, 1, 0, -2, -2, -2, -1, -1, 0, 1, 2, 2, 3, 4, 2, 1, 0, 0, 1, 1, 1, -1, -2, -2, -2, -2, -1, 0, 2, 1, 3, 3, 2, 1, -1, -1, -3, -3, -3, 0, 2, 2, 1, 2, 3, 3, 1, 0, 0, 0, 2, 1, 0, 0, -1, -3, -3, -1, 0, 0, 1, 2, 2, 2, 1, 0, 0, -3, -3, -3, 0, 0, 2, 2, 2, 2, 3, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 1, 1, 1, 2, 1, 0, -2, -2, -3, -2, -1, 1, 1, 3, 1, 2, 2, 2, 2, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, 0, 1, 1, 2, 1, 1, 0, -1, -2, -4, -3, -3, -1, 0, 0, 1, 2, 2, 2, 3, 2, 2, 0, -1, -1, 0, -1, -1, -1, -1, 0, -1, 1, 1, 1, 0, 0, 0, 0, -1, -4, -5, -5, -2, -1, 0, 0, 0, 1, 1, 3, 4, 4, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, -5, -5, -5, -3, 0, 0, 0, 0, 0, 0, 2, 3, 3, 2, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, -2, -5, -4, -4, -2, 0, 0, 0, 0, 0, 1, 3, 4, 5, 1, 0, -2, -1, 0, 0, 0, 0, 1, 2, 2, 2, 0, 0, 0, 0, -1, 0, -1, -3, -3, -1, 0, 0, 2, 2, 1, 0, 2, 4, 3, 4, 0, 0, -2, -2, 0, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 3, 2, 3, 1, 2, 3, 3, 2, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 1, 1, 2, 2, 0, 1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -3, 0, -1, -2, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, -2, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -2, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, -2, -1, 0, -2, -2, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, -2, -1, 0, -1, -1, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 1, 0, -1, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 1, 2, 2, 1, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 2, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 2, 1, 0, 1, 1, 1, -1, -1, 0, 0, -2, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 2, 2, 0, 2, 0, 1, 0, 0, -1, -1, 0, -2, 0, 0, 0, -1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 2, 1, 0, 0, 1, 2, 2, 3, 1, 2, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, -2, 0, 0, 0, 1, 2, 1, 0, 1, 1, 2, 2, 2, 1, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 2, 0, -2, -1, 0, 0, 0, 2, 0, 1, 2, 2, 2, 2, 2, 2, 1, 1, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, -2, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 2, 0, 0, 0, 1, 1, 3, 3, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 2, 2, 1, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 1, -2, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 2, 2, 2, 1, 1, 1, -1, 0, 0, 0, -1, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, -3, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 2, 2, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -2, 0, -1, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 2, 1, 0, 2, 2, 1, 1, 1, 1, 1, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 1, 1, 1, 0, 0, 0, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 0, 0, 0, 0, -1, -1, -2, -1, 0, -1, 0, -1, -1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 1, 1, 0, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 0, 0, -2, 0, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 1, 0, 1, 1, 0, 0, -1, 0, -2, -1, 0, 0, 0, 0, -1, 1, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, -1, 0, 1, 1, 0, 0, -1, -2, -2, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, 0, 1, 1, 1, 1, 0, 0, -2, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, -3, 0, -1, -1, -1, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, -1, 0, -3, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, -1, -1, -1, -2, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 0, 0, 0, 2, 0, -1, 0, -2, -2, -2, -2, -2, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 3, 1, 3, 4, 1, 1, 2, 2, 1, 2, 0, 0, -1, -3, -2, -3, -2, -1, -1, -2, -2, 0, 0, -1, 0, 0, -1, 0, 0, 1, 2, 2, 4, 3, 3, 3, 1, 3, 3, 1, 2, 4, 2, 2, 0, -2, -2, -2, -1, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, -1, 0, 0, 2, 2, 3, 3, 5, 2, 2, 3, 4, 2, 2, 4, 2, 3, 2, -1, -1, 0, -1, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 2, 4, 3, 3, 3, 2, 4, 4, 3, 1, 2, 3, 3, 2, 0, 1, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 1, 0, -1, 0, 2, 1, 2, 3, 2, 2, 3, 3, 3, 4, 3, 2, 2, 1, 3, 3, 1, 1, 2, 1, 1, 0, -1, 0, 0, -2, 1, 0, 1, 0, 0, 0, 2, 1, 2, 2, 2, 1, 2, 2, 4, 2, 1, 3, 1, 1, 4, 2, 1, 1, 2, 2, 2, 0, 0, 0, 0, -3, 0, 2, 1, 0, -1, 1, 1, 1, 3, 2, 1, 2, 1, 2, 4, 2, 0, 1, 2, 0, 2, 3, 0, 1, 1, 2, 1, 0, -1, 0, 0, -3, 0, 2, 1, 0, 0, 1, 3, 2, 3, 3, 2, 2, 2, 3, 3, 3, 0, 2, 3, 2, 2, 2, 0, 1, 3, 1, 0, 1, 0, 0, 0, -3, -1, 0, 1, 0, 2, 1, 3, 3, 5, 2, 2, 2, 1, 3, 4, 2, 0, 0, 0, 2, 1, 1, 0, 0, 2, 1, 1, 0, -2, 0, 0, -1, 0, 2, 1, 1, 1, 2, 2, 3, 3, 3, 2, 4, 3, 2, 4, 0, 0, 0, -1, 1, 0, 0, 0, 1, 2, 3, 1, 1, -3, 0, 0, -1, 0, 1, 0, 0, 3, 1, 2, 3, 3, 5, 4, 4, 4, 4, 3, 0, -1, -1, -1, 0, 0, 2, 0, 1, 3, 3, 1, 0, -3, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 3, 4, 4, 4, 4, 4, 4, 4, 0, 0, 0, 0, -1, 0, 1, 0, 0, 4, 3, 1, 0, -3, 0, 0, 1, 0, 0, -1, 0, 1, 2, 3, 3, 3, 4, 3, 2, 4, 5, 4, 1, 0, 0, 0, -2, -1, 1, 0, 1, 3, 3, 2, 1, -2, -1, 0, 1, 0, 0, 0, -1, 0, 1, 3, 3, 3, 4, 5, 3, 4, 4, 4, 2, 1, 2, 1, -1, 0, 0, 0, 1, 2, 2, 1, 1, -2, -2, 0, 1, 0, -1, 0, 0, 0, 2, 4, 3, 5, 3, 4, 4, 2, 1, 1, 2, 1, 2, 1, 0, -1, 0, 0, 0, 1, 2, 1, 0, -4, -3, 0, 0, -1, 0, 0, 0, 1, 1, 4, 4, 4, 3, 3, 3, 2, 1, 1, 1, 0, 1, 1, -1, 0, 0, 0, 0, 2, 2, 0, -1, -3, -2, 0, 0, -1, 0, 0, 2, 1, 1, 4, 5, 4, 2, 3, 2, 3, 0, 2, 1, 1, 2, 0, 0, 1, 0, 0, 1, 2, 1, 0, 0, -3, -2, 0, 1, -2, 0, 1, 2, 1, 0, 3, 4, 4, 2, 3, 3, 1, 0, 2, 2, 0, 1, 2, 0, 0, 0, 0, 0, 2, 1, 1, 0, -3, -1, 0, 0, -1, 0, 0, 0, 0, 0, 2, 4, 4, 3, 3, 3, 2, 0, 2, 1, 0, 1, 1, 0, 2, 0, 0, 1, 1, 1, 0, 0, -1, -1, 0, -1, -2, 0, 1, 1, 0, 0, 2, 2, 2, 1, 0, 4, 1, 1, 3, 2, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, 2, 1, 0, 1, 3, 2, 2, 2, 0, 3, 2, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, -2, -1, 0, 0, 0, 0, 1, 1, 0, 0, 2, 2, 3, 1, 0, 2, 3, 0, 1, 0, 0, 0, 0, 2, 1, 0, -1, 1, 0, -1, 0, 0, -2, -2, 0, -1, 0, 0, 2, 1, 0, 0, 1, 2, 0, 0, 1, 2, 3, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -2, 0, 0, 0, 2, 1, 0, 0, -2, 0, 0, 0, 1, 1, 3, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, 0, -1, 0, -2, -2, 0, 0, 0, 1, 1, 1, 0, -2, -1, 0, 0, 1, 1, 3, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 2, 2, 3, 4, 3, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, -2, 0, 3, 3, 4, 3, 1, 1, 2, 2, 2, 2, 1, 0, 0, 0, -1, -2, -1, -1, -2, 0, -2, 0, 0, -1, 0, 0, 0, 2, 0, 0, 0, 0, 2, 2, 3, 2, 1, 2, 1, 2, 0, 1, 1, 0, -1, -1, 0, -1, 0, -1, -1, 0, -3, 0, -1, -1, 0, 0, 1, 0, 1, 0, -1, 0, 1, 1, 1, 0, 0, 1, 1, 0, 1, 1, 0, -1, 0, 0, -1, -1, 0, -1, -2, 0, -2, 0, -2, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, 0, -3, -1, -2, -2, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 2, 3, 4, 4, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -2, -2, -1, -1, 0, -1, -1, -2, -1, -1, 0, 0, 1, 2, 2, 2, 3, 2, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, -2, -2, -1, 0, 0, 0, 1, 1, 1, 2, 1, 1, 0, 0, 2, 0, 0, 0, 1, 3, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, -2, 0, -1, 0, 0, 1, 0, 1, 2, 0, 2, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, -2, -2, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, -1, -1, -1, -3, -2, -1, -1, 0, 0, 1, 0, 0, 0, -2, -2, -1, 0, 0, 0, 1, 1, 0, 1, 1, 3, 2, 1, 2, 2, 2, 0, 0, 0, -1, -1, -2, -2, -2, 0, 0, 0, 0, 0, 1, 0, -1, -2, -1, 0, 0, -1, 0, 1, 0, 1, 1, 1, 2, 0, 2, 4, 4, 1, 1, 0, 0, -2, -2, -4, -3, -1, 0, 0, 1, 0, 0, -1, -1, -2, -3, -1, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 2, 3, 2, 1, 0, 0, 0, -2, -3, -4, -5, -3, -1, 0, 0, 0, 0, 0, 0, -1, -3, -2, -2, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 3, 0, 0, 0, 0, 0, -1, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 0, 0, 0, 0, -1, -1, -2, -2, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -3, -3, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, -1, -1, -1, -1, -2, -4, -2, -1, 0, 1, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -2, -2, -2, -2, -2, -2, -1, -1, 0, 1, 2, 1, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, -1, -2, -1, -2, -1, -4, -4, -2, -2, -3, -1, -1, 0, 1, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -2, -2, -3, -2, -3, -2, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, -1, 0, -1, -1, 0, 0, 1, 1, -1, -1, 0, 0, 0, 0, -1, -2, -2, -2, -3, -3, -2, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -2, -3, -2, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 1, 1, 0, 1, 0, 0, 1, 0, -1, -2, -2, -1, -2, -2, -1, -1, -1, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 1, 1, 0, -1, -2, -1, -2, -2, -1, -1, 0, 0, -1, 0, -2, -2, -1, -1, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 0, 1, 0, -1, -3, -2, -2, -2, -2, -1, -1, 0, -1, 0, 0, -1, 0, -2, -1, -2, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 2, 1, 0, 0, 0, -1, -3, -4, -3, -2, -2, -2, -2, -1, -2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 1, 0, -1, 0, -1, -2, -2, -3, -2, -2, -1, -1, -1, -2, -1, 0, 0, 0, -2, -2, 0, -1, 0, 1, 2, 0, 1, 0, 2, 0, 1, 0, 0, 0, 0, -2, -2, -3, -2, -3, -1, 0, 0, -2, -1, -1, 0, -1, -1, -3, -3, -2, -2, 0, 0, 0, 2, 2, 2, 2, 1, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -2, -3, -2, -3, -2, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, -1, -1, -3, -3, -4, -2, -1, -2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, -3, -3, -3, -2, -2, -1, -2, -1, -2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 0, 0, 0, 0, 0, 0, -1, -2, -2, -3, -2, -2, -1, -1, -2, -1, 0, 1, 2, 1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -2, -2, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 2, 1, 1, 1, 0, 0, 2, 1, 1, 0, 2, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 2, 2, 1, 1, 2, 1, 1, 2, 2, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 1, 1, 2, 2, 0, 1, 2, 1, 2, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, 0, 0, 1, 2, 1, 1, 2, 1, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 2, 1, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 1, 1, 2, 1, 1, 1, 1, 0, 0, 2, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 1, 0, 1, 0, 2, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -2, -1, 0, 0, 0, 1, 3, 1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 1, 0, -1, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 1, 2, 2, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 1, 0, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -2, 0, -2, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 0, 2, 2, 0, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 3, 1, 2, 1, 1, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, -2, 0, 0, -1, -1, -1, 0, 1, 2, 2, 1, 2, 3, 3, 2, 2, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 2, 1, 2, 2, 3, 2, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 2, 3, 2, 2, 3, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 0, 2, 2, 2, 1, 1, 1, 3, 3, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 2, 1, 1, 2, 2, 2, 1, 2, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 1, 1, 2, 3, 2, 2, 2, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 3, 2, 2, 0, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, 1, 2, 1, 3, 2, 2, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 3, 1, 1, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, -2, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -2, 0, 1, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 2, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 2, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -1, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, -1, -2, -1, -1, -2, -2, 0, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 2, 2, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, -3, -2, 0, 0, 0, 0, 1, 0, 1, 2, 2, 1, 1, 0, 1, 1, 0, 0, 1, 1, 2, 3, 4, 5, 5, 5, 5, 4, 3, 1, 0, 0, 0, 0, 0, 1, 2, 2, 2, 3, 4, 3, 2, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 3, 4, 3, 3, 1, 1, 0, 0, 1, 0, 1, 2, 3, 3, 3, 3, 2, 1, 0, -1, -1, 0, -1, 0, -1, -2, 0, -1, -1, -1, 0, 0, 1, 2, 3, 3, 1, 0, 0, 0, 2, 2, 1, 2, 3, 3, 1, 1, 0, 0, 0, -1, -1, 0, -1, -2, -2, -4, -2, -2, -3, -2, 0, 0, 1, 2, 3, 4, 1, 0, 1, 2, 0, 1, 0, 2, 1, 3, 2, 1, 1, 0, 1, 0, 0, 0, 0, -4, -5, -5, -3, -2, -2, -3, -1, 0, 0, 1, 2, 3, 2, 0, 0, 1, 1, 0, -1, 0, 1, 1, 1, 1, 0, 1, 2, 2, 0, 0, 0, -1, -2, -3, -4, -1, -1, 0, 0, 1, 0, 2, 4, 4, 2, 1, 1, 1, 0, 0, 0, -1, 0, -1, -1, -2, 0, 2, 2, 1, 2, 1, 1, -1, -3, -1, -3, -1, -1, -1, 0, 1, 1, 0, 2, 3, 2, 0, 2, 2, 2, 1, 0, -1, 0, -3, -3, -2, 0, 1, 2, 3, 3, 3, 2, -1, -3, -4, -2, -3, -2, -1, 0, 1, 0, 0, 1, 3, 2, 1, 2, 4, 3, 3, 0, 0, -2, -3, -4, -4, -2, 0, 2, 4, 3, 4, 1, -1, -3, -3, -4, -5, -2, -3, -1, 0, 0, 0, 1, 1, 0, 2, 2, 4, 2, 3, 1, 0, -2, -2, -4, -4, -4, 0, 0, 1, 3, 4, 1, 0, -1, -2, -4, -3, -4, -2, -1, 0, 0, -1, 0, 1, 1, 2, 2, 2, 3, 1, 1, 0, -2, -3, -4, -4, -3, -1, 0, 2, 2, 2, 1, 1, 0, -1, -2, -2, -3, -3, 0, -1, 0, -1, 0, 1, 2, 1, 2, 3, 1, 1, 0, 0, -1, -3, -4, -5, -3, -1, 0, 0, 1, 2, 2, 2, 1, 0, -1, -2, -3, -1, -1, -1, 0, -2, -1, 0, 2, 1, 1, 1, 0, 0, -1, -2, -1, -3, -6, -5, -3, 0, 0, 3, 3, 5, 3, 3, 2, 0, -1, 0, -2, -1, -3, -1, -1, -2, 0, 0, 1, 0, 0, 0, 0, -1, -2, -1, -2, -4, -6, -5, -3, 0, 2, 4, 5, 5, 4, 3, 1, 0, -2, -1, -2, -2, -2, -2, -1, -2, 0, 1, 0, 0, 0, 0, -2, -3, -3, -2, -2, -5, -5, -6, -4, 0, 0, 2, 3, 6, 3, 3, 1, 0, -2, -1, -3, -3, -2, -2, -2, -1, 0, 0, 0, 0, 0, -1, 0, -2, -1, -2, -4, -7, -7, -5, -3, -1, 0, 1, 3, 3, 3, 1, 0, 0, -3, -3, -2, -2, -2, -3, -1, -1, 0, 1, 0, 1, 0, -2, -1, -1, -2, -3, -5, -7, -6, -5, -5, -2, 1, 2, 2, 4, 3, 1, 0, 0, -2, -3, -2, -3, -3, -3, -2, -3, 0, 1, 0, 0, 0, -1, 0, -1, -1, -3, -4, -5, -5, -5, -4, -2, 0, 3, 4, 4, 2, 0, 1, 0, -2, -2, -2, -3, -5, -2, -3, -3, 0, 1, 0, 0, 0, 0, -1, 0, -1, -2, -5, -6, -5, -5, -4, -1, 0, 2, 4, 4, 2, 0, 1, 0, -2, -2, -3, -3, -5, -4, -3, -2, 0, 1, 2, 0, 0, 0, 0, 0, 0, -2, -3, -4, -4, -4, -5, -3, 0, 0, 1, 3, 1, 0, -1, -2, -3, -2, -3, -5, -5, -3, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, -1, -3, -5, -6, -5, -4, -2, 0, 0, 1, 2, 0, -1, 0, -1, -3, -3, -5, -4, -3, -1, 0, 0, 0, 2, 2, 2, 1, 2, 2, 1, 0, -1, -3, -6, -4, -5, -4, -3, 0, 2, 2, 2, 1, 0, 0, -3, -3, -3, -5, -3, -3, 0, 1, 1, 2, 2, 2, 2, 2, 3, 3, 1, 0, -1, -3, -4, -5, -3, -3, 0, 0, 1, 1, 1, 0, 0, 0, -3, -3, -5, -3, -3, -1, 0, 1, 2, 2, 3, 1, 0, 2, 3, 2, 1, 0, -1, -4, -4, -3, -4, -1, 0, 1, 0, 1, 0, -1, 0, -2, -4, -3, -3, -3, -3, -1, 0, 2, 2, 3, 3, 1, 0, 1, 2, 0, 0, -2, -3, -4, -3, -4, -2, 0, 0, 1, 1, 1, 0, 0, -2, -4, -4, -4, -5, -4, -3, 0, 0, 2, 2, 2, 4, 1, 0, 0, 1, 0, 0, -2, -2, -2, -2, -2, 0, 0, 2, 1, 2, 0, 0, -2, -4, -5, -6, -6, -5, -3, -2, -2, 0, 0, 1, 3, 3, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 1, 0, -1, -2, -5, -5, -7, -7, -5, -4, -3, -1, -1, 0, 0, 3, 3, 2, 0, 1, 1, 1, 1, 1, 0, 0, 1, 0, 2, 2, 2, 2, 1, -1, 0, -1, -5, -7, -7, -7, -5, -4, -3, -2, -1, -1, 0, 3, 4, 1, 1, 0, 0, 0, 1, 0, 1, 2, 2, 2, 2, 3, 1, 0, 0, -1, -1, -2, -3, -5, -5, -5, -3, -2, 0, -1, -1, 0, 1, 4, 4, 2, 0, -1, -1, 0, 0, 0, 0, 1, 2, 2, 2, 2, 1, 0, 0, -2, -2, -2, -2, -1, -1, -1, 1, 0, 1, 1, 2, 3, 4, 4, 4, 1, 0, -2, 0, 0, 0, 0, 0, 1, 3, 3, 3, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 3, 2, 3, 3, 3, 3, 4, 3, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -3, -2, -2, -1, -2, -1, -2, -3, -2, -2, -2, -4, -3, -4, -2, -2, -3, -3, -2, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, -2, -1, -1, -1, -2, -3, -2, -4, -3, -4, -2, -1, -3, -1, -2, -2, -3, -3, -2, -2, -2, -1, 0, 0, 0, -2, 0, -1, 0, -2, -3, -3, -1, -2, -1, 0, 0, -2, 0, -2, -4, -3, -2, -1, 0, -1, -1, 0, -3, -2, -2, -2, -2, -1, 0, 0, -2, -2, 0, -1, -1, -1, -2, -3, -3, -1, 0, 0, 0, 0, 0, -1, -3, 0, -1, 0, 1, 1, 1, 0, -1, 0, -2, -2, -2, -2, -1, 0, -1, -1, 0, -1, -2, -1, -1, -3, -2, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 3, 2, 1, 0, 0, -1, -2, 0, 0, 0, 0, -2, 0, 0, -2, -1, 0, -1, 0, -1, 0, 0, 2, 1, 1, 0, 0, 0, 1, 0, 0, 1, 2, 3, 2, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, -1, 0, 1, 2, 1, 2, 1, 0, 2, 2, 0, 1, 1, 2, 3, 2, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 2, 1, 1, 2, 0, 1, 0, 1, 0, 1, 1, 3, 2, 0, 0, 0, -1, -1, 0, 0, 0, -2, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 2, 2, 2, 1, 2, 3, 1, 0, 1, 0, 2, 2, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 2, 1, 2, 1, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, -2, -1, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 2, 2, 3, 3, 1, 1, 1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, -1, -2, -2, 0, -2, -1, 0, 0, 0, -1, 0, 0, 0, 2, 2, 3, 2, 3, 3, 1, 1, 0, 0, 0, 0, 2, 1, 1, 0, 1, 0, 0, -1, -2, -2, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 2, 3, 4, 5, 4, 3, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, -1, -2, -1, 0, 0, -1, -1, 0, 0, 0, 0, 2, 1, 3, 4, 4, 4, 5, 2, 0, -1, -1, -1, -2, 0, 0, 1, 1, 2, 0, 0, -2, -2, -1, -1, 0, 1, 0, -1, 0, 1, 1, 2, 2, 3, 2, 3, 3, 2, 4, 2, 0, -1, -1, 0, -2, -1, 0, 0, 0, 1, 1, 1, 0, -1, -2, -1, 0, 0, 0, -1, 0, 0, 2, 2, 3, 2, 4, 2, 3, 2, 3, 4, 0, 0, -1, 0, -1, -1, 0, 1, 0, 0, 1, 0, 0, -1, -2, 0, 0, 1, -1, -1, 1, 0, 2, 3, 3, 3, 3, 4, 3, 3, 3, 3, 1, 0, 0, 0, -1, 0, 1, 1, 1, 0, 1, 0, -1, -2, -2, -2, 0, 0, 0, 0, 0, 1, 3, 4, 3, 4, 2, 3, 2, 4, 3, 3, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, -1, -1, -3, 0, 0, 0, -2, 0, 0, 1, 1, 3, 2, 4, 1, 1, 2, 3, 3, 2, 1, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -2, -2, 0, 0, -1, -1, 0, 1, 2, 1, 2, 2, 3, 1, 1, 3, 3, 2, 3, 1, -1, 0, 1, 0, 0, 1, 0, 1, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 2, 1, 2, 2, 2, 2, 1, 3, 3, 2, 3, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, -2, 0, 2, 1, 1, 2, 2, 1, 1, 1, 1, 2, 2, 1, 1, -1, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 1, 1, 1, 2, 1, 1, 1, 1, 1, 3, 1, 1, 1, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 2, 2, 4, 3, 2, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 2, 2, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -1, -2, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 2, 4, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, -1, -2, -2, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 2, 2, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, -1, -2, -3, -3, -1, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 1, 0, 1, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, -2, -2, -3, -2, -1, 0, 0, -1, -1, 0, 0, -2, -1, 0, -3, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, -1, -2, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -2, -1, 0, 0, 0, -1, -2, -2, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -3, -2, -1, -2, 0, -1, 0, 0, 0, 1, 0, -1, -2, -4, -4, -4, -4, -4, -3, -3, -2, -1, 0, 0, 1, 1, 1, 0, 0, 0, -2, -1, -3, -4, -1, 0, 0, 0, 0, 1, 1, 2, 1, -2, -3, -5, -3, -5, -2, -1, -2, -2, -1, -1, 1, 0, 1, 0, 0, 2, 1, 0, -1, 0, -2, -3, -2, -1, 0, 0, 1, 2, 3, 3, 2, 0, -2, -1, -1, -1, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 2, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -2, -2, 0, 0, 0, 0, 1, 2, 3, 2, 2, 1, 3, 2, 1, 0, 1, 2, 0, 0, 1, 1, 0, -1, 0, 1, 2, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 3, 4, 3, 4, 2, 1, 0, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 2, 5, 4, 4, 5, 4, 3, 1, 1, 1, 2, 2, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 2, 2, 0, 0, -1, 0, 0, -2, -1, 0, 2, 4, 4, 5, 6, 4, 3, 3, 1, 2, 3, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 3, 1, 0, 0, 0, 0, -1, -1, 0, 3, 4, 3, 5, 5, 5, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 3, 1, 0, -1, 0, -1, -1, 0, 1, 2, 2, 5, 5, 4, 2, 2, 1, 1, 2, 2, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, -1, -1, 0, 0, 0, 3, 4, 5, 5, 6, 4, 3, 2, 2, 1, 1, 1, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 2, 2, 4, 6, 6, 4, 3, 3, 2, 2, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -2, 0, 0, 0, 1, 3, 3, 4, 5, 7, 7, 4, 3, 3, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 2, 3, 3, 4, 5, 5, 7, 6, 5, 4, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, -2, -3, -1, 0, 1, 2, 3, 3, 4, 5, 5, 7, 6, 4, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -2, -2, -2, 0, -1, 0, 1, 2, 4, 3, 5, 5, 6, 6, 5, 4, 3, 3, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -2, -1, -1, -1, -1, 0, 1, 2, 3, 3, 3, 5, 4, 6, 5, 3, 3, 2, 2, 0, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 1, 2, 2, 5, 4, 7, 6, 4, 3, 3, 3, 1, 1, 2, 0, 0, -1, -2, -1, 1, 2, 0, 0, 0, -2, -2, -1, 0, 0, -1, 0, 0, 1, 1, 3, 3, 5, 5, 5, 5, 3, 3, 3, 1, 1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 1, 1, 2, 2, 3, 4, 5, 3, 3, 3, 2, 2, 2, 0, 0, -1, -1, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, 0, 1, 1, 3, 4, 3, 4, 3, 1, 3, 2, 1, 2, 0, 0, 0, -1, -2, 0, 0, 1, 1, 0, 0, 1, 0, 1, 1, 1, 0, -1, -2, 0, 0, 2, 3, 4, 3, 1, 1, 1, 3, 1, 2, 2, 0, 0, -1, -1, -1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -2, -1, 1, 2, 4, 3, 2, 3, 2, 1, 3, 3, 1, 1, 1, 0, 0, -1, -1, 0, 2, 2, 1, 0, 0, 0, 1, 1, 1, 0, -1, 0, -1, 0, 0, 3, 4, 3, 2, 3, 3, 2, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 2, 3, 4, 3, 2, 4, 3, 2, 1, 0, 0, 0, -1, -1, -1, -2, -1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, -2, -2, -1, 0, 1, 2, 3, 2, 3, 2, 3, 2, 1, -1, 0, -1, 0, -2, -2, -1, -2, -1, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 3, 1, 2, 1, 2, 2, 0, 0, 0, -1, -1, -2, -1, -2, -3, -2, 0, 0, 2, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, -2, -2, 0, 1, 1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, 1, 1, 3, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, 0, 1, 0, -1, 0, -2, -3, -2, -3, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, -3, -1, -2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 1, 1, 2, 1, 1, 1, 1, 1, 1, 3, 2, 2, 2, 2, 2, 2, 1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 1, 2, 1, 1, 1, 1, 0, 1, 2, 2, 1, 2, 3, 3, 3, 2, 3, 2, 3, 3, 3, 3, 0, 0, 0, 0, -1, 0, 0, 1, 0, 2, 1, 1, 2, 1, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 3, 4, 2, 4, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 2, 0, 1, 0, 0, 0, 0, -2, -2, -2, -2, -2, -2, -1, 0, -1, 0, 0, 1, 2, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, -1, -2, -3, -3, -4, -2, -3, -1, 0, 0, 0, 0, 1, 1, 2, 2, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, -1, -2, -3, -3, -5, -2, -2, 0, -1, 0, 0, 0, 0, 2, 3, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, -1, -2, -3, -3, -3, -1, 0, 0, 0, 0, 1, 0, 3, 3, 2, 0, 0, 1, 0, -1, -1, 0, 0, -1, -1, 0, 0, 1, 1, 1, 2, 0, -1, -2, -3, -1, -1, -1, -1, 0, 0, 1, 2, 2, 2, 2, 2, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 1, 1, 1, 2, 0, 0, -1, -1, -3, -1, 0, -1, 0, 1, 2, 0, 1, 1, 2, 2, 0, 1, 1, 0, 1, 0, 0, -1, -1, -1, -2, 0, 0, 0, 2, 3, 1, 0, -1, -1, -2, -1, 0, -1, -1, 1, 1, 1, 0, 1, 2, 1, 0, 1, 1, 0, 1, 1, 0, -1, -1, -2, -2, -1, 1, 1, 2, 2, 2, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 3, 2, 0, 1, 1, 0, 1, 1, 1, 0, -2, -1, -1, -1, 0, 2, 1, 1, 0, 1, 0, -1, -2, 0, -1, -1, -1, -1, 0, 0, 0, 2, 2, 2, 0, 1, 0, 0, 1, 1, 0, 0, -1, -2, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -1, 0, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, 0, 3, 2, 0, 0, 1, 0, 1, 0, 0, 0, -1, -3, -3, -1, 0, 1, 2, 2, 1, 0, 0, -1, 0, 0, 0, -1, -1, -1, -2, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -3, -1, 0, 1, 2, 2, 0, 0, -1, 0, 0, 0, 0, -1, -2, -2, -1, -1, 0, 0, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, -2, -3, -2, -2, -1, 0, 2, 3, 0, 0, -1, -1, 0, 0, 0, -1, -1, -3, -1, -1, -1, 0, 2, 1, 0, -1, 0, 0, 1, -1, 0, -1, -1, -1, -4, -3, -1, 0, 2, 3, 2, 0, 0, 0, 0, -1, 0, -1, -1, -3, -3, -1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -3, 0, 1, 1, 3, 3, 1, 0, 0, 0, -1, -1, -2, -2, -3, -2, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, -3, 0, 0, 2, 3, 2, 0, 0, 0, 0, -1, 0, -1, -3, -3, -2, 0, 0, 2, 2, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 1, 3, 3, 2, 0, 0, 0, 0, -1, 0, -2, -2, -1, -1, 0, 0, 3, 4, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -2, 0, 0, 1, 2, 2, 0, 0, 0, -2, -3, -1, -2, -1, -1, 0, 1, 2, 2, 4, 2, 0, 0, 1, 1, 1, 1, 0, -1, -1, -1, -1, -1, 0, 1, 1, 1, 1, 1, 0, -1, -3, -3, -3, -2, -1, 0, 0, 0, 2, 3, 3, 2, 0, 1, 1, 1, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 0, 0, 0, -2, -2, -2, -3, -2, -1, 0, 0, 1, 1, 2, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -3, -2, -1, -1, 0, 0, 0, 1, 2, 3, 3, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, -1, -3, -4, -4, -4, -2, 0, 0, 0, 0, 1, 3, 3, 4, 2, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -3, -4, -4, -4, -3, -2, 0, 0, 0, 0, 2, 2, 4, 4, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -3, -4, -4, -5, -3, -1, 0, 0, 0, 1, 2, 2, 3, 4, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -4, -4, -4, -3, -2, -1, 0, 1, 1, 2, 4, 3, 3, 2, 0, -1, 0, -2, 0, 0, 1, 1, 0, 1, 1, 1, 2, 2, 0, 1, 0, -1, -3, -3, -2, -1, 0, 0, 0, 0, 2, 2, 3, 4, 2, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 1, 1, 1, 1, 2, 3, 2, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, -2, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 2, 0, 0, -1, 0, -1, -1, -3, -1, -2, -2, -2, -3, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 1, 0, 1, 1, 0, 3, 1, 0, -1, -1, 0, 0, 0, -1, -1, -3, -3, -1, -2, -1, -1, -2, -2, 0, -1, -2, 1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 2, 5, 3, 0, 0, 1, 0, 1, 0, 0, 1, -1, -2, 0, 0, -1, 0, -2, -2, 0, 0, -1, 2, 1, -1, -1, -1, 0, 1, 1, 2, 3, 4, 4, 3, 1, 3, 1, 1, 2, 3, 1, 2, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 2, 0, 4, 3, 4, 4, 3, 2, 4, 3, 2, 2, 3, 2, 2, 2, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 2, 2, 3, 3, 2, 4, 2, 1, 4, 3, 1, 0, 2, 2, 4, 4, 0, 3, 2, 1, 0, 0, 1, 0, 0, 0, 3, 1, 0, 0, 0, 0, 0, 2, 3, 1, 2, 2, 2, 3, 3, 1, 0, 2, 2, 3, 4, 4, 0, 2, 3, 0, 1, -1, 1, 0, 0, 0, 2, 3, 1, 1, 0, 2, 0, 2, 1, 1, 3, 2, 1, 3, 3, 3, 0, 2, 0, 1, 4, 1, 0, 1, 2, 2, 0, 0, 0, 1, 0, -2, 3, 4, 3, 1, 1, 2, 3, 3, 3, 2, 3, 2, 2, 4, 3, 2, 0, 2, 0, 1, 2, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 3, 2, 1, 1, 1, 1, 3, 3, 3, 4, 2, 2, 4, 3, 2, 0, -1, 0, 2, 3, 1, 0, 1, 2, 1, 1, -1, -2, 0, 0, -1, 1, 2, 2, 1, 2, 2, 2, 2, 2, 4, 5, 3, 3, 4, 3, 1, 0, -1, 0, 1, 2, 1, 1, 2, 3, 2, 1, 0, -1, 0, 0, 0, 3, 1, 2, 1, 2, 1, 2, 3, 3, 4, 5, 4, 5, 4, 1, 0, 0, -1, -1, 0, 1, 1, 0, 2, 4, 3, 1, 0, -1, 0, 1, 2, 4, 0, 0, 2, 1, 1, 3, 2, 3, 4, 5, 5, 5, 5, 2, 0, 1, 0, 0, 0, 0, 2, 0, 2, 4, 4, 2, 0, 0, 0, 1, 2, 3, 0, -1, 0, 2, 1, 2, 2, 3, 4, 4, 4, 6, 7, 3, 0, 0, 1, -1, -2, 0, 0, 0, 1, 4, 3, 3, 1, -2, 0, 0, 3, 3, 0, 0, 0, 1, 2, 1, 2, 3, 4, 5, 3, 5, 4, 2, 1, 1, 1, -1, -3, 0, 0, 0, 1, 4, 4, 0, 0, -1, 0, 0, 2, 1, -1, 1, 1, 1, 1, 2, 3, 5, 4, 4, 4, 4, 4, 2, 1, 0, 2, 0, 0, -1, 0, 1, 2, 4, 4, 0, 0, -1, 0, 0, 2, 0, 0, 0, 2, 0, 1, 2, 3, 4, 3, 4, 3, 4, 3, 2, 2, 2, 3, 0, 0, 0, 0, 1, 2, 4, 2, 1, 0, -1, 0, 1, 0, 1, 0, 2, 3, 0, 1, 2, 3, 4, 2, 4, 3, 2, 3, 3, 1, 1, 2, 0, 1, 0, 1, 0, 1, 2, 3, 0, -1, -1, 0, 0, 1, 0, 1, 2, 1, 0, 1, 3, 3, 3, 2, 3, 3, 1, 3, 4, 1, 0, 2, 1, 0, 2, 1, 2, 2, 2, 1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 2, 1, 1, 4, 3, 3, 2, 3, 4, 3, 3, 3, 1, 0, 2, 1, 0, 1, 1, 1, 3, 2, 1, 2, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 0, 3, 2, 2, 2, 1, 4, 2, 2, 4, 0, 0, 0, 0, 0, 0, 1, 0, 3, 2, 0, 1, 0, 1, 0, 0, 0, 1, 3, 2, 2, 0, 0, 2, 1, 0, 0, 1, 4, 3, 2, 2, 0, 0, 0, 0, 1, 1, 1, 1, 3, 1, 0, 1, 0, 0, 0, 1, 0, 1, 3, 3, 3, 1, 1, 2, 2, 0, 1, 3, 5, 3, 1, 0, 0, 0, 1, 2, 2, 1, 0, 2, 2, 0, 0, 0, 0, -1, 0, 0, 0, 2, 3, 2, 2, 0, 0, 2, 2, 1, 1, 2, 4, 1, 0, 0, 0, 0, 0, 1, 2, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 3, 1, 2, 0, -1, 1, 1, 1, 1, 3, 4, 1, 0, 1, 0, 1, 1, 0, 1, 2, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, -1, 0, 2, 1, 2, 5, 1, 1, 2, 1, 1, 1, 0, 1, 2, 2, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 3, 2, 5, 3, 0, 0, 1, 1, 0, 1, 2, 1, 2, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 2, 0, 0, 0, 3, 3, 3, 4, 1, 0, 1, 0, 2, 2, 2, 0, 0, 1, 0, 0, 0, -1, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 0, -1, 0, 2, 2, 3, 2, 1, 0, 0, 2, 1, 0, 1, -1, -1, -1, 0, 0, -1, -1, -2, 0, 0, 0, 0, -3, 0, 0, -1, 0, 1, 0, 0, 0, 1, 2, 2, 2, 0, 0, 1, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, -1, 0, 0, 0, 1, 1, 1, 2, 1, 1, 1, 2, 1, 1, 0, 1, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 2, 1, 1, 2, 1, 2, 3, 6, 6, 6, 5, 3, 0, 0, 0, -1, 1, 2, 0, 0, 1, 0, -2, -2, -1, 0, 0, 0, 1, 0, 0, 1, 2, 2, 0, 0, 0, 1, 2, 4, 4, 5, 6, 6, 2, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 1, 2, 1, 0, 1, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, -1, 1, 1, 0, 0, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, 0, 0, 2, 2, 1, 0, 0, 1, 0, -1, 0, 0, 0, -1, -1, -1, -2, -3, -3, -1, -2, -1, 0, -1, -1, -2, -2, -1, 0, -1, 0, 0, 0, 0, 2, 2, 1, 0, 1, 0, 0, 0, 0, 2, 0, 0, 0, -2, -2, -4, -4, -3, -3, -2, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, -4, -5, -4, -2, 0, 0, 1, 0, 1, -1, 0, 1, 0, 1, 0, 0, 1, 2, 1, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -3, -4, -2, -2, 0, 1, 1, 2, 0, 0, 0, 1, 1, 1, 0, 0, 2, 2, 2, 0, 0, 0, -1, -2, -1, -2, 0, 0, -1, 0, 0, -1, -3, -3, -4, -3, -3, 0, -1, 0, 0, 0, 0, -1, 1, 1, 0, 0, 1, 3, 2, 1, 1, 1, -1, -1, -1, -3, -2, -2, -2, 0, 0, 0, -1, -2, -3, -3, -4, -3, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 1, 0, 0, -1, -2, -2, -2, -3, -3, -3, -1, -2, -1, -3, -3, -3, -5, -3, -3, -2, -1, 0, 0, 0, -2, 0, 1, 0, 0, 0, 2, 1, 0, 0, -1, -2, -3, -2, -3, -2, -2, -2, -2, -3, -3, -4, -4, -4, -4, -1, -2, 0, 0, 0, 1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -3, -4, -4, -2, -3, -1, -1, -3, -4, -3, -3, -2, -1, -2, -1, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -3, -3, -3, -3, -2, 0, 0, 0, -1, -2, -3, -1, -1, -1, -2, -1, -1, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -2, -3, -3, -3, -3, -3, -2, -1, 0, 0, -2, -2, -1, -2, -2, 0, -1, -2, 0, 0, 0, 0, 0, -2, -1, 0, 0, 1, 1, 0, 0, 0, -1, -3, -4, -4, -3, -4, -5, -4, -1, 0, -1, -2, -2, -3, -1, 0, 0, 0, 0, -1, 0, -1, 0, -2, -2, 0, 0, 2, 1, 0, 0, 0, -2, -2, -3, -3, -3, -4, -4, -3, -4, -2, -2, -2, -2, -3, -3, -1, -1, -2, -2, -1, -1, 0, 0, 0, -2, 0, 0, 0, 2, 0, 0, -1, -1, -1, -1, -3, -2, -3, -1, -2, -4, -4, -2, -2, -1, 0, 0, 0, 0, -1, -2, -2, -1, -1, -1, -2, -2, -1, 0, 1, 2, 1, 0, 0, -1, -1, -1, -2, -2, -2, -3, -1, -2, -3, -2, -2, -1, 0, 1, 0, -1, -1, -1, -1, -1, -2, -2, -2, -2, -1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, -1, -1, -2, -2, -3, -2, -3, -3, -1, 0, 0, 0, -2, -2, -2, -1, -3, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -3, -2, -3, -2, -2, -1, -1, -1, -1, -2, -2, -2, -2, -1, -1, -1, -2, 0, 0, 2, 1, 0, 1, 0, -1, 0, 1, 1, 0, 1, 0, 0, -1, -1, -3, -2, -2, -3, -4, -3, -2, -3, -3, -2, -2, -1, 0, -1, -1, 0, 0, 3, 1, 1, 2, 0, 0, 0, 0, 1, 0, -1, -1, -1, -1, -2, -3, -2, -2, -3, -3, -3, -4, -4, -3, -3, -2, -2, -1, -2, -1, 0, 0, 2, 2, 2, 1, 1, 1, 1, 1, 0, 0, 0, -2, -3, -3, -3, -3, -3, -1, -2, -2, -3, -4, -3, -3, -3, -1, -2, -2, -1, -2, 0, 2, 2, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, -3, -3, -4, -2, -1, -2, -2, -3, -1, -1, 0, 0, 0, -1, -1, -2, 0, 1, 2, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 1, 0, -1, -2, 0, -1, -1, -2, -3, -2, -2, 0, 1, 0, 0, -1, -2, 0, 0, 3, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 1, 2, 2, 2, 0, -1, 0, 0, -1, -1, -2, -3, -2, -1, 0, 0, 0, -2, -1, 0, 1, 2, 3, 1, 0, 0, 0, 0, 0, 0, 0, 2, 4, 5, 4, 4, 2, 1, -1, -1, -2, -2, -2, -4, -4, -3, -2, -1, -1, -1, -3, 0, 1, 3, 2, 2, 2, 2, 2, 1, 2, 2, 1, 2, 4, 5, 5, 5, 3, 3, 0, -1, -4, -5, -4, -5, -4, -3, -4, -2, -2, -1, -1, -1, 0, 0, 2, 2, 1, 2, 1, 0, 1, 2, 1, 1, 1, 1, 1, 0, 0, -1, -2, -2, -4, -4, -5, -5, -5, -5, -3, -2, 0, 0, 0, 0, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, -1, -1, -1, 0, 0, 1, 2, 1, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -3, -3, -2, -1, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, -1, -2, -1, -2, 0, -2, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -2, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 2, 3, 1, 0, 0, -1, 0, 0, -2, -2, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, -2, -2, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 0, 0, -1, 0, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, -1, -1, -2, -2, -1, 0, 0, -1, 0, 0, 0, 0, 1, 2, 0, 1, 1, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, 0, -1, -2, -2, -1, -2, 0, -1, -1, 0, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, -1, 0, 0, -2, -2, -2, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -2, -2, -1, 0, 0, 0, -1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 1, 1, 0, 0, 0, -1, -1, -2, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, -1, -2, -3, -2, -1, -2, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -2, -3, -2, -2, -1, -1, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 1, 1, -1, 0, 0, 0, 1, 1, 1, 2, 0, 1, 0, -1, -1, -2, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, -2, 0, -1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 3, 2, 1, 3, 2, 2, 2, 3, 4, 4, 3, 3, 3, 3, 3, 4, 3, 3, 3, 1, 0, 0, -2, -2, 0, 0, 0, 1, 0, 1, 2, 3, 2, 2, 3, 2, 2, 3, 3, 2, 3, 4, 3, 3, 3, 3, 4, 4, 5, 4, 4, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 2, 0, 2, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 2, 3, 4, 4, 3, 0, -1, -2, 0, 0, 0, 0, 2, 2, 2, 1, 0, 1, 0, 0, 0, -1, -3, -3, -3, -3, -3, -2, -1, -1, -1, 0, 1, 3, 4, 3, 3, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, -1, -3, -3, -5, -4, -3, -2, -2, 0, 0, 0, 0, 0, 3, 3, 2, 0, 0, -2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, -1, -1, -4, -4, -4, -3, -3, -2, 0, 0, 0, 1, 0, 3, 3, 4, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 3, 2, 1, 0, -1, -2, -2, -3, -2, -2, -1, 0, 0, 0, 2, 3, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 2, 1, -2, -1, -2, -1, -2, -1, 0, 0, 1, 1, 2, 2, 3, 1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, 0, 1, 3, 2, 2, 2, 1, 0, 0, -1, -3, -3, -2, 0, 0, 0, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 2, 3, 3, 1, 2, 1, 0, 0, -1, -1, -2, -3, 0, 0, 0, 1, 1, 3, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, 0, 0, 2, 2, 2, 2, 3, 1, 1, 0, 0, -2, -2, -2, 0, 0, 0, 0, 2, 3, 3, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 1, 3, 3, 3, 2, 2, 1, 0, 0, 0, -1, -1, -2, -1, -1, 0, 2, 3, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 2, 1, 3, 3, 4, 3, 3, 2, 0, 0, -1, -4, -3, -2, -2, -1, 1, 3, 3, 1, 1, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 3, 2, 3, 3, 2, 4, 3, 3, 1, 0, -3, -3, -3, -3, -3, -2, 1, 2, 2, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, -1, -1, 0, 2, 3, 2, 3, 2, 3, 2, 2, 0, 0, -3, -4, -4, -4, -3, -1, 0, 2, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, -1, 2, 3, 2, 2, 3, 3, 1, 1, 1, 0, 0, -2, -3, -4, -4, -2, -1, 1, 2, 2, 0, 0, 0, 1, 1, 0, 1, 0, -1, -3, -1, 0, 1, 2, 3, 3, 2, 2, 1, 1, 2, 2, 0, -1, -3, -4, -3, -3, -2, 1, 1, 3, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, 0, 2, 3, 2, 3, 2, 1, 2, 1, 1, 1, 0, -1, -3, -4, -4, -2, -1, 2, 1, 3, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -2, 0, 1, 2, 4, 3, 2, 2, 3, 1, 2, 1, 0, -2, -4, -3, -3, -1, 0, 2, 2, 2, 0, -1, 0, 0, -1, 0, 0, 0, -1, -2, -2, -1, 0, 3, 4, 2, 3, 4, 2, 1, 1, 0, 0, -3, -3, -3, -2, 0, 0, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, 0, 1, 4, 3, 4, 2, 2, 0, 0, 0, -2, -4, -4, -2, -2, 0, 1, 2, 2, 2, 0, 0, 1, 0, 1, 0, 0, 0, -3, -2, -1, -1, 0, 1, 3, 2, 3, 4, 1, 1, 0, -1, -1, -2, -3, -2, 0, 0, 2, 3, 2, 3, 0, 0, 1, 2, 1, 1, 0, -1, -2, -2, -1, 0, -1, 2, 2, 2, 4, 2, 2, 0, 0, -1, -1, -3, -2, -1, 0, 0, 2, 2, 3, 3, 1, 0, 0, 1, 1, 0, 0, -1, -1, -2, -2, 0, 0, 2, 3, 2, 2, 3, 0, 0, -2, -2, -3, -2, -1, -1, 0, 0, 1, 3, 2, 2, 0, 0, -1, 1, 0, 0, 0, -1, -2, -2, 0, 0, 0, 1, 2, 3, 2, 0, 0, 0, 0, -2, -1, -2, -1, -1, 0, 1, 3, 3, 3, 2, 0, -1, -1, -1, -1, -1, 0, -1, 0, -2, -2, 0, -1, 0, 3, 2, 0, -1, -1, -2, -3, -2, -3, -1, 0, 0, 0, 1, 3, 5, 2, 3, 0, 0, -1, -1, 0, 0, 0, -1, 0, -2, -2, 0, 0, 1, 0, 0, 0, -2, -4, -3, -2, -3, -1, -2, -1, 0, 1, 1, 3, 4, 2, 2, 0, 0, -2, -1, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 1, 0, -1, -3, -4, -2, -3, -2, -1, 0, 0, 1, 2, 3, 3, 4, 4, 2, -1, 0, -3, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -2, -2, -2, -3, -1, 0, 0, 1, 1, 3, 2, 3, 3, 6, 3, 3, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 1, 2, 2, 4, 4, 5, 4, 5, 4, 3, 3, -1, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 2, 3, 4, 4, 5, 4, 3, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, -2, -1, -1, -2, -1, -1, -1, -3, -1, -2, -3, -3, -4, -4, -5, -4, -3, -3, -3, -4, -4, -4, -4, -2, -2, -3, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, -2, -1, -2, -1, -3, -2, -2, -3, -5, -5, -4, -3, -2, -3, -2, -3, -4, -3, -4, -4, -3, -2, -3, -2, 0, -1, 0, 0, 0, 0, -2, -1, -1, -1, -2, 0, -2, -2, -2, -3, -3, -4, -3, -2, 0, -1, -1, -1, -2, -2, -2, -3, -3, -2, -4, 0, 0, -1, 0, 0, 0, -1, -3, -1, -2, -2, 0, -1, -1, -2, 1, 0, 0, -2, -2, 0, 0, 0, 0, 1, 1, 0, 0, -1, -2, -2, -4, -1, 0, -2, -1, 0, 0, -1, -3, -1, -2, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 2, 0, 0, 0, -1, -1, -2, -1, 0, -2, 0, 0, -1, -1, -2, -3, -2, -1, 0, 0, 0, 0, 2, 1, 0, 0, 2, 0, 0, 2, 2, 3, 3, 1, 0, 1, 0, -1, -1, -1, -1, -1, -1, 1, -1, -2, -1, -1, -2, -1, 0, 0, 1, 1, 3, 0, 0, 3, 2, 2, 1, 2, 1, 4, 3, 2, 0, 0, 1, -1, -1, -1, -1, -1, -1, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 2, 1, 1, 0, 2, 2, 2, 0, 1, 1, 5, 4, 2, 1, 0, 1, 0, -1, -1, 0, -1, -2, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 3, 1, 1, 0, 1, 2, 0, 1, 2, 2, 5, 3, 1, 1, 0, 0, 0, -1, -1, -1, -2, -1, -1, -1, 0, 0, 0, 1, 0, 0, 1, 1, 3, 3, 2, 3, 1, 2, 0, 0, 1, 2, 4, 3, 2, 2, 2, 0, 1, -2, -2, 0, -1, -1, -1, -1, -1, -1, 0, 1, 0, 0, 2, 1, 3, 4, 2, 2, 2, 1, 0, 0, -1, 3, 3, 1, 1, 2, 3, 1, 0, -1, -2, 0, -1, -1, 0, 0, 0, 0, 1, 1, -1, 0, 0, 2, 3, 4, 4, 3, 1, 0, 0, 0, 0, 1, 2, 2, 1, 2, 3, 3, 0, -2, -4, 0, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 3, 4, 3, 3, 3, 1, 0, 0, -1, -2, 0, 1, 1, 1, 2, 5, 3, 0, -2, -2, -1, 0, 1, 1, -1, -1, 0, 2, 1, 1, 2, 2, 3, 4, 2, 3, 4, 1, 0, 0, -1, -3, 0, 1, 2, 2, 4, 5, 3, 0, -1, -3, 0, -1, 1, 0, -1, 0, 0, 1, 2, 3, 3, 1, 2, 4, 1, 2, 3, 0, -2, -2, 0, 0, -3, 0, 2, 3, 3, 4, 4, 0, -1, -3, -1, 0, 1, 2, -1, 0, 1, 3, 4, 3, 3, 1, 3, 3, 0, 2, 3, 0, 0, 0, 0, 0, -2, 0, 2, 3, 3, 4, 2, 1, -1, -3, -1, 0, 3, 0, -1, 0, 2, 3, 3, 5, 2, 2, 4, 3, 1, 2, 4, 1, 0, 0, 0, 0, -1, 1, 2, 2, 4, 3, 3, 1, -1, -3, -1, 0, 1, 0, 0, 1, 1, 3, 4, 3, 2, 3, 1, 4, 2, 2, 3, 0, 0, 0, 0, 0, -1, 1, 2, 1, 3, 4, 4, 0, 0, -1, 0, 0, 2, 0, 0, 0, 2, 3, 3, 3, 1, 3, 1, 2, 2, 3, 3, 1, 0, -1, 1, 0, -1, 1, 2, 2, 3, 3, 1, 1, 0, -1, -1, 0, 1, 0, -1, 0, 3, 2, 1, 3, 2, 2, 0, 1, 1, 2, 3, 2, -2, -2, 1, 0, 0, 3, 2, 2, 3, 3, 0, 0, -1, 0, -1, 0, 0, -1, -1, 1, 1, 2, 1, 2, 1, 2, 2, 2, 2, 2, 2, 2, 0, -1, 2, 1, 1, 1, 1, 1, 3, 0, 0, 0, -1, 0, 0, 0, -1, -2, -1, 1, 1, 1, 2, 2, 2, 2, 1, 1, 2, 2, 2, 3, 0, -1, 1, 0, 0, 1, 1, 1, 1, 1, 0, 0, -2, 0, 0, 0, 0, 0, -1, 0, 1, 2, 0, 3, 1, 0, 0, 2, 3, 1, 2, 0, 0, 0, 1, 1, 0, 2, 2, 1, 2, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 2, 0, 2, 0, 0, 0, 1, 3, 3, 2, 1, -1, -1, 0, 0, 0, 2, 2, 1, 0, 0, -1, -1, -3, -1, 0, -1, 0, 1, 0, 1, 0, 0, 0, 1, 1, 1, 1, 2, 3, 1, 2, 0, 0, 0, 0, 1, 0, 1, 1, 2, 0, 0, -1, -1, -2, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 3, 1, 1, 2, 2, 1, 0, 0, 1, 3, 2, 2, 0, -1, -1, -3, -3, -1, 0, -1, 0, 0, 0, -1, 1, 1, -1, -2, -1, 0, 1, 1, 2, 1, 1, 3, 2, 1, 0, -1, 0, 2, 1, 2, 0, 0, -3, -3, -2, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, -1, 0, -2, -3, -3, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, -3, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, -2, -2, -2, -3, 0, 0, -1, -1, 0, -1, -2, 0, 0, 0, -1, -2, -1, 0, -2, -1, -1, -2, -2, -1, -3, -2, 0, 0, 0, 0, -1, -2, -1, -4, -3, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -2, -2, -2, -1, -4, -2, -2, 0, -1, -2, -2, -3, -2, -2, -3, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -2, -1, 0, -2, -2, -2, -3, -3, -3, -3, -3, -3, -1, -2, -3, -2, -3, -1, -3, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -2, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -2, -3, -2, -1, 0, 0, 0, 1, 0, -1, -2, -4, -5, -5, -5, -4, -4, -3, -2, -1, 0, 1, 0, 0, 1, 2, 2, 1, -1, -2, -2, -2, -2, -2, -1, 0, -1, -1, 1, 1, 1, 0, -3, -4, -4, -4, -4, -4, -4, -2, -2, -1, -1, 0, 0, 0, 1, 0, 1, 1, 0, -2, -2, -2, -3, -2, -1, -1, 0, 0, 1, 2, 1, 1, 0, -1, -1, -1, -2, -1, -1, 0, 0, -2, -2, -1, 0, 0, -1, 0, 1, 1, -1, 0, 0, 0, -2, 0, -1, 0, 0, 0, 1, 1, 2, 2, 2, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, -1, -1, 0, 0, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 3, 2, 3, 2, 2, 2, 3, 2, 0, 0, 1, 0, 0, -1, 0, -2, -1, -1, 1, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 2, 2, 3, 3, 3, 4, 4, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 1, 2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 4, 4, 2, 4, 5, 2, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 1, 0, 0, 0, 2, 1, 1, 0, 1, 0, 0, -1, -1, 1, 3, 3, 4, 3, 4, 3, 2, 1, 0, -1, 0, 1, -1, -2, 0, 0, -1, 0, 0, 1, 0, 1, 2, 2, 1, 0, 0, 1, 0, -2, -1, 0, 1, 2, 2, 3, 3, 2, 2, 1, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 1, 1, 3, 2, 0, 1, 0, 0, 0, 0, 0, 2, 3, 3, 3, 2, 2, 1, 1, 1, 2, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 1, 0, 1, 0, 1, 3, 3, 4, 4, 2, 3, 2, 0, 1, 2, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 2, 2, 4, 4, 5, 2, 1, 2, 2, 2, 0, 0, 1, 0, -1, -2, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 3, 3, 3, 4, 4, 5, 6, 3, 3, 3, 2, 2, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, -2, -1, 0, 2, 2, 2, 3, 2, 3, 4, 6, 4, 3, 2, 2, 2, -1, 0, 0, 0, -1, -1, -1, -2, -1, -1, -1, 0, 0, 0, -2, -2, -2, 0, 0, 3, 3, 2, 3, 3, 5, 4, 6, 4, 4, 1, 2, 0, -1, 0, -1, 0, 0, 0, -1, -1, -2, -2, 0, 0, 0, 0, -2, -2, -1, 0, 0, 2, 1, 3, 2, 3, 3, 4, 4, 5, 2, 2, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, 0, 0, -2, -2, -1, 1, 0, 1, 2, 1, 1, 2, 2, 5, 5, 3, 4, 3, 1, 0, 1, 0, 1, 2, 0, -1, -1, -2, -2, 0, 0, 0, 0, 0, -2, -1, -1, 2, 2, 2, 2, 1, 2, 1, 1, 2, 3, 3, 4, 2, 2, 1, 1, 0, 0, 2, 1, 0, -2, -2, -2, 0, 0, 1, 0, 0, -2, -1, 0, 0, 2, 1, 1, 0, 1, 0, 1, 2, 2, 5, 3, 3, 2, 2, 2, 1, 1, 1, 0, -2, -1, -2, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 2, 0, 0, 0, 0, 1, 1, 1, 3, 4, 4, 2, 2, 2, 2, 2, 0, 0, -1, -1, -2, -2, -1, 0, 2, 2, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, -1, -1, 1, 0, 2, 1, 2, 0, 2, 2, 1, 0, 0, -1, -2, -1, -1, -2, 0, 1, 2, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -3, -2, 0, 0, 1, 2, 0, 1, 0, 2, 3, 2, 0, 0, -1, -2, -1, 0, 0, 1, 1, 3, 2, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -2, 0, 2, 2, 2, 2, 1, 2, 2, 3, 3, 1, 0, 0, 0, 0, -1, 0, 0, 1, 3, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -2, 0, 2, 2, 2, 3, 1, 2, 2, 1, 0, 0, 0, 0, -2, -2, -1, 0, 1, 2, 3, 1, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 1, 2, 3, 2, 3, 3, 1, 0, -1, -1, -1, -1, -2, -2, -3, -2, 0, 1, 2, 2, 0, 0, 0, 0, -1, -1, -1, -2, -2, 0, 0, 2, 1, 3, 2, 2, 2, 2, 2, 0, -3, -2, -2, -1, -3, -3, -4, -4, -2, 1, 1, 2, 0, 0, 0, 0, -1, -1, 0, -2, -1, 0, 0, 2, 1, 1, 0, 0, 1, 1, 1, 0, -2, -2, -1, -1, -2, -2, -4, -4, -2, 0, 1, 1, 0, 0, -1, -1, -1, -1, -2, -2, -2, -1, 0, 2, 0, 0, -2, -2, 0, 0, 0, -1, -2, -2, -2, 0, -1, -3, -2, -2, 0, 2, 3, 1, 0, -1, -1, -1, -1, -1, -1, -1, -2, -1, 0, 0, 0, -1, -3, -3, -3, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 4, 4, 3, 0, 0, 0, -2, -1, 0, 0, -1, -1, -2, 0, -1, -1, -1, -1, -2, -2, -2, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 2, 3, 4, 2, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, -1, -2, 0, 0, 0, 2, 2, 2, 1, 1, 2, 1, 2, 2, 2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 2, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 1, 1, 2, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 2, 2, 1, 2, 2, 1, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 1, 1, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 2, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 2, 1, 0, 0, 1, 1, 1, 1, 1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 2, 2, 1, 0, -1, 0, 0, 0, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, -1, -1, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 2, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 2, 0, 0, 2, 1, 2, 1, 2, 1, 2, 3, 3, 2, 3, 2, 2, 3, 3, 3, 3, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 1, 2, 2, 2, 2, 2, 3, 4, 4, 3, 2, 2, 2, 2, 3, 3, 2, 2, 2, 3, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 1, 2, 1, 2, 1, 3, 3, 2, 2, 2, 1, 0, 0, 0, 1, 1, 2, 3, 4, 3, 2, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 0, 1, 0, 2, 1, 2, 1, 0, 0, 0, -1, 0, -1, -1, -1, -2, -2, -2, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 2, 3, 3, 1, 0, 1, 1, 3, 1, 2, 1, 1, -2, -3, -3, -2, -2, -2, -2, -1, -2, -2, 0, 1, 2, 1, 0, 0, 1, 2, 1, 0, 1, 2, 1, 1, 0, 0, 1, 3, 3, 3, 1, 0, -2, -5, -4, -3, -4, -3, -3, -2, -1, -3, -2, 0, 0, 1, 0, 0, 1, 2, 0, 1, 1, 2, 1, 1, 0, 1, 3, 3, 3, 2, 1, 0, -2, -4, -5, -4, -3, -3, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 2, 1, 0, 0, 0, 1, 1, 0, -1, 0, 1, 4, 3, 2, 2, 0, -2, -2, -3, -4, -2, -3, -1, 0, 0, 0, 0, 2, 2, 2, 1, 0, 2, 2, 1, 0, 0, 0, 0, -1, -1, 0, 0, 3, 2, 3, 2, 1, -1, -2, -4, -3, -3, -1, -1, 0, 0, 0, 1, 1, 2, 3, 1, 0, 3, 2, 0, 0, 2, 0, 0, 0, -2, -2, 0, 1, 2, 2, 1, 1, -1, -3, -2, -4, -4, -3, -3, -1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 1, 2, 0, -2, -2, -1, -1, 0, 1, 0, 1, 1, 0, -2, -3, -4, -4, -4, -3, -3, -1, 0, 0, -1, 1, 1, 1, 0, 2, 2, 0, 0, 1, 1, -1, -3, -3, -2, -2, 0, 0, 1, 2, 1, 0, -1, -1, -4, -5, -3, -4, -3, -2, 0, -2, -1, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, -3, -4, -3, -1, 0, 0, 1, 0, 2, 0, -1, -2, -3, -3, -3, -3, -4, -3, -1, -2, -2, 0, 1, 1, 2, 1, 1, 0, 0, 1, 0, 0, -3, -4, -4, -2, 0, 1, 0, 2, 0, 0, -2, -2, -2, -2, -2, -4, -3, -3, -3, -3, -2, -1, 1, 0, 1, 1, 0, 0, 0, 1, 0, -1, -3, -4, -4, -3, -1, 0, 2, 1, 0, 0, -2, -2, -2, -2, -3, -3, -5, -5, -4, -3, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -3, -4, -5, -4, -3, -1, 0, 1, 3, 2, -1, -2, -2, -2, -1, -2, -4, -4, -4, -5, -3, -2, -1, 0, 0, 1, 0, 1, 1, 1, 0, 0, -3, -4, -5, -4, -4, -2, 0, 1, 1, 2, 0, -2, -2, -3, -3, -2, -4, -4, -4, -4, -3, -2, -1, 0, 0, 0, 0, 1, 2, 1, 0, -1, -2, -3, -4, -3, -4, -3, 0, 0, 1, 0, 0, 0, -3, -3, -2, -1, -3, -4, -5, -5, -3, -2, -2, 0, 0, 1, 0, 1, 2, 2, 0, -2, -2, -3, -2, -3, -3, -1, -2, 0, 0, 0, 0, 0, -1, -2, -1, -1, -2, -4, -5, -4, -3, -1, 0, 0, 0, 1, 0, 2, 1, 1, 0, 0, -2, -1, 0, -2, -2, -1, 0, 0, 1, 0, 0, -1, -1, -1, -1, -1, -2, -3, -4, -4, -3, -1, 0, 1, 0, 0, 1, 1, 2, 1, 0, 0, -2, -1, -1, 0, -1, -1, 0, 0, 2, 0, -1, 0, -1, -2, -1, -1, -4, -5, -3, -3, -2, -1, 0, 1, 1, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 0, 0, -1, -2, -4, -2, -3, -5, -4, -3, -3, -1, -1, 0, 0, 1, 0, 2, 1, 0, 1, 0, 0, 0, -1, 0, 1, 1, 1, 3, 1, 2, 1, -1, -1, -3, -3, -4, -5, -5, -5, -3, -2, -1, 0, 1, 0, 0, 1, 2, 2, 0, 0, 2, 0, 0, 0, 0, 0, 1, 1, 3, 2, 2, 0, 0, -2, -3, -5, -5, -6, -5, -4, -3, -1, -1, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 1, 1, 1, 1, 1, 2, 0, 0, -1, -3, -4, -4, -5, -4, -5, -3, -4, -2, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 3, 1, 1, 0, 0, -4, -5, -5, -4, -4, -3, -3, -3, -2, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 1, 1, 3, 2, 2, 3, 1, 1, -2, -5, -4, -4, -3, -3, -2, -3, -2, -1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 4, 3, 3, 1, -1, -4, -5, -5, -3, -3, -2, -3, -2, 0, 0, 0, 3, 2, 0, 0, 1, 1, 1, 0, 1, 0, 1, 1, 2, 1, 1, 2, 3, 5, 4, 2, 0, -3, -5, -5, -4, -4, -3, -4, -3, -1, 0, 0, 2, 0, 0, 0, 0, 2, 2, 1, 2, 0, 2, 3, 3, 3, 2, 2, 3, 3, 3, 4, 0, -1, -2, -2, -2, -3, -3, -2, -3, -2, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 2, 3, 3, 4, 2, 3, 2, 4, 4, 3, 3, 1, 0, -1, -2, -3, -3, -1, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 2, 1, 2, 2, 0, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 3, 2, 2, 3, 2, 2, 1, 1, 2, 1, 1, 0, -1, 0, -1, -2, -3, -2, -2, -2, -1, -1, -1, -3, -2, -3, -4, -1, -2, 0, 1, 2, 4, 2, 3, 3, 1, 1, 2, 2, 2, 1, 0, -1, 0, -2, -3, -3, -3, -4, -2, -1, -2, 0, 0, -1, -2, -3, -3, -1, 0, -1, 0, 2, 3, 2, 2, 2, 1, 0, 0, 0, 2, 0, 0, -1, -1, 0, 0, -1, -4, -3, -3, 0, 0, 1, 4, 2, 1, 1, -1, -2, 0, -1, 2, 3, 3, 3, 2, 1, 1, 0, 0, 1, 2, 0, 0, -1, -1, 0, -1, -1, -2, -3, -1, 0, 0, 1, 2, 3, 4, 3, 0, 0, -1, 0, 1, 1, 2, 2, 1, 1, 0, 0, 0, 1, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 3, 1, 1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 2, 2, 0, 0, 0, -1, 0, 0, 2, 1, 0, 2, 2, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 2, 1, 1, 2, 1, 1, 0, 0, 1, 2, 1, 1, 0, 0, 0, -1, 0, 2, 0, 0, 2, 4, 1, 1, 0, 2, 1, 0, 0, 0, 0, 1, 3, 2, 1, 1, 1, 1, 0, -1, 0, 1, 0, 0, 0, 1, -1, 0, 0, 1, 2, 1, 1, 5, 4, 2, 3, 3, 0, 0, 0, 0, 0, 0, 2, 2, 1, 1, 0, 1, 0, -1, 0, 0, 0, 1, 1, 0, -1, -2, -1, 0, 1, 0, 1, 4, 4, 3, 3, 1, 2, 0, 0, 1, 0, 1, 3, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -2, -2, 0, 0, 1, 3, 6, 4, 3, 1, 2, 2, 1, 1, 0, 1, 3, 3, 3, 1, 0, 0, 0, 0, 1, 0, -1, -2, 0, -1, -1, 0, -2, -2, -2, -2, 1, 3, 5, 5, 3, 1, 1, 3, 3, 1, 0, 0, 2, 3, 2, 3, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, -2, -2, -3, -2, -2, -2, 0, 2, 3, 4, 2, 1, 2, 4, 3, 2, 0, 0, 2, 1, 3, 2, 0, 0, -1, 1, 1, 0, -2, 0, 0, 0, -3, -3, -3, -2, -2, -1, 0, 1, 4, 4, 3, 2, 1, 4, 4, 3, 1, 0, 2, 1, 1, 2, 0, -2, -1, 1, 1, 0, -1, -2, 0, -1, -4, -6, -4, -1, 0, -1, 0, 1, 2, 2, 2, 3, 1, 3, 5, 3, 1, -1, 0, 2, 1, 3, 0, -1, -1, 0, 0, 0, -1, -2, 0, 0, -5, -4, -2, -2, 0, -1, -2, 0, 1, 2, 2, 3, 3, 2, 3, 2, 0, 0, 0, 0, 1, 3, 0, -1, -1, 0, 0, 0, -2, 0, 0, 0, -2, -4, -4, -2, -3, -1, -2, -1, 0, 1, 2, 5, 4, 3, 2, 2, 0, 0, 0, 1, 2, 2, 0, -2, 0, 0, 0, -1, -3, -2, 0, 1, -2, -2, -3, -3, -3, 0, 0, 0, 0, 2, 4, 5, 5, 4, 3, 2, 0, 0, 0, 0, 1, 3, 1, -1, 0, 0, 0, -1, -3, -3, -2, 0, -2, -1, -2, -2, -2, 0, 1, 1, 2, 3, 2, 4, 6, 4, 3, 3, 0, 0, 2, 0, 0, 0, 1, 0, -1, 0, -1, -1, -1, -3, -2, -1, -1, 0, -1, -4, -3, 0, 2, 2, 1, 3, 3, 3, 4, 5, 1, 1, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -2, 0, 0, -1, 0, 0, 3, 5, 3, 3, 3, 2, 3, 3, 1, 1, 1, 0, 1, 2, 1, 0, -1, 1, 0, -1, -1, -1, -2, -1, -1, -3, -1, 0, 0, -1, 0, 1, 5, 6, 3, 4, 2, 1, 3, 2, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, -1, -1, 0, -1, 0, 0, -2, -3, 0, 0, 0, 1, 2, 4, 4, 2, 3, 2, 1, 3, 3, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, -1, -3, 0, 0, 1, 2, 1, 3, 2, 4, 4, 3, 4, 3, 2, 0, 0, 0, 0, 1, 2, 1, 0, -1, -1, 0, 0, -1, -1, 0, -1, -1, -2, -2, 0, 1, 0, 1, 0, 0, 1, 3, 3, 4, 3, 2, 2, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 2, 0, 0, 0, 1, 1, 1, 2, 2, 1, 1, 0, -1, -1, 0, 1, 0, 1, 0, -1, 0, 0, 1, 1, 0, 0, -1, 0, -1, -1, 1, 1, 2, 0, 0, -1, 0, 0, 2, 1, 1, 2, 1, -1, 0, 0, 0, 1, 0, 1, 0, -1, 0, 1, 1, 0, 1, 0, -1, 0, -2, 0, 1, 1, 2, 1, -1, -1, 0, 0, 2, 3, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 1, 0, 2, 1, 0, -1, -2, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 2, 2, 0, 0, 0, 0, 0, 1, 1, 0, -1, -2, -1, 0, 0, -1, 0, -2, -2, -3, -2, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 1, 0, 0, 0, 0, -1, -2, -3, -4, -4, -4, -3, -4, -3, -4, -4, -5, -3, -2, 0, 2, 2, 1, 1, 0, 0, 0, 1, 0, 3, 3, 3, 3, 1, 0, 0, 1, 0, -3, -6, -7, -6, -5, -5, -6, -6, -7, -7, -6, -4, -1, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -5, -5, -5, -5, -5, -5, -5, -5, -5, -4, -4, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -2, -2, -1, -1, -1, -2, -1, -1, 0, -1, -1, -2, -2, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, -1, -2, -2, -2, 0, -1, 0, 0, -1, -2, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -1, 0, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -2, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -2, -1, -2, -1, -1, 0, -1, -1, -1, -1, -2, -1, -1, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -2, -2, -1, -2, -1, 0, -2, -1, 0, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 3, 0, -2, 0, 0, 1, 0, 0, -2, -4, -4, -4, -4, -3, -1, -2, -3, 0, 0, -2, 1, 0, 0, -2, 0, 0, 0, 2, 2, 3, 2, 5, 3, 1, 1, 0, 2, 3, 2, 2, 0, -2, -3, -2, -3, -2, 0, -4, -4, 0, 0, -1, 1, 0, -2, -1, 0, -1, 1, 1, 3, 4, 3, 7, 4, 4, 4, 2, 1, 3, 4, 4, 4, 3, 0, 0, 0, -1, 0, -4, -4, 0, 0, -1, 1, 0, -2, 0, -1, -1, 0, 2, 3, 4, 6, 7, 4, 4, 5, 5, 2, 3, 5, 5, 7, 3, 1, 4, 2, 0, 1, -3, -3, 0, -1, 0, 2, 0, 0, -1, -3, -1, 0, 0, 4, 5, 5, 6, 3, 5, 6, 5, 4, 4, 6, 5, 6, 5, 1, 3, 4, 1, 0, -3, 0, 0, 0, 0, 4, 1, 0, 0, -2, 0, 1, 1, 3, 3, 4, 5, 5, 5, 7, 5, 5, 4, 4, 6, 8, 5, 2, 3, 5, 3, 1, -3, -1, 0, -2, -1, 3, 2, 1, 0, -1, 1, 0, 2, 2, 3, 5, 5, 5, 6, 8, 5, 3, 5, 4, 5, 9, 6, 3, 2, 4, 2, 2, -1, -2, 1, 0, -3, 3, 3, 2, -1, 0, 1, 2, 3, 3, 4, 4, 3, 5, 6, 9, 5, 4, 5, 6, 3, 7, 5, 2, 2, 3, 3, 2, -1, -2, 0, -1, -3, 2, 3, 3, 0, 0, 0, 1, 3, 4, 3, 5, 4, 5, 8, 9, 3, 1, 1, 3, 6, 6, 2, 2, 4, 4, 4, 2, -1, -4, 0, 0, -2, 2, 3, 1, 1, 1, 0, 0, 1, 4, 5, 7, 6, 6, 8, 6, 2, 0, 0, 1, 5, 6, 1, 2, 4, 6, 5, 3, -2, -4, 0, 0, 0, 3, 2, 0, 1, 1, -1, 0, 0, 4, 6, 7, 8, 7, 9, 4, 2, 2, -1, 0, 5, 4, 3, 1, 3, 7, 5, 3, -1, -4, 0, 0, 1, 3, 0, -2, 0, 0, 0, 0, 0, 2, 5, 7, 7, 8, 10, 4, 0, 0, 0, -1, 2, 4, 2, 0, 3, 7, 7, 4, 0, -3, 1, 2, 3, 2, -2, -3, 0, 0, 0, 2, 3, 2, 6, 6, 5, 9, 10, 5, 2, 1, 1, -2, -1, 2, 4, 2, 3, 6, 7, 4, -1, -5, 0, 0, 3, 2, -2, -3, -1, 0, 1, 2, 2, 5, 7, 7, 5, 8, 10, 6, 2, 2, 3, -1, -1, 0, 2, 2, 3, 6, 6, 4, -1, -4, 0, 1, 3, 2, -1, -1, -1, 0, 0, 2, 2, 4, 6, 6, 5, 7, 8, 5, 3, 4, 3, 1, -2, 1, 2, 2, 2, 6, 6, 3, 0, -6, 0, 2, 3, 2, -1, 0, -1, 0, 0, 3, 3, 5, 7, 9, 4, 6, 5, 5, 4, 4, 5, 2, 0, 0, 2, 2, 3, 5, 5, 1, -2, -6, 0, 3, 3, 0, 0, 0, 1, 0, 0, 3, 4, 4, 4, 7, 5, 6, 5, 4, 3, 3, 6, 3, 1, 1, 2, 2, 3, 6, 4, 1, -2, -4, 0, 2, 2, 2, 0, 0, 0, 0, 0, 3, 4, 4, 4, 6, 5, 4, 5, 3, 2, 2, 7, 2, 2, 3, 0, 2, 4, 5, 3, 3, -3, -3, 0, 2, 0, 0, 0, 2, 1, 0, 0, 4, 5, 5, 4, 4, 7, 4, 5, 6, 1, 3, 6, 2, 2, 4, 0, 1, 4, 4, 4, 3, -3, -3, 0, 2, 1, 0, 0, 3, 1, -1, -1, 3, 3, 3, 4, 3, 7, 5, 5, 6, 3, 2, 5, 2, 3, 4, 2, 0, 4, 2, 1, 3, -3, -2, 0, 1, 0, 0, 1, 3, 2, 0, 0, 5, 3, 1, 1, 3, 7, 6, 5, 6, 2, 2, 2, 3, 3, 2, 2, 0, 4, 1, 0, 1, -2, -1, 0, 0, 0, 1, 1, 3, 2, 0, 0, 5, 2, 1, 1, 5, 8, 5, 4, 4, 0, 0, 3, 2, 2, 2, 1, 1, 4, 1, -1, 1, -2, -2, 0, 0, 0, 2, 3, 4, 2, 0, -1, 5, 4, 1, 2, 4, 7, 5, 4, 3, 0, 0, 0, 1, 3, 2, 3, 3, 3, 0, -1, 1, -4, -3, 0, 0, 0, 2, 3, 2, 2, -1, 0, 3, 3, 3, 2, 4, 7, 3, 2, 2, 1, 0, 1, 1, 1, 2, 4, 3, 3, 0, -3, 0, -4, -2, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 2, 4, 5, 7, 4, 0, 2, 3, 3, 1, 0, 2, 3, 3, 2, 0, -1, -3, -1, -3, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, 0, 4, 4, 6, 7, 3, 1, 3, 3, 4, 2, 1, 2, 1, 3, 2, 0, 0, -1, 0, -4, -1, 0, 0, 0, 1, -1, 0, 2, 1, 0, -2, 0, 4, 5, 5, 7, 2, 2, 2, 3, 3, 2, 1, 2, 1, 0, 1, 0, -1, -2, -1, -4, -2, 0, 0, 0, 1, -1, 0, 2, 2, 1, 0, 0, 3, 4, 5, 5, 2, 3, 4, 3, 3, 3, 2, 1, 1, 0, 0, 0, 0, -2, -2, -4, -2, 0, 0, -1, 2, 0, 0, 1, 3, 3, 0, 0, 3, 2, 3, 3, 1, 1, 2, 3, 1, 0, 1, 0, 0, -1, 0, 0, 0, -2, -2, -2, -2, 0, 0, 0, 2, 0, 0, 2, 3, 3, 2, 0, 2, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, -2, -1, -2, 0, 0, -2, -1, -1, -2, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, -1, -2, 0, -2, 0, -2, -1, 0, -1, -2, -2, -1, -1, -1, -1, 0, -1, 0, 0, -1, 0, -2, -3, -3, -2, -2, -2, -2, -1, -1, -1, 0, 1, 0, 2, 0, 2, 0, 1, 0, -1, -1, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, -3, -3, -3, -1, -1, -1, -1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 2, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, -2, -2, 0, 1, 0, 2, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 2, 2, 1, 0, 0, -1, -1, 0, -1, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 2, 1, 1, 2, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 2, 2, 3, 2, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 1, 0, -1, 0, 0, 2, 3, 3, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 2, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 3, 2, 3, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 3, 2, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, -2, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 3, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, -1, -2, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -2, -1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 2, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -2, -1, 0, 1, 0, 0, 2, 1, 0, 1, 1, 0, 0, 0, -1, -1, 0, -1, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 1, 2, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 2, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, -2, -2, -1, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -2, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 3, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 2, 0, 1, 2, 1, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -3, -2, -3, -1, -2, -2, -1, -2, -2, -2, -2, -3, -3, -4, -4, -4, -4, -2, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -1, -3, -1, -2, -1, -2, 0, 0, -1, -2, -2, -5, -5, -6, -4, -4, -3, -2, -3, -3, -3, -1, -1, -1, 0, 0, 0, 1, -1, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, -3, -3, -5, -4, -3, -2, -1, -1, 0, 0, -2, -2, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, -1, 0, -1, -1, -1, -1, -2, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 2, 0, 0, -1, -1, -1, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 1, 0, 0, 0, 1, 2, 2, 3, 2, 2, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 2, 2, 2, 1, 1, 2, 1, 2, 0, 1, 2, 4, 3, 2, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 2, 2, 3, 0, 1, 2, 2, 1, 1, 0, 3, 3, 3, 2, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, -2, 0, 0, 0, -1, 0, 0, 3, 3, 2, 2, 1, 0, 1, 2, 1, 2, 2, 2, 2, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 2, 3, 2, 0, 1, 1, 0, 1, 1, 2, 3, 2, 1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 3, 2, 1, 1, 0, 0, 0, 1, 2, 2, 1, 1, 1, 2, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, -1, -1, 0, 2, 4, 4, 4, 2, 2, 1, 1, 0, 0, 1, 2, 2, 2, 0, 0, 1, 1, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 1, 3, 4, 4, 4, 2, 1, 0, 0, 0, 0, 0, 3, 1, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, -1, -2, -2, 0, 0, 0, 0, 1, 2, 3, 4, 4, 3, 2, 0, 0, -1, -1, 0, 0, 2, 2, 1, 1, 2, 2, 0, -1, 0, -2, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 2, 3, 4, 3, 1, -1, 0, 0, 0, 0, 0, 2, 1, 1, 2, 2, 0, -1, -2, -1, -2, 0, 0, -1, -1, 0, 1, 0, 2, 0, 2, 3, 4, 3, 4, 3, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, -1, -1, -1, -2, 0, 0, -2, 0, 0, 1, 1, 2, 2, 2, 4, 2, 3, 3, 3, 1, 0, -1, 0, 0, 1, 1, 1, 1, 2, 2, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 3, 1, 2, 2, 3, 3, 4, 3, 2, 0, 0, 1, 1, 1, 2, 2, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 1, 1, 1, 3, 1, 2, 1, 3, 4, 4, 3, 3, 0, 0, 0, 0, 1, 1, 1, 1, 2, 2, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 1, 0, 0, 0, 2, 1, 1, 2, 2, 3, 5, 2, 0, 1, 3, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 2, 2, 2, 3, 2, 0, 1, 2, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 1, 1, 1, 0, 0, 1, 0, 3, 3, 1, 1, 2, 1, 0, 0, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 1, 3, 2, 1, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 2, 0, 1, 1, 1, 2, 1, 1, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 2, 1, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 2, 1, 1, 2, 2, 2, 1, 0, 0, 0, 0, -1, -1, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 2, 1, 0, 0, 0, 0, 0, -1, -2, -2, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -2, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, -2, 0, 0, 0, -1, 0, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 1, 1, 3, 2, 4, 4, 3, 2, 1, 0, -1, 0, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 2, 2, 1, 1, 1, 3, 2, 2, 3, 4, 2, 0, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 1, 2, 0, -1, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -2, -1, -2, -2, -1, -1, 0, -1, -2, -1, -1, -1, 1, 2, 3, 0, -1, -2, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, -3, -3, -2, -2, -1, -1, -1, 0, -2, -1, 0, 1, 2, 0, 0, -1, -1, -2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 1, 0, -1, -2, -2, -1, -1, 0, 0, 0, -1, 0, 0, 1, 2, 0, 0, -1, 0, -1, -1, 0, -1, 0, -2, -2, -2, 0, 1, 1, 1, 1, 2, 1, 0, -1, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, 2, 0, -1, -1, 0, 0, -1, 0, 0, -1, -3, -2, -2, -1, 0, 2, 2, 1, 2, 0, 0, -1, -1, -4, -3, -3, -3, -2, -1, -2, 0, 0, 0, 0, -1, 0, 1, 1, 0, -1, 0, -1, -3, -3, -4, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -4, -3, -3, -2, -1, -2, -2, -1, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, -2, -2, -3, -1, 0, 1, 0, 1, 1, 1, 0, 0, 0, -2, -2, -2, -2, -1, -2, -2, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, 0, 0, 0, 1, 2, 1, 2, 1, 0, 0, -1, -2, -1, -1, -3, -2, -1, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, 0, 1, 0, 1, 2, 3, 2, 1, 0, 0, -1, -3, -3, -3, -2, -2, 0, 1, 0, 0, -2, -1, -1, 0, 0, 1, 1, 0, -1, -2, -2, 0, 0, 2, 1, 0, 2, 3, 1, 1, 0, 0, -1, -3, -3, -4, -2, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -2, 0, 0, 0, 1, 2, 1, 1, 3, 2, 0, 0, -1, -2, -2, -3, -4, -4, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -2, -2, -1, 0, 0, 0, 2, 0, 1, 2, 2, 0, -1, 0, 0, -2, -3, -4, -3, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 0, 0, -1, -2, -2, -2, -3, -2, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 2, 1, 1, 1, 0, 0, -2, -3, -5, -3, -2, -1, 1, 0, 0, 0, 0, 0, 2, 2, 1, 1, 0, 0, -1, 0, 0, 1, 0, 2, 2, 1, 1, 1, 2, 1, 0, -1, -4, -5, -5, -3, -2, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 2, 1, 0, -1, -1, -3, -3, -4, -3, -1, 0, 1, 0, 0, -1, 0, 0, 0, 2, 1, 0, 0, 0, 0, -1, 0, 1, 0, 2, 0, 1, 0, 1, 0, -1, -2, -2, -2, -3, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -2, -2, -1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 1, -1, -1, -3, -3, -2, -2, 0, -1, 0, 1, 0, 0, 0, 0, 1, 1, 1, -1, -2, -3, -2, -2, -2, 0, 0, 0, 1, 0, 2, 1, 0, 0, -1, -2, -4, -3, -2, -2, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 1, -1, -1, -1, -2, -1, -2, 0, 0, 1, 1, 2, 2, 0, 0, 0, -2, -3, -3, -4, -3, -2, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, -2, -1, -2, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -2, -3, -3, -2, -3, -2, 0, 0, 0, 1, 0, -1, -1, -1, 0, -1, -1, -1, -1, -2, -2, 0, 0, 0, 0, 1, 1, 1, 0, -2, -1, -1, -3, -3, -3, -3, -1, -1, 0, 0, 0, 2, 0, 0, -1, -2, 0, -1, 0, -1, -2, -1, 0, 0, -1, 0, 1, 1, 1, 0, -1, -2, -3, -3, -1, -2, -2, -2, -2, -1, 0, 0, 0, 2, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, 0, -1, -1, -2, -1, -2, -2, -3, -2, -4, -3, -1, 0, 0, 1, 0, -1, -2, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, -1, -2, -2, -1, -1, -1, -2, -1, -1, -1, 0, 2, 1, 3, -1, -2, -2, -2, -1, 0, 0, -2, -1, -2, -1, -1, -2, -3, -2, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 2, 2, 2, 3, 3, 0, -2, -3, -2, -1, -2, -2, -3, -2, -2, -2, -2, -2, -3, -1, -2, -1, 0, 0, 1, 2, 3, 3, 4, 4, 5, 4, 4, 4, 4, 2, 3, 0, -1, -3, -2, -3, -1, -1, 0, -1, -2, -2, -1, -2, -1, -1, -1, 0, 0, 1, 2, 1, 2, 4, 3, 4, 3, 4, 3, 3, 2, 1, 2, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, -2, -1, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 2, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 2, 1, 0, 1, 1, 0, -1, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, 0, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, -1, -1, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, -2, 0, -2, -2, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 1, -1, 0, -1, -2, 0, -1, -3, 1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, -1, 0, 0, 1, 0, -1, 0, -1, 0, 1, 0, 1, 0, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 1, 1, 3, 2, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 1, 0, 0, 1, 2, 0, 2, 0, 2, 3, 2, 1, 1, 3, 2, 1, 0, 1, 1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 3, 1, 2, 3, 2, 1, 2, 3, 3, 2, 3, 1, 2, 2, 0, 0, 2, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 2, 2, 3, 3, 4, 2, 1, 2, 3, 4, 3, 2, 1, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 3, 3, 2, 3, 4, 4, 2, 2, 2, 2, 3, 2, 2, 1, 1, 2, 1, 0, 0, 0, -1, -1, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 3, 4, 2, 1, 3, 1, 1, 2, 2, 2, 2, 1, 1, 1, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 3, 3, 1, 4, 3, 2, 1, 3, 0, 0, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, -2, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 2, 2, 3, 3, 2, 2, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 1, 2, 2, 3, 2, 1, 0, 0, 1, 1, 1, 0, 1, 2, 1, -1, 0, 0, 0, -2, -1, 0, -1, 0, 1, 0, -1, -1, 0, 1, 1, 2, 2, 2, 5, 3, 3, 2, 0, 1, 0, 0, 0, 2, 1, 2, 2, 0, 1, 0, 0, -1, -1, 0, 0, 0, 1, 0, -1, -1, 0, 0, 1, 2, 1, 4, 6, 3, 2, 3, 1, 0, 0, 0, 0, 2, 2, 2, 2, 1, 0, 0, 0, -2, -2, 0, -1, 0, 1, 0, 0, -1, 1, 2, 1, 1, 2, 4, 6, 4, 3, 3, 2, 0, 0, 1, 1, 1, 2, 1, 0, 1, 0, -1, 0, -1, -2, 0, 0, 0, 1, 0, 0, 0, 0, 2, 1, 1, 0, 3, 4, 4, 3, 3, 2, 0, 0, 1, 0, 0, 1, 1, 2, 2, 0, -1, 0, -2, -2, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 1, 0, 0, 4, 5, 3, 3, 1, 0, 0, 2, 1, 0, 1, 1, 1, 1, 1, 0, 0, -1, -2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 2, 4, 4, 2, 4, 3, 0, 0, 2, 1, 1, 1, 1, 0, 1, 1, 0, 0, -2, -1, 1, 0, 1, -1, 0, 0, 0, 2, 1, 0, 2, 2, 2, 4, 4, 4, 5, 3, 0, 2, 2, 1, 1, 2, 1, 1, 1, 2, 0, -1, -1, -2, 1, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 1, 3, 5, 3, 4, 5, 3, 1, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, -1, 0, 0, 0, 2, 1, 0, 2, 1, 3, 5, 4, 5, 5, 3, 0, 1, 1, 1, 2, 2, 0, 0, 0, 1, 0, 0, -1, -1, 1, 0, 0, -1, -2, 0, 0, 2, 2, 2, 2, 3, 3, 5, 3, 4, 3, 1, 1, 2, 1, 1, 2, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 2, 2, 2, 2, 2, 4, 2, 3, 3, 1, 2, 0, 1, 1, 1, 1, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 3, 2, 2, 3, 3, 3, 3, 3, 2, 1, 0, 1, 2, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 3, 2, 3, 3, 2, 2, 2, 2, 2, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, -1, -1, 0, 1, 1, 4, 2, 3, 3, 3, 2, 1, 2, 3, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, 0, -1, -1, 0, 1, 2, 2, 2, 2, 3, 3, 1, 2, 2, 3, 1, 1, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, -2, 1, 0, 0, 0, -1, 0, -1, 1, 2, 1, 1, 2, 2, 2, 2, 2, 1, 2, 1, 1, 2, 0, -1, -2, -1, 1, 1, 1, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 2, 1, 1, 2, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, -2, -2, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, -1, -2, -2, -2, -1, 0, -1, 0, -3, -1, -2, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, -1, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 2, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 2, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 2, 2, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 2, 3, 2, 1, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 2, 2, 2, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 2, 2, 1, 0, -1, 0, 0, 2, 1, 0, 0, 1, 1, 0, 0, 0, -1, 1, 0, 0, 1, 2, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 2, 1, 1, -1, 0, 0, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 1, 2, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, -1, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 2, 2, 0, 0, 0, 0, 0, -1, -1, -1, -1, -3, -2, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 1, 1, 1, 1, 0, 0, -2, -4, -4, -3, -3, -1, -2, -2, -1, -1, 0, 2, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 1, 2, 2, 2, 1, 1, 0, 0, 0, -2, -3, -3, -3, -2, -2, -2, 0, -1, 0, 1, 2, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 2, 3, 3, 3, 2, 0, 1, 0, 1, 0, 0, -2, -1, -1, -1, -1, -2, -2, 0, 1, 2, 2, 1, 0, 0, 0, -1, -1, -2, 0, 1, 2, 3, 3, 4, 3, 2, 1, 1, 1, 0, 2, 1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 2, 2, 0, 0, 0, -1, -2, -2, -3, -1, 0, 0, 1, 4, 4, 4, 3, 3, 2, 2, 2, 1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 2, 1, 1, -1, 0, -2, -2, -3, -3, -2, -3, -1, 1, 2, 4, 4, 3, 3, 2, 1, 0, 0, -1, -1, -2, -1, -2, -1, -2, -1, 0, 2, 2, 1, 0, 0, 0, 0, -3, -2, -3, -3, -3, -2, 0, 2, 3, 4, 2, 1, 1, 0, 0, 0, -2, -2, -2, -1, -3, -3, -2, -2, 0, 0, 1, 2, 0, 0, -1, -1, -2, -5, -4, -4, -3, -3, -1, 0, 2, 2, 2, 1, 1, 0, 0, -1, -1, -1, -1, -1, -2, -3, -3, -1, 0, 2, 2, 1, -1, -2, -1, -2, -4, -4, -5, -4, -5, -3, 0, 1, 3, 2, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, -3, -3, -2, 0, -1, 1, 2, 0, -1, -1, -2, -2, -5, -6, -6, -7, -4, -3, -1, 1, 3, 3, 2, 2, 1, 1, 1, 2, 0, 0, -1, -1, -2, -3, -2, -2, 0, 1, 0, -1, -2, -2, -3, -2, -4, -6, -6, -6, -5, -3, 0, 1, 4, 3, 3, 3, 2, 2, 1, 1, 0, -1, -1, -2, -1, -2, -2, -2, 0, 1, 0, -1, -3, -2, -3, -4, -6, -6, -7, -8, -6, -2, 0, 3, 4, 2, 2, 1, 2, 1, 0, 1, 0, 0, 0, 0, -2, -1, -3, -1, -1, 0, 0, -1, -2, -2, -2, -3, -6, -8, -8, -6, -5, -4, -1, 1, 3, 4, 3, 1, 2, 2, 1, 1, 0, -1, -2, 0, -2, -2, -1, -3, 0, 0, 1, 0, -1, -2, -4, -5, -6, -6, -7, -5, -5, -4, -1, 1, 3, 3, 1, 2, 2, 1, 2, 2, 1, -1, -1, -2, -1, -1, -1, -2, -1, 0, 1, 0, -1, -2, -4, -3, -5, -5, -6, -5, -4, -3, 0, 0, 3, 2, 1, 2, 3, 1, 3, 2, 1, -1, -3, -2, -1, -2, -2, -1, -1, 1, 0, 0, 0, -2, -2, -4, -5, -5, -5, -5, -4, -2, -1, 1, 3, 3, 2, 3, 3, 3, 4, 3, 0, -1, -2, -2, -1, -1, -1, -2, -1, 0, 1, 0, 0, -2, -3, -2, -5, -5, -4, -3, -3, -1, -1, 1, 3, 3, 2, 4, 4, 4, 4, 2, 0, 0, -2, -2, 0, -2, -2, -1, -1, 0, 1, 0, 0, -1, -2, -3, -4, -3, -2, -3, -2, -1, 0, 2, 3, 3, 3, 3, 3, 3, 3, 2, 0, -1, -2, -1, -1, -1, -1, -2, -2, 1, 0, 1, 0, -1, -1, -3, -3, -4, -2, -2, 0, 0, 0, 3, 4, 3, 2, 3, 3, 2, 3, 1, 0, 0, -2, -2, -2, 0, -1, -1, -1, 0, 2, 0, 0, 0, -1, -2, -4, -4, -3, -1, 0, 1, 2, 3, 5, 4, 4, 2, 2, 0, 2, 0, -2, 0, -2, -1, -2, -1, -1, -2, -1, 1, 0, 0, 0, 0, -2, -3, -2, -4, -1, -1, 0, 1, 3, 2, 3, 3, 2, 2, 1, 1, 0, 0, -1, -1, -1, -2, -3, -2, 0, -1, 0, 1, 0, 0, -1, -1, -2, -3, -3, -3, -1, 0, 0, 1, 2, 3, 3, 2, 2, 3, 1, 2, 0, 0, 0, -3, -2, -3, -2, -1, -1, -1, 0, 0, 1, 0, 0, -1, -1, -1, -3, -3, 0, 0, 0, 2, 3, 2, 2, 2, 1, 0, 1, 1, 1, 0, -2, -3, -3, -1, -1, -1, -1, 0, -1, 0, 0, 0, -1, -1, -2, -1, -2, -1, 0, 1, 3, 2, 3, 1, 1, 2, 2, 0, 1, 0, 0, -1, -2, -1, -3, -1, -1, -1, 0, 0, 0, 1, 1, 1, 0, -1, 0, -1, -1, -1, 1, 1, 2, 2, 2, 2, 2, 2, 1, 1, 0, 0, 0, -2, -2, -3, -2, -3, -2, 0, 0, 0, -1, 1, 1, 2, 1, -1, 1, 0, 0, 1, 0, 2, 3, 2, 2, 2, 1, 1, 1, 0, 0, -1, -2, -3, -4, -2, -4, -3, -3, -1, -1, -1, -1, 0, 1, 1, 1, 1, 2, 0, 2, 1, 1, 2, 3, 1, 1, 2, 0, 0, 0, 0, -2, -2, -2, -3, -3, -4, -4, -4, -2, -2, -1, -1, 0, -1, 0, 0, 1, 0, 1, 1, 2, 2, 2, 1, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, 0, -2, -2, -2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -2, -1, 0, -1, -1, -1, 0, 0, 1, 1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, -2, 0, -1, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 1, 1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, -1, -2, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, -1, -1, 0, 1, 0, 0, 1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -2, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, -2, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, -2, -1, 0, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -2, -2, -1, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 2, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 2, 2, 1, 0, 2, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, -1, 1, 1, 0, 1, 1, 1, 1, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 1, 0, 2, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 2, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, -1, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -2, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, -1, 0, 1, 1, 1, 0, 1, 1, 1, 1, 1, 0, 0, -1, -2, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, -1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, -2, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, -1, -1, -1, -1, -3, -2, -1, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -3, -1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, -2, -2, -1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, -1, -2, -2, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, -1, -2, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, -1, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, -2, -1, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -2, -1, 0, -1, -1, 0, 0, 1, 0, 1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -2, -1, -1, -1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 2, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 2, 2, 2, 1, 2, 1, 2, 3, 3, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 1, 0, 1, 1, 1, 1, 1, 2, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 2, 2, 3, 4, 4, 4, 4, 2, 4, 5, 5, 6, 5, 5, 4, 3, 3, 1, 0, 1, 1, 1, 1, 2, 0, 0, -2, -3, -3, 0, -1, 0, 2, 3, 5, 5, 4, 5, 4, 5, 5, 7, 8, 6, 6, 6, 5, 4, 2, 1, -1, 0, 2, 1, 3, 4, 2, 0, 1, -3, -2, -1, 0, 0, 1, 3, 3, 4, 4, 2, 1, 3, 4, 6, 7, 7, 5, 3, 3, 3, 1, 0, -1, -2, -1, 0, 0, 2, 4, 5, 4, 1, 0, 0, 0, 0, 2, 3, 3, 3, 2, 1, 0, 3, 3, 6, 5, 5, 4, 1, 0, 0, -1, -1, -3, -2, -3, -2, -2, 0, 0, 3, 4, 3, 1, 1, 0, 1, 3, 2, 3, 4, 2, 0, 0, 3, 5, 7, 6, 5, 4, -2, -3, -2, -2, -3, -2, -3, 0, -2, -3, -3, -2, 1, 3, 1, 0, 0, 1, 1, 2, 1, 3, 3, 2, 2, 1, 3, 8, 9, 6, 5, 4, -1, -5, -4, -4, -3, -3, 0, 1, 1, -1, -1, -1, 0, 2, 0, 1, 0, 1, 1, 1, 0, 2, 3, 2, 2, 3, 5, 8, 9, 7, 5, 2, -1, -4, -5, -3, -4, -5, -2, 1, 2, 1, -1, 0, 1, 0, 0, 0, 1, 1, 1, 1, 1, 2, 2, 2, 2, 2, 4, 7, 7, 5, 6, 2, -2, -4, -3, -4, -4, -4, -2, 0, 3, 4, 0, 0, 2, 1, 1, 1, 1, 2, 2, 1, 3, 4, 3, 2, 2, 2, 3, 4, 4, 4, 5, 2, -1, -4, -5, -5, -6, -5, -2, 0, 3, 4, 1, 0, 2, 4, 2, 2, 1, 2, 2, 3, 4, 5, 3, 2, 1, 1, 3, 3, 5, 4, 4, 1, 0, -2, -4, -5, -6, -7, -3, 0, 2, 3, 0, 0, 0, 3, 4, 4, 1, 1, 1, 2, 4, 7, 5, 2, 1, 1, 3, 3, 3, 3, 4, 2, 1, -1, -5, -5, -7, -8, -5, -2, -1, 1, 0, -3, 0, 3, 5, 4, 3, 0, 2, 4, 6, 6, 6, 2, 0, 0, 3, 2, 2, 4, 4, 2, 2, -2, -6, -5, -6, -8, -6, -5, -4, -1, -3, -3, -1, 2, 4, 4, 2, 0, 1, 2, 5, 6, 5, 0, 0, 1, 4, 5, 2, 3, 3, 3, 1, -3, -5, -6, -5, -7, -6, -4, -4, -3, -5, -4, -2, 1, 3, 4, 1, 0, 0, 1, 3, 5, 3, 0, 0, 1, 2, 3, 4, 4, 4, 4, 1, -4, -6, -6, -5, -6, -7, -6, -5, -5, -6, -6, -2, -2, 1, 4, 2, -1, 0, 1, 1, 5, 2, -1, -1, 0, 1, 2, 4, 3, 4, 5, 0, -4, -6, -5, -5, -5, -8, -6, -7, -8, -7, -7, -3, -3, 0, 2, 2, 0, 0, 0, 1, 3, 3, 0, -1, 0, 0, 1, 4, 3, 3, 5, 2, -4, -7, -6, -5, -4, -6, -7, -7, -9, -6, -4, -2, -2, 0, 3, 2, 0, 1, 1, 2, 3, 2, 0, -1, 0, 0, 0, 2, 1, 1, 2, 1, -3, -5, -7, -7, -6, -6, -7, -7, -9, -7, -4, -2, -3, 0, 2, 1, 0, 2, 2, 1, 1, 3, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, -3, -5, -7, -7, -6, -5, -6, -6, -9, -7, -5, -2, -1, 0, 2, 1, 1, 3, 4, 1, 0, 0, 2, 1, 1, 0, 0, -1, 0, 0, 0, 0, -2, -4, -7, -7, -6, -4, -4, -6, -8, -5, -4, -2, -1, 0, 1, 2, 0, 1, 3, 2, 0, 0, 2, 3, 2, 0, 0, 0, 0, 1, 0, -1, -3, -3, -6, -5, -5, -3, -2, -4, -5, -3, -4, -2, -1, 0, 0, 0, 0, 1, 2, 2, 1, 2, 2, 2, 2, 1, 0, 1, 1, 1, 1, 0, -2, -3, -4, -5, -5, -3, -2, -4, -3, -1, -2, -3, 0, 1, 1, 0, 0, 1, 1, 3, 3, 2, 3, 3, 3, 3, 0, 2, 2, 3, 0, -2, -4, -3, -4, -5, -6, -5, -4, -3, -1, -1, 0, 0, 1, 1, 0, 0, 1, 0, 3, 2, 4, 2, 2, 3, 3, 4, 2, 2, 4, 4, 1, -2, -3, -5, -5, -7, -5, -7, -4, -3, -2, 0, 0, 0, 1, 2, 1, 0, 0, 0, 2, 3, 3, 4, 3, 2, 4, 5, 4, 5, 3, 2, 2, -1, -3, -3, -5, -6, -6, -6, -5, -4, -1, -1, 0, 0, 1, 1, 1, 0, -1, 0, 0, 2, 3, 2, 2, 2, 4, 6, 5, 3, 2, 3, 0, -1, -4, -6, -6, -5, -6, -5, -6, -3, -2, -3, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 5, 4, 6, 6, 4, 2, 0, -2, -5, -7, -6, -4, -5, -6, -4, -4, -4, -1, 1, 0, 2, 2, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 3, 5, 5, 7, 5, 5, 1, -1, -5, -6, -6, -4, -3, -4, -5, -3, -2, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, -1, -2, 0, -1, 0, 3, 4, 6, 9, 9, 6, 4, 0, -4, -7, -7, -5, -4, -4, -5, -3, -3, 0, 1, 1, 0, -1, -2, -1, 0, 0, 0, -1, 0, -1, 0, 1, 3, 3, 5, 8, 9, 9, 5, 2, -1, -6, -7, -5, -7, -5, -6, -4, -4, -3, -2, 0, -1, -3, -4, -1, 0, 1, 0, 1, 0, 1, 1, 2, 3, 4, 5, 8, 9, 11, 10, 5, 3, -1, -5, -4, -6, -6, -8, -4, -6, -6, -4, -4, -4, -5, -3, -1, 0, 1, 0, 0, 0, 2, 2, 4, 3, 2, 5, 6, 10, 11, 9, 7, 4, 1, -1, -2, -4, -5, -6, -5, -3, -4, -4, -4, -4, -5, -5, -3, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 2, 3, 4, 5, 5, 5, 2, 2, 0, 0, 0, -3, -3, -1, -2, -1, -3, -2, -1, -3, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, -1, -2, -1, -3, -2, -1, -2, -1, 0, 2, 2, 3, 2, 1, 3, 1, 2, 0, 0, -1, -1, 0, 0, 1, 1, 1, 2, 2, 2, 0, 0, -2, -4, -4, -5, -4, -4, -3, -2, -1, -2, 0, 1, 2, 4, 1, 2, 2, 2, -1, -1, -1, -2, -1, 0, 1, 1, 1, 1, 3, 3, 2, 0, -2, -4, -5, -5, -4, -4, -3, -2, -3, -3, -1, 1, 2, 1, 2, 2, 2, 1, 0, 0, 0, -1, 0, 0, 1, 2, 2, 1, 3, 1, 2, 0, -2, -3, -3, -2, -2, -3, -3, -2, -3, -2, -1, 0, 0, 0, 1, 2, 1, 3, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 2, 1, 1, 0, 0, -1, 0, -1, -1, -3, -3, -2, -2, -2, -1, 0, 0, 0, 0, 1, 3, 3, 0, 1, 1, 0, 0, 0, 1, 2, 1, 0, 1, 2, 2, 1, 1, 1, 2, 2, 0, -2, -2, -1, -2, -1, 0, 0, 1, 0, 0, 2, 4, 4, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 3, 3, 3, 2, 2, 1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 3, 0, 1, 3, 2, 0, 0, 0, 0, -2, -3, -3, -2, 1, 3, 3, 6, 6, 4, 2, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 3, 3, 0, 3, 5, 3, 2, 0, 0, -1, -4, -4, -4, -3, 0, 2, 3, 7, 6, 5, 2, 0, -2, -1, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 3, 6, 6, 3, 0, 0, -1, -3, -4, -5, -3, 0, 1, 3, 4, 5, 4, 0, -1, -2, -2, -1, -2, -2, 0, 0, 0, 0, 1, 1, 1, 1, 3, 6, 5, 4, 1, -1, -1, -2, -3, -3, -3, -2, 1, 2, 4, 4, 3, 2, 0, -1, -1, -1, -2, -1, 0, 0, 0, -1, 0, 0, 0, 1, 3, 4, 3, 2, 0, -1, -1, -2, -2, -2, -1, 0, 1, 3, 4, 5, 4, 2, 1, 0, 0, 0, -1, -1, -2, -1, -1, -1, -1, 0, 1, 0, 3, 4, 3, 0, 0, -1, -1, -1, -2, -3, 0, 2, 3, 4, 3, 6, 4, 5, 3, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 1, 1, 0, -1, -2, -2, 0, 0, -3, -2, 0, 3, 5, 6, 7, 5, 4, 4, 2, 0, 0, -1, -1, -1, -2, -1, -1, -2, 0, 0, 0, 0, 0, 0, -2, -3, -2, -1, 0, -1, -2, -1, 0, 2, 5, 5, 8, 6, 5, 4, 1, 0, -2, -1, 0, -2, -2, 0, -1, -1, -1, 0, 0, 0, -1, -1, -3, -3, -3, -1, -1, -3, -3, -2, 0, 1, 4, 5, 6, 5, 5, 2, 1, 0, -1, -2, -2, -2, -1, 0, -1, -1, 0, 0, 0, 0, -1, -3, -3, -2, -1, -3, -2, -4, -2, -2, 0, 0, 4, 4, 4, 5, 4, 3, 0, 0, -1, -2, 0, -1, -1, -2, -3, -2, 0, 0, 0, 0, -1, -2, -2, -1, 0, -2, -3, -3, -2, -1, 0, 1, 2, 3, 4, 5, 3, 2, 1, 2, -1, -1, 0, -1, -2, -2, -3, -1, 0, 0, 1, 0, -1, -2, -2, 0, 0, -2, -2, -3, -1, 0, 0, 0, 3, 4, 5, 5, 4, 3, 3, 2, 0, 0, -1, -1, -3, -3, -2, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -3, -3, -2, -1, -1, 0, 2, 2, 4, 4, 2, 0, 1, 1, 0, 0, 0, -3, -2, -3, -1, -1, 0, 1, 1, 0, 0, 0, 1, 0, 1, -2, -3, -2, -2, -2, 0, 0, 0, 2, 2, 3, 1, 0, 0, 0, 0, 0, 0, -2, -1, -2, -1, -1, 0, 2, 2, 0, 0, 0, 1, 1, 2, 0, -4, -5, -4, -3, -2, 0, 0, 2, 3, 3, 2, 1, 2, 0, 0, 0, 0, -2, 0, -1, 0, 0, 1, 2, 3, 1, 2, 2, 1, 1, 1, 0, -4, -4, -5, -5, -2, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, -1, -1, -2, 0, 0, 1, 1, 1, 3, 1, 1, 2, 2, 2, 1, 1, -1, -3, -4, -6, -5, -2, 0, 1, 0, 0, 0, 1, 2, 2, 0, -1, -1, -1, -1, 0, 1, 2, 2, 2, 3, 2, 2, 3, 3, 1, 0, -1, -2, -3, -4, -5, -4, -2, 0, 2, 1, 1, 1, 1, 0, 1, -2, -1, -1, -3, -2, 0, 2, 2, 2, 3, 4, 3, 1, 2, 2, 1, -1, -1, -1, -3, -3, -3, -1, 0, 2, 2, 2, 1, 2, 2, 0, -1, -2, -2, -3, -3, -2, -1, 1, 0, 2, 2, 4, 1, 1, 1, 2, 1, 0, 0, -1, -2, -1, 0, 0, 2, 2, 2, 3, 3, 3, 1, 0, -1, -4, -5, -5, -3, -3, -2, -1, -1, 0, 2, 2, 3, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 3, 3, 3, 2, 2, 0, 0, 1, 0, -3, -5, -6, -4, -3, -4, -2, -3, -3, -1, 0, 2, 1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 2, 4, 3, 3, 0, 0, -1, 0, 0, -3, -4, -5, -4, -3, -2, -3, -3, -2, -2, 0, 2, 3, 2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 2, 4, 2, 0, 0, -2, -3, -1, -1, -3, -3, -4, -1, 0, -1, -1, -2, -2, 0, 1, 2, 4, 3, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 3, 2, 0, 0, -3, -2, -2, -2, -2, -2, -1, 0, 1, 1, 0, 1, 1, 1, 2, 4, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, -3, -2, -3, -2, -3, -2, -1, 0, 0, 0, 2, 2, 2, 1, 1, 0, 0, 0, -2, -1, 0, 0, 0, 1, 1, 1, 1, 1, 1, -1, -3, -4, -4, -5, -4, -3, -2, -3, -3, -2, 0, 0, 0, 2, 1, 0, 1, 1, -1, -1, -2, -2, -1, 0, 1, 0, 1, 1, 1, 0, 1, 0, -3, -3, -3, -4, -3, -2, -3, -2, -2, -2, -1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, -2, -1, 1, 2, 1, 0, 1, 1, 1, 0, -3, -3, -2, -1, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 3, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -2, -1, -1, 1, 0, 2, 3, 2, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 1, 2, 2, 1, 2, 1, 2, 0, 0, 0, -1, -1, -3, -3, -1, 0, 1, 2, 3, 4, 2, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 3, 3, 4, 2, 1, 0, -1, -3, -4, -3, -1, -1, 2, 2, 4, 3, 1, 1, -1, -1, -1, -2, -2, -1, 0, -1, 0, 0, 0, 0, 1, 1, 2, 4, 3, 1, 0, 0, 0, -2, -2, -3, -3, -1, 0, 1, 3, 2, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 3, 3, 1, 0, 0, -1, -2, 0, -1, -2, -1, 1, 1, 3, 2, 0, 1, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 4, 4, 2, 2, 0, 0, -1, 0, -1, -1, 0, 2, 1, 2, 0, 0, 2, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 3, 1, 1, 0, -1, -1, 0, 0, -1, 0, 1, 2, 3, 2, 2, 2, 2, 1, 1, 0, 0, 0, 0, -2, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, -2, -2, -2, -1, 0, 0, 0, 0, 2, 2, 3, 6, 5, 3, 2, 3, 0, -1, 0, 0, -1, -1, -1, 0, 0, -2, -1, 0, 0, 0, 0, -2, -1, -2, -3, -1, 0, 0, -1, 0, 1, 2, 2, 4, 4, 3, 3, 2, 0, 0, -1, -2, -2, -2, 0, 0, 0, -1, 0, -1, 0, 0, 0, -2, -3, -3, -2, -1, -1, 0, -1, 0, 0, 2, 1, 4, 3, 3, 2, 1, 1, 0, -1, -2, -2, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, -2, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, 2, 3, 2, 3, 2, 0, 1, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, -1, -2, -1, -1, 0, 0, 1, 1, 2, 2, 2, 1, 1, 1, 0, 0, -1, 0, 0, -1, -1, -2, -1, 0, 0, 1, 0, 0, -2, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 4, 1, 2, 0, 0, 1, 0, 0, 0, 0, -2, -2, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 1, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 2, 1, -1, 0, -1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 2, 2, 0, -1, -1, -4, -2, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 1, 0, 2, 1, 1, 0, 1, 2, 0, 1, 0, -1, -2, -3, -3, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -2, 0, 0, 1, 1, 1, 1, 2, 1, 0, 2, 1, 1, 0, 0, -1, -1, -3, -4, -2, -2, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 2, 3, 0, 0, 2, 1, 1, -1, -1, -2, -2, -1, -3, -1, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, -2, -2, -2, -2, 0, 0, 1, 1, 1, 2, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, -2, 0, 1, 2, 2, 0, 0, 1, 2, 0, -1, -3, -3, -3, -1, -2, -1, 0, 0, 0, 1, 1, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 2, 3, 2, 3, 0, 0, 2, 0, 0, -2, -3, -3, -3, -2, -2, -1, -2, -1, 0, 0, 2, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 2, 3, 3, 2, 2, 1, 0, 1, 0, -1, -2, -4, -3, -2, -2, -1, -2, -2, -2, 0, 0, 2, 1, 0, 0, 1, 1, 1, 0, 0, 1, 1, 2, 3, 3, 3, 1, 0, -1, 0, -1, -1, -2, -2, -1, 0, 0, 0, -2, -2, -2, 0, 0, 2, 1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 3, 2, 0, 0, -2, 0, 0, 0, -1, -1, 0, -1, 0, 1, 0, 0, -1, 0, 1, 2, 3, 1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 2, 2, 0, 1, 2, 2, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 1, 0, 1, 1, 1, 2, 0, 0, 0, 0, -1, 0, -2, -2, -2, -2, -2, -2, -1, -2, -1, -3, -3, -2, -4, -2, -2, -1, 0, 1, 0, 2, 1, 1, 1, 0, 0, 0, 1, 1, 1, 0, -1, -1, 0, -1, -2, -2, -2, -1, 0, 0, 0, -1, -2, -1, -2, -2, -2, -2, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -2, 0, -1, -1, -2, -2, 0, 0, 1, 1, 0, 0, 1, 0, 0, -2, -2, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, 0, 0, 0, 1, 2, 2, 2, 0, -1, -1, -1, -1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 2, 2, 1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 0, 0, 1, 2, 2, 1, 0, -1, 0, 0, 0, 0, 1, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 1, 1, 2, 0, 1, 0, 0, -1, 0, -1, 0, 1, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 3, 3, 3, 2, 2, 1, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 4, 4, 2, 2, 2, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 3, 2, 0, 0, 3, 1, 1, -1, 0, 0, 0, 0, 1, 0, -1, -1, 0, -1, -1, -1, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 3, 3, 3, 1, 0, 2, 2, 2, 0, -1, 0, 1, 0, 0, 0, -1, -1, 0, 0, -1, -2, -2, -2, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 4, 4, 1, 1, 3, 2, 3, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, -1, -1, -1, -1, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 2, 3, 3, 2, 2, 3, 2, 0, -1, -1, 0, 1, 2, 1, 0, -1, 0, 0, -1, -2, -2, 0, 0, 0, -2, 0, 0, -1, -1, 0, 0, 1, 1, 1, 3, 2, 3, 3, 3, 1, -2, 0, 0, 1, 2, 0, 0, -1, 0, 1, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 3, 3, 2, 0, -2, 0, 0, 1, 1, 1, -1, 0, 0, 1, 0, -2, -2, 0, 1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 2, 3, 3, 2, 3, 1, 1, 0, 0, 0, 1, 3, 0, -1, -1, 0, -1, 0, -2, -1, -2, 0, 0, -1, 0, 0, -1, -1, 0, 1, 0, 1, 2, 3, 3, 3, 4, 3, 0, -1, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, -2, -1, 0, 0, 1, 1, 1, 3, 4, 5, 3, 1, 0, -1, 0, 0, 1, 2, 1, 0, 0, -1, -1, -1, -1, -1, -2, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 1, 2, 1, 2, 5, 4, 2, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 2, 3, 3, 3, 2, 3, 3, 3, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -1, -1, -1, 0, 1, 1, 0, 0, 2, 3, 2, 3, 3, 2, 2, 2, 1, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 2, 3, 3, 2, 3, 2, 3, 2, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 2, 3, 3, 2, 2, 2, 1, 1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 3, 4, 2, 0, 0, 0, -2, -2, -1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 2, 2, 3, 2, 2, 0, 0, 0, -2, 0, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, 0, 1, 2, 1, 2, 1, 0, -1, -2, -2, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 2, 1, 0, 1, 0, 0, 1, 3, 1, 0, 0, -1, -1, -1, -1, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 1, 0, 1, 0, 1, 1, 2, 0, 0, 0, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -2, -3, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -2, 0, -2, -2, -2, -2, -3, -4, -2, -2, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -3, -3, -4, -3, -2, -4, -5, -4, -5, -4, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -3, -2, -4, -3, -2, -3, -4, -2, -4, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 0, 0, -1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 2, 2, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 3, 3, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -2, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 1, 1, 3, 1, 0, 0, 0, -2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, -1, -1, -1, 0, 0, 1, 2, 2, 1, 1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, -1, 1, 1, 0, -1, 1, 0, 0, -1, 0, 0, -2, -1, 0, 0, 0, 1, 2, 3, 2, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 2, 2, 3, 1, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 3, 2, 3, 1, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 1, 2, 3, 1, 0, 0, 0, -1, -1, 0, -1, -2, -1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 1, 3, 3, 1, 0, 1, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 2, 2, 1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, 0, 0, 0, 2, 2, 2, 2, 1, 1, 1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 1, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 2, 0, 2, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, -2, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 2, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -3, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 2, 2, 1, 1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 1, 1, 1, 2, 1, 1, -1, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 2, 2, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 1, 0, 0, 2, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, 1, 2, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 0, -1, 0, 0, 2, 0, 0, -1, 0, 0, 0, -1, 0, 1, 3, 2, 3, 3, 2, 0, 0, 0, 1, 0, 0, 1, 3, 2, 0, 1, 1, 2, 0, 0, 0, 0, 2, 1, 1, 0, -1, 0, 0, 0, 0, 1, 2, 3, 2, 3, 3, 0, 0, 0, 0, 0, 1, 1, 3, 2, 1, 0, 1, 1, 2, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, 0, 1, 1, 2, 3, 3, 3, 0, 0, -1, 0, 0, 0, 1, 1, 2, 2, 1, 0, 2, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, -1, 0, 1, 2, 2, 3, 3, 3, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 2, 2, 2, 3, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 2, 0, 0, -1, 0, 1, 0, 0, 1, 0, -1, 0, 0, 1, 0, 1, 2, 2, 2, 1, 0, -1, -1, -1, -1, -1, 0, 1, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 2, 2, 1, 3, 3, 1, 0, 0, 0, -2, -2, -1, 0, 0, 1, 0, 1, 1, 0, 1, 0, -2, -1, 0, -1, 0, 0, 0, -2, -1, 0, 1, 2, 2, 3, 5, 3, 2, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -2, 0, 0, 1, 1, 2, 2, 4, 4, 1, 1, 0, -1, -1, -1, 0, -1, 0, 1, 1, 0, 1, 1, 0, 0, -2, 0, 0, -1, 0, -1, -2, -2, -1, 0, 0, 0, 1, 1, 2, 3, 2, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, -2, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 3, 3, 2, 1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 1, 1, 3, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, -1, 0, 1, 0, -1, -2, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 1, 1, 0, 0, 0, 1, 0, 1, 1, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 2, 2, 0, 1, 2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 3, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 2, 2, 2, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 1, 1, 0, 0, -1, -1, 0, -1, 0, 0, -2, -1, 0, 0, 1, 1, 0, 0, 0, 0, 2, 2, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 2, 1, 1, 0, -1, 0, 0, -1, -2, 0, -2, -3, -2, 0, 1, 1, 0, -2, 0, -1, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, -1, -1, 0, -1, -2, -2, -2, -2, -1, -1, 0, -1, -1, 0, -2, 1, 1, 0, 0, 1, 0, 1, 2, 0, 1, 0, 0, 0, -1, 0, -2, -1, 0, 0, -1, -1, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -3, -3, -3, -1, -1, -2, -1, -2, -2, -3, -2, -2, -3, -2, -2, 0, 0, 0, -1, 0, 0, -1, -1, -2, -2, -1, -1, -1, 0, -1, -1, -2, -3, -3, -3, -4, -2, -2, -2, -1, -3, -3, -2, -1, -3, -2, -4, -1, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, 0, -1, 0, -1, -1, 0, -2, -2, -4, -2, -1, -1, 0, 0, -1, 0, -1, -1, -1, -2, -3, -3, 0, -1, 0, 0, 0, -2, -2, -2, -2, 0, 1, -1, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 1, 3, 1, 0, 0, 0, -1, -1, -2, -2, 0, 0, -1, 0, 0, -2, -2, -3, -2, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, 1, 0, 2, 2, 5, 4, 2, 2, 1, 0, -1, -1, -1, 0, 0, 0, 1, 0, -2, -2, -2, 0, -1, 0, 0, 0, 0, 1, 2, 2, 3, 3, 2, 3, 3, 3, 5, 5, 3, 2, 2, 1, 0, -2, -1, 0, -1, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 1, 1, 3, 2, 2, 2, 3, 3, 4, 3, 4, 7, 6, 4, 4, 1, 1, 0, -2, -2, 0, -1, -1, 2, 1, 0, -1, -3, -1, 0, 0, 0, 0, 2, 3, 2, 2, 3, 3, 2, 4, 5, 4, 6, 6, 4, 3, 1, 1, 1, -1, -2, 1, 0, -1, 1, 1, 0, -1, -2, 0, 0, 0, 1, 1, 4, 3, 3, 4, 4, 3, 3, 4, 3, 4, 5, 5, 3, 3, 2, 0, 1, 0, -2, 1, -1, 0, 1, 1, 0, 0, -2, -2, 0, 1, 1, 1, 4, 5, 3, 4, 4, 2, 0, 2, 2, 5, 6, 5, 4, 2, 2, 1, 1, 0, -3, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 3, 4, 5, 5, 3, 4, 2, 1, 1, 1, 4, 5, 4, 2, 2, 4, 3, 2, -2, -2, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 3, 5, 4, 4, 5, 3, 1, 2, 1, 0, 2, 6, 4, 3, 3, 3, 2, 2, -1, -2, 0, 0, 0, 1, 0, -2, -2, -1, 0, 0, 0, 0, 2, 4, 4, 5, 5, 3, 0, 0, 0, 0, 2, 5, 5, 3, 2, 4, 5, 2, -1, -3, 0, 0, 1, 1, -1, -3, -3, 0, 0, -1, 0, 0, 1, 4, 3, 5, 5, 4, 1, 0, 0, 0, 0, 2, 3, 4, 4, 4, 4, 2, 0, -3, 0, 0, 2, 0, 0, -2, -1, -1, 0, 0, 0, 1, 1, 4, 3, 3, 4, 4, 0, 0, 0, 1, 1, 2, 2, 3, 3, 6, 4, 3, 0, -3, 0, 0, 2, 1, -1, -2, -2, 0, 0, 0, 1, 0, 3, 4, 3, 3, 4, 4, 0, 1, 2, 3, 1, 0, 4, 2, 3, 5, 5, 3, 0, -3, 0, 0, 2, 0, -2, -1, 0, 0, 0, 1, 0, 0, 1, 3, 3, 3, 4, 4, 2, 1, 2, 3, 0, 2, 4, 2, 3, 5, 4, 1, -1, -2, 0, 0, 2, 0, -1, -1, 0, 0, 0, 0, 1, 1, 2, 2, 2, 3, 3, 4, 2, 0, 3, 3, 1, 3, 3, 2, 3, 5, 3, 0, 0, -2, 0, 0, 2, 0, -1, 0, 0, 1, 0, 2, 1, 2, 2, 2, 3, 2, 4, 4, 2, 1, 3, 4, 3, 3, 4, 3, 4, 5, 4, 0, -1, -1, 0, 1, 2, 1, -1, 0, 0, -1, 0, 0, 1, 1, 2, 3, 4, 3, 3, 4, 0, 1, 4, 5, 3, 4, 3, 3, 3, 4, 2, 1, 0, -2, 0, 1, 1, 1, -1, 0, 1, 0, 0, 1, 0, 0, 1, 3, 4, 3, 5, 4, 2, 0, 3, 3, 3, 4, 3, 2, 3, 3, 2, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 2, 5, 5, 4, 3, 1, 0, 4, 3, 3, 3, 3, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 2, 0, 0, 0, 3, 5, 4, 4, 3, 0, 0, 1, 3, 3, 3, 3, 2, 3, 1, 0, -1, -2, -1, 0, 0, 0, 1, 1, 2, 0, 0, 0, 1, 1, 0, 0, 2, 4, 4, 4, 4, 2, 0, 1, 3, 2, 3, 3, 3, 1, 0, -1, 0, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 3, 2, 2, 3, 3, 2, 1, 1, 2, 4, 4, 3, 2, 0, 0, -1, -2, -1, 0, 0, 1, 0, 0, 0, 0, 2, 0, 0, 0, 2, 1, 1, 4, 3, 3, 4, 3, 2, 1, 2, 3, 3, 3, 2, 1, 0, -1, -2, -3, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 2, 2, 1, 2, 1, 2, 3, 3, 2, 4, 3, 1, 3, 3, 2, 1, 0, -1, -2, -4, -1, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 3, 0, 2, 1, 1, 3, 2, 3, 3, 2, 2, 2, 1, 1, 1, 0, 0, -3, -4, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 2, 2, 2, 2, 1, 1, 1, 2, 1, 0, 0, 0, -1, -3, -3, -2, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -2, -2, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 2, 1, 1, 2, 2, 3, 1, 2, 1, 2, 2, 1, 2, 2, 2, 1, 2, 1, 1, 0, 0, 0, 1, 0, 1, 2, 2, 1, 2, 2, 2, 3, 2, 2, 3, 4, 3, 3, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 0, 0, 1, 3, 2, 2, 3, 1, 2, 2, 3, 4, 3, 2, 2, 2, 2, 1, 1, 0, 0, 0, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 1, 1, 2, 2, 3, 2, 1, 2, 1, 0, -1, -1, -2, -1, -2, -2, -3, -2, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 2, 0, 1, 0, 3, 2, 3, 2, 0, 0, -1, -3, -2, -2, -2, -1, -3, -1, -2, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 0, 1, 1, 1, 1, 3, 2, 2, 3, 2, 0, -1, -2, -2, -4, -1, -1, -1, -2, -1, -1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 2, 2, 3, 1, 0, 1, 0, -2, -1, -3, -2, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, -2, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 2, 2, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -2, -1, -2, -2, -2, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -3, -2, -2, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, -2, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -2, -3, -3, -3, -2, -1, 0, 2, 1, 0, 0, 0, 0, 1, 0, 0, -1, -2, 0, -1, -1, -1, 0, 0, 1, 2, 0, 0, 0, 0, -1, -1, -2, -3, -2, -4, -1, -2, 0, 1, 0, 0, 1, 0, 1, 1, 0, -1, -2, -2, -1, -1, -2, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, -1, -2, -2, -4, -2, -2, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, -3, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -4, -4, -3, -2, -1, -1, 1, 0, 1, 0, 1, 0, 1, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -5, -4, -3, -3, -2, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, -2, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -3, -4, -5, -4, -3, -1, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, 0, -1, -2, -3, -2, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, -3, -4, -2, -3, -3, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -2, -2, -3, -3, -2, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -2, -2, -2, -2, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 1, 2, 0, 1, 0, -1, 0, -1, -2, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 2, 1, 2, 1, 0, 0, 0, -1, -1, -2, -2, -2, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 1, 0, 1, 0, 0, 0, 2, 1, 0, 0, -1, -2, -2, -1, -1, -2, -1, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, -1, -1, -1, -2, -2, -2, 0, -2, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 0, 1, 0, -1, -3, -2, -2, -1, -1, 0, -1, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, -3, -2, -3, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 2, 1, 0, 0, -2, -3, -3, -3, -2, 0, -1, -1, 0, -1, 0, 1, 1, 1, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, -2, -2, -3, -3, -1, -2, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 1, 2, 1, 0, 1, 0, 0, 0, 2, 0, 0, -2, -1, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 1, 2, 2, 2, 1, 2, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, -2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 3, 3, 1, 1, 1, 2, 3, 1, 1, 1, 3, 3, 3, 5, 4, 2, 2, 3, 2, 0, -2, -2, 0, -1, 0, 0, 1, 2, 3, 2, 4, 4, 3, 2, 1, 2, 3, 3, 3, 2, 1, 1, 2, 2, 0, 0, 1, 2, 3, 3, 2, 0, -1, 0, 0, 0, 0, 1, 2, 2, 2, 2, 3, 3, 2, 0, 0, 2, 1, 0, 0, 0, -1, 0, -2, 0, -1, -1, 0, 1, 2, 2, 1, 0, -1, 0, 0, 0, 0, 1, 3, 3, 2, 0, 0, 0, 0, 0, 2, 1, 0, -2, -3, -3, -2, -3, -4, -3, -1, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, -1, 0, 1, 2, 1, 2, 1, 0, 1, 2, 1, 2, 1, 0, -4, -5, -6, -4, -5, -3, -2, -1, -1, 0, 0, 1, 2, 2, 0, 0, 0, 0, -1, 0, 1, 2, 1, 1, 0, 0, 1, 2, 2, 2, 0, 0, -3, -5, -5, -4, -2, -2, 0, 0, 0, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 2, 2, 1, 1, 1, 0, -2, -3, -4, -3, -1, -2, 0, 1, 0, 0, 0, 3, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -2, 0, 1, 2, 1, 2, 0, 0, -1, -3, -3, -3, -1, -2, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -3, -1, -1, 0, 0, 2, 1, 0, 0, -1, -2, -4, -3, -3, -2, -2, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -2, -2, 0, 0, 0, 2, 2, 0, -1, -1, -3, -2, -2, -3, -2, -2, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, -1, -3, 0, -1, 0, 1, 3, 1, 0, 0, -1, -1, -2, -2, -2, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 2, 1, -1, -1, -1, 0, 0, 1, 2, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 2, 2, 0, 0, 0, 1, 0, 1, 1, 0, 0, -2, -2, -1, 0, 0, 2, 2, 1, 2, 0, 1, 0, -1, -1, -2, -2, 0, 0, 0, -2, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -1, -1, 1, 1, 3, 2, 1, 0, 0, -1, -1, -1, -2, -1, 0, -1, -2, -1, -1, 0, 2, 1, -1, -1, 0, 1, 0, 0, 0, -1, -2, -4, -3, -1, 0, 2, 2, 2, 1, 0, 0, -1, -1, -1, -2, -2, 0, 0, -2, 0, 0, 1, 1, 0, -2, -2, 0, 0, 0, 0, -1, -2, -3, -4, -3, -1, 1, 1, 0, 2, 1, -1, -1, -1, -2, 0, 0, -1, -1, 0, -2, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -3, -3, -4, -3, 0, 0, 1, 2, 3, 0, -1, -2, 0, -1, 0, -1, -1, -3, -2, -2, 0, 1, 2, 1, 0, -2, 0, 0, 1, 1, 0, -2, -3, -2, -3, -3, -1, -1, 2, 3, 3, 0, 0, 0, 0, 0, -1, -1, -1, -2, -3, -2, 0, 0, 2, 1, 0, -2, -2, 0, 1, 0, -1, -1, -3, -2, -2, -2, -2, 0, 3, 4, 4, 1, -1, 0, -1, -1, 0, -2, -2, -3, -1, 0, 0, 0, 3, 3, 0, -2, -1, -1, 0, 0, -1, -2, -2, -2, -3, -3, -3, 0, 2, 4, 3, 1, 0, 0, -1, -2, -2, -3, -2, -1, 0, 1, 2, 2, 4, 3, 0, -1, -1, 0, 0, 0, 0, -2, -2, -2, -3, -3, -1, 0, 3, 4, 3, 0, 0, 0, -2, -2, -1, -4, -2, 0, 0, 2, 1, 2, 3, 3, 0, 0, 0, 2, 1, 1, 0, -1, -2, -4, -3, -4, -1, 0, 1, 4, 2, 1, 0, 0, -3, -3, -2, -2, -2, 0, 1, 2, 3, 4, 4, 2, 0, 0, 0, 2, 1, 0, 0, -2, -1, -3, -3, -2, -1, 1, 2, 1, 1, 2, 0, -1, -3, -4, -3, -3, 0, 1, 1, 2, 2, 3, 5, 3, 0, 0, 0, 1, 1, 1, 0, -1, -2, -1, -1, -1, 0, 2, 1, 1, 1, 1, 0, -1, -2, -3, -3, -2, 0, 1, 1, 3, 3, 3, 5, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 2, 1, 0, -2, -2, -3, -4, -3, -1, 0, 0, 2, 3, 3, 3, 5, 1, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 2, 1, 2, 1, 1, -1, -4, -6, -6, -3, -1, 0, 1, 2, 1, 2, 2, 4, 4, 2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, -5, -6, -5, -3, -2, 0, 1, 1, 1, 1, 3, 4, 4, 3, 0, -2, -2, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -3, -4, -6, -4, -2, 0, 0, 1, 0, 0, 1, 3, 4, 4, 3, 1, -2, -1, -2, -1, 0, 0, 1, 0, 1, 2, 1, 0, -1, 0, -1, -1, -2, -5, -4, -3, 0, 1, 0, 1, 1, 1, 3, 5, 5, 4, 2, 0, -4, -2, -2, -2, 0, 0, 0, 1, 2, 1, 1, 0, 0, -2, 0, -1, -2, -2, -2, 0, 2, 4, 3, 4, 2, 2, 4, 5, 5, 4, 2, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 3, 5, 5, 4, 4, 3, 5, 4, 4, 3, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 1, 1, 1, 2, 2, 2, 4, 4, 3, 3, 4, 4, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, -2, -3, -2, -2, -1, 0, 0, 0, 0, 1, 2, 2, 3, 2, 3, 3, 5, 5, 4, 4, 2, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, 2, 2, 3, 1, 3, 2, 4, 3, 3, 3, 0, 1, -1, -1, -2, -3, -1, -2, -1, -1, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 2, 2, 0, 0, 2, 3, 3, 3, 2, 0, 0, -1, -2, -3, -3, -4, -3, -3, -3, -3, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 2, 2, 4, 2, 2, 0, 0, -3, -2, -3, -4, -4, -2, -3, -2, -2, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 2, 1, 0, 1, 3, 3, 3, 2, 2, 0, -1, -2, -4, -3, -4, -2, -2, -1, -1, 0, -1, -2, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 2, 2, 4, 1, 1, 0, -2, -3, -3, -2, -3, -1, -2, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 3, 3, 0, 0, 0, -1, -2, -3, -2, -1, -1, -3, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 2, 1, 2, 0, 0, -1, 0, -3, -1, -2, -2, -1, -3, -1, 0, 1, 0, 0, -1, 0, 1, 2, 0, 0, 0, 1, 2, 2, 1, 1, 1, 1, 3, 1, 1, 1, 0, 0, -2, -2, -1, -1, -3, -2, -1, -2, 0, 0, 0, -2, -1, 0, 2, 1, 0, 0, 0, 1, 3, 3, 3, 2, 1, 1, 3, 3, 1, 2, 0, 0, -1, -1, -1, -3, -2, -2, -3, -1, -2, -1, -1, -4, -1, 0, 2, 3, 1, 0, 0, 2, 2, 5, 4, 0, 0, 1, 3, 3, 2, 2, 1, 1, -2, -2, -3, -1, -2, -2, -3, -3, -3, -2, -4, -4, -2, 0, 2, 2, 1, 0, 1, 1, 2, 3, 3, 1, 0, 2, 4, 3, 3, 1, 0, 1, -2, -3, -2, -1, 0, -2, -2, -2, -4, -4, -4, -5, -2, -1, 1, 3, 1, 0, 0, 1, 2, 3, 2, 1, 2, 3, 3, 3, 3, 3, 0, 1, -1, -4, -4, -1, -1, -1, -1, -3, -4, -4, -5, -4, -3, -2, 0, 1, 0, 0, 0, 0, 0, 3, 3, 0, 1, 3, 3, 2, 3, 2, 1, 1, -1, -3, -4, -1, -1, 0, -1, -2, -3, -6, -6, -5, -4, -3, 0, 3, 2, 0, 0, 0, 0, 1, 1, 0, 2, 3, 2, 2, 3, 1, 1, 1, 0, -3, -3, -2, 0, 0, 0, -3, -5, -5, -5, -5, -4, -2, 0, 2, 1, 0, 0, 0, 0, 1, 2, 0, 0, 2, 1, 1, 1, 0, 0, 0, -2, -4, -3, -3, -2, -1, 0, -2, -4, -6, -7, -4, -4, -2, 0, 2, 1, 0, 1, 0, 0, 0, 2, 2, 2, 3, 2, 1, 1, 0, 0, 0, -1, -3, -2, -3, -1, -1, -1, -2, -4, -6, -5, -5, -4, -2, 0, 2, 1, -1, 0, 0, 0, 0, 1, 1, 3, 1, 0, 0, 0, 0, 1, 0, -2, -3, -3, -2, -1, -1, -1, -1, -3, -3, -3, -5, -4, -1, 0, 1, 1, 0, -1, 0, 0, 0, 0, 1, 3, 3, 0, 1, 0, 1, 1, 0, -1, -3, -2, -1, -1, -2, -1, -1, -1, -2, -2, -3, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 3, 2, 1, 1, 1, 1, 0, 0, 0, -2, -1, -2, -2, -3, -1, 0, -1, -1, -1, -1, -2, -1, 0, 0, 0, -1, 0, 0, 1, 1, 2, 2, 3, 2, 2, 1, 1, 1, 2, 0, -1, -2, -2, -3, -2, -3, -2, -2, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 2, 3, 4, 2, 3, 3, 1, 2, 1, 1, 1, 0, 0, -1, -2, -1, -2, -2, -1, -1, -2, 0, 0, 0, 1, 0, 0, 1, -1, -1, -1, 0, 2, 2, 3, 2, 2, 2, 2, 3, 3, 1, 0, -1, -2, -2, -1, -2, -2, -1, 0, -2, -1, -2, -1, 1, 1, 0, 0, 0, 0, -2, -2, 0, 0, 2, 0, 2, 2, 2, 3, 3, 2, 0, 0, -1, -2, -1, -2, -2, -2, 0, -1, -1, 0, -1, -1, 0, 1, 1, 0, 0, -1, -1, -1, -1, 0, 0, 1, 1, 2, 3, 3, 3, 3, 1, 0, 0, -2, -3, -3, -3, -2, -1, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 3, 2, 2, 3, 1, 1, 0, -1, -3, -3, -4, -1, -2, -1, 0, 0, -1, 0, 2, 2, 0, -1, -1, -1, -1, -1, -2, -2, -1, -1, 0, 0, 1, 2, 1, 3, 2, 1, 0, -2, -4, -4, -5, -3, -3, -3, -2, -1, 0, 0, 1, 1, 0, 0, -1, -2, -1, -2, -1, -1, 0, -1, 0, 0, 1, 2, 2, 2, 2, 3, 1, 0, -2, -4, -4, -5, -4, -3, -2, 0, -1, -1, -1, 0, 0, -1, -2, -3, -2, -3, -3, -2, -2, 0, 0, 0, 0, 0, 2, 3, 3, 3, 4, 3, 0, -2, -3, -2, -3, -3, -1, 0, 0, 0, -2, -2, -1, -4, -4, -3, -2, -2, -2, -2, 0, -1, 0, 0, 0, 0, 2, 3, 5, 4, 5, 4, 1, 0, 0, -1, -1, -3, -1, -1, 0, -1, -2, -3, -2, -4, -3, -3, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 2, 2, 2, 3, 3, 3, 2, 1, 0, -1, -1, -2, 0, -1, 0, -1, -2, -2, -1, -2, -1, -2,
    -- filter=0 channel=2
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 2, 2, 0, 2, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 2, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 2, 1, 1, 0, 1, 2, 0, 1, 0, 1, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 1, 1, 0, 2, 1, 2, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 2, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 1, 0, 0, 0, 2, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, -1, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 2, 0, 1, 0, 0, -2, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -2, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -2, 0, -2, -1, 0, -2, 0, 0, 0, -1, 1, 1, 0, 0, 1, 0, 0, 0, 0, -2, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, -1, -1, -2, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, -1, 0, -1, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, -1, -1, -1, -2, -1, -2, 0, -1, 0, 0, 0, 0, 1, 2, 1, 1, 2, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -1, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 2, 1, 0, -2, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, -1, -1, -1, 0, 0, 1, 1, 1, 1, 1, 1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 1, 1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 2, 0, 1, 0, 0, -1, 0, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 1, 1, 0, -1, 0, -2, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 2, 1, 1, 2, 2, 0, 1, 1, 0, 1, 2, 1, 0, 0, 1, 0, 0, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 2, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, -2, -2, -2, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, -2, -2, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -2, 0, -1, -2, -1, 0, 0, 0, 1, 0, 1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 2, 1, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 2, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 2, 1, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 1, 1, 0, 0, 1, 2, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 2, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 1, 2, 2, 1, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, -1, -2, 0, -1, -2, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 1, 0, 1, 1, 2, 1, 1, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, -2, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, -2, -1, -2, -2, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -3, -2, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 2, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 1, 2, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 2, 0, 1, 2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 2, 0, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 1, 2, 1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 2, 3, 2, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 1, 1, 0, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, 1, 1, 1, 2, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 1, 2, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 2, 2, 1, 1, 1, 1, 1, 1, -1, -1, -2, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 2, 1, 0, 1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, -1, 0, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -2, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, -1, -2, -1, -2, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, 1, 1, 1, 1, 2, 1, 2, 1, 1, 0, 0, -1, -1, -1, 0, 0, 0, -1, -2, -1, 0, 1, 2, 2, 1, 1, 0, 1, 0, 0, 0, 0, 2, 3, 3, 2, 3, 4, 3, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 3, 3, 3, 1, 0, 0, 2, 3, 3, 4, 4, 2, 2, 2, 3, 1, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 2, 1, 1, 2, 3, 1, 0, 1, 1, 3, 4, 5, 4, 2, 2, 2, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 2, 2, 1, 1, 1, 2, 0, 0, 1, 2, 4, 3, 3, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 1, 1, 1, 2, 1, 2, 3, 2, 3, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 2, 2, 1, 2, 1, 1, 2, 2, 2, 3, 3, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 1, 2, 2, 1, 1, 3, 2, 2, 2, 2, 3, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 1, 1, 0, 2, 3, 2, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, 0, 1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 2, 1, 2, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, -1, -1, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 1, 2, 1, 0, 0, 0, 1, 0, 1, 2, 2, 2, 2, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 3, 1, 0, 1, 0, 1, 1, 2, 2, 1, 1, 1, 1, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 2, 2, 0, 0, 1, 1, 2, 1, 2, 2, 1, 1, 1, 1, 2, 0, 1, 0, 2, 2, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 0, 1, 2, 1, 0, 1, 1, 2, 1, 2, 1, 3, 1, 2, 2, 1, 1, 1, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 2, 2, 0, 2, 2, 2, 2, 1, 1, 1, 1, 0, 1, 0, 0, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, 1, 2, 1, 2, 2, 3, 3, 2, 2, 2, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 2, 1, 3, 4, 3, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 1, 2, 2, 2, 2, 2, 1, 1, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 2, 2, 2, 1, 1, 1, 1, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 1, 2, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 2, 2, 2, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 2, 1, 0, 1, 0, 1, 1, 1, 0, 1, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 2, 1, 2, 1, 2, 3, 1, 1, 2, 0, 1, 1, 1, 0, 0, 1, 2, 1, 1, 1, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 2, 3, 1, 3, 1, 1, 0, 1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 2, 1, 2, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -2, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, -3, -2, -2, -2, -2, -1, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, -2, 0, 0, -1, -2, -1, -3, -4, -3, -2, -2, 0, -1, -1, -1, -2, -1, -1, 0, -2, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, -1, -1, -1, -2, -2, -1, -2, -2, -1, -2, -2, 0, -1, -1, -1, -1, -1, -1, -2, 0, -1, -1, 0, 0, 0, 0, -1, -2, -1, -2, -2, -2, -2, -1, -2, -1, -3, 0, -2, -3, 0, -1, -1, -1, -1, -1, 0, -1, -2, -1, -2, -2, -1, -2, -1, -2, -2, -2, -1, -1, 0, 0, -1, -1, -1, -1, -1, -1, -2, 0, 0, -2, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, -2, 0, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 2, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, -1, -2, -1, 0, -1, 0, 1, 1, 3, 2, 2, 1, 1, 1, 0, 0, 1, 1, 2, 1, 1, 0, 2, 3, 2, 1, 2, 0, 0, 2, 1, 0, 0, -1, -2, -1, 0, 1, 0, 1, 3, 4, 3, 4, 1, 2, 1, 1, 1, 2, 3, 2, 2, 2, 2, 3, 2, 1, 1, 1, 3, 3, 1, 0, 0, -1, -2, 0, 0, 1, 1, 1, 3, 3, 5, 4, 2, 1, 3, 2, 3, 3, 4, 2, 2, 4, 3, 4, 4, 2, 2, 2, 4, 3, 1, 0, 0, -2, -2, 0, 0, 1, 1, 1, 3, 3, 4, 4, 3, 1, 3, 2, 2, 3, 5, 3, 4, 5, 3, 3, 4, 2, 2, 4, 5, 3, 2, 1, 0, -1, 0, 0, 0, 0, 1, 2, 2, 2, 3, 3, 1, 2, 3, 2, 4, 5, 4, 4, 3, 4, 4, 4, 4, 4, 3, 5, 4, 4, 2, 0, 0, -2, 0, 0, 0, 1, 0, 2, 0, 2, 2, 1, 1, 2, 3, 3, 5, 6, 4, 3, 2, 2, 3, 3, 4, 5, 3, 4, 3, 3, 3, 1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 1, 3, 6, 6, 6, 5, 5, 3, 4, 3, 3, 3, 5, 4, 3, 4, 3, 2, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 2, 2, 2, 4, 5, 5, 7, 6, 5, 4, 4, 3, 3, 3, 3, 4, 4, 3, 3, 2, 1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 2, 2, 4, 4, 6, 7, 6, 6, 4, 4, 3, 2, 1, 1, 2, 2, 2, 2, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 3, 2, 4, 4, 4, 4, 5, 4, 3, 3, 2, 3, 2, 2, 2, 1, 2, 2, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 3, 2, 4, 3, 2, 3, 2, 2, 2, 3, 2, 2, 1, 0, 2, 2, 2, 0, -1, 0, -1, -2, -1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 2, 2, 3, 2, 1, 2, 2, 3, 2, 3, 3, 1, 2, 1, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 1, 2, 2, 1, 2, 1, 3, 2, 2, 3, 2, 4, 3, 3, 3, 2, 3, 3, 4, 3, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 3, 3, 3, 3, 4, 3, 3, 2, 4, 5, 5, 3, 2, 2, 3, 4, 3, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 1, 0, 1, 2, 2, 2, 5, 4, 6, 4, 4, 3, 4, 5, 4, 5, 2, 3, 4, 4, 4, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 3, 4, 5, 5, 3, 3, 2, 3, 4, 5, 4, 2, 3, 3, 2, 2, 1, 0, 0, -1, -1, 0, 0, 1, -1, -1, -1, -1, 0, 0, 0, 1, 0, 2, 3, 2, 3, 2, 2, 2, 3, 3, 4, 2, 1, 1, 2, 1, 1, 0, 0, -2, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 1, 2, 1, 1, 2, 3, 1, 2, 3, 2, 1, 0, 0, 0, 1, 0, 0, 0, -2, -2, -1, 0, -1, -2, -2, -1, -3, -3, 0, -1, -1, -2, 0, 0, 1, 1, 1, 1, 1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, -2, -3, -3, -3, -1, -1, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, -2, 0, -1, -2, -1, 0, -1, -2, 0, -1, -2, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, 0, -2, -2, 0, 0, -2, -1, -1, -1, 0, -2, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -2, -2, 0, -2, -2, 0, 0, -2, 0, -2, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -2, 0, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, -2, 0, 1, 1, 0, 0, 0, 2, 1, 0, 1, 0, 0, -1, 0, 0, -1, -1, -1, 0, -2, -2, -2, -1, 0, -1, 0, -2, -1, -2, -2, 0, 0, 1, 0, 3, 2, 1, 2, 2, 2, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -2, -2, -1, -2, -2, -2, -2, -1, -2, -2, -2, 0, 1, 3, 4, 3, 3, 3, 3, 1, 2, 1, 1, 1, 2, 0, 1, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, -1, -1, -1, -1, 0, 1, 3, 3, 2, 1, 2, 2, 3, 1, 2, 0, 1, 3, 2, 3, 2, 3, 3, 3, 4, 4, 3, 2, 2, 2, 1, 0, -1, -2, -1, 0, 0, 0, 2, 1, 1, 1, 1, 2, 3, 4, 3, 3, 4, 4, 5, 5, 4, 4, 4, 5, 4, 4, 4, 4, 3, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 2, 1, 1, 2, 1, 2, 3, 3, 2, 2, 5, 5, 4, 6, 4, 4, 4, 5, 5, 5, 4, 3, 1, 1, 1, 0, -1, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 2, 2, 2, 3, 5, 5, 6, 4, 4, 3, 5, 4, 4, 5, 3, 2, 0, 1, -1, -2, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 2, 0, 2, 2, 3, 4, 5, 4, 2, 2, 4, 4, 6, 5, 5, 3, 2, 1, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, -2, -1, 0, 1, 1, 2, 2, 4, 4, 3, 3, 2, 0, 1, 1, 4, 3, 4, 4, 4, 2, 0, -1, -3, -1, 0, 0, -2, -2, -1, -1, -2, -3, -1, 0, 1, 2, 3, 4, 5, 4, 2, 2, 0, -1, 0, 0, 3, 4, 4, 4, 2, 0, 0, -2, -3, -2, -1, -1, -2, -1, -1, -1, -3, -3, -2, 0, 0, 2, 1, 3, 4, 2, 0, -1, -1, -1, 0, 0, 1, 2, 3, 2, 3, 0, 0, -2, -4, -3, -2, -1, -2, 0, -1, -1, -2, -2, -2, 0, 0, 0, 0, 1, 2, 0, -2, -2, -1, -1, -1, 0, 0, 2, 2, 2, 2, 0, -2, -4, -5, -3, -1, 0, 0, 0, -1, 0, 0, -2, -2, 0, 0, 0, 0, 0, -1, -3, -4, -3, -2, -2, -1, 0, 0, 1, 1, 2, 1, 0, -1, -4, -5, -4, -1, -2, -2, -1, -1, 0, -1, -2, -1, 0, -2, -2, -1, -3, -5, -5, -5, -4, -4, -4, -1, -2, -1, 0, 1, 1, 0, 0, -3, -5, -6, -4, -2, 0, -2, -1, -1, -2, -1, -1, 0, -2, -2, -3, -5, -4, -6, -6, -6, -6, -4, -2, -2, -2, -3, -1, 0, 0, 0, -1, -3, -5, -4, -4, -2, -2, -2, -1, -3, -3, -4, -2, -1, -2, -3, -4, -7, -8, -6, -6, -7, -7, -4, -3, -2, -2, -2, 0, 0, 0, 0, -1, -2, -4, -5, -3, -2, 0, -2, -2, -2, -3, -2, -3, -1, -2, -3, -6, -6, -8, -7, -6, -6, -5, -3, -1, 0, 0, 0, 0, 0, 1, 1, 0, -2, -3, -6, -4, -1, 0, -2, 0, -1, -2, -1, 0, 0, 0, -4, -6, -6, -7, -6, -6, -5, -4, -2, 0, 0, 0, 0, 0, 1, 2, 1, 0, -2, -5, -6, -3, -2, -1, 0, 0, -1, -1, -1, 0, 0, 0, -3, -4, -5, -6, -7, -6, -5, -3, -1, 0, 0, 0, 0, 1, 2, 1, 2, 0, -2, -4, -5, -3, -3, 0, -2, 0, 0, 0, 0, 0, 0, -2, -1, -4, -4, -5, -5, -3, -3, -4, -2, -2, -1, 1, 0, 2, 3, 3, 2, 0, -1, -5, -6, -2, -2, 0, -2, 0, 0, -1, -2, -1, -2, -2, -2, -3, -3, -2, -2, -2, -2, -3, -2, -2, 0, 1, 3, 2, 3, 3, 1, 0, 0, -3, -5, -4, -2, -1, 0, 0, 0, -2, -2, -2, -2, 0, 0, 0, 1, 0, 0, 0, -1, -3, -2, -3, 0, 0, 2, 4, 4, 3, 3, 1, 0, -3, -4, -4, -2, -1, 0, 0, -1, -2, -3, -2, -2, 0, 0, 0, 1, 2, 2, 2, 0, -1, -3, -2, -1, 1, 3, 5, 5, 3, 2, 1, 0, -2, -3, -3, 0, 0, 0, -2, -2, -2, -3, -2, -2, 0, 2, 2, 3, 4, 3, 3, 1, 1, 0, 0, 1, 3, 5, 5, 4, 3, 3, 2, 0, -3, -3, -2, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, 2, 3, 3, 5, 4, 3, 4, 2, 2, 2, 3, 4, 3, 3, 3, 1, 1, 2, 0, -1, -2, -1, 0, -1, -1, 0, -1, -2, 0, 0, 0, 1, 1, 3, 3, 3, 3, 4, 2, 3, 2, 2, 4, 3, 4, 4, 2, 2, 0, 0, -1, -2, -3, -2, 0, 0, -1, 0, -1, 0, 0, 0, 2, 2, 3, 1, 2, 2, 1, 3, 3, 3, 3, 2, 2, 4, 2, 2, 3, 3, 1, 0, -1, -3, -3, -1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 3, 2, 2, 2, 0, 2, 2, 1, 2, 3, 2, 3, 2, 4, 3, 2, 2, 2, 0, -1, -3, -4, -2, 0, 1, 0, 2, 2, 0, 3, 3, 3, 2, 3, 2, 1, 0, 2, 2, 2, 2, 1, 1, 2, 1, 1, 2, 2, 2, 1, 0, -1, -4, -3, -1, 0, 0, 1, 2, 3, 2, 3, 3, 3, 4, 3, 2, 2, 2, 0, 2, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, -1, -3, -3, -3, -1, 0, 1, 0, 2, 0, 1, 1, 1, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -3, -3, -2, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 2, 1, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -2, -2, -1, -1, -2, -2, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -2, -2, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, -1, -1, -1, -2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 1, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 1, 0, -2, -1, -1, -1, -1, -1, 0, 0, -1, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -2, -2, -2, 0, -1, -1, -1, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -2, -3, -4, -1, -1, -1, 0, -2, -1, -1, 1, 0, -1, -1, -1, 0, 0, -1, 0, -1, -1, -2, -2, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, -3, -2, -2, 0, 0, 0, 0, 0, 0, 1, 0, -2, -2, -2, -1, 0, -1, 0, 0, -1, -1, -3, -2, -1, 0, -1, 0, 1, 1, 1, 0, 0, -2, -1, -2, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, -2, 0, -1, -1, 0, -1, -2, -3, -4, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, -2, -2, -1, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, 0, 0, -2, -2, 0, -1, -1, -3, -3, -2, -2, -1, -2, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, -1, -1, 0, 1, 0, -1, -2, -2, 0, -1, -1, -1, -2, -2, -2, -3, -3, -3, -2, -1, -2, -1, 0, 1, 1, 0, 0, -2, -1, -2, 0, 0, -2, -1, 0, 0, 1, 0, -1, -1, 0, 0, -1, -1, -1, -1, -2, -2, -3, -2, 0, -2, -1, -1, 0, 1, 2, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, -2, -1, -2, -2, -2, -2, -1, 0, -1, -2, -2, -3, 0, 1, 1, 0, 0, 0, -1, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -2, -1, -2, -2, 0, 0, 0, -2, -3, -2, -1, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, 0, 0, -1, -1, 0, 0, -1, -2, -1, 0, -2, -1, -3, -2, -2, 0, 0, 0, -2, -1, 0, -2, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 2, 0, 0, -2, -1, 0, -1, -1, -1, 0, 0, -1, -2, -1, -2, 0, 0, 0, -1, -1, 0, -1, 0, -2, -1, -2, -1, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, -2, 0, -1, 0, -2, -1, 0, 0, -1, -1, -1, -1, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -3, -2, 0, 0, -1, -1, -1, -1, -2, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -3, -3, -2, 0, 0, -1, -1, -1, -2, -2, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -3, -1, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -1, 0, -1, -1, 0, -2, -1, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, -1, -2, -2, -2, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, -1, -1, -1, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 3, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 2, 3, 2, 2, 1, 1, 1, 0, 1, 1, 0, 0, -2, -1, -1, 0, 1, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 2, 2, 0, 0, 1, 2, 2, 1, 3, 1, 1, 2, 2, 1, 1, 2, 0, 0, 0, 0, 1, 0, 1, 1, 0, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 2, 2, 1, 1, 1, 1, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 1, 1, 1, 0, 0, 1, 0, 1, 0, 2, 2, 2, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 2, 1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 2, 2, 1, 1, 0, 1, 1, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, 2, 0, 1, 1, 0, 1, 1, 2, 1, 1, 1, 1, 2, 1, 2, 1, 1, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 0, 0, 2, 2, 1, 0, 1, 2, 2, 1, 0, 1, 1, 1, 1, 2, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 1, 2, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 1, 1, 0, 1, 2, 2, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 2, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -2, -1, -3, -3, -1, -2, -1, 0, 0, 1, 2, 0, 0, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -3, -2, -2, -2, -1, 0, -1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -3, -3, -3, -3, -3, -2, -3, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, -1, -1, 0, 0, 0, 0, -1, -2, -3, -3, -4, -4, -3, -1, -1, -1, -2, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, -1, -2, -2, -2, -4, -4, -3, -2, -1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 0, -2, -2, -2, -2, -3, -3, -2, -2, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -2, -1, -1, -2, -2, -4, -2, -2, -1, 0, 0, 0, 2, 0, 1, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, -1, 0, -2, -2, -3, -3, -1, -1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -2, -2, -2, -1, -1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -3, -2, -1, -1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 1, 1, 2, 2, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 1, 2, 1, 0, -1, -1, -1, 0, 2, 1, 1, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 1, 2, 0, 0, 0, -1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 1, -1, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 2, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, -1, -1, -1, -1, 0, 0, 1, 2, 1, 1, 1, 2, 2, 2, 2, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 1, 0, 1, 1, 2, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, -1, -2, -2, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -2, -3, -2, -2, -1, -3, -4, -4, -4, -5, -3, -4, -3, -2, -3, -2, -2, 0, -1, -2, 0, 1, 1, 1, 0, 0, 0, 0, -1, -1, -1, -1, -3, -3, -2, -3, -2, -2, -3, -3, -2, -2, -3, -2, -1, -2, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -3, -2, -3, -3, -3, -3, -2, -2, -3, -2, -2, -3, -2, -2, -1, -1, -1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -3, -1, -2, -2, -2, -3, -3, -2, -1, -2, -3, -1, -3, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, -2, -2, -3, -3, -3, -2, -2, -2, -3, -3, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, 0, 1, 0, 0, 0, 0, 2, 0, 0, 0, -1, -3, -3, -2, -3, -4, -2, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, -2, -2, 0, -1, -1, -1, -2, -3, -1, -1, 0, 0, 2, 1, 2, 1, 0, -3, -3, -4, -4, -4, -1, 0, 0, 0, 2, 1, 1, -1, 0, -1, -1, -1, -1, 0, 0, -2, -1, -2, -2, -1, 0, 1, 3, 3, 2, 1, 0, 0, -2, -3, -2, -1, 0, 0, 0, 1, 1, 3, 1, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 2, 3, 3, 1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 1, 2, 3, 4, 2, 0, -1, -1, -2, -1, -3, -1, -1, 0, 0, 2, 1, 1, 2, 3, 2, 2, 0, -1, 0, -1, 0, -1, -1, -2, -1, 0, 1, 1, 2, 4, 2, 0, 0, -2, -3, -2, -3, -2, -1, 0, 1, 2, 3, 4, 4, 4, 2, 1, -1, 0, -1, -1, 0, -1, 0, -1, -1, -1, 1, 2, 3, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 3, 2, 2, 1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 2, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 1, 1, 0, 0, 0, 0, 1, 2, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, -3, -2, -1, 0, -1, 0, 0, 0, 2, 3, 3, 2, 0, -1, -2, -1, -1, 0, -1, 1, 0, 2, 3, 2, 3, 0, 0, 0, 0, 1, 0, 0, -3, -4, -3, -3, -2, -1, 0, 2, 4, 4, 2, 1, 0, 0, -2, -2, -1, 0, 0, 1, 1, 2, 2, 2, 1, 0, 1, 0, -1, 0, 0, -3, -3, -3, -2, -3, -2, -3, -2, 0, 3, 3, 2, 1, 0, -2, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -2, -3, -2, -1, -2, -3, -1, 0, 1, 2, 1, 1, -1, 0, 0, 0, 0, 0, 1, 2, 3, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -2, -2, -1, 0, 2, 2, 3, 0, -1, 0, -1, -1, 0, 1, 2, 2, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -3, -4, -3, -2, -2, -1, 0, 1, 1, 3, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, -1, -2, -1, -2, -1, -2, -1, -3, -2, -3, -1, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -2, -3, -2, -3, -2, -3, -1, -1, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -2, -1, 0, 0, -1, 0, -1, -1, -2, -1, -2, -2, -3, -3, -1, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, -1, -2, -1, 0, -1, -1, -1, -2, 0, -1, -1, -2, -1, -1, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -2, -2, -2, -3, -2, -3, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, -1, 0, -1, -3, -2, -3, -4, -3, -4, -2, -4, -2, -2, 0, 0, 0, 2, 2, 1, 0, -1, 0, 0, -1, -2, 0, 0, -2, -1, 0, 0, 0, 0, -2, -2, -2, -2, -3, -5, -3, -4, -2, -3, -2, -2, -1, -1, -1, 0, 2, 1, 0, 1, 0, 0, -1, -1, 0, 0, -1, -2, -2, -1, -3, -2, -4, -2, -2, -1, -3, -3, -3, -2, -2, -2, 0, -2, -1, 0, 0, 0, 2, 1, 0, 3, 2, 2, 0, 1, 0, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 3, 1, 0, 0, 2, 2, 2, 1, 2, 1, 1, 2, 1, 0, 0, 0, 1, 0, 0, 1, 2, 3, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 1, 1, 1, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, -1, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 2, 1, 0, 0, 0, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 0, 1, 1, 0, 1, 1, 2, 1, 0, 0, -1, -1, -2, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 2, 2, 1, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 1, 0, 0, 1, 1, 1, 1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 2, 0, 1, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 2, 2, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 2, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 2, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 1, 2, 1, 1, 2, 1, 1, 0, 1, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 1, 1, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 1, 0, 1, 0, 1, 0, 0, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 1, 1, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -2, -2, 0, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, -1, -1, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -2, -1, -1, -1, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, -1, -2, -1, -1, -2, -1, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -2, -1, -2, -2, -1, 0, -1, -1, 0, 1, 2, 2, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -2, -1, -2, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -2, 0, -2, -2, -2, -1, 0, 0, -1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -2, -2, -1, -2, -2, -2, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -3, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 2, 0, 0, 0, 2, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 1, 2, 2, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 2, 2, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, -1, -1, 0, 0, -1, -1, 0, 0, 1, 2, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -2, -1, 0, 0, -1, 0, -1, -2, -1, -3, -2, -2, 0, 1, 2, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 2, 1, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 3, 2, 0, 1, 1, 1, 1, 2, 1, 1, 1, 2, 2, 2, 2, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 2, 2, 1, 2, 0, 1, 1, 1, 1, 2, 0, 3, 3, 2, 3, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 2, 1, 1, 2, 1, 1, 2, 2, 2, 3, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 2, 0, 0, 0, 1, 2, 1, 2, 1, 0, 1, 1, 3, 1, 3, 2, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 1, 2, 1, 3, 3, 1, 0, -1, 0, 0, 0, -2, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 3, 2, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 3, 0, 0, 0, 0, -1, 0, 0, 2, 2, 1, 0, 0, -1, 0, -1, -1, -3, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, 2, -1, -1, -1, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -3, -4, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 1, 1, 1, 0, 0, -1, -1, -2, -3, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -2, -2, -1, -2, -2, -1, -1, -2, -2, 0, 0, 0, 1, 1, 0, 0, 0, -3, -2, -2, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -2, -2, -3, -3, -2, -3, -2, -2, -1, -1, -1, -2, -1, 0, 1, 0, 0, 0, -2, -2, -3, -3, -1, 0, 0, 0, 0, -1, -2, -1, 0, -1, -1, -2, -4, -3, -3, -3, -2, -3, -2, -1, 0, -1, -2, -1, 0, 1, 0, 0, -1, -1, -2, -2, -3, 0, 0, 0, 0, -2, -1, -1, 0, 0, -2, -4, -4, -3, -4, -3, -4, -3, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, -2, -3, -3, -3, 0, 0, 0, 0, 0, 0, 0, 1, 0, -3, -3, -3, -2, -2, -3, -4, -2, -1, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, -1, -2, -3, -2, 0, 0, 1, 0, 0, 0, 0, 1, 0, -2, -3, -4, -1, -1, -1, -2, -2, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, -3, -2, -4, -3, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -2, -1, -2, -1, -1, -2, -3, -2, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, -2, -4, -3, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -2, -1, -1, -2, -2, -2, -1, 0, 0, 1, 2, 1, 2, 1, 0, 0, 0, -1, -3, -4, -2, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 1, 1, 0, 0, -2, -1, -1, 0, 1, 3, 2, 3, 1, 1, 0, 0, -1, -3, -3, -2, 0, 0, 0, -1, -1, -2, -2, -1, 0, 1, 1, 0, 2, 1, 0, 1, 0, -1, 0, 0, 1, 3, 3, 2, 2, 0, 1, 0, 0, -1, -3, -2, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 2, 2, 2, 1, 0, 0, 0, 0, 3, 2, 4, 1, 1, 1, 0, 0, 0, -2, -3, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 2, 2, 2, 2, 0, 1, 0, 1, 1, 2, 2, 1, 1, 0, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 2, 1, 1, 1, 2, 1, 2, 1, 2, 2, 2, 0, 0, -1, 0, -1, -1, -3, -2, 0, 0, 0, 0, 0, 0, -1, 1, 1, 1, 0, 2, 0, 2, 1, 1, 1, 1, 1, 2, 1, 2, 1, 2, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 0, 1, 1, 1, 0, 0, 1, 1, 2, 2, 1, 0, 2, 2, 2, 0, -1, -1, -1, -2, -2, -1, 0, 1, 1, 0, 0, 0, 0, 2, 2, 1, 1, 1, 0, 0, 0, 1, 1, 1, 2, 1, 0, 2, 2, 1, 2, 0, -1, -1, -1, -2, -1, -1, 0, 0, 1, 1, 1, 0, 2, 2, 2, 1, 2, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, -1, -1, -2, -2, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, -2, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, -1, 0, 1, 1, 0, 0, -1, 0, 0, 1, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 0, 1, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, -2, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, -1, -1, -2, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -2, 0, -2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, -2, 0, 0, 1, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, -2, -1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 1, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, 0, -1, -1, -1, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -2, -1, -1, -1, -3, -3, -2, -1, -2, -2, -2, -3, -2, -2, -3, -1, -1, 0, -1, -1, -1, -2, 0, 0, 0, 0, -2, 0, 1, 0, -2, 0, -1, -1, -2, -2, -2, -3, -3, -2, -1, -2, -3, -3, -3, -3, -2, -2, -2, 0, 0, 0, 0, -2, -1, 0, 0, 0, -2, 0, 2, 0, -2, 0, -1, -1, 0, -2, -1, -3, -3, -2, -2, -3, -3, -3, -2, -4, -4, -3, -1, 0, -1, -1, 0, -1, -1, -1, 0, 0, -2, 0, 2, 0, -2, 0, -2, -2, -1, -1, -1, -1, -3, -2, -3, -4, -2, -2, -3, -3, -2, -3, -1, 0, 0, -2, -2, -1, -1, -2, 0, 0, -2, -1, 1, 0, 0, 0, -2, -2, -2, -1, 0, -1, -3, -3, -2, -3, -2, -3, -3, -3, -2, -2, -3, -1, -2, -1, -1, 0, 0, -1, -1, 0, 0, -1, 0, 1, 0, 0, -1, -2, 0, -1, 0, -3, -4, -1, -2, -3, -3, -2, -4, -2, -1, 0, -1, 0, -1, -3, 0, -2, 0, -2, -2, -1, -1, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, -2, -2, -1, -3, -2, -3, -3, -6, -4, -2, -1, -1, 1, 0, -1, -1, 0, -2, -3, -2, -1, -2, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -2, -2, -1, -2, -2, -1, -4, -5, -3, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, -3, -3, -1, 1, 1, 0, 0, 0, -1, -2, 0, -1, -2, -2, -1, -2, -2, -3, -4, -3, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -3, -1, 0, 2, 0, 0, 0, 1, -1, -1, 0, 0, -1, -2, -2, -2, -1, -2, -2, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, -1, -3, -1, 0, 1, 0, 0, 0, 1, 0, -1, -1, -1, 0, -2, -2, 0, -2, -3, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, -3, -2, 0, 0, 0, -1, 0, -1, 1, 0, -1, -1, 0, 0, -1, -1, -1, -1, -2, 0, 1, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, -1, 0, -1, -3, -2, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 1, -1, -3, -4, -1, 1, 0, 1, 0, 0, -1, -2, 0, -2, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, -1, -2, -3, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -2, -4, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 2, -1, 0, -1, 0, 0, -1, -4, -3, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 2, 0, -1, 0, 0, -2, -2, 0, 1, -1, 0, -1, -1, 0, 0, -2, -1, -2, 1, 0, 0, -1, -1, 0, -1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, -3, -2, -2, -1, -1, -2, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, -2, -1, -1, -1, 1, 2, 0, -1, -1, 0, 0, -1, 0, 1, 0, 0, -2, -1, -2, -1, 0, -1, -4, -3, -1, 0, -1, -1, 1, 2, 0, 0, -2, -2, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, -2, -1, -2, 0, -2, -3, -3, -3, -2, -2, -2, 0, 1, 0, 0, -2, -2, 0, -1, 0, 1, -1, -1, -1, 0, -1, 0, 0, 1, 0, 0, -2, -2, -2, -2, 0, -2, -3, -3, -4, -3, -2, -2, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, -3, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, -1, -3, -3, -4, -3, -2, -3, -2, 0, 0, 0, 1, 1, 0, -2, -2, 0, -1, -1, -1, -1, -2, 0, 0, 1, 2, 0, 0, -2, -2, 0, 0, -2, -2, -3, -4, -4, -3, -4, -2, -1, -2, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, -2, -2, 0, 1, 1, 1, 0, -1, -2, 0, 0, -2, -3, -3, -3, -4, -3, -3, -2, -2, -1, -1, 0, 0, 0, 0, -2, -2, -1, -1, -1, 0, 0, 0, -1, 0, 2, 2, 0, -1, -1, 0, -1, -2, -3, -2, -3, -3, -4, -3, -3, -3, -4, -3, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -4, -2, -2, -2, -2, -4, -3, -3, -4, -4, -4, -1, 0, -1, 0, -2, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, -1, -1, -4, -3, -2, -3, -1, -3, -2, -3, -2, -3, -3, -3, -2, -1, -2, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 0, -1, -1, 0, -1, -2, -3, -3, -2, -3, -3, -3, -1, -2, -3, -3, -3, -1, -1, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, -1, -1, -1, -2, -2, 0, -2, -3, -3, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, -1, -1, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 3, 1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, -2, -1, 0, 0, 1, 0, 0, 1, 2, 2, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, -1, 0, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, 0, -1, -2, -1, -2, -2, -2, -1, -1, -1, -1, 0, -1, -1, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, -2, -2, -2, -2, -2, -2, -2, -2, -2, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, -2, -2, -2, -3, -2, -3, -1, -1, -2, -1, -2, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -2, -4, -3, -2, -2, -1, -3, -1, -1, -2, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, -1, -3, -2, -2, -3, -3, -3, -2, -2, -1, -1, -2, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, -2, -1, -2, -1, -2, -1, 0, 0, -1, -1, -2, -2, -1, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -1, -2, -1, -1, -1, 0, 0, -2, -2, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, -1, -2, -1, -1, -3, -1, -1, -1, -1, -1, -2, 0, 0, -1, -1, -1, 0, 0, -2, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -2, -2, -2, -2, -2, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, -3, -2, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, -2, -3, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 1, 2, 0, 1, 1, 1, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 2, 0, 0, 0, 0, 1, 0, 0, 2, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 2, 1, 2, 1, 1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 1, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 1, 1, 2, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 1, 1, 3, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 2, 1, 1, 1, 1, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 2, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 2, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 3, 3, 3, 2, 2, 1, 1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 1, 2, 2, 2, 1, 2, 2, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 2, 2, 2, 2, 2, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 2, 2, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -2, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, -2, -2, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, 2, 0, 2, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, -1, -1, -2, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 2, 1, 2, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 2, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, -1, -1, -1, 0, -2, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, -1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 1, 0, 1, 1, 3, 3, 2, 1, 2, 1, 0, 0, 0, 0, 1, 0, -1, -2, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 0, 2, 1, 1, 1, 2, 1, 0, 1, 2, 0, 2, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 2, 1, 1, 1, 1, 0, 1, 0, 2, 1, 2, 3, 1, 2, 2, 3, 1, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 2, 1, 1, 4, 4, 4, 2, 3, 4, 3, 3, 3, 1, 1, 2, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 3, 2, 3, 4, 4, 3, 3, 2, 2, 3, 2, 1, 1, 2, 1, 2, 1, 0, 0, -1, 0, -1, 0, 0, 1, 0, 1, 0, 1, 1, 0, 3, 2, 3, 2, 4, 3, 3, 3, 2, 1, 3, 2, 3, 2, 3, 2, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 3, 4, 4, 2, 3, 3, 1, 3, 3, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 2, 0, 2, 2, 2, 3, 3, 2, 0, 1, 2, 2, 1, 3, 3, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 1, 2, 2, 2, 1, 2, 1, 0, 0, 0, 0, 1, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 3, 0, 1, 0, 0, 0, -1, -1, 0, 1, 1, 2, 2, 1, 0, 1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 0, -2, -3, -2, -1, -1, -1, 0, 0, 1, 1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, -1, 0, 0, -1, -2, -3, -3, -3, -1, -1, 0, 1, 2, 0, 0, 0, -1, -3, -2, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -2, 0, -1, -2, -3, -3, -3, -4, -4, -3, -2, -2, -1, 1, 0, 1, 0, -1, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -5, -5, -5, -4, -3, -4, -3, -3, -2, -2, 0, 0, 0, 0, -1, -1, -2, -1, -3, -2, -1, -2, 0, 0, 0, -1, 0, 0, -1, -2, -2, -4, -4, -6, -5, -4, -4, -3, -1, -2, -3, -3, -2, 0, 0, 0, 0, -1, -2, -1, -2, -1, -1, -2, -1, -1, 0, -1, -1, 0, 0, -1, -3, -4, -6, -5, -4, -5, -5, -4, -3, -2, -2, -3, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, -3, -5, -4, -3, -4, -3, -3, -2, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, -4, -4, -4, -5, -4, -4, -4, -3, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, -2, -1, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, -3, -3, -3, -3, -5, -4, -3, -3, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, -1, -1, -1, 0, -1, 0, 0, 1, -1, 0, -1, -1, -1, -1, -3, -3, -2, -3, -4, -3, -2, -2, -1, 0, 0, 1, 1, 0, 1, 0, -1, -1, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -2, -2, -1, -2, -2, -3, -2, -2, -1, 0, 0, 1, 1, 0, 1, 0, 0, -1, -2, -3, -2, -1, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -3, -3, -1, 0, 2, 2, 1, 2, 2, 0, 0, 0, -2, -1, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 1, 2, 2, 0, 0, -1, -2, -2, 0, 1, 3, 3, 3, 1, 1, 0, 0, 0, -1, -1, -1, 0, -2, 0, 0, -1, -1, -1, -1, 0, 1, 1, 3, 2, 2, 2, 1, 0, 0, 0, 1, 1, 2, 4, 2, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 3, 4, 3, 3, 2, 1, 0, 2, 1, 1, 2, 3, 3, 2, 2, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 1, 1, 2, 3, 2, 3, 2, 3, 1, 1, 1, 1, 2, 1, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 2, 2, 1, 2, 2, 2, 2, 2, 2, 3, 3, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 2, 0, 1, 1, 2, 2, 1, 2, 2, 2, 3, 3, 3, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 2, 2, 2, 2, 2, 0, 2, 1, 0, 1, 1, 2, 1, 1, 2, 1, 2, 2, 3, 1, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 1, 1, 3, 2, 4, 2, 2, 0, 1, 1, 0, 1, 0, 0, 1, 2, 2, 2, 1, 2, 1, 1, 0, -1, -1, -2, -2, 0, 0, 0, 1, 0, 0, 1, 1, 2, 1, 0, 1, 1, 0, 1, 0, 0, 0, 1, 2, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 2, 1, 2, 2, 1, 0, 0, 1, 0, 2, 3, 2, 2, 2, 2, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 3, 2, 1, 1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 2, 1, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 3, 1, 1, 2, 1, 1, 1, 1, 3, 2, 3, 2, 1, 1, 1, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 1, 1, 1, 3, 2, 2, 1, 3, 1, 2, 2, 2, 1, 1, 2, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 1, 1, 0, 2, 2, 1, 3, 2, 2, 2, 2, 2, 1, 1, 1, 2, 1, 1, 2, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 3, 2, 3, 3, 2, 3, 3, 3, 2, 3, 1, 1, 2, 0, 0, 2, 1, 1, 2, 2, 2, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 2, 3, 3, 3, 1, 3, 4, 3, 3, 1, 3, 1, 1, 2, 1, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 3, 2, 3, 3, 3, 3, 2, 2, 1, 1, 1, 1, 0, 0, 0, 1, 0, 2, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 3, 3, 4, 2, 2, 1, 2, 2, 2, 2, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 2, 2, 2, 2, 2, 2, 1, 2, 1, 2, 1, 1, 1, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 3, 1, 1, 2, 2, 2, 1, 1, 1, 1, 1, 2, 2, 1, 1, 1, 0, 2, 2, 2, 2, 0, 0, 0, -1, 0, 0, 0, 1, -1, -1, 1, 1, 2, 2, 1, 3, 2, 2, 1, 1, 1, 1, 2, 2, 1, 0, 0, 0, 2, 2, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 3, 1, 2, 1, 3, 3, 0, 2, 1, 0, 2, 2, 2, 0, 0, 0, 1, 2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 2, 4, 2, 3, 2, 1, 1, 1, 1, 1, 0, 0, 0, 2, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 2, 2, 3, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 3, 3, 1, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 2, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, -1, -1, 0, -1, -1, -1, -1, -1, -1, -2, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, -2, -2, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -2, -2, -1, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 1, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 2, 1, 0, 1, 1, 1, 2, 1, 2, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 1, 1, 1, 0, 1, 0, 1, 1, 0, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 2, 1, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 2, 1, 2, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 1, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 2, 1, 0, 0, 0, 0, 1, 2, 2, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 2, 1, 2, 0, 1, 1, 1, 3, 1, 3, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 1, 2, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 2, 2, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 1, 2, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -2, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 2, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, -2, -2, 0, -1, -2, 0, -1, -1, -1, -2, -1, -1, 0, 0, 1, 1, 2, 2, 3, 1, 3, 1, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, 0, 0, 0, 1, 1, 1, 1, 2, 3, 3, 2, 2, 1, 1, 0, 1, 1, 1, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, -3, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 0, 1, 0, 1, 1, 0, 2, 1, 2, 2, 4, 3, 3, 1, 1, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 1, 1, 0, 1, 1, 2, 2, 2, 0, 1, 0, 2, 2, 2, 1, 3, 2, 4, 4, 3, 3, 1, 1, 1, 1, 0, -2, -2, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 0, 0, 1, 1, 0, 1, 2, 1, 3, 2, 3, 2, 4, 3, 3, 1, 1, 0, 0, 0, -1, -1, 0, 1, 1, 1, 0, -1, 0, 0, 1, 1, 1, 1, 0, 0, 2, 2, 2, 1, 2, 0, 2, 3, 3, 3, 1, 1, 1, 1, 0, -1, -3, -1, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 1, 2, 0, 0, 1, 3, 1, 1, 1, 2, 1, 2, 2, 3, 1, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 2, 3, 2, 0, 1, 1, 0, 0, 1, 2, 1, 2, 1, 1, 0, 0, -2, -4, -2, 0, 0, 0, 0, -2, -1, -1, 0, -1, 0, 1, 1, 2, 2, 2, 1, 1, 0, 0, 0, 1, 1, 1, 2, 2, 1, 1, 0, 0, -2, -3, -2, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 1, 2, 2, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 1, 0, 0, -1, -4, -5, -1, 0, -1, 0, -2, -1, -2, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, -1, -2, -1, 0, 0, 1, 0, 1, 2, 0, 0, 0, 0, -2, -4, -3, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, -2, 0, 0, -2, -1, -2, -2, -1, -2, 0, 0, 0, 2, 0, 2, 0, 0, -2, -4, -5, -2, 0, 0, 0, -1, -1, -2, 0, 0, -1, -1, -2, -2, -1, -2, -3, -1, -3, -2, -1, -2, -1, -1, 0, 0, 1, 1, 0, -1, -2, -4, -5, -1, 0, -1, -1, -1, -1, -2, 0, -1, -1, -3, -2, -4, -3, -3, -3, -2, -2, -2, -1, -2, 0, 0, 0, 0, 1, 1, 0, 0, -2, -5, -5, -3, 0, -1, 0, -1, -1, -2, -1, -1, -1, -2, -3, -4, -3, -2, -3, -2, -2, -1, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, -2, -3, -4, -2, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, -2, -3, -3, -3, -3, -3, -2, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -3, -4, -4, -2, 0, -1, 0, 0, -1, -1, -1, 0, 0, -1, -1, -2, -2, -3, -2, -2, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, -3, -4, -6, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -2, -2, 0, -2, -2, -2, -1, -1, 1, 1, 0, 1, 0, 2, 1, 1, 0, 0, -2, -3, -4, -2, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 2, 3, 2, 2, 3, 1, 0, 0, -3, -4, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 1, 1, 2, 1, 2, 3, 1, 0, 0, -3, -4, -2, 0, 0, 0, 0, -2, -2, -2, -1, 0, 0, 1, 0, 2, 1, 1, 0, 0, 0, -1, 0, 1, 2, 2, 2, 2, 2, 1, 1, 0, -3, -3, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 1, 1, 2, 0, 1, 0, 0, 0, 1, 1, 1, 2, 1, 1, 1, 1, -1, -3, -4, -1, 0, 0, 0, 0, 0, -1, -2, 0, 0, 1, 1, 0, 2, 2, 2, 3, 1, 2, 0, 2, 1, 2, 2, 1, 1, 1, 0, 0, 0, -2, -3, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 2, 2, 1, 1, 2, 3, 2, 1, 1, 1, 3, 3, 2, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 1, 0, 1, 2, 0, 1, 1, 2, 2, 2, 1, 2, 2, 2, 1, 0, 0, 0, 0, -2, -2, -1, 0, 0, 1, 0, 0, 0, 1, 2, 1, 1, 0, 0, 1, 0, 0, 2, 2, 2, 3, 3, 2, 3, 2, 1, 2, 1, 0, 0, -1, -2, -3, -1, 0, 0, 2, 0, 0, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, 1, 0, 1, 2, 1, 2, 1, 2, 2, 1, 0, 0, -1, 0, -1, -1, -1, 0, 2, 3, 1, 2, 1, 1, 1, 1, 2, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -2, -2, -2, -2, -3, 0, 0, 1, 2, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -2, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -1, -2, -2, -2, -1, -2, -2, -3, -2, -2, -1, -2, -2, -1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 1, -2, 0, 0, -1, -2, -1, -2, -2, -1, -2, -1, -2, -3, -1, -2, -1, -2, -3, -2, 0, 0, 0, 0, -2, -1, 0, 0, 0, -1, 0, 0, 2, -2, 0, 0, -2, -2, 0, -2, -1, -2, -2, -2, -1, -3, -2, -1, -1, -2, -1, -2, -1, 0, -1, -1, -1, -1, -1, 0, 0, -1, 0, 1, 0, -1, 0, 0, -1, -2, -1, 0, -1, -2, -2, -1, -1, -2, -1, -2, -1, -1, -2, -1, -1, 0, -1, 0, -1, -1, 0, 0, -1, 0, -1, 0, 1, -1, 0, 0, -1, 0, 0, -1, 0, -2, -2, -2, -1, -1, -2, 0, -2, -2, -1, -1, -1, 0, 0, -1, -1, -2, -1, -1, 0, -1, -2, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, -2, -3, 0, -1, -2, -1, -2, -3, -2, -1, -2, -1, 0, -1, -1, -1, -1, 0, -2, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, -2, -1, -2, -2, 0, -2, -4, -2, 0, 0, 0, 1, -1, -1, 0, -1, -1, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -2, -1, 0, -1, -4, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 1, 0, 0, -2, 0, 0, 0, 0, 0, -2, -2, 0, -1, -1, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, -2, 0, -1, 1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -2, 0, 0, 0, 0, -1, -1, -1, 0, 1, 1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, -1, -2, -1, 1, 2, 1, 2, 2, 0, -2, 0, -1, -1, -1, 0, 1, 0, 0, 1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -3, 0, 2, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, -3, -2, 0, 1, 2, 1, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, 1, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, -2, -1, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 2, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -2, -2, 0, -1, 0, 0, -2, 0, 0, -1, 0, 0, 0, 1, 0, 0, -2, -2, -1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -3, -1, 0, 0, 0, -1, -3, -2, 0, 0, 0, 0, 0, 1, 0, 0, -3, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -4, -1, -1, 0, 1, -1, -3, -2, -1, -2, 0, -1, 1, 0, 0, 0, -2, -3, -1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, -1, -3, -1, -1, 0, 0, -1, -3, -2, -2, -1, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, -2, -1, -1, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, -2, -3, -2, -2, -2, -2, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -2, -1, 0, 1, 2, 1, 0, 0, -1, 0, 0, 0, 0, -3, -2, -3, -3, -2, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -2, 0, -1, 0, 1, 1, 0, 0, -2, 0, 0, 0, -1, -2, -2, -2, -2, -2, -3, -2, -3, -1, -2, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, 2, 1, 0, 0, -1, 0, 0, 0, -1, -1, -2, 0, -2, -3, -2, -2, -3, -3, -2, -1, 0, -1, 0, 0, -2, 0, -1, 0, 0, 0, -1, 0, 1, 1, 0, -1, 0, 0, 0, -1, -1, -1, -1, -2, -2, -4, -3, -3, -2, -3, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, -2, -3, -2, -1, -1, -2, -2, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -2, -2, -1, -1, -2, -2, -2, -1, 0, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -2, -1, 0, 0, -2, -2, -1, -2, 0, -2, -2, -1, -1, -1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, 1, -2, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -3, -1, -1, -2, 0, -2, 0, 0, 0, 2, 2, 1, 1, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, -2, -2, -1, -1, -2, -3, -2, -2, -1, -2, -2, -1, 0, 1, 2, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 2, 1, 0, -1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 2, 2, 2, 1, 1, 1, 1, 0, -1, 0, -1, -1, 0, 0, 0, -2, -2, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, -1, -3, -3, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 2, 2, 2, 1, 2, 2, 1, 0, -2, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 1, 0, 0, 0, 0, -1, -1, 0, 1, 2, 2, 2, 2, 1, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 2, 1, 2, 0, 0, 0, -1, -1, 0, 1, 0, 1, 0, 0, 0, -2, -2, -3, -1, -2, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, -2, -1, -1, 0, 1, 2, 1, 0, 0, 0, -1, -2, -2, -2, -1, -2, -2, -1, 0, 0, 1, 0, 1, -1, 0, -1, 0, 1, 0, 1, 0, 0, 0, -2, -2, -1, 0, 0, 1, 0, 0, 1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 2, 2, 1, 1, 0, -1, -1, 0, -1, -1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -2, 0, 0, -1, -1, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, 0, -2, 0, 0, 0, -2, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, -1, -2, 0, -1, -1, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, -1, -1, -2, -2, -2, -2, 0, 0, 1, 2, 1, 2, 0, 1, 0, -1, -1, -2, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, -1, 1, 0, 0, -2, -2, -2, -2, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, -2, -1, -1, 0, 1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -2, -1, 0, 0, 1, 0, -1, -2, 0, -2, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, -1, -2, -2, -2, -1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, -2, -1, -2, -3, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, -1, 0, 0, 1, 1, 0, 0, 1, 2, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -2, -1, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 2, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -3, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 2, 2, 2, 1, 2, 1, 1, 2, 1, 0, 1, 1, 1, 0, 0, 0, 1, 2, 1, 0, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 1, 1, 0, 0, 0, -1, -1, -2, -1, -1, -1, -2, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, -1, -1, -2, -2, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, -1, 0, -1, -2, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, -1, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, -1, -2, 0, -1, -1, -1, -1, -1, -1, -1, -2, -2, -2, -2, -3, -1, -1, -1, -2, 0, -1, 1, 0, 1, 1, 1, 1, 2, 0, 1, 0, 0, 0, 0, -2, 0, -1, -2, -2, -1, 0, -1, 0, 0, -1, -2, -2, -1, -2, -1, -2, -1, 0, 1, 0, 1, 2, 1, 3, 2, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 1, 3, 3, 3, 2, 2, 2, 0, 1, 0, 1, 0, 1, 1, 1, 3, 2, 2, 2, 2, 1, 0, 1, 0, -1, -2, -1, -2, 0, 0, 1, 1, 2, 2, 1, 1, 1, 1, 1, 1, 0, 0, 2, 1, 3, 3, 3, 4, 4, 4, 3, 2, 2, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 2, 3, 3, 3, 3, 4, 3, 5, 4, 4, 2, 1, 2, 1, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 2, 0, 0, 1, 2, 3, 2, 4, 3, 1, 4, 5, 4, 3, 4, 2, 2, 0, 1, 0, -2, -2, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 1, 0, 2, 2, 2, 2, 3, 2, 1, 1, 3, 4, 3, 4, 4, 2, 1, 1, -1, -3, -2, -2, 0, 0, -1, -1, -1, 0, -1, -1, 0, 2, 2, 2, 2, 3, 4, 3, 2, 1, 0, 0, 1, 2, 3, 4, 3, 3, 1, 1, -1, -3, -3, -1, 0, 0, -1, -1, -1, -1, -1, -1, 0, 1, 2, 4, 3, 4, 3, 1, 1, 1, 1, 1, 0, 1, 3, 2, 2, 2, 0, 0, -2, -4, -3, -2, 0, 0, -2, -3, -2, -1, -1, 0, 0, 1, 2, 4, 3, 4, 4, 0, 0, 0, 0, 1, 0, 0, 1, 2, 2, 1, 1, -1, -3, -4, -3, -3, -1, -1, -2, -1, -1, -1, -1, -1, 0, 0, 0, 2, 3, 3, 2, 0, -1, 0, 0, 0, 1, 1, 1, 1, 2, 2, 0, -1, -4, -5, -3, -3, 0, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 1, 0, 0, 1, 2, 1, 1, 0, -1, -3, -5, -3, -3, 0, -2, -2, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -4, -6, -4, -3, 0, -2, -1, -2, -2, -2, -3, -1, -1, -1, -2, -2, -3, -2, -4, -2, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -4, -6, -3, -2, -1, -1, -3, -2, -2, -3, -3, -2, 0, -2, -4, -5, -4, -2, -4, -3, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -3, -4, -6, -4, -3, 0, -1, -2, -1, -2, -3, -2, -2, -1, -3, -4, -5, -5, -3, -2, -3, -3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -4, -6, -3, -2, 0, -1, -1, 0, 0, -1, -1, 0, 0, -2, -2, -4, -5, -3, -1, -1, -1, 0, 0, 0, 1, 1, 1, 1, 1, 2, 1, -2, -4, -5, -5, -4, 0, 0, -1, 0, 0, 0, -1, -1, 0, -2, -2, -4, -3, -1, -2, 0, -1, -1, 0, 0, 0, 0, 1, 2, 2, 2, 1, -1, -6, -6, -3, -3, 0, -1, 0, -1, 0, -1, -1, 0, -1, -2, -1, -1, -3, -1, -1, -1, 0, 0, 0, 0, 1, 1, 2, 4, 3, 2, 1, -1, -4, -5, -4, -3, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 4, 3, 2, 1, -1, -4, -4, -2, -3, 0, -1, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, -1, 0, 1, 2, 3, 3, 4, 2, 1, -1, -2, -5, -2, -3, 0, 0, 0, -2, -1, -2, -3, -1, 0, 0, 1, 1, 1, 2, 2, 2, 1, 0, -1, 0, 2, 2, 2, 3, 3, 3, 1, 0, -2, -3, -3, -2, 0, 0, -1, -1, -2, -1, -2, 0, 0, 1, 0, 1, 2, 2, 1, 1, 0, 0, 0, 1, 1, 2, 1, 2, 3, 2, 1, -1, -2, -5, -2, -2, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 2, 1, 3, 2, 2, 3, 2, 0, 1, 1, 2, 0, 2, 2, 0, -2, -2, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 1, 2, 2, 2, 2, 1, 1, 3, 1, 1, 2, 0, 0, 0, -1, -3, -3, -1, -1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 1, 1, 1, 1, 2, 2, 2, 3, 2, 2, 2, 2, 0, 0, 0, 1, 0, -1, -3, -3, -2, 0, 1, 0, 1, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 3, 2, 1, 2, 1, 1, 0, 0, -2, -2, -4, -1, -2, 2, 1, 0, 1, 1, 1, 2, 1, 1, 2, 1, 0, 0, 1, 0, 1, 2, 0, 1, 2, 2, 1, 0, 2, 0, 1, -1, -2, -4, -4, -2, -1, 1, 1, 1, 2, 2, 2, 2, 1, 2, 2, 0, 0, -1, 0, 1, 0, 1, 0, 1, 1, 1, 1, -1, -1, 0, -1, -1, -3, -2, -3, -1, -2, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -2, -2, -1, -2, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, 0, 0, -1, -1, 0, 0, -1, -2, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 2, 1, 2, 2, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 3, 0, 0, 0, 0, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 3, 1, 0, -1, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 1, 0, 0, 1, 1, 0, 2, 1, 1, 0, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 3, 2, 1, 1, 0, 0, 2, 1, 1, 1, 2, 2, 2, 1, 0, 0, 0, 1, 2, 1, 1, 0, -1, 0, 1, 0, 0, 0, 2, 0, 1, 1, 2, 1, 1, 2, 1, 1, 1, 1, 1, 1, 2, 2, 2, 1, 1, 0, 1, 0, 1, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 1, 3, 2, 2, 3, 2, 1, 1, 1, 1, 1, 2, 1, 0, 0, 2, 3, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 2, 0, 1, 2, 2, 1, 1, 2, 2, 1, 1, 1, 1, 1, 1, 0, 0, 2, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 1, 1, 3, 2, 2, 2, 2, 3, 1, 2, 1, 0, 1, 2, 0, 1, 1, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 3, 3, 3, 2, 2, 4, 2, 3, 3, 2, 1, 1, 1, 1, 0, 1, 2, 1, 1, 1, 3, 2, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 2, 3, 3, 3, 3, 2, 3, 2, 3, 3, 2, 1, 1, 2, 1, 1, 1, 1, 0, 0, 2, 0, 0, 0, -2, 0, 0, -1, 0, 0, 1, 1, 1, 3, 1, 2, 2, 3, 2, 2, 2, 0, 1, 0, 0, 2, 1, 0, 1, 1, 0, 0, 1, 1, 0, -1, -2, 0, 0, -1, 0, 0, 0, 0, 2, 1, 1, 3, 3, 2, 3, 2, 1, 2, 0, 1, 0, 1, 1, 1, 0, 1, 1, 1, 1, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 1, 2, 3, 2, 1, 3, 3, 2, 2, 2, 1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 2, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 2, 1, 4, 4, 4, 2, 0, 1, 0, 0, 0, 2, 1, 0, 0, 0, 1, 1, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 2, 2, 1, 3, 4, 2, 3, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 1, 2, 3, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 2, 1, 1, 2, 3, 2, 2, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 3, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 2, 2, 1, 1, 0, 2, 1, 0, 0, 0, 0, 1, 3, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 2, 2, 1, 0, 0, 1, 0, 1, 0, 1, 1, 1, 2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 2, 1, 0, 0, 1, 1, 1, 0, 1, 0, 2, 0, 0, 0, -1, -1, -1, 0, -2, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 2, 2, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 2, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, -1, -2, 0, -1, 0, -1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, -1, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, 2, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 1, 1, 0, 1, 1, 1, 3, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 2, 1, 1, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, -1, -1, 0, 0, 1, 1, 2, 2, 2, 0, 0, 1, 0, -1, 0, 1, 0, 1, 1, 0, -1, 0, 0, 0, 0, 1, 2, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 1, 2, 1, 2, 0, 1, 0, 0, -1, 0, 0, 2, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, -1, -1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, -2, 0, -1, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 1, 1, 1, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 1, 1, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 2, 1, 3, 2, 0, 0, 0, 2, 3, 4, 1, 1, 1, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 2, 3, 2, 3, 2, 1, 0, 0, 1, 3, 2, 1, 2, 2, 1, 1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 1, 2, 1, 3, 2, 2, 0, 1, 1, 2, 2, 2, 3, 2, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, 2, 1, 0, 0, 0, 1, 2, 3, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 1, 2, 2, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 2, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 1, 2, 0, -1, -1, 0, -2, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 1, 0, 1, 1, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 1, 0, -1, -1, -1, -1, -1, 0, 0, 0, -1, 1, 0, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -2, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, -2, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, -1, 0, -2, -2, 0, -1, -1, -2, 0, -2, -1, -1, 0, 0, 0, 3, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, 0, 0, -1, -1, -2, -1, -2, -1, -1, -1, -2, -3, -1, -1, 0, 0, 0, 0, 1, 2, 2, 1, 1, 1, 1, 3, 2, 1, 0, -1, -1, 0, 0, 2, 1, 0, -1, -2, -1, 0, 0, 0, 0, -1, -2, -1, -2, -2, 0, 0, 2, 3, 2, 2, 3, 1, 2, 3, 2, 3, 2, 1, 0, 0, 0, 2, 3, 1, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 2, 3, 3, 2, 2, 1, 4, 3, 1, 1, 0, 0, 0, 0, 1, 2, 0, 1, 2, 1, 1, 1, 1, 0, 1, 1, 0, 0, -1, 0, 0, 1, 1, 1, 2, 1, 0, 1, 2, 3, 2, 1, 0, 0, 1, 0, 0, 2, 0, 2, 2, 3, 3, 2, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 2, 2, 1, 1, 0, 1, 1, 1, 0, 1, 0, 1, 2, 3, 3, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 1, 0, 1, 1, 1, 0, 0, 1, 1, 0, 1, 0, 1, 1, 2, 2, 2, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 2, 3, 2, 2, 1, 0, 0, 0, 1, 1, 0, 0, -2, 0, 1, 2, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 2, 3, 2, 3, 3, 3, 0, 1, 1, 0, 1, 0, 0, -2, 0, 1, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 4, 3, 3, 2, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, -2, -2, 0, 0, 0, 0, 0, -1, 0, -2, 0, 1, 3, 3, 3, 2, 2, 1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, -1, -2, -2, -1, -2, -1, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 3, 3, 3, 3, 2, 0, 0, 0, -1, 0, -2, 0, 1, 1, 0, 0, -2, 0, -1, -1, -1, -3, -2, -2, 0, -2, -2, -1, -2, -1, 0, 0, 2, 4, 4, 3, 2, 1, 1, 0, 0, -1, -2, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -2, -2, -2, -2, -1, -2, -1, -2, -1, -2, 0, 2, 3, 4, 2, 2, 2, 1, 0, 0, -2, -2, -1, 0, 0, 0, -2, 0, -1, -1, -1, 0, -3, -1, -2, -3, -3, -3, -1, -1, -1, -1, 0, 1, 1, 3, 2, 3, 2, 1, 1, 0, -2, -2, -1, 0, 1, 0, -2, -1, 0, 0, -1, 0, -1, -3, -2, -3, -3, -4, -2, -1, 0, -1, 0, 0, 1, 2, 1, 2, 2, 1, 1, 0, -1, 0, -2, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, -1, -2, -2, -4, -2, 0, 0, 0, -1, 1, 1, 1, 2, 1, 1, 2, 1, 0, -1, -1, -1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, -2, 0, -2, -3, -3, -3, 0, 0, 0, 0, 1, 1, 2, 0, 2, 1, 1, 2, 0, 0, -2, -1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, -2, -2, -3, -3, -2, 0, 0, 1, 2, 1, 0, 0, 1, 2, 1, 0, 0, 0, -1, -1, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, -3, -3, -2, 0, 1, 1, 1, 1, 0, 1, 1, 3, 2, 2, 0, -1, 0, -1, 0, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, -3, -2, 0, 1, 2, 2, 2, 1, 1, 1, 1, 2, 2, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, 1, 2, 1, 0, 0, 0, 1, 2, 2, 1, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, -2, -1, 0, 0, 2, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 1, 2, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 1, 2, 1, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 2, 3, 1, 2, 1, 0, 1, 2, 1, 1, 3, 2, 2, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 2, 1, 0, 1, 1, 1, 2, 2, 2, 1, 1, 1, 0, 2, 2, 2, 3, 2, 2, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 1, 1, 0, 1, 2, 2, 1, 2, 1, 0, 0, 0, 0, 2, 1, 1, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 3, 2, 2, 2, 3, 1, 0, 0, 0, -1, 0, 1, 1, 1, 1, 2, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, 1, 3, 4, 4, 2, 3, 3, 4, 1, 2, 1, 1, -1, 0, -1, 0, 1, 2, 0, 1, 1, 1, 1, 2, 0, 0, 0, 0, 0, 1, 1, 0, 2, 3, 4, 4, 2, 3, 3, 2, 2, 1, 1, 1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 2, 2, 3, 2, 1, 3, 2, 1, 2, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 0, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 1, 1, 2, 0, 0, 0, 1, 1, 0, 0, 0, -3, -3, -3, -3, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, -2, -4, -2, -4, -4, -3, -3, -2, -1, -1, -1, -1, 0, 0, 0, -2, 0, -1, -1, 0, -1, -2, -2, -2, -1, -1, -2, 0, -1, 0, 0, 3, 0, -2, -2, -3, -2, -2, -3, -3, -2, -1, -2, -1, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -3, -2, -2, -1, -1, 0, -2, 0, 0, 2, 0, -2, -3, -2, -2, -1, 0, -1, -1, -2, 0, -1, 0, -1, -1, -2, -1, 0, -1, 0, -2, -2, -1, -1, -2, -1, -1, 0, 0, 0, 0, 1, -1, -2, -1, -3, -2, -1, -1, -1, -3, -2, -2, -1, -1, -1, 0, -2, -2, -1, 0, -1, -2, -1, -2, -1, -2, -1, -1, 0, -1, 0, 0, 1, -2, -1, 0, -2, -2, 0, 0, -1, -1, -2, 0, -1, -2, 0, 0, -1, -2, -1, -2, 0, -1, -2, -3, -2, -1, 0, 0, -1, -1, 0, 0, 2, -1, -2, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, -2, -1, -2, -1, 0, -2, -2, -2, -2, -2, -1, -1, -1, -1, 1, 2, -1, -2, -1, -1, 0, -1, 0, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -2, -3, -3, -1, -2, 0, -2, 0, 0, 1, 3, -1, -2, -3, 0, 0, 0, -1, -1, -2, -2, -3, -3, 0, -1, -2, -1, 0, -1, 0, 0, -2, -2, -3, -4, -3, -1, 0, 0, -1, 0, 1, 1, -1, -3, -3, -1, 0, 0, -1, -1, -2, -1, -3, -4, -2, -2, -1, -1, 0, 0, 0, -1, 0, -1, -2, -3, -3, 0, 0, 0, -1, 0, 0, 2, -1, -2, -1, -1, -1, -2, -2, -1, 0, -2, -3, -6, -3, -3, -1, -1, 0, 0, 1, 0, 0, -2, -2, -3, -2, 0, 0, -1, -1, 0, 0, 2, -1, -3, -3, -1, 0, -1, -3, -2, -1, -1, -3, -4, -3, -1, -1, 0, -1, -1, 0, 0, -1, -2, -2, -3, -2, -2, 0, 0, 0, -1, 0, 1, 0, -3, -3, -2, 0, 0, -1, -1, 0, 0, -1, -2, -1, 0, 0, -2, -2, -3, -1, -1, -2, -2, -3, -1, -1, -3, -1, 0, -2, 0, 0, 1, 0, -1, -1, -2, 0, 0, -1, -1, 0, -1, 0, -2, -2, 0, -1, -1, -2, -2, -1, 0, 0, -2, -2, -2, -2, -3, -2, -2, -3, -1, 0, 2, 0, -1, -1, -1, 0, 0, -2, -1, 0, -1, -2, -1, -2, 0, 1, 0, -3, -3, -2, 0, -1, -2, -2, -2, -3, -2, -2, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -2, -1, -2, -1, 0, 0, 0, 1, -1, -1, 0, -2, -2, -2, -2, -1, -2, -2, -1, -2, 0, 0, 0, 1, 0, -2, 0, 0, 0, 0, -1, 0, -1, -2, -1, 0, 0, 0, 2, 1, 0, 0, -1, 0, -1, -3, -3, -2, -1, -1, -1, -2, -2, 0, 1, 2, 0, -2, -2, 0, 0, -1, -1, -1, 0, 0, -2, 0, 0, -1, 2, 2, 0, 0, 0, -2, -1, -3, -3, -2, -2, -1, 0, 0, 0, 0, 0, 2, -1, -1, -2, -1, -1, 0, -1, -1, 0, 0, -1, -2, 0, 0, 0, 2, 1, 0, -1, -1, -3, -3, -4, -3, -1, -2, 0, -1, -1, 0, 0, 3, -1, -1, -2, -1, 1, 0, -1, 0, 0, 0, -1, -1, -1, -2, 0, 2, 0, -1, 0, -3, -3, -2, -4, -3, -1, -2, -2, -2, -1, -1, 0, 2, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, 1, 2, 1, 0, -2, -2, -2, -3, -3, -1, -1, -1, -2, 0, 0, 0, 2, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 1, 1, 0, 0, -1, -1, -2, -1, 0, 0, 0, -1, -1, -1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, -3, -3, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, -1, -2, -1, 0, 0, 0, 0, 1, 1, 0, -1, -1, -1, -2, -1, -1, -3, -1, -1, -1, -2, -2, 0, 1, 0, 1, 0, -1, 1, 0, 3, -1, 0, 0, -1, 0, -1, -2, -1, 0, 0, 0, -1, -1, 0, -2, -2, -2, -2, -3, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -2, -1, -1, 0, 0, -2, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -2, -2, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 2, 0, 0, -1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 3, 0, -1, -2, -2, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 3, 0, 0, -1, -2, 0, -2, -3, -2, -2, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 3, 1, 0, 0, -1, 0, -1, -2, -1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 1, 0, 1, 1, 2, 0, 0, 1, 1, 3, 3, 1, 2, 1, 2, 2, 1, 1, 2, 2, 2, 1, 1, 1, 1, 0, 0, 0, 0, 2, 1, 1, 1, 0, 1, 3, 2, 1, 1, 1, 1, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 1, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 1, 1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 2, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, -1, -2, -1, 0, -1, -2, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, -2, 0, 0, 0, 0, -1, 0, 1, 2, -2, 0, 0, -1, -2, -2, -3, -2, -3, -4, -2, -1, -2, -3, -2, -2, -3, -1, -2, 0, 0, 0, 0, -1, -3, -1, 0, 0, 0, 0, 0, 2, -4, 0, 0, -4, -3, -1, -2, -3, -2, -3, -2, -2, -3, -4, -1, -1, -3, -2, -4, -1, 0, -1, -1, -1, -3, -2, 0, 0, -1, 0, 0, 1, -2, 0, 0, -3, -2, -1, -2, -2, -2, -2, -1, -2, -2, -3, -2, -3, -2, -3, -4, -1, -1, 0, -2, -2, -2, -1, -2, -1, -3, -1, 0, 2, -1, 0, 0, -4, -2, -2, -2, -1, -2, -3, -3, -2, -3, -2, -1, -3, -3, -2, -2, -1, 0, 0, -1, -1, -1, -2, -1, -1, -1, -1, 0, 1, -1, 0, -1, -3, -1, -1, -1, -2, -3, -3, -1, -3, -3, -1, -2, -4, -3, -1, -3, -2, -1, -1, -3, 0, -2, -1, -3, -1, -1, -2, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, -4, -3, -2, -1, -2, -2, -3, -6, -4, -2, -1, -1, 0, -1, -1, -1, -2, -2, -2, -1, 0, -2, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, -3, -3, -1, -1, 0, -1, -2, -5, -4, -3, 0, 0, 1, 0, -2, 0, -2, -2, -2, -2, -2, -2, -1, 0, 2, -1, -1, -1, 0, -1, 0, 0, -1, -3, 0, -1, 0, 0, -1, -6, -3, -2, -1, 0, 1, 0, -1, 0, -2, -3, -3, -3, -1, -2, 0, 1, 2, 0, -1, 0, 1, 0, 0, 0, -2, -2, -2, 0, 0, 0, -1, -5, -2, -1, -2, -1, -1, 0, 0, -1, 0, -1, -2, -2, -2, -2, 0, 1, 1, 0, 0, -2, 0, 0, 0, 0, -1, -3, -3, 0, 0, -2, -3, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, -3, -3, -2, -1, 1, 0, 0, -2, -2, 0, 0, 2, 0, 0, 0, -2, -1, 0, -1, -2, -1, -1, -2, -1, -1, 0, -1, 1, 0, 0, 0, 0, -1, -2, -3, 0, 1, 0, 0, -1, -3, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, -3, -2, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, -1, 0, 1, 0, 0, 0, -3, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, -3, -1, -1, -2, -2, 0, 0, 0, 0, 2, 0, -1, 0, 0, -1, -1, -1, 1, 0, 0, 0, -2, 0, -1, -3, -2, 0, 2, 2, 1, 2, 0, -1, -1, -1, -3, -1, -1, 0, -1, 0, 0, 1, -2, -2, 0, -1, -1, -2, 1, 1, 0, 0, -3, 0, 0, -3, -4, 0, 1, 2, 2, 2, 0, 0, 0, -2, -1, -1, -1, 0, 0, 0, 1, 0, 0, -2, 0, 0, -2, -2, 0, 2, 0, -1, -3, 0, -1, -3, -3, -1, 1, 2, 3, 1, -1, 0, -1, -1, -1, -1, -3, -2, 0, -1, 1, 1, 0, 0, -1, -1, -2, -1, 1, 1, 0, -1, -3, -1, 0, -1, -1, 0, 0, 1, 2, 1, 0, 0, 0, -1, -1, -1, -2, -1, 0, 0, 0, 1, 0, 0, -1, -1, -2, 0, 1, 0, 0, 0, -2, 0, -1, 0, 0, -1, -2, 0, 2, 0, 0, 1, 2, 0, 0, -1, -2, -3, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 2, 0, 0, -1, -3, -2, 0, 1, 1, 0, -3, -1, 0, 0, 0, 3, 3, 1, 1, -1, -3, -4, -3, -1, 0, 2, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -4, -2, -2, 0, 1, 0, -3, -2, -1, 0, 0, 1, 3, 2, 1, 0, -4, -3, -1, -2, 0, 0, 0, -2, -2, 0, 0, 0, 3, 1, 0, -1, -5, -1, 0, 0, 2, -1, -4, -4, -5, -3, -1, 0, 2, 2, 2, 1, -1, -2, -2, -1, 0, -1, -1, -2, -3, 0, 0, 1, 2, 1, 0, 0, -3, -2, -1, 0, 0, -1, -3, -4, -4, -2, -2, -1, 0, 1, 1, 1, 0, 0, -1, 0, 0, -1, 0, -1, -3, -1, 0, 0, 3, 1, 0, -1, -2, -2, 0, 0, 0, -3, -3, -5, -4, -2, -2, -1, -1, 0, 0, 1, 1, 0, -1, -1, 0, 0, 0, 0, -3, -2, 0, 0, 2, 2, 0, -1, -2, 0, 0, 0, 0, -3, -2, -3, -5, -4, -4, -2, -3, -2, 0, 0, 2, 0, 0, -1, -1, 0, 0, 0, -1, -2, 0, -1, 2, 2, 0, 0, -1, -1, -1, -1, -1, -3, -1, -2, -5, -4, -5, -5, -5, -3, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -2, -1, 0, 2, 2, 0, 0, -1, 0, 0, -2, -2, -2, -2, -2, -4, -5, -4, -4, -5, -4, -3, -1, -1, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, 1, 2, 0, 0, 0, 0, -1, -2, -4, -2, -3, -2, -2, -4, -3, -3, -3, -5, -4, -2, -1, -2, 0, -1, -2, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -3, -4, -2, -1, -1, -3, -5, -3, -2, -2, -3, -4, -1, -1, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -4, -1, 0, -1, -3, -3, -1, -2, -2, -2, -2, -1, -1, -1, -3, -1, -2, -1, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -2, -2, 0, 0, -1, -1, -2, 0, -1, -1, -3, -1, 0, -1, -1, -1, 0, 0, 1, 1, 0, 1, 0, 0, 1, -1, 0, 0, -1, -1, 0, 0, -1, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 1, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 2, 0, 0, 0, 0, 1, 2, 1, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 1, 0, 0, 0, 0, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 2, 2, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 2, 2, 2, 1, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 1, 1, 0, 2, 1, 1, 1, 3, 2, 0, 2, 1, 2, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 2, 3, 3, 2, 1, 2, 2, 3, 3, 2, 1, 1, 2, 3, 1, 2, 0, 1, 1, 1, 2, 2, 1, 1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 1, 2, 2, 2, 1, 3, 3, 1, 1, 2, 1, 1, 1, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 2, 0, 1, 1, 1, 1, 1, 1, 3, 2, 3, 2, 2, 3, 2, 3, 2, 2, 2, 2, 2, 3, 2, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 2, 2, 2, 2, 2, 2, 3, 1, 1, 2, 3, 2, 2, 3, 2, 2, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 1, 2, 3, 2, 4, 3, 2, 2, 1, 2, 2, 1, 2, 1, 1, 2, 2, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 3, 3, 2, 4, 3, 3, 1, 2, 2, 1, 2, 1, 1, 1, 1, 1, 2, 2, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 2, 2, 2, 3, 4, 3, 2, 4, 2, 1, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 3, 2, 3, 3, 2, 3, 2, 1, 1, 1, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 2, 2, 3, 2, 3, 3, 3, 2, 1, 0, 1, 1, 1, 0, 1, 0, 0, 1, 1, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 3, 3, 3, 2, 3, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 2, 3, 3, 3, 3, 3, 2, 1, 2, 1, 2, 2, 2, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 2, 3, 4, 2, 4, 3, 2, 0, 1, 0, 2, 1, 1, 0, 0, 1, 2, 2, 2, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 3, 4, 3, 3, 2, 1, 1, 2, 2, 0, 0, 1, 1, 3, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 3, 3, 4, 3, 3, 1, 1, 1, 2, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 2, 1, 2, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 2, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, 0, 0, -1, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -2, -1, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, 0, 0, 0, -1, 0, -1, -2, -1, -1, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, -1, -1, 0, -2, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, -2, -1, 0, -1, -1, -2, -1, -2, 1, 1, 2, 2, 3, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, -1, -2, 0, -1, -2, -1, 1, 0, 1, 1, 2, 1, 1, 1, 0, 1, 0, 1, 1, 0, 1, 0, 0, 1, 1, 0, 1, 2, 2, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 3, 1, 1, 2, 2, 1, 0, 2, 1, 0, 1, 1, 1, 1, 2, 2, 0, 1, 0, 0, -1, -2, -2, -1, -1, 0, 0, 1, 1, 2, 1, 2, 3, 3, 3, 2, 1, 1, 3, 1, 2, 2, 0, 1, 2, 3, 2, 2, 2, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 1, 1, 2, 2, 2, 3, 2, 2, 1, 0, 0, 1, 2, 3, 3, 1, 2, 1, 2, 2, 3, 2, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 1, 1, 2, 1, 2, 1, 0, 0, 1, 3, 3, 4, 3, 2, 0, 2, 1, 3, 3, 2, 2, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 2, 2, 1, 3, 2, 3, 3, 2, 1, 1, 1, 2, 3, 4, 2, 2, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 3, 3, 2, 3, 2, 3, 3, 3, 1, 1, 0, 0, 2, 2, 3, 2, 2, 0, 0, -1, 0, -2, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, 2, 3, 5, 5, 3, 4, 2, 1, 2, 0, 0, 0, 1, 1, 2, 2, 2, 1, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 4, 3, 4, 3, 2, 1, 2, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, -2, -2, -2, -2, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 2, 3, 3, 2, 1, 0, 0, 0, -1, 0, -1, -1, 1, 0, 1, 1, 1, 0, -1, -3, -2, -2, 0, 0, 1, 0, 0, 1, 1, 1, 3, 2, 1, 2, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, -1, -1, -2, -2, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -2, -1, 0, -1, 0, -1, -1, -2, 0, -1, -1, 0, -1, -1, -2, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, -2, -2, -2, -2, -1, 0, -1, -1, -1, -2, -1, -1, -1, 0, -2, -3, -4, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, -2, -1, -2, -1, -1, 0, -1, -1, 0, 0, -2, -2, -3, -4, -5, -4, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -3, -2, -1, -2, -2, -1, -2, 0, 0, -1, 0, 0, 0, -1, -1, -2, -3, -4, -3, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, -1, -1, -3, -4, -3, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -1, 0, 0, 0, 0, 1, 2, 0, 0, -1, -2, -4, -2, -2, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 1, 1, 2, 1, 1, 1, 0, -1, -2, -2, -2, 0, -1, -1, 0, -2, -1, -1, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 1, 0, -2, -2, -3, -2, -1, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 2, 3, 1, 2, 2, 2, 0, 0, 0, 0, 1, 1, 3, 2, 1, 0, 0, -1, -2, -2, -1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 2, 1, 3, 2, 4, 3, 3, 2, 1, 0, 0, 1, 0, 1, 0, 0, -1, -2, -3, -3, -3, -1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 2, 1, 3, 1, 3, 3, 2, 3, 1, 0, 0, 0, 1, 1, 0, -1, -1, -2, -3, -3, -2, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 2, 2, 2, 1, 2, 1, 0, 0, 0, 0, -1, -1, -2, -2, -3, -2, -1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 3, 2, 2, 0, 0, 0, 0, 0, 0, -1, -3, -4, -4, -3, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, -1, -2, -3, -4, -3, -2, 0, 0, 1, 1, 0, 0, 1, 1, 0, 1, 2, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -3, -4, -1, -2, 0, 0, 1, 1, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -2, -2, 0, -1, 0, -2, -3, -4, -3, -2, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -2, -2, -2, -1, -2, -2, -2, -2, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 1, 2, 2, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 1, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -2, -2, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, -2, -2, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -2, -2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -3, -2, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 1, 0, 1, -1, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, -2, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -2, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, -1, 0, -2, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, 2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -2, -2, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, -2, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, -1, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, -2, -1, 0, -1, -2, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, -1, 0, 1, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, -1, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, -2, -1, -1, 0, 0, 1, 1, 0, 1, 1, 2, 1, 0, 0, 0, 0, -1, -1, -2, -2, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 2, 1, 0, 0, 2, 2, 0, 0, -1, -2, 0, -1, 0, -1, -2, -1, -2, -1, -1, -1, -1, -1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 2, 2, 1, 1, 0, 0, 0, 0, 0, -2, 0, -1, 0, -1, -2, -2, -2, -3, -2, -1, -1, -2, -1, -1, 0, 0, 0, 1, -1, 0, -1, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -2, -1, -2, -2, -2, -1, -2, -1, -2, -2, -2, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -2, -2, -2, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -2, -3, -3, -2, -1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, -1, -3, -3, -2, -2, -3, -1, -3, -2, -2, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -2, -2, -1, -2, -2, -2, -2, 0, 0, 0, 0, 1, 1, 1, 0, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, -2, -2, -3, -2, -1, -2, -1, -1, -1, 0, -1, 0, 1, 0, 0, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, -2, -2, -2, -1, -2, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, -1, -2, -2, -3, -1, -1, -1, -1, 0, -1, -1, -1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, -1, -2, -2, -3, -3, -2, -2, 0, -1, -1, 0, 0, 0, 0, 0, 1, 2, 1, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, -2, -3, -3, -3, -2, -2, -1, 0, 0, 0, -2, -2, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -4, -2, -3, -2, -1, 0, 0, -1, -2, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -3, -3, -2, -1, 0, 0, 0, -1, -2, -2, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -3, -3, -2, -2, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -2, -2, -2, -1, 0, -1, 0, 0, -2, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, -1, -1, 0, 0, -1, 0, -2, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 2, 1, 1, 1, 2, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 2, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 2, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 2, 1, 2, 2, 0, 0, 1, 0, 1, 0, 1, 2, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 1, 1, 1, 1, 1, 2, 2, 1, 1, 2, 1, 1, 1, 2, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 1, 0, 1, 1, 1, 0, 1, 2, 2, 1, 2, 1, 1, 2, 1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 1, 1, 1, 0, 1, 0, 1, 1, 0, 1, 1, 1, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 2, 1, 2, 1, 1, 1, 0, 0, 1, 0, 1, 2, 1, 1, 0, 0, 0, -1, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 1, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -2, -2, -3, -2, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -3, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, -2, -1, -2, -2, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -3, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -2, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -2, -1, 0, -2, -1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 1, 0, 1, 2, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 2, 1, 1, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, -2, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 1, 0, 2, 2, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, 0, 1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -2, 0, 0, 2, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, -1, -2, 0, -2, 0, 0, 0, 0, 0, 4, 2, 1, 0, 0, 0, 0, 1, 0, -2, -1, -1, 0, 0, 1, 1, 0, 0, -2, 0, 0, 0, 0, -1, -2, -3, -2, -1, 0, 0, 0, 0, 5, 5, 2, 2, 1, 0, 2, 2, 2, 1, -1, -1, -1, 0, 3, 3, 1, 0, -1, 0, 1, 0, 0, -2, -2, -3, -2, 0, 0, 0, 0, 0, 5, 5, 4, 2, 2, 1, 3, 5, 4, 1, 0, -1, -2, 0, 2, 3, 2, 0, 0, 2, 2, 1, 0, 0, 0, -1, -1, 0, -1, -2, -1, 0, 4, 6, 4, 3, 1, 1, 4, 5, 5, 1, 0, 0, -1, 0, 1, 3, 2, 1, 1, 4, 3, 2, 2, 1, 0, 1, 1, 1, -1, -1, -1, -1, 4, 6, 3, 3, 0, 1, 3, 4, 4, 0, 0, 0, 0, -1, 0, 2, 1, 1, 3, 4, 5, 3, 1, 0, 0, 3, 2, 0, 0, -2, -1, 0, 4, 4, 2, 1, 1, 0, 2, 3, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 3, 3, 4, 5, 1, 0, 1, 2, 1, 1, 0, -1, -3, -1, 3, 5, 1, 0, 0, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 2, 3, 2, 1, 0, 0, 0, 2, 1, -1, -2, -2, 0, 2, 3, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 4, 3, 4, 2, 0, 0, 0, 1, 2, 0, -4, -1, 0, 2, 2, 0, -1, -1, 0, 1, 0, 0, 1, 2, 0, -2, -3, -1, 0, 0, 0, 2, 4, 4, 4, 3, 1, -1, 0, 0, 0, -1, -3, -2, 0, 1, 1, 0, -1, -3, -1, 0, -1, 0, 1, 2, 1, -3, -4, -2, 0, 0, 0, 2, 5, 6, 4, 2, 0, -1, -1, -1, 0, -2, -3, -2, -1, 2, 1, -1, -2, -2, 0, 0, 0, -1, 0, 1, 2, -2, -4, -4, -1, -3, 0, 2, 3, 5, 6, 2, 0, -1, -1, 0, 0, -1, -3, -2, 0, 1, 0, -2, -2, -3, 0, 0, -2, -4, -2, 0, 0, -1, -3, -3, -3, -2, -2, 0, 1, 3, 6, 4, 1, 0, 0, -1, -2, -3, -4, -4, -2, 2, 0, 0, -3, -2, 0, 0, 0, -4, -2, -1, -1, -3, -4, -1, -2, -3, -2, -1, 1, 3, 6, 6, 3, 2, 0, 0, -2, -5, -6, -3, -1, 1, 0, -1, -3, -1, 0, 0, -1, -3, -4, -3, -2, -4, -3, -2, 0, -2, -3, -4, -1, 1, 4, 6, 4, 2, 0, 0, -1, -4, -6, -5, -1, 0, 0, -2, -1, -1, 0, 0, -1, -2, -4, -3, -3, -3, -3, -2, 0, 1, -2, -2, -3, 0, 2, 3, 2, 3, 1, 0, 0, -3, -4, -3, 0, 1, 1, -1, -2, -1, 0, 1, -2, -4, -4, -1, -3, -4, -6, -4, 0, 2, 0, -3, -1, -1, 1, 2, 2, 1, 0, 0, 0, -1, -4, -3, 0, 2, 1, 0, -1, 0, 0, 0, -1, -3, -2, -2, -2, -3, -5, -5, -1, 2, 1, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, -1, -3, -3, -1, 2, 2, 0, -1, -1, 0, 1, -2, -3, -2, -1, 0, -1, -5, -6, -4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4, -3, -1, 3, 4, 2, -2, 0, 2, 1, 0, 0, -1, 0, 1, -1, -3, -5, -5, 0, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, -2, -4, -3, -2, 3, 4, 2, 0, 0, 0, 3, 0, 0, 0, 1, 1, 1, -1, -4, -5, 0, 1, 2, 3, 2, 1, 1, 0, 1, 2, 1, 0, 0, -3, -3, -1, 3, 4, 2, 0, 0, 1, 2, 2, 0, 1, 1, 3, 3, 0, -2, -4, -1, 1, 3, 3, 3, 1, 1, 1, 1, 2, 3, 3, -1, -2, -1, 0, 2, 3, 3, 1, 0, 0, 1, 2, 0, 1, 4, 2, 3, 2, 0, -2, 0, 3, 5, 4, 2, 0, 1, 0, 1, 3, 3, 4, 0, -1, -1, 0, 3, 3, 2, 1, 0, 1, 2, 2, 2, 1, 3, 3, 3, 1, 0, -1, 0, 3, 4, 4, 2, 1, 0, 0, 1, 3, 4, 2, 0, 0, 0, 0, 2, 4, 3, 1, 0, 1, 3, 2, 2, 1, 1, 2, 3, 2, 2, 2, 1, 3, 3, 3, 3, 1, 0, 0, 0, 3, 3, 3, 1, -1, -1, 1, 4, 3, 4, 2, 1, 3, 3, 3, 4, 1, 2, 2, 2, 3, 2, 3, 4, 5, 3, 3, 3, 1, 1, 0, 0, 2, 3, 3, 0, 0, 0, 0, 5, 5, 3, 2, 2, 3, 5, 4, 3, 1, 1, 2, 2, 3, 4, 6, 7, 5, 4, 4, 4, 4, 2, 0, 0, 1, 3, 3, 1, 0, 0, 1, 4, 5, 5, 2, 3, 4, 5, 4, 1, 2, 2, 2, 1, 0, 1, 6, 6, 6, 4, 3, 4, 5, 3, 1, 0, 1, 2, 2, 2, 2, 1, 0, 6, 6, 5, 3, 3, 4, 6, 5, 3, 1, 2, 2, 0, 0, 1, 5, 5, 4, 2, 2, 4, 5, 4, 2, 2, 0, 1, 3, 3, 5, 1, 0, 6, 7, 5, 5, 4, 5, 6, 4, 2, 3, 1, 1, 0, -2, 0, 2, 4, 4, 2, 3, 4, 4, 4, 3, 0, 0, 1, 3, 5, 4, 3, 1, 7, 8, 7, 6, 5, 5, 5, 5, 5, 5, 4, 1, 0, -2, -1, 2, 4, 1, 0, 1, 3, 5, 4, 2, 0, -1, 0, 0, 2, 4, 3, 2, 3, 4, 5, 3, 4, 2, 4, 3, 1, 1, 2, 1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -2, -1, 0, 0, 0, 0, 1, 1, 2, 1, 2, 2, 2, 1, 1, 2, 2, 2, 2, 1, 1, 0, 0, 1, 0, 1, 1, 0, 0, -1, -2, -1, -2, -1, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 3, 2, 1, 3, 2, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -2, -3, -1, -1, -1, -1, 0, -1, 0, 1, 1, 2, 2, 3, 3, 3, 1, 1, 2, 2, 1, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, -1, -1, -2, -2, -1, -1, -2, 0, 0, 0, 0, 1, 2, 3, 4, 2, 2, 3, 1, 2, 1, 2, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -2, -2, -2, 0, 1, 0, 2, 1, 1, 3, 3, 3, 1, 2, 2, 2, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -2, -1, 0, 0, 1, 1, 1, 2, 2, 3, 1, 2, 1, 0, 0, 1, 1, 2, 2, 1, 1, 0, -1, 0, 0, -1, 0, -1, 0, 1, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 2, 1, 1, 0, 0, 0, 0, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 1, 0, 0, 0, 0, 0, 2, 2, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 1, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -2, -1, -2, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -2, -3, -2, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, -2, -1, 0, 0, 0, 1, 1, 2, 1, 0, 1, 0, 0, 0, -1, -1, -2, -2, -4, -4, -3, -2, -1, -2, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 2, 2, 1, 1, 0, 1, 0, -1, -1, -2, -3, -2, -3, -3, -2, -2, -4, -3, -1, -1, -1, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, -2, -4, -4, -3, -4, -3, -2, -2, -3, -3, -2, -2, -1, 0, -1, 0, -1, -1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 2, 1, 2, 0, -1, -2, -4, -3, -3, -2, -2, -2, -1, -2, -2, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 1, 0, 1, 1, 0, 0, 0, -3, -3, -2, -2, -3, -4, -2, -1, -1, -2, -3, -3, -3, -2, -2, -2, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, 1, 1, 2, 1, 0, -2, -2, -3, -2, -2, -3, -3, -1, 0, -2, -1, -2, 0, -1, -1, -1, 0, 0, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, 2, 2, 1, -1, 0, -1, -1, -3, -2, -3, -2, -2, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, -1, -2, -2, -1, -1, -1, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, -1, -2, -3, -4, -5, -2, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -2, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -3, -4, -4, -4, -3, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, -2, -2, -4, -3, -1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, -1, 0, -1, -2, -1, 0, -1, 0, -2, -2, 0, 1, 1, 2, 2, 2, 1, 0, 0, -2, -3, -1, 0, 2, 3, 2, 2, 2, 2, 2, 1, 0, 0, 0, -1, -2, -2, 0, -1, 0, -2, -1, -1, 1, 1, 3, 2, 3, 3, 3, 1, 0, -1, 0, 1, 3, 3, 3, 2, 1, 2, 2, 1, 1, 1, 0, -1, -2, -2, 0, 0, 0, 0, 0, 1, 0, 1, 3, 3, 2, 2, 2, 1, 1, 0, 0, 2, 2, 3, 3, 3, 1, 2, 2, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 2, 3, 3, 2, 1, 1, 1, 1, 0, 0, 1, 3, 5, 4, 2, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 1, 1, 0, 1, 1, 0, 1, 1, 2, 4, 5, 3, 3, 1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 2, 1, 1, 0, 2, 1, 1, 0, 2, 2, 4, 5, 4, 3, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 1, 0, 2, 2, 1, 2, 3, 2, 3, 3, 2, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 2, 1, 1, 2, 2, 1, 1, 1, 1, 2, 2, 2, 2, 3, 2, 3, 1, 0, -1, 0, -1, -2, -1, 0, -1, 0, -1, -1, -1, 0, 0, 1, 0, 1, 2, 1, 1, 2, 0, 0, 1, 2, 1, 2, 2, 1, 1, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, -2, -2, 0, 0, 0, 0, 1, 2, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -2, -1, -1, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, -3, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, -2, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, -1, 0, -1, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, -1, -2, 0, -2, -1, -1, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 2, 0, 2, 1, 0, 1, 0, 0, -1, -1, -1, -1, 0, -1, -2, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, -1, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, -1, -1, -1, -1, -2, -1, -1, -1, 0, 0, 1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, -1, -1, -1, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 1, 0, 1, 0, 0, 0, -1, -2, -2, -2, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, -2, -1, -2, -2, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, 1, 1, 2, 1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 1, 0, 1, 1, 1, 2, 2, 1, 0, -1, 0, 0, -1, -1, 0, 0, -2, 0, 0, 1, 1, 2, 3, 2, 1, 0, 1, 0, -1, -1, 0, 1, 2, 1, 2, 2, 2, 2, 2, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, -1, 1, 1, 1, 1, 1, 2, 2, 2, 0, 0, 0, 1, 2, 3, 3, 1, 0, 1, 2, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 3, 1, 1, 2, 0, 1, 1, 0, 1, 2, 3, 3, 1, 1, 2, 2, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 1, 2, 2, 2, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 2, 1, 1, 1, 1, 0, 0, 1, 2, 2, 3, 3, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 3, 3, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 2, 2, 2, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 2, 1, 3, 1, 0, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 2, 0, 0, -1, -2, -2, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, -2, -3, -3, -2, -2, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, -1, -2, -3, -2, -1, -2, -2, -1, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, -3, -1, -2, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, 1, 0, 0, -1, -2, -2, -1, -1, -1, -1, -1, -1, -1, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, -1, 0, 0, -1, -2, 0, -1, 0, 0, 1, 1, -1, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, -2, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, -2, -1, -1, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, 1, 0, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, -1, -2, 0, -1, 0, -1, -2, -1, 0, 1, 0, 1, -2, -2, 0, 0, 0, -1, 0, -1, -1, 0, -2, 0, 0, -1, -2, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 2, 0, -2, -1, 0, -1, -1, 0, 0, 0, -1, -2, -1, -2, -1, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, -1, 0, -1, -1, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, -1, 0, 1, 1, -1, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, -2, -1, -2, 0, -1, 0, -1, 0, 0, 1, 1, -2, -1, -2, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, -1, -1, -1, 0, -2, 0, 0, 0, -1, 0, 1, 0, -1, -1, -2, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, -1, -1, 0, -1, -1, -1, 0, -1, -1, 0, 2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -2, -2, -2, -2, -1, -2, 0, -1, -1, -2, -1, -1, 0, 0, 2, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, -2, -2, -2, -1, -2, -1, 0, -1, -1, -1, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, -2, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 2, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 2, 1, 0, -1, -2, -1, -3, -2, -1, -1, 0, -1, 0, 0, 0, 2, 0, 0, -2, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 2, 2, 0, 0, -1, -2, -1, -2, -2, -2, -1, 0, 0, -1, 0, 1, 1, 1, -2, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 2, 1, 0, 0, -1, -2, -3, -1, -2, -1, -2, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, -1, -1, -1, 0, -1, 0, 0, 1, 0, 0, -1, -2, -1, -1, -2, 0, -1, -2, -1, -2, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -2, 0, 0, -1, 0, -1, 0, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, -1, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, -2, -2, 0, 0, -1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, -2, -1, -2, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, -2, -2, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, -1, -1, -2, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 1, 2, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, -1, -1, -1, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 2, 1, 1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 2, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 2, 1, 1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, -1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -2, -1, 0, 0, -1, -1, -2, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 1, 0, -1, -2, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, -1, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, -2, -1, 0, 0, -1, 0, 0, 0, -2, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, -1, -1, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 2, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, -1, -2, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 2, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, 0, -2, 0, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, -2, -1, -2, -2, -1, -2, -2, 0, -1, -1, -2, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, -2, -2, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, 0, -2, -1, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -2, -1, -2, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 2, 1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -2, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 1, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 2, 0, 1, 0, 0, 0, 1, 3, 2, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 2, 0, 0, 0, 1, 1, 0, 2, 1, 0, 1, 2, 2, 0, 0, -1, 0, 0, -1, -1, 0, 0, 1, 1, 2, 2, 1, 1, 0, 0, 0, 0, 1, 1, 0, 1, 2, 0, 0, 1, 0, 0, 0, 3, 2, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 1, 2, 2, 1, 2, 2, 0, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 1, 2, 2, 0, 0, -2, -1, 0, 0, -1, 0, 0, 2, 3, 2, 2, 1, 3, 3, 1, 0, 1, 0, 1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 2, 1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 2, 3, 3, 2, 2, 3, 1, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 2, 1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 2, 3, 2, 4, 3, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 3, 2, 0, 0, -1, -2, 0, 0, 0, 1, 0, 1, 2, 2, 3, 2, 3, 3, 2, 1, 0, 0, 0, 0, 0, 2, 1, 0, -1, 0, 1, 2, 2, 1, 0, 0, -2, -2, 0, 0, 1, 1, 0, 0, 0, 2, 2, 2, 3, 2, 3, 2, 1, -1, 1, 0, 0, 1, 1, 0, 0, 0, 1, 2, 4, 3, 0, 0, -2, 0, 0, 0, 1, 0, -1, -1, 0, 0, 2, 2, 3, 2, 2, 2, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 3, 2, 0, 0, -2, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 3, 3, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 1, 2, 2, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 1, 0, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, -1, -2, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -2, 0, -1, 0, -2, -1, 0, -1, -1, -3, -2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, -1, -2, -2, 0, -1, -1, -2, 0, -1, -1, -2, -2, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, 0, -1, -2, -2, -2, -2, -1, -2, 0, -2, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, -2, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -2, -1, 0, 0, -1, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 1, 1, 1, 2, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 2, 2, 2, 1, 1, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 0, 0, 2, 1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, 1, 1, 0, 0, -1, -1, 0, 0, 2, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 2, 1, 0, 1, 1, 1, 1, 0, 0, -1, -1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, 0, -1, -2, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, -2, -1, 0, 0, 0, -1, 0, -2, 0, 0, -1, -1, -1, 0, 0, -1, -1, -2, -2, -1, 0, 0, 1, 2, 2, 1, 1, 1, 0, 0, -1, 0, -1, 0, 1, 0, 0, -1, 0, -2, -1, 0, -1, -1, 0, -1, -1, -1, -2, -1, -1, 0, 0, 0, 0, 2, 2, 0, 1, 1, 0, 0, -1, -1, -2, -1, 0, 0, -1, 0, -2, -3, -2, -1, -2, -1, -2, -2, -1, -2, -2, -1, -1, -1, 0, 0, 1, 1, 2, 1, 2, 1, 0, 0, 0, -1, -2, -1, 0, 1, 0, -1, -1, -1, -1, -1, -1, -3, -2, -2, -2, -1, -1, -2, -2, -1, 0, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, -1, -1, 0, 0, -2, -1, -2, -1, -1, -2, -2, -1, 0, 0, 0, 0, 1, 3, 1, 1, 2, 2, 1, 1, 0, -1, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, -1, -2, -1, -1, -1, -2, -3, -1, 0, 0, 0, 0, 1, 3, 2, 3, 1, 1, 2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -2, -1, -3, -1, 0, 0, 0, 0, 0, 1, 2, 2, 2, 1, 2, 0, 0, 0, -1, -1, 1, 0, 0, 1, 0, 0, -1, -1, -1, -1, -2, -1, -1, -1, -1, -2, -1, -1, 0, 0, 1, 2, 2, 2, 2, 2, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, -1, 0, 1, 1, 1, 1, 0, 1, 2, 1, 0, 0, 0, -2, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 2, 2, 1, 2, 1, -1, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 2, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 1, 1, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 2, 1, 2, 0, 1, 1, 0, 0, 0, -1, 1, 0, 0, -1, -1, 0, 0, 1, 2, 2, 1, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 1, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 3, 1, 1, 0, 1, 2, 3, 1, 1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 3, 3, 2, 2, 2, 2, 2, 3, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 3, 4, 2, 2, 2, 2, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 2, 3, 2, 1, 2, 1, 2, 1, 1, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, -1, -1, 0, -1, -2, -1, -1, -2, -1, 0, 1, 2, 1, 1, 1, 2, 2, 2, 1, 0, 0, 0, -1, 0, -1, 0, 1, 0, -1, -2, -1, 0, 0, 0, 0, 0, -1, -2, -1, -1, -2, 0, 1, 1, 2, 1, 1, 2, 2, 0, 1, 0, 0, 0, -1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 1, 2, 1, 1, 1, 0, 2, 1, 1, 2, 2, 1, 3, 3, 3, 2, 1, 0, 0, 0, 0, -2, 0, 0, 0, 1, 1, 1, 1, 0, 1, 2, 3, 3, 1, 2, 0, 0, 1, 2, 3, 2, 1, 3, 4, 4, 3, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, -1, 0, 1, 3, 2, 1, 0, 2, 2, 3, 3, 2, 1, 2, 3, 2, 4, 3, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 2, 3, 1, 2, 2, 1, 2, 3, 2, 3, 1, 1, 0, 0, -1, 0, -1, 0, 0, 1, 2, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 1, 2, 2, 3, 4, 3, 3, 2, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, -1, -1, -1, 1, 0, 0, 1, 2, 1, 2, 1, 0, 0, 0, 0, 0, 2, 2, 3, 3, 2, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, -2, 0, 0, 0, 0, 1, 3, 4, 2, 2, 0, 0, 0, -1, 0, 1, 2, 3, 3, 1, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 2, 2, 0, 1, -1, -1, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, -1, -2, -2, -2, 0, 0, 0, 0, -1, -2, 0, 0, 0, -1, 0, 0, 2, 1, 0, -1, -2, 0, -1, 0, -1, 0, 1, 1, 2, 0, 0, 0, -2, -3, -5, -3, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -3, -1, -2, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, -3, -4, -2, 0, 0, 0, 0, 0, -2, -1, 0, 0, -1, -1, -1, -2, -3, -3, -3, -3, -2, -2, -1, 0, -1, -1, 0, 1, 0, 0, -1, -1, -3, -3, -2, 0, 0, -1, -2, -2, -3, -2, 0, -2, -1, -2, -3, -2, -3, -3, -3, -4, -3, -2, -1, -2, 0, -1, 0, 0, 0, 0, 0, -2, -2, -3, -2, 0, 0, -1, -2, -2, -3, -1, -1, -2, -2, -2, -3, -3, -2, -3, -3, -2, -1, -1, -1, -1, 0, -1, 1, 1, 0, 0, 0, -1, -1, -3, -2, 0, 0, 0, 0, -1, -3, -1, 0, -1, -3, -3, -3, -4, -3, -4, -3, -2, -2, 0, 0, 0, 0, 0, 1, 1, 3, 1, 0, -2, -3, -4, -2, 0, -1, 0, -1, 0, -1, 0, 0, 0, -2, -3, -3, -4, -2, -3, -2, -1, -1, 0, 0, 0, 1, 2, 2, 1, 2, 1, -1, -2, -4, -4, -3, 0, -1, -1, 0, -1, 0, 0, 0, 0, -2, -2, -4, -4, -3, -2, -3, -1, 0, 0, 0, 1, 2, 2, 3, 2, 2, 0, 0, -1, -2, -4, -3, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -3, -2, -1, -1, -1, -3, -1, -2, 0, 0, 0, 2, 2, 2, 1, 3, 0, 0, -1, -4, -4, -2, -1, 0, 0, 0, 0, -1, -2, -2, -1, -1, -1, -1, 0, 0, 0, -1, -2, -1, 0, 0, 1, 3, 2, 1, 1, 1, 0, 0, -2, -2, -3, -3, 0, 0, 0, 0, 0, -2, -3, -2, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, -2, 0, 1, 2, 3, 3, 1, 1, 1, 0, -1, -1, -3, -3, 0, 0, 0, 0, -2, -3, -2, -1, 0, 1, 0, 0, 1, 2, 3, 0, 0, -1, 0, 1, 1, 3, 3, 3, 2, 0, 0, 1, 0, -2, -2, -1, 0, -1, 0, 0, 0, -2, -2, -1, 0, 2, 2, 2, 2, 3, 3, 2, 0, 0, 0, 1, 2, 3, 3, 2, 2, 0, 0, 0, 0, -2, -3, -2, -1, 0, 0, 0, -1, -2, 0, 0, 2, 2, 2, 2, 3, 2, 2, 1, 0, 2, 0, 2, 3, 3, 1, 2, 0, -1, 0, 0, 0, -1, -2, -3, 0, 0, 0, 0, 0, -1, -1, 1, 1, 1, 1, 2, 2, 1, 1, 2, 2, 2, 3, 2, 2, 1, 1, 1, 0, -1, 0, -1, -1, -3, -3, -1, 0, 0, 0, 1, 0, 0, -1, 1, 2, 1, 1, 1, 2, 0, 1, 1, 2, 1, 2, 1, 1, 1, 1, 2, 0, 0, -1, -2, -2, -1, -3, -2, 0, 1, 0, 1, 0, 0, 0, 2, 2, 3, 2, 1, 2, 1, 0, 0, 0, 2, 1, 1, 0, 1, 2, 1, 1, 1, -1, -1, -1, -3, -3, -2, 0, 1, 1, 1, 1, 1, 2, 2, 4, 2, 2, 2, 2, 1, 1, 0, 1, 1, 2, 1, 0, 0, 0, 1, 0, 0, -2, -3, -3, -1, -2, -1, 0, 1, 1, 0, 0, 1, 2, 3, 4, 2, 2, 2, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, -3, -2, -4, -2, -3, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, -1, -2, -1, -2, -2, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 2, 2, 0, -1, -1, 0, 1, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 1, 3, 3, 0, -1, 0, 0, 2, 0, 0, -1, -1, -1, -1, 0, 1, 1, 0, 0, 0, -1, 0, 1, 1, -1, 0, -1, 0, 1, 0, 0, 1, 1, 3, 1, 0, 0, 0, 2, 3, 2, 2, 1, 0, 0, 0, 0, 2, 3, 3, 1, 0, 1, 1, 2, 1, 0, 1, 0, 0, 1, 2, 0, 2, 0, 2, 3, 0, 2, 0, 1, 3, 4, 3, 0, 0, 0, 0, 0, 2, 4, 3, 2, 1, 2, 3, 3, 2, 0, 0, 1, 0, 1, 0, 0, 1, 1, 3, 3, 1, 2, 1, 1, 3, 4, 3, 1, 0, 0, -1, 0, 0, 1, 1, 2, 1, 3, 4, 4, 2, 1, 0, 0, 1, 0, 1, -1, 0, 0, 3, 2, 1, 0, 0, 1, 2, 3, 2, 0, -1, 0, 0, 0, 1, 0, 2, 2, 2, 4, 4, 3, 2, 1, 2, 1, 2, 2, 0, 0, 0, 0, 3, 2, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 3, 3, 3, 3, 1, 1, 3, 2, 1, 0, -1, 0, 0, 1, 2, 1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 3, 4, 3, 1, 1, 2, 4, 2, 0, -2, -2, -2, 3, 3, 0, 0, 0, 1, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 3, 3, 1, 2, 1, 3, 2, 0, -1, -2, -2, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 2, 2, 0, 0, 0, 0, 0, 1, 1, 2, 3, 2, 1, 1, 0, 1, 1, 0, -1, -3, -1, -2, 2, 0, -1, -2, -1, -1, -1, -1, 0, 1, 2, 2, 0, 0, 0, 0, 0, 1, 0, 1, 2, 3, 3, 2, 1, 0, 1, 0, -2, -3, -2, 0, 1, 1, 0, -2, -1, -1, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 2, 2, 3, 2, 2, 1, 0, -1, 0, -2, -4, -4, 0, 1, 1, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 2, 2, 3, 4, 2, 2, 0, -1, -1, -2, -4, -3, 0, 1, 0, -1, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 2, 3, 2, 3, 2, 1, 0, 0, -3, -5, -4, -1, 0, 0, -1, -1, -1, -1, 0, 0, -3, -2, -1, -1, 0, -1, -1, 0, -1, -1, -2, 0, 1, 1, 2, 1, 1, 2, 0, -2, -3, -5, -3, -3, 1, 0, -1, -1, -2, 0, 0, 0, -2, -2, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 2, 1, 0, 0, -3, -3, -4, -1, 1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -2, -1, -1, -1, 0, 1, 0, -1, 0, 1, 2, 1, 1, 0, 0, 0, 0, -2, -4, -4, -2, 1, 1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, -2, -4, -3, -2, 2, 2, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -2, -3, -3, -2, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -2, -4, -3, -1, 1, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, -4, -4, -2, 1, 1, 1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -2, -2, -1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 0, -3, -3, -3, -2, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 0, 0, -2, 0, 1, 0, 1, 1, 0, 1, 1, 2, 2, 2, 0, -1, -2, -2, -1, 2, 1, 1, 0, 0, 0, 1, 1, 1, 1, 2, 2, 3, 3, 2, 1, 1, 1, 2, 0, 0, 1, 0, 0, 1, 1, 3, 1, 0, -1, -2, 0, 1, 3, 1, 0, 0, 0, 2, 2, 1, 1, 1, 2, 4, 3, 2, 1, 1, 1, 2, 1, 1, 0, 0, 0, 2, 1, 3, 2, 0, -2, 0, 0, 2, 2, 1, 1, 1, 1, 2, 2, 2, 1, 2, 2, 3, 2, 2, 2, 4, 3, 4, 2, 1, 0, 1, 1, 0, 1, 1, 2, 0, -1, 0, 0, 2, 2, 2, 1, 1, 3, 2, 3, 3, 1, 1, 1, 2, 1, 2, 4, 4, 4, 3, 1, 2, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 2, 3, 2, 2, 2, 2, 3, 3, 3, 0, 2, 2, 2, 2, 3, 4, 4, 5, 4, 3, 2, 1, 2, 0, 0, 2, 2, 0, 0, 0, 1, 1, 4, 5, 3, 2, 2, 2, 3, 3, 2, 2, 1, 2, 2, 1, 2, 3, 5, 4, 4, 4, 3, 5, 3, 3, 1, 2, 1, 1, 1, 1, 0, 1, 3, 5, 3, 3, 2, 2, 4, 3, 2, 3, 2, 2, 1, 1, 3, 4, 5, 5, 4, 4, 4, 4, 4, 3, 1, 1, 1, 2, 1, 2, 1, 1, 5, 5, 5, 4, 3, 2, 4, 4, 2, 2, 2, 1, 2, 1, 1, 2, 5, 3, 2, 3, 4, 5, 4, 2, 1, 1, 1, 1, 2, 2, 2, 1, 4, 5, 4, 4, 2, 3, 2, 3, 3, 2, 3, 1, 1, 0, 0, 1, 3, 2, 0, 1, 1, 2, 1, 0, 1, 0, 1, 2, 1, 2, 3, 2, 0, 2, 2, 2, 1, 1, 1, 2, 1, 0, 1, 1, 0, 0, 0, 1, 2, 1, 0, 0, 2, 1, 0, 1, 0, 1, 0, 0, 1, 0, 1, 2,
    -- filter=0 channel=3
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, -2, -2, -1, -1, -1, -2, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, -2, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 2, 0, 1, 1, -1, 0, 0, 0, 0, 0, -1, -1, -1, -2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, -1, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 2, 1, 2, 1, 3, 3, 2, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 1, 1, 0, 1, 2, 1, 2, 0, 0, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 2, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, -1, -1, -1, -1, -1, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, -2, 0, 0, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -2, -3, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, -1, -2, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 0, 1, 1, 0, 1, 1, 1, 0, 1, 1, 1, 0, 2, 1, 0, 1, 0, 1, 0, 2, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 2, 1, 2, 2, 2, 1, 1, 2, 0, 1, 2, 1, 0, 0, 1, 1, 2, 1, 1, 1, 1, 1, 0, 1, 1, 1, 0, 1, 1, 1, 2, 1, 1, 1, 1, 0, 1, 1, 1, 0, 1, 2, 2, 0, 1, 1, 1, 1, 1, 1, 1, 2, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 2, 1, 1, 2, 1, 0, 1, 0, 1, 1, 1, 0, 1, 2, 0, 2, 1, 1, 1, 2, 2, 0, 0, 0, 1, 2, 1, 1, 1, 1, 1, 1, 2, 1, 2, 2, 2, 0, 1, 0, 1, 1, 1, 1, 1, 1, 0, 2, 1, 0, 0, 0, 0, 1, 1, 0, 1, 2, 0, 1, 2, 2, 0, 2, 2, 2, 1, 1, 1, 1, 0, 1, 0, 1, 1, 0, 0, 1, 1, 1, 1, 2, 2, 0, 0, 1, 0, 1, 1, 1, 2, 2, 1, 1, 1, 1, 0, 1, 1, 0, 1, 1, 1, 0, 1, 2, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 2, 0, 2, 2, 1, 1, 1, 2, 1, 0, 0, 0, 1, 1, 1, 1, 1, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 2, 1, 2, 1, 2, 1, 1, 2, 1, 1, 2, 1, 1, 1, 2, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 3, 3, 1, 2, 2, 1, 1, 2, 1, 1, 1, 0, 2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, 2, 1, 2, 3, 1, 0, 0, 1, 0, 1, 1, 2, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 1, 0, 0, 2, 1, 2, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 1, 1, 1, 1, 2, 1, 2, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 1, 1, 0, 1, 1, 1, 2, 1, 1, 1, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, 0, 0, 0, 0, 0, 2, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 2, 2, 0, 1, 1, 0, 2, 0, 1, 1, 2, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 2, 1, 2, 2, 1, 1, 0, 1, 2, 1, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 1, 1, 1, 1, 1, 2, 1, 0, 2, 1, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 2, 2, 2, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 2, 0, 1, 1, 2, 2, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 2, 2, 2, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 2, 1, 1, 1, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 2, 1, 2, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 2, 2, 2, 2, 1, 1, 1, 2, 0, 2, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 1, 2, 2, 1, 0, 1, 0, 1, 1, 1, 1, 2, 2, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 2, 1, 0, 1, 0, 1, 0, 0, 1, 1, 1, 2, 1, 1, 0, 1, 2, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 1, 1, 2, 2, 1, 0, 1, 2, 0, 1, 2, 1, 1, 1, 2, 2, 2, 2, 1, 0, 0, 1, 0, 1, 0, 1, 1, 2, 1, 0, 1, 2, 2, 1, 2, 2, 2, 2, 2, 2, 1, 2, 2, 0, 1, 1, 2, 2, 1, 3, 3, 0, 0, 2, 0, 0, 1, 0, 1, 1, 0, 1, 0, 1, 0, 1, 2, 1, 1, 2, 2, 1, 1, 1, 2, 2, 3, 2, 1, 3, 3, 3, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 2, 2, 2, 1, 2, 2, 2, 3, 2, 3, 3, 3, 3, 2, 3, 2, 1, 0, 1, 1, 0, 0, 1, 1, 1, 0, 2, 1, 0, 0, 0, 1, 1, 0, 1, 2, 1, 2, 2, 2, 2, 1, 2, 1, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -2, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, -1, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -2, -1, 0, -1, 0, 0, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 1, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 3, 2, 2, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 3, 2, 1, 2, 1, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 1, 2, 1, 2, 2, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 1, 2, 0, 1, 0, 0, 0, 0, -1, 1, 1, 0, 1, 1, 1, 2, 2, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 2, 1, 1, 0, 1, 0, -1, 0, -2, -2, -2, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 2, 2, 0, 0, 0, 0, -1, 0, 1, 1, 1, 3, 1, 0, 0, -1, -2, -1, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 0, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, -1, -1, 1, 1, 1, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -2, -1, -2, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 2, 2, 2, 0, 0, -2, -2, 0, 0, -1, -1, -1, 0, -2, -1, -2, -2, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, -1, -1, -2, -1, -2, -1, -2, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 2, 2, 0, 0, -2, -1, 0, -1, -3, -2, -1, -3, -1, -2, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, -1, 0, -1, -2, -2, -3, -1, -2, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 2, 2, 0, -1, -1, 0, 0, 0, -3, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, -2, -1, -2, -3, -3, 0, -1, 0, 0, 0, 0, 2, 0, 1, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 2, 0, 1, 1, 2, 0, 0, 0, -2, -2, -1, -3, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 1, 2, 1, 2, 2, 0, 0, 0, -1, -1, -1, -3, -2, -2, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 2, 2, 2, 2, 1, 1, 2, 2, 1, 0, 0, 0, 0, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 1, 2, 3, 1, 0, 1, 0, 2, 0, 0, 0, -1, -2, -1, -2, -2, -1, -1, 0, 0, 0, -1, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 2, 0, -1, -1, 0, -1, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 1, 0, 0, -1, 0, -1, -2, -1, -2, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -2, -2, -2, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 1, 0, -1, -1, -2, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 2, 0, 1, 1, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 2, 1, 0, 0, 0, 2, 1, 1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 1, 0, 2, 1, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 2, 1, 0, 1, 1, 0, 1, 1, 1, 2, 1, 1, 0, 1, 1, 0, 0, -1, 0, -1, 0, 0, -1, -1, -2, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 2, 2, 1, 0, 0, 1, 2, 1, 1, 0, 2, 0, 1, 1, 0, 1, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 2, 3, 3, 4, 3, 3, 2, 1, 3, 2, 2, 2, 2, 2, 3, 1, 3, 1, 2, 2, 1, 3, 1, 1, 0, -2, -2, 0, 0, 0, 0, 1, 3, 4, 4, 4, 4, 4, 4, 3, 3, 3, 1, 2, 2, 1, 2, 3, 4, 3, 2, 2, 2, 2, 1, 1, 0, -2, -1, 0, 0, 1, 1, 2, 2, 2, 4, 4, 3, 4, 4, 4, 1, 1, 0, 0, 0, 2, 1, 3, 2, 3, 3, 3, 2, 1, 0, 0, -1, -3, -2, -1, 0, 0, 0, 0, 0, 2, 1, 3, 2, 2, 3, 3, 0, 0, -1, 0, 0, 1, 1, 1, 3, 3, 1, 1, 2, 2, 2, 0, -2, -1, -2, -3, -2, -1, 0, 0, 0, 1, 2, 2, 1, 1, 1, 0, -1, 0, -1, 0, 0, 0, 0, 2, 1, 2, 2, 1, 2, 2, 1, 1, 0, -3, -2, -2, -1, 0, 0, 1, 0, 0, 1, 0, 0, -1, -2, -2, -2, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 2, 2, 0, -1, -2, -3, -2, -2, 0, 0, 0, 1, 2, 0, 0, -1, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 2, 1, 2, 0, -2, -2, -3, -2, 0, 0, 0, 1, 0, 0, 0, -2, -4, -3, -2, -2, -1, -1, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 1, 2, 1, 0, -2, -2, -3, -2, -1, -1, -1, -1, 0, -1, -2, -2, -3, -4, -3, -1, -1, -2, -1, -1, 0, -1, 0, -1, -2, -1, -1, 0, 1, 3, 2, -1, -3, -2, -2, -1, -3, -3, -3, -3, -1, -2, -2, -3, -3, -3, -4, -1, -3, -1, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 2, 2, 2, -2, -3, -2, -3, -4, -3, -4, -5, -2, -3, -2, -2, -3, -2, -2, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 2, -1, -2, -3, -3, -2, -4, -4, -5, -3, -2, -2, -3, -3, -2, -2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, -2, -1, -1, -2, -3, -3, -4, -4, -3, -3, -3, -2, 0, -1, 0, 0, 0, 0, 0, 1, 2, 3, 1, 0, 0, 0, -1, 0, -1, 1, 2, 0, -2, -1, -1, -1, -2, -3, -4, -2, -3, -3, -3, 0, 0, 0, 0, 1, 2, 1, 0, 1, 3, 2, 1, 2, 0, -1, 0, 0, 0, 1, 1, 0, -3, -2, 0, -2, -2, -3, -4, -4, -3, -3, -3, -1, -1, 1, 0, 0, 1, 1, 1, 0, 2, 1, 2, 0, -1, -1, -1, 0, 0, 0, 2, -2, -2, 0, -1, -1, -4, -4, -4, -3, -2, -2, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 1, 0, -1, 0, 0, 1, 1, 1, 1, -1, -2, 0, 0, -3, -3, -4, -3, -4, -2, -2, -2, -2, 0, 0, 0, 0, -1, 0, 1, 2, 2, 1, 0, 0, 1, 0, 2, 3, 3, 2, 1, -1, -1, 0, -1, -2, -3, -3, -3, -4, -2, -3, -2, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 3, 2, 2, 2, 1, 2, -1, -2, -2, -1, -3, -2, -3, -3, -3, -4, -3, -3, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 3, 3, 2, 2, 0, 1, 0, 0, 0, -1, -2, -3, -4, -3, -2, -3, -3, -2, -1, 0, 0, 0, 0, -1, -2, -1, -1, 0, -2, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, -3, -4, -3, -5, -4, -4, -2, -3, -2, 0, 0, -1, 0, -2, -2, -2, -3, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -3, -2, -3, -2, -2, -2, -1, -1, -1, 0, 0, -1, -2, -4, -2, -2, 0, -2, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, -2, -3, -4, -3, 0, -1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, -2, 0, 0, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, -1, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, -1, -1, 0, -1, 1, 1, 1, 2, 2, 2, 1, 2, 1, 2, 0, 1, 1, 0, 1, 1, 2, 2, 1, 1, 0, 1, 2, 1, 1, 1, 1, 0, -2, -2, 0, 0, 2, 3, 3, 3, 4, 2, 3, 2, 3, 2, 2, 3, 2, 1, 1, 1, 2, 2, 2, 2, 3, 2, 2, 2, 1, 2, 1, 0, -1, -1, 0, 0, 3, 3, 4, 4, 5, 3, 2, 1, 1, 3, 3, 3, 3, 3, 3, 1, 1, 2, 2, 1, 2, 3, 2, 2, 0, 1, 1, 0, 0, -1, 0, 0, 0, 2, 2, 3, 3, 3, 3, 2, 2, 3, 2, 2, 2, 2, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 1, 1, 1, 0, 0, 1, 2, 0, 0, 1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 2, 1, 2, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 2, 1, 2, 1, 3, 3, 1, 3, 3, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 2, 1, 0, 0, 1, 1, 2, 2, 2, 1, 2, 2, 2, 3, 3, 2, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 2, 1, 0, 0, 0, 0, 1, 1, 1, 1, 2, 1, 1, 2, 2, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, 1, 2, 0, 0, 1, 3, 2, -1, 0, 0, 0, 1, 0, 2, 2, 1, 0, 1, 1, 1, 1, 1, 2, 1, 1, 0, -1, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 2, 2, -1, -1, 0, -1, 0, 1, 0, 0, 0, 1, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -2, 0, 0, 0, 1, 1, 0, 1, 3, 2, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 1, 0, 0, 0, 1, 0, -1, -2, -1, -1, 0, 0, 0, 1, 0, 2, 2, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 1, 1, 2, 2, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -2, -1, -1, -1, -2, -2, -1, 0, -1, -1, -1, -1, 0, 0, 0, 1, 1, 3, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -3, -2, -2, -3, -1, -1, -1, -1, 0, -1, 0, 0, -2, -1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, -1, -1, 0, -3, -2, -1, -2, -1, -2, -2, -2, -3, -3, -2, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -2, -1, -2, -2, -2, -2, -1, -3, -2, -2, 0, 0, 0, 0, 1, 1, 0, -1, -1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -2, -1, -1, -1, -1, -1, -2, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, -1, -1, -2, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, -1, -1, 0, 0, 1, 0, -1, 0, -2, -1, -3, -1, -1, -2, -2, -2, -2, -2, -2, 0, 0, 1, 2, 0, 0, 1, 1, 0, 1, 2, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, -2, -1, -3, -1, -2, -3, -2, -1, -2, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 0, -1, 0, 1, 1, 0, -1, -1, -1, 0, -1, -2, -2, -2, -1, -2, -2, -3, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -2, -1, -1, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, -1, -1, 0, 1, 0, 0, -1, 0, 0, 0, -1, -2, -1, 0, -2, -3, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -2, -2, -1, -2, -1, -2, -2, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, 0, -1, 0, 0, 0, -1, -1, -1, -2, -1, -1, -1, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, -2, 0, 0, 1, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -2, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, -2, 0, -2, -1, 0, 1, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 2, 1, 1, 2, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 1, 2, 1, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 1, 2, 2, 3, 3, 1, 2, 2, 1, 1, 2, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, -1, -2, 0, 0, 1, 2, 2, 5, 4, 6, 5, 5, 6, 4, 5, 5, 3, 3, 4, 2, 3, 2, 1, 2, 2, 2, 3, 1, 1, 0, 1, 0, 0, -3, -2, 0, 1, 3, 3, 5, 6, 6, 7, 6, 6, 6, 6, 6, 5, 3, 3, 3, 2, 2, 2, 1, 3, 2, 3, 1, 1, 1, 1, 1, -1, -2, -1, -1, 0, 3, 4, 3, 5, 4, 5, 7, 6, 7, 6, 6, 6, 2, 2, 1, 2, 2, 1, 3, 3, 4, 1, 2, 1, 1, 0, 2, -2, -3, -3, -1, 0, 1, 2, 2, 3, 3, 4, 4, 5, 4, 4, 4, 4, 1, 1, 0, 0, 2, 2, 2, 2, 2, 2, 1, 2, 2, 2, 2, 0, -3, -3, -2, -3, 0, 0, 1, 1, 1, 2, 2, 3, 2, 1, 2, 1, 1, 0, 0, 1, 1, 0, 1, 3, 2, 3, 2, 1, 3, 1, 2, -1, -2, -5, -4, -3, -2, 1, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 1, 2, 3, 1, 0, -2, -3, -4, -5, -2, 0, 0, 0, 1, 0, 0, -2, -1, -2, -1, -1, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 2, 0, -3, -5, -3, -3, -4, -1, -1, -2, -1, -1, -2, -4, -3, -3, -4, -2, -2, -1, -1, 0, -1, -1, 0, -2, -1, 0, -1, 0, 0, 1, 3, 0, -2, -4, -3, -4, -4, -4, -4, -4, -2, -4, -3, -5, -6, -6, -4, -5, -3, -4, -2, -1, -1, -1, 0, -2, -1, -3, -3, -2, 0, 2, 3, 0, -3, -3, -2, -2, -4, -4, -5, -4, -3, -5, -4, -4, -5, -5, -5, -5, -5, -4, -4, -2, 0, -1, 0, 0, -2, -3, -4, -2, 0, 2, 3, 0, -2, -1, -2, -1, -5, -6, -6, -6, -5, -4, -4, -4, -5, -6, -6, -5, -4, -4, -2, -1, 0, 0, 1, 0, 0, -2, -2, 0, 0, 1, 3, 0, 0, -2, 0, -2, -3, -5, -6, -5, -5, -6, -5, -6, -6, -5, -5, -4, -4, -3, -3, -2, 0, 0, 2, 0, 0, -1, -1, -1, 0, 2, 3, -1, 0, -1, 0, -1, -2, -5, -6, -5, -5, -4, -5, -5, -4, -5, -5, -4, -4, -3, -2, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 2, 2, -1, -3, -2, -1, -1, -3, -4, -5, -6, -4, -6, -6, -5, -5, -5, -4, -3, -4, -3, -3, -1, 0, 2, 3, 2, 0, -1, 0, 0, 0, 1, 1, 0, -1, -2, 0, -1, -3, -6, -6, -5, -5, -6, -6, -6, -5, -5, -4, -4, -2, -2, -2, -1, 1, 1, 2, 0, 0, 0, 0, 0, 1, 3, 2, -1, -1, -2, 0, -1, -4, -6, -6, -6, -5, -6, -7, -6, -5, -3, -4, -3, -3, -1, -1, 0, 0, 2, 1, 0, 0, 0, 0, 1, 3, 3, 4, -1, -2, -3, -1, -3, -3, -4, -6, -6, -6, -5, -6, -5, -4, -3, -3, -3, -3, -2, 0, -1, 0, 1, 1, 0, 1, 1, 2, 2, 3, 2, 2, -1, -2, -1, -1, -2, -3, -5, -5, -5, -6, -6, -6, -5, -3, -2, -3, -4, -3, -1, -1, 0, 0, 0, 1, 0, 2, 3, 2, 3, 2, 1, 2, 0, -1, -1, -1, -2, -3, -4, -5, -6, -5, -5, -6, -4, -4, -3, -3, -1, -2, -1, 0, 0, 0, 0, 1, 0, 0, 1, 3, 2, 0, 0, 0, 0, -1, -1, -2, -2, -3, -4, -4, -5, -6, -6, -5, -5, -4, -2, -2, -1, -3, -2, -2, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -1, -3, -3, -3, -5, -4, -5, -5, -4, -5, -4, -2, -2, -2, -3, -4, -3, -1, -1, -2, -2, -1, -1, 0, 0, 0, -1, -2, 0, 0, -3, -2, -3, -3, -2, -3, -3, -3, -4, -2, -4, -2, -1, 0, -1, -3, -4, -4, -3, -1, -2, -1, 0, -1, 0, -1, -1, -1, -1, -1, -1, -1, -3, -4, -2, -2, -1, -1, -1, -1, -1, -2, -2, 0, 0, 0, -2, -2, -2, -3, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -3, -4, -3, -2, -1, -1, 0, -1, 0, -2, 0, 0, 0, 0, -1, -3, -1, 0, 1, 2, 0, 0, 0, 0, -1, -1, -1, 0, -1, -2, 0, -1, -2, -4, -2, -2, -1, 0, 0, 1, 0, 0, 0, 1, 0, -1, -1, -2, -2, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -3, -2, -1, -1, 0, 0, 1, 2, 2, 1, 1, 1, 1, 0, 0, -1, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, -1, -2, -3, 0, 0, 0, 1, 2, 2, 2, 1, 2, 2, 0, 2, 1, 1, 1, 0, 1, 0, 1, 1, 0, 0, 2, 1, 3, 2, 0, 0, 0, -1, -2, -3, -1, 0, 1, 1, 3, 3, 5, 4, 2, 2, 0, 1, 1, 1, 1, 1, 2, 1, 2, 2, 1, 1, 1, 1, 2, 2, 1, 0, 0, 0, -2, -1, 0, 0, 0, 1, 4, 4, 4, 5, 4, 3, 2, 1, 1, 2, 1, 2, 2, 1, 1, 1, 1, 1, 1, 2, 2, 2, 0, 0, 0, 0, -1, -1, 0, 0, 0, 2, 3, 4, 4, 3, 4, 2, 1, 1, 1, 1, 1, 2, 2, 1, 0, 1, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 2, 1, 2, 1, 3, 3, 2, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 1, 1, 2, 2, 1, 2, 1, 1, 2, 1, 1, 0, -1, -1, 0, -1, -1, -1, -2, -2, -2, -1, -1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 3, 1, 2, 1, 1, 0, 0, 0, -2, -3, -4, -4, -3, -2, -4, -3, -5, -5, -3, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 3, 2, 2, 1, 1, 0, 0, -1, -2, -3, -4, -3, -2, -3, -5, -4, -3, -5, -3, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 2, 2, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, -2, -3, -3, -4, -4, -3, -2, 0, 1, 0, 0, 0, 1, 0, 1, 0, -1, 0, 1, 1, 1, -1, 0, -1, -2, -2, -1, -2, 0, -1, -1, 0, -1, -2, -3, -4, -3, -3, -1, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 1, 0, 1, 0, -2, -3, -2, -3, -3, -2, -1, 0, 1, 1, 0, 0, -1, -2, -3, -2, -1, 0, 0, 0, 0, 2, 1, 2, 1, 0, 3, 3, 3, 1, 1, 0, 0, -2, -3, -3, -2, -2, 0, 0, 0, 1, 0, 0, 0, -2, -2, -2, -2, 0, 1, 0, 1, 3, 2, 2, 1, 1, 4, 4, 4, 3, 3, 0, 0, -1, -2, -3, -1, -1, 0, 1, 0, 0, -1, 0, -1, -1, -3, -1, 0, 0, 1, 0, 0, 2, 1, 0, 0, 2, 2, 3, 4, 3, 3, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -2, -1, 0, 1, 2, -1, 0, 0, 0, 0, 0, 1, 1, 2, 4, 2, 1, 1, 0, 0, -1, 0, 1, 1, -1, -2, -2, -1, -3, -1, -2, 0, -1, 0, 0, 0, 1, -1, 0, -1, -1, -3, -2, -2, 0, 0, 0, 2, 1, 0, -1, -2, 0, 0, 0, 0, -2, -1, -3, -3, -1, -3, 0, -1, -1, 0, 0, 0, 1, 0, -1, -1, -2, -3, -3, -3, -3, -1, 0, 0, 0, -1, -1, -2, -1, 0, 1, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, -1, -2, -4, -5, -5, -4, -2, -2, 0, 0, 0, 0, 0, -1, 0, 0, 2, 1, 0, 1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, -2, -2, -3, -5, -5, -6, -5, -3, -3, -2, 0, 1, 1, 3, 0, 1, 1, 1, 2, 1, 1, 1, 2, 2, 3, 2, 3, 2, 0, 0, 1, 0, 0, 0, -2, -4, -6, -7, -7, -5, -3, -1, 1, 1, 1, 3, 2, 3, 2, 3, 0, 0, 0, 2, 3, 2, 2, 3, 2, 1, 0, 1, 0, 0, 0, 0, 0, -4, -4, -6, -7, -4, -2, -1, 0, 1, 2, 2, 2, 3, 2, 3, 1, 0, 0, 2, 2, 3, 3, 2, 2, 2, 1, 2, 1, -1, 0, 0, -1, -4, -6, -7, -8, -4, -2, -1, 0, 1, 0, 2, 3, 3, 2, 2, 0, 1, 0, 1, 3, 3, 3, 3, 3, 4, 2, 2, 1, 0, 0, 1, -1, -4, -4, -5, -5, -6, -3, -2, 0, 0, 0, 1, 2, 1, 2, 0, 0, 0, 1, 2, 3, 4, 4, 3, 3, 4, 2, 2, 1, 0, 0, 1, -1, -4, -4, -4, -3, -4, -2, 0, 0, 0, 0, 1, 1, 2, 1, -1, 0, 1, 1, 2, 3, 5, 4, 3, 2, 3, 1, 1, 0, 1, 1, 0, 0, -2, -4, -2, -2, -2, -1, 0, 1, 0, 1, 1, 1, 0, 0, 0, -1, 0, 1, 2, 2, 3, 3, 1, 1, 2, 0, 1, 0, 0, 1, 1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, 0, 1, 1, 2, 3, 3, 1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 2, 1, 2, 3, 3, 4, 4, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 4, 2, 2, 1, 3, 2, 1, 1, 2, 4, 4, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 5, 4, 3, 4, 4, 3, 3, 4, 2, 2, 3, 0, 0, -1, -2, 0, 0, 2, 1, -1, 0, 1, 0, 1, 0, 1, 1, 0, 0, 1, 0, 1, 5, 5, 3, 5, 4, 5, 4, 3, 3, 1, 0, 0, 0, -1, -1, 0, 1, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 1, 2, 4, 4, 3, 3, 4, 4, 4, 3, 3, 1, 1, 1, 1, 0, 0, 0, 0, 2, 1, 2, 2, 1, 1, 0, -1, -1, -2, -1, 0, 1, 1, 1, 3, 3, 2, 2, 3, 4, 3, 2, 2, 2, 2, 1, 2, 2, 0, 0, 0, 2, 2, 1, 2, 0, 0, -1, -1, -3, -1, -1, -2, 0, 0, 0, 2, 1, 1, 1, 1, 2, 1, 2, 2, 2, 3, 2, 2, 2, 0, -1, 0, 0, 0, 1, 0, -1, -1, -2, -4, -4, -4, -3, -3, 0, 1, 0, 2, 0, 1, 1, 1, 0, 0, 0, 1, 2, 2, 3, 2, 0, 0, -1, -2, -1, 0, -1, -1, -3, -4, -4, -6, -7, -6, -4, -3, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, -1, 0, -2, -3, -3, -2, -3, -5, -5, -6, -6, -6, -4, -3, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 2, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 2, 1, 1, 1, 0, 0, 1, 2, 1, 0, 0, 2, 2, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 2, 0, 1, 1, 0, 0, 2, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, 1, 1, 2, 0, 1, 0, 0, 1, 1, 1, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -3, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -2, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 1, 0, 0, 0, 0, 2, 1, 2, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 2, 2, 3, 3, 3, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 2, -1, 0, 0, 1, 1, 1, 2, 3, 2, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 2, 0, -1, -1, 0, 2, 3, 2, 2, 2, 3, 2, 0, 0, -1, -2, -1, 0, 0, -2, -2, -1, -1, -2, -1, -1, 1, 0, 0, -1, -1, 1, 1, 0, -1, -1, 0, 2, 3, 2, 1, 1, 3, 3, 1, 0, 0, 0, 0, 0, 0, -1, -2, -3, -4, -2, 0, -1, 0, 1, 1, 0, 0, 1, 0, 0, -1, 0, 0, 1, 1, 3, 2, 1, 2, 2, 1, 0, 0, 0, -1, -1, 0, -1, -2, -3, -2, -2, -1, 0, 0, 1, 1, 0, 0, 0, 2, 0, 0, 0, 1, 0, 1, 2, 1, 1, 1, 1, 2, 1, 0, -1, -1, -2, -2, -3, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 1, 3, 3, 1, 1, 2, 3, 2, 1, 0, 0, 0, -1, -3, -3, -3, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 2, 3, 3, 4, 3, 3, 3, 1, 1, 0, 0, 0, -1, -1, -2, -2, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 1, 0, 2, 4, 4, 3, 3, 3, 3, 1, 1, 0, 0, -1, -2, -3, -3, -3, -1, -1, -1, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 1, 2, 2, 3, 2, 1, 2, 3, 3, 0, 0, 0, 0, 0, -2, -3, -3, 0, -1, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 2, 3, 1, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, -3, -4, -3, -2, 0, -1, -2, 0, 1, 1, 1, 0, 0, 1, 0, -1, 0, 1, 0, 1, 1, 0, 1, 0, 0, 1, 0, -1, -2, -2, -2, -3, -2, -3, -2, -1, 0, -1, 0, -2, 0, 0, 2, 1, 0, 0, 0, 0, 0, 2, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, -1, -2, -3, -1, -3, -3, -2, -2, 0, -2, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -3, -1, -2, -3, -2, -2, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 2, 2, 3, 2, 2, 0, 0, 1, 2, 0, 0, 0, -2, -2, -1, 0, -2, -2, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 2, 1, 1, 2, 1, 0, 0, 0, 2, 0, 0, 0, 0, -1, 0, -1, 0, -2, -2, -1, -2, -2, -1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, -2, -1, -1, -1, -1, -1, 0, 0, 1, 0, 1, 0, 0, 3, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 3, 3, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 1, 0, 0, -1, 0, -1, 0, 0, 0, 2, 1, 0, 0, 1, 0, 2, 3, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 0, 1, 2, 2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 2, 1, 1, 1, 2, 1, 2, 1, 1, 0, 1, 2, 0, 2, 2, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 0, 1, 1, 0, -1, 0, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 1, 1, 1, 1, 1, 0, 0, 0, -1, -1, 0, -1, -2, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 1, 0, 1, 0, 0, -1, -2, -1, -1, 0, 0, -2, -1, -1, 0, -3, -1, 0, 1, 1, 1, 0, 1, 0, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, -1, -1, 0, 0, 0, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 1, 0, 1, 0, 1, 1, 1, 0, -1, 0, 0, -1, -1, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 1, 2, 1, 1, 1, 2, 1, 1, 0, 0, -1, -1, -2, -2, -2, -2, 0, -2, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 2, 0, 0, 1, 0, 0, 3, 2, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 2, 1, 1, 1, 2, 2, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 1, 2, 2, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 1, 1, 0, 0, 0, -2, -1, -2, -1, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 2, 1, 2, 1, 1, 0, 0, 0, -1, 0, -1, -1, -2, -2, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 1, 2, 1, 1, 1, 0, 1, 1, 2, 1, 3, 2, 1, 0, 0, 0, 0, 0, -1, -2, -3, -2, -2, -1, 0, 1, 1, 1, 1, 2, 1, 1, 1, 0, 0, 0, 0, 2, 2, 2, 3, 2, 1, 3, 1, 0, 0, 0, 0, 0, 0, -2, -2, -2, 0, 0, 1, 1, 2, 0, 0, 1, 1, 2, 1, 2, 0, 0, 1, 1, 2, 2, 1, 1, 2, 3, 1, 0, 0, 0, 0, -1, -2, -2, -2, -1, 0, 0, 0, 1, 2, 1, 0, 2, 2, 2, 0, 1, 0, 2, 2, 2, 3, 2, 2, 2, 3, 3, 1, 1, 2, 1, 0, -1, -1, -2, -2, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 1, 1, 2, 1, 2, 3, 3, 3, 2, 3, 1, 1, 2, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 2, 1, 3, 2, 1, 0, 1, 2, 1, 1, 2, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 2, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 0, 0, 0, 1, 0, 0, 0, 1, 0, 2, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 1, 0, 2, 4, 1, 2, 2, 2, 2, 1, 1, 1, 1, 1, 2, 2, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 3, 1, 1, 2, 1, 2, 0, 1, 2, 2, 3, 2, 1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 3, 3, 2, 3, 4, 3, 2, 1, 2, 2, 3, 2, 1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 2, 0, 0, 0, 1, 1, 1, 3, 3, 2, 2, 4, 3, 3, 1, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 1, -1, 0, 0, 0, 1, 4, 3, 2, 2, 2, 3, 1, 2, 1, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 3, 3, 2, 2, 2, 1, 1, 0, 2, 2, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 2, 2, 2, 2, 2, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, -1, -1, 0, -1, 0, 0, -1, -1, -2, -3, -3, -2, -3, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -2, -3, -1, -4, -3, -1, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -2, -2, -1, -1, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 2, 1, 1, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 4, 6, 5, 3, 3, 3, 3, 3, 2, 3, 3, 3, 3, 1, 1, 2, 2, 4, 3, 2, 2, 1, 0, 0, 0, 0, 0, 2, 3, 0, -1, 0, 2, 3, 3, 2, 1, 2, 3, 4, 4, 5, 3, 4, 4, 3, 3, 3, 4, 4, 2, 3, 2, 1, 1, 0, 0, 1, 1, 3, 4, 0, 0, 0, 1, 2, 2, 2, 2, 1, 3, 4, 4, 3, 3, 4, 3, 4, 3, 3, 3, 2, 0, 1, 0, 0, 1, 0, 0, 1, 3, 2, 2, 1, 0, 0, 0, 2, 3, 4, 3, 2, 2, 1, 0, 2, 1, 3, 2, 3, 3, 3, 1, 1, 0, -1, 0, 1, 0, 1, 0, 1, 3, 3, 2, 2, 0, 0, 2, 3, 3, 3, 3, 1, 0, 0, 1, 1, 0, 0, 1, 1, 2, 0, 0, 0, 0, -1, 0, 1, 1, 2, 1, 2, 2, 2, 3, 2, 1, 1, 2, 3, 3, 4, 4, 3, 2, 2, 2, 1, -1, -1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 2, 1, 2, 0, 0, 0, 2, 1, 0, 0, 1, 4, 4, 5, 5, 6, 3, 4, 3, 4, 2, 1, 1, 1, 1, 0, -1, 0, 0, 0, 0, 2, 3, 3, 3, 2, 0, 1, 1, 0, -1, -1, 1, 4, 6, 4, 5, 6, 5, 4, 2, 1, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 1, 1, 0, 1, 2, 1, 0, 0, 1, 0, 0, 0, 1, 4, 4, 3, 3, 4, 4, 4, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -2, 0, 0, 0, 0, 1, 4, 3, 3, 4, 2, 3, 4, 2, 0, 0, 0, 1, 0, 1, 0, 0, -1, -1, -2, -2, -2, -2, 0, -1, 0, -1, 0, 0, 2, 3, 0, 1, 3, 4, 3, 3, 1, 1, 3, 4, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, -2, -1, -1, -2, -2, 0, 0, -1, 0, 1, 2, 1, 0, 0, 0, 2, 2, 2, 3, 1, 1, 3, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, -2, -2, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 1, 2, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, -1, -3, -1, -2, -1, -3, -1, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 2, 0, 0, 0, 0, 2, 1, 1, 2, 1, 2, 1, 1, 0, 0, 1, 1, 1, 0, -1, 0, -1, 0, 1, 1, 0, 0, 2, 4, 4, 3, 2, 3, 1, 0, 0, 1, 2, 4, 2, 2, 2, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 3, 5, 4, 3, 3, 3, 4, 2, 1, 2, 2, 2, 4, 4, 3, 2, 2, 2, 3, 1, 1, 0, -1, -2, -2, -2, -1, 0, 1, 1, 0, 1, 2, 3, 2, 1, 0, 0, 1, 2, 2, 0, 1, 1, 0, 0, 1, 2, 3, 2, 0, 0, 0, 0, -1, 0, 0, 0, 2, 1, 2, 1, 0, 1, 2, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 1, 0, 0, 2, 1, 2, 1, 0, 1, 1, 3, 1, 0, 2, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 2, 0, 1, 2, 0, 0, 1, 1, 0, 1, 1, 2, 2, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, 0, 1, 0, 1, 1, 1, 0, 0, 1, 1, 3, 2, 3, 1, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, -2, -2, 0, 0, 1, -1, 0, 0, 0, 1, 2, 4, 3, 2, 2, 2, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, -2, -1, -2, -1, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 4, 3, 4, 4, 3, 3, 2, 2, 0, 0, 1, 1, 1, 2, 2, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 4, 3, 3, 3, 3, 3, 2, 2, 2, 2, 3, 3, 2, 1, 0, 1, 0, 1, -1, -1, -2, -1, -1, -1, 0, 1, 1, 2, 2, 2, 0, 1, 5, 3, 3, 2, 2, 3, 3, 2, 2, 3, 2, 1, 2, 0, 0, 0, 0, 0, 0, -2, -2, -1, -2, 0, 0, 1, 2, 4, 1, 2, 1, 2, 6, 6, 3, 4, 3, 4, 3, 1, 1, 1, 0, 1, 0, 0, 2, 1, 0, 0, 0, -1, -1, 0, 0, -1, 1, 1, 3, 3, 4, 3, 2, 0, 4, 5, 3, 3, 2, 2, 2, 2, 0, 0, 0, 0, 1, 1, 2, 2, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 3, 4, 3, 3, 2, 1, 1, 2, 2, 2, 1, 1, 3, 2, 1, 2, 1, 1, 1, 3, 2, 3, 2, 0, 0, 1, 1, 1, 2, 2, 3, 3, 4, 4, 3, 2, 2, 0, 1, 1, 0, 0, 2, 2, 1, 1, 3, 2, 3, 1, 1, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 2, 1, 0, 0, 0, 0, -1, 0, 0, 3, 3, 2, 1, 0, 1, 1, 2, 1, 3, 4, 4, 3, 3, 2, 0, 0, 0, -1, -1, -2, -3, -3, -2, -3, -3, -3, -2, -3, -3, -2, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 1, 1, 2, 2, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 2, 2, 0, 2, 2, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 2, 1, 0, 1, 1, 2, 1, 2, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 3, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 1, 1, 0, 1, 0, 0, 1, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 1, 0, 1, 1, 1, 0, 0, 1, 2, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 1, 1, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, -1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 2, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 1, 0, 1, 2, 2, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 1, 0, 2, 1, 1, 1, 1, 0, 1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 1, 2, 2, 2, 1, 1, 1, 2, 1, 0, -1, -1, -1, -2, -1, -1, -1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 1, 2, 0, 0, 0, 2, 0, 0, 2, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 1, 0, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 2, 1, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 1, 2, 2, 2, 1, 1, 1, 3, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -1, 0, 0, -1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, -1, 0, -1, 0, 0, 2, 1, 0, 1, 1, 1, 0, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 2, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, -2, 0, -1, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 2, 2, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -2, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 2, 2, 1, 2, 1, 2, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 2, 2, 2, 1, 2, 3, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 2, 3, 2, 2, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, -1, 0, 0, 1, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 2, 0, 1, 1, 1, 1, 1, 1, 0, 1, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 0, 2, 1, 1, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 1, 0, 1, 0, 1, 1, 2, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 2, 2, 2, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 3, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 2, 1, 1, 2, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 2, 2, 3, 2, 0, 1, 1, 0, 1, 0, 2, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 2, 3, 2, 2, 2, 1, 3, 1, 1, 0, 1, 1, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 2, 3, 3, 3, 3, 3, 3, 2, 2, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 3, 3, 2, 3, 2, 2, 2, 1, 2, 1, 1, 2, 3, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 3, 2, 2, 1, 3, 1, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 3, 1, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 1, 1, 1, 2, 1, 0, 1, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -2, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -2, 0, -1, 0, 1, 2, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, -2, -1, -2, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -2, -1, -2, -1, -1, -2, -1, -2, -1, -2, -1, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -1, -1, -3, 0, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -2, 0, -2, -2, -2, -1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -2, -2, -1, -1, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, -1, -1, -2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -3, -2, 0, -1, -1, 0, 0, 0, -1, -1, -3, -1, -1, 0, -1, -2, 0, 0, 2, 0, 0, 0, 0, 1, 0, 0, 1, 1, -1, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, -2, -2, -1, 0, 0, -2, 0, 0, 2, 1, 0, 0, 0, 0, 1, 0, 2, 0, -1, 0, -2, 0, -1, 0, -1, 0, -1, -1, 0, -1, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, -2, 0, -2, -1, 0, 0, -1, 0, -1, -1, -3, -2, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, -1, -2, 0, 2, 0, 1, 0, -1, -2, -1, 0, 0, -1, -2, 0, 0, -1, -2, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -3, -1, -1, 0, -2, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -3, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -3, -2, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -2, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 1, -1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, -2, -4, -3, -1, -1, 0, 2, 1, 1, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 1, 0, 1, 0, -1, -2, -3, -3, -3, -2, -1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 2, 0, 0, 0, 0, 1, -1, -2, -3, -4, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 2, 2, 1, 1, 2, 2, 0, 0, 0, 1, 1, -1, -3, -3, -3, -3, -3, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, 1, 1, 2, 1, 2, 1, 1, 1, 1, 0, 1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, 0, 1, 2, 1, 1, 2, 1, 0, 0, 1, 0, 2, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -2, -1, -1, 0, 0, 1, 1, 1, 0, 1, 0, -1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, -1, -2, -3, 0, 0, 0, -1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, -2, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 1, 1, 0, 1, 0, 2, 1, 2, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 1, 0, 2, 2, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, -2, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 3, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 3, 3, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 3, 3, 1, 2, 1, 2, 1, 1, 1, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 2, 2, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -1, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -1, 0, 1, 0, 0, 0, -1, -1, -2, -1, -1, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -2, -1, -2, -3, 0, -2, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -1, 0, -1, -2, -1, -3, -2, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -2, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 2, 2, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, -1, 0, 1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, -1, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 2, 0, -1, -1, -2, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, -2, -1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 0, -1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, -1, 0, 0, 0, 1, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 2, -1, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, -1, 1, 0, 0, 1, 0, -2, 0, -1, 0, 0, 0, -2, -1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, -1, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, -1, -2, -1, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, -1, -1, 0, 0, 0, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, -1, -2, 0, 0, -1, -1, -1, -1, 0, -1, 0, -2, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -2, -1, -1, 0, 1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -2, 0, 0, 0, 0, -1, -2, -1, -1, -3, -1, -1, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -3, -2, 0, 1, -1, -1, -2, -2, -3, -3, -2, -2, 0, 0, -1, 0, 0, 2, 1, 0, 0, 1, 0, -1, 0, 0, 1, -1, -1, 0, 0, -2, -4, -1, 0, 0, -1, -2, -2, -1, -3, -4, -4, -3, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, -1, -1, 0, 0, -4, -3, -2, -1, 0, -2, -2, -2, -1, -3, -3, -4, -2, -1, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, -2, -2, -2, 0, -1, -3, -3, -2, -1, -1, -3, -3, -2, -2, -1, -2, -3, -3, -1, 0, 0, 0, 1, 2, 0, 0, 0, 1, 0, 0, -1, -1, -1, -3, -2, -1, 0, -3, -4, -2, 0, -2, -3, -2, -2, -2, -2, -2, -1, -2, -2, 0, -1, 0, 2, 2, 1, 0, 0, 1, -1, 0, 0, 0, -2, -3, -3, -1, 0, -3, -4, -2, -2, -2, -4, -3, -3, -3, -1, 0, -1, -1, -1, 0, 0, -1, 1, 0, 1, 1, 0, 1, -1, -1, 0, 0, -2, -3, -3, -3, -4, -4, -2, -2, -1, -2, -3, -3, -2, -2, -2, -1, 0, -1, -2, -1, 0, 0, 1, 0, 2, 2, 0, 0, 0, -1, 0, 1, 0, -2, -2, -3, -4, -3, -3, -2, -3, -2, -2, -3, -2, -3, -2, -1, 0, 0, -1, -1, -1, 0, 2, 1, 1, 3, 0, 1, 0, -1, 0, 0, 0, -1, -2, -3, -4, -4, -2, -1, -3, -1, -1, -3, -2, -1, -2, -1, 0, 0, -2, -1, -1, 1, 2, 0, 2, 3, 0, 2, 0, -2, -1, 0, 0, -1, -2, -3, -6, -3, -2, -2, -2, -2, -3, -3, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, 2, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -4, -4, -5, -2, 0, -2, -3, -4, -2, -3, -3, -3, -1, -1, 0, 0, 0, 0, 0, 3, 2, 1, 3, 0, 0, 1, 0, 0, 1, 0, 0, -2, -3, -4, -3, -2, 0, 0, -4, -4, -3, -2, -2, -1, -1, 0, 1, 0, -1, 0, 0, 1, 0, 2, 2, 0, -2, 1, 1, 0, 0, 0, -1, -1, -3, -3, -2, -1, 0, -1, -4, -5, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 0, -1, 1, 1, 0, 1, -1, 0, -1, -3, -1, -3, 0, 0, 0, -4, -5, -2, -2, -1, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 2, 2, 0, 0, 2, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, 0, -1, -3, -3, -3, -3, 0, -1, -3, -2, 0, -2, 0, 0, 0, 0, 0, 1, 3, 0, 0, 1, 0, 0, 1, 0, -2, -2, -1, 0, -2, -1, -1, -1, -4, -1, -1, -2, -1, -2, -3, -2, 0, -2, -1, 0, 0, 0, 0, 1, 3, 0, 0, 2, 0, 0, 0, 0, 0, -3, -2, -1, -2, -3, 0, -3, -3, -2, -2, -2, -1, -3, -1, -1, 0, -3, -1, 0, 0, -1, 0, 2, 1, 0, 0, 1, 0, -1, 0, -1, -1, -1, -3, -1, -3, -3, -1, -2, -3, -1, -1, -2, -2, -2, -2, 0, -2, -2, -1, 0, 0, 0, 0, 1, 2, 0, 1, 3, 0, -1, -1, 0, 0, -2, -3, -3, -2, -3, -2, -2, -2, -2, -3, -3, -2, -2, -3, -1, -2, -2, -1, 0, 0, 0, 0, 1, 2, 0, 0, 2, 0, -2, 0, -1, -1, -2, -1, -2, -1, -1, 0, -3, -1, -3, -3, -3, -4, -3, -2, -3, -3, -2, 0, 0, 0, 0, 0, 1, 3, 0, 0, 3, 0, -2, 0, 0, -1, -2, -3, -2, -1, -1, 0, -3, -1, -3, -3, -3, -2, -3, -3, -3, -4, -2, 0, 0, 0, 0, 0, 0, 3, 0, 0, 3, 0, -2, 0, 0, 0, -2, -2, -2, 0, 0, 0, -2, -1, -1, -2, -3, -3, -1, -2, -3, -4, -4, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, -2, -2, 0, -1, -1, 0, -2, -2, -1, -2, -1, -4, -2, -2, -2, -2, -2, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, -2, -2, 0, 0, -1, -2, -1, 0, -2, -2, -2, -1, 0, 0, 0, -1, -3, -2, -2, -2, -2, -1, 1, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, -2, -2, -1, -1, -1, 0, -1, -1, -1, 0, -1, -2, -2, -1, 0, 0, 0, 2, 0, 1, 0, 1, -1, 1, 0, 1, 0, 0, -2, -1, -1, -2, -2, -2, -1, -1, -2, 0, -1, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 3, 1, 0, 1, 1, -2, -1, 0, 1, 1, 0, -2, -2, -1, -2, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 2, -3, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 2, 1, 1, 0, 1, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 1, 2, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 2, 1, 2, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, -2, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 2, 3, 2, 4, 3, 2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 3, 4, 3, 2, 0, 1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 2, 2, 3, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, -1, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 1, 2, 2, -1, -2, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, -1, -1, 0, -1, 0, -1, -2, 0, 0, 0, 0, 0, 2, 1, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, -2, -2, -1, -2, -2, -1, 0, 1, 2, 2, 1, 1, 3, 3, 2, 2, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, 1, 2, 2, 3, 3, 3, 2, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, -1, -1, -1, -1, -2, -1, 1, 0, 1, 3, 2, 3, 2, 4, 2, 1, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 2, -1, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 2, 3, 2, 1, 2, 2, 2, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, -1, -1, 0, -1, -1, 0, -1, -2, -1, 0, 0, 0, 1, 2, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 2, 2, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 2, 2, 2, 1, 0, 0, 1, 0, 1, -1, 0, 1, 0, -1, -1, 0, -2, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, -1, 1, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, -1, -2, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, -1, 0, -1, 0, 0, 0, -1, 0, 1, 1, 1, 2, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, -2, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, -1, 0, -2, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 1, -1, 0, 1, 0, 0, 1, 0, 1, 1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 0, 2, 2, 2, 2, 1, 0, 0, 1, 2, 1, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 2, 1, 2, 1, 1, 2, 1, 2, 2, 2, 1, 1, 0, 0, 0, 2, 1, 2, 0, 0, 0, 0, 0, 0, 1, -1, 0, 1, 1, 0, 1, 0, 1, 1, 0, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, 0, -1, -1, -2, -2, -2, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, -2, -1, -2, -1, -2, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, -2, -1, -2, -2, -1, -2, -2, -2, -1, -2, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, -2, -2, -3, -2, -1, -2, -3, -2, -2, -1, -2, -1, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, -2, -2, -2, -1, -2, -2, -2, -1, -3, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -3, -3, -1, -2, -2, -2, -2, -2, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, -2, -1, -3, -2, -1, -1, -1, -1, -1, 0, -2, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -1, -1, -2, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -2, -1, -2, -1, -2, -1, -2, -1, -2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, -2, -1, -2, -1, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, -1, 0, -2, -2, -2, -1, -1, -2, -2, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -2, -1, -2, -1, -2, -1, -2, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -2, -2, -2, -1, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -2, -1, 0, -1, -1, -1, -2, -2, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, -1, -2, -2, -2, 0, -1, 0, -1, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -2, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 1, 1, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, -2, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, -2, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, -2, 0, 0, 0, -1, -1, -1, -2, -1, -1, -2, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -2, 0, 0, 0, -1, 0, -2, -2, 0, 0, 0, -1, -1, -1, -1, -1, -2, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, -2, -1, -2, -1, -1, 0, -1, -2, -1, 0, 0, 0, 0, -1, -1, -1, -2, -2, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, -1, 0, -1, -2, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -2, -1, -1, -1, -1, 0, -1, -1, -2, 0, -2, 0, 0, 0, 0, 0, -1, -1, -2, 0, -2, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, 0, -1, -1, 0, -1, -1, 0, -2, -1, -1, 0, -1, -1, 0, 0, -1, 0, -2, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -2, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -2, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, -1, -1, -1, 0, -1, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -2, -1, -1, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, -2, -2, 0, 0, 0, -2, -1, -1, -1, 0, -2, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -2, -1, -2, 0, -1, -2, 0, 0, -1, -1, -1, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 2, 2, 2, 1, 1, 0, 1, 0, 0, -1, -2, -1, -2, -1, -2, -1, -1, -3, -2, -1, -2, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 1, 1, 2, 3, 3, 3, 1, 0, 1, 0, 0, 0, -1, -1, -2, -1, -1, -1, -1, -1, -2, -1, 0, 1, 1, 0, 1, 1, 1, 1, 0, 0, 1, 1, 2, 3, 2, 1, 1, 0, 0, 0, 0, -2, -2, -1, 0, -1, -1, -2, -1, -2, 0, -1, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 1, 2, 1, 2, 1, 1, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, -2, -2, -1, 0, -2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, -1, -1, -1, -2, -2, 0, 0, 0, 0, 0, 1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 0, 1, 1, 2, 1, -1, -1, -1, -2, -3, -1, -1, -2, 0, 0, 0, 0, 0, -1, -2, -2, -1, 0, 0, 0, 1, 1, 1, 1, 2, 2, 4, 3, 4, 4, 2, 1, -1, -1, -3, -2, -3, -2, -1, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, 0, 0, 1, 0, 2, 2, 0, 1, 3, 3, 4, 4, 3, 2, 2, 0, 0, -3, -2, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -2, 0, 1, 2, 1, 0, 0, 0, 0, 2, 1, 2, 3, 3, 3, 1, 1, -1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 3, -1, 0, 0, -1, -1, 0, 1, 1, 2, 2, 2, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 3, 2, 0, -1, -2, -2, -1, -1, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 2, 3, 3, 0, -1, -2, -3, 0, -2, -2, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 1, 2, 0, -1, -2, -2, -2, -3, -4, -4, -1, -2, 0, -1, 0, 0, 0, 0, 2, 2, 2, 1, 1, 1, 2, 1, 1, 1, 0, 0, 2, 1, 0, 0, -1, -1, -3, -2, -2, -4, -4, -4, -3, -1, -1, 0, 1, 2, 1, 2, 2, 3, 2, 2, 1, 2, 2, 3, 2, 2, 1, 2, 2, 1, 0, 0, 0, -1, 0, 0, -3, -3, -4, -4, -3, -1, -1, 0, 0, 2, 3, 3, 3, 2, 3, 1, 2, 2, 2, 3, 3, 3, 1, 1, 2, 2, 1, 1, 0, -1, 0, 0, -2, -3, -5, -5, -3, -1, 0, 0, 0, 2, 2, 2, 2, 4, 3, 2, 1, 3, 3, 2, 3, 2, 1, 1, 1, 2, 1, 2, 0, 0, 0, -1, -3, -3, -3, -3, -1, -1, 0, 0, 1, 1, 2, 2, 3, 4, 2, 3, 1, 2, 3, 2, 2, 2, 3, 3, 4, 3, 1, 2, 0, 0, 0, 0, -3, -2, -3, -4, -2, -1, 0, 0, 1, 2, 2, 2, 2, 2, 2, 1, 2, 3, 1, 3, 4, 4, 4, 4, 3, 2, 1, 3, 0, 0, 0, -1, -2, -3, -2, -2, -1, -1, 0, 0, 1, 1, 2, 2, 2, 1, 0, 0, 1, 2, 3, 3, 4, 3, 3, 2, 3, 1, 1, 1, 0, 0, 1, 0, -3, -2, -1, -1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, -1, 0, 2, 0, 1, 2, 2, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 2, 2, 1, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 1, 1, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 1, 0, 2, 1, 2, 1, 3, 3, 1, 3, 2, -1, -2, -1, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 2, 0, 1, 3, 2, 1, 2, 1, 2, 3, 2, 4, 3, 2, 1, 0, -1, -2, -2, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 2, 4, 3, 3, 1, 4, 3, 3, 3, 3, 2, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 2, 0, 2, 4, 4, 2, 3, 4, 3, 2, 2, 1, 2, 1, 0, 0, 0, -1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 3, 2, 2, 4, 4, 4, 3, 2, 3, 3, 2, 2, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, 0, -1, 0, 1, 1, 1, 2, 1, 3, 2, 4, 3, 3, 3, 3, 2, 2, 2, 3, 1, 1, 1, 0, 0, 0, 2, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 2, 1, 1, 2, 3, 3, 1, 2, 2, 3, 3, 1, 3, 3, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -3, -3, -1, -2, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 1, 1, -1, -1, -2, 0, -1, -1, -3, -4, -3, -4, -5, -5, -2, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -2, -2, -1, -4, -4, -4, -4, -4, -4, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 1, 2, 1, 1, 3, 2, 3, 2, 1, 1, 1, 1, 0, 2, 1, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 2, 2, 1, 3, 2, 2, 1, 3, 2, 0, 2, 0, 0, 0, 1, 1, 1, 0, 0, 2, 2, 1, 0, 2, 2, 0, 2, 0, -1, 0, 1, 1, 2, 1, 0, 1, 1, 1, 2, 3, 2, 2, 2, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 2, -1, -1, 0, 0, 1, 1, 1, 2, 1, 1, 2, 0, 1, 2, 1, 2, 1, 1, 1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 2, 2, 1, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 1, 1, 3, 1, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 1, 2, 1, 0, -2, 0, -1, -1, -1, 0, -1, -1, 0, 0, -1, -1, -2, -1, -1, -2, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 1, 1, 0, -1, -1, -1, -1, 0, -1, -1, -1, 0, -1, -1, -3, -1, -1, -2, -1, -1, 0, 0, 0, 0, -1, 0, -2, -1, -1, 0, 0, 1, 1, 3, 0, -1, -1, -2, -2, -1, -2, -2, -2, -1, -2, -2, -1, -3, -2, -1, -2, -3, -2, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 2, 2, 0, -1, -1, -1, -1, -1, -1, -2, -2, -1, -1, -2, 0, -1, -3, -2, -2, -4, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 0, 0, -1, -1, 0, 0, -1, -1, -1, -1, -1, -3, -1, -2, -3, -2, -2, -2, -2, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 3, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -2, -2, -2, -2, -2, -2, -2, -1, -2, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 3, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -1, -3, -1, -1, -2, -3, -2, -2, -1, -1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -3, -1, -2, -2, -3, -3, -2, 0, -1, 0, 1, 1, 0, 0, 1, 0, 0, 1, 2, 2, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, -2, -2, -2, -1, -2, -2, -1, -1, -2, 0, 0, 1, 1, 0, 0, 0, 0, 1, 2, 2, 2, 0, 0, 0, 1, 1, -1, -2, -1, 0, -1, 0, -1, -1, -1, -2, -3, -2, -3, -1, -2, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 3, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, -2, 0, 0, -1, -3, -1, -1, 0, -1, 0, 0, 2, 0, 0, 0, 0, 1, 2, 1, 2, -1, -1, 0, 0, 1, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, -2, -2, -1, -1, -1, -1, 0, 0, 1, 0, -1, 0, 0, 0, 2, 1, 2, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, -1, -1, 0, 1, 0, 0, -1, 0, 0, 0, -2, -1, -2, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, -2, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, -2, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, -1, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, -1, -1, -2, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, -1, -2, -3, -2, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -2, -1, -1, -2, -1, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, -1, -1, -2, -2, -1, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, -2, -1, -1, -1, -1, 0, 1, 1, 2, 1, 1, 2, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 2, 0, 0, 1, 1, 1, 2, 1, 2, 0, 1, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 2, 2, 0, 0, 1, 2, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 1, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 2, 1, 1, 1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, -2, -1, 0, 0, 0, 1, 2, 1, 1, 3, 3, 2, 2, 2, 1, 1, 1, 1, 1, 0, 2, 0, 1, 1, 2, 2, 2, 2, 2, 2, 0, -1, -2, -2, 0, 0, 0, 1, 2, 3, 2, 4, 3, 3, 3, 2, 1, 2, 1, 1, 0, 1, 0, 1, 2, 1, 2, 1, 2, 2, 1, 2, 0, 0, -2, -1, -1, 0, 0, 0, 1, 2, 1, 1, 2, 2, 3, 2, 2, 2, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 1, 0, 1, 1, 1, 0, -1, -3, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 1, 1, 1, -1, -1, -2, -2, -2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 2, 3, 2, -1, -2, -4, -3, -2, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 2, 1, 2, 0, -1, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, -2, -2, -1, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 2, 0, -3, -3, -4, -3, -1, -1, 0, 0, 0, 0, -1, -1, -2, -2, -1, -2, -3, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, -1, -2, -2, -3, -3, -2, -3, -2, -2, -1, -1, -2, -3, -4, -3, -3, -1, -3, -2, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 2, -1, -1, -2, -3, -1, -2, -3, -2, -1, -2, -2, -3, -3, -2, -2, -3, -3, -2, -3, -2, 0, -1, 0, 0, 0, 0, -2, -1, 0, 0, 2, 3, 0, -2, -2, -1, -2, -2, -4, -3, -3, -1, -2, -2, -3, -3, -2, -3, -2, -2, -1, -2, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 1, 1, 0, -1, -2, -2, -1, -3, -3, -2, -3, -3, -3, -2, -3, -2, -1, -1, -2, -1, -2, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, -2, -2, -1, -1, -2, -2, -4, -2, -2, -3, -4, -3, -3, -3, -2, -1, -2, -1, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 0, -3, -2, -1, -1, -1, -2, -4, -2, -2, -2, -3, -2, -2, -3, -2, -1, -2, 0, 0, 0, 0, 1, 1, 1, -1, -1, -1, 0, 0, 1, 0, -2, -2, 0, 0, 0, -2, -3, -2, -2, -2, -3, -3, -2, -2, -1, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 2, 2, -2, -2, -1, 0, -1, -2, -3, -4, -2, -2, -1, -3, -2, -1, -1, -2, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 1, 0, -1, 0, 0, -1, -3, -4, -2, -3, -2, -3, -2, -3, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 2, 1, -1, -1, -1, 0, -1, -2, -3, -4, -3, -3, -1, -2, -1, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 1, 1, 0, -1, -1, -1, 0, -3, -4, -4, -3, -3, -2, -2, -2, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, -1, -2, -1, -2, -3, -4, -2, -3, -3, -1, -2, -1, -1, -1, -2, 0, 0, 0, -1, -1, -1, -1, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, -2, -2, -2, -3, -3, -2, -2, -2, -2, -1, -1, 0, 0, -1, -1, -3, -2, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, -2, -2, -1, -2, -3, -3, -2, -2, -2, -1, -1, -1, -1, -1, 0, -2, -2, -2, -1, -2, 0, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, -2, -2, -2, -1, -2, -1, -2, -1, -1, 0, 0, 0, -1, 0, -1, -2, -1, 0, -1, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -3, -2, -2, -2, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, -1, -1, -1, -1, 0, 1, 2, 2, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 2, 1, 0, 2, 0, -1, -2, 0, 0, 0, 0, 0, 2, 2, 1, 1, 2, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 1, 1, 2, 2, 1, 1, 2, 0, 0, -1, 0, 0, 0, 0, 0, 1, 3, 3, 2, 2, 1, 0, 0, 1, 0, 1, 2, 1, 1, 0, 0, 0, 1, 1, 1, 0, 2, 0, 1, 0, 0, -1, 0, -1, -1, 1, 0, 2, 1, 1, 1, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -2, -2, -3, -2, -1, -2, -2, -3, -2, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -3, -2, -2, -2, -4, -3, -4, -3, -2, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -2, -2, -3, -1, -3, -2, -3, -4, -4, -4, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, -2, -2, -2, -3, -3, -2, -3, -2, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -2, -1, -3, -2, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, -2, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, -1, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 3, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 2, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, -2, 0, 0, 0, 0, -1, 0, 1, -2, 0, -1, -2, -2, 0, 0, 2, 2, 2, 2, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -2, -1, -2, -2, -1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, -2, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -2, -3, -2, -2, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -3, -2, -3, -2, -1, 0, 1, 2, 1, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, -1, -3, -4, -4, -3, -2, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 2, 2, 1, 0, -1, 0, 0, 1, 0, -1, -2, -2, -3, -4, -3, -2, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 1, 2, 1, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, -2, -2, -3, -3, -2, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 1, 2, 2, 2, 1, 2, 1, 1, 0, -1, 0, 1, 0, -1, 0, -3, -3, -2, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 1, 2, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 1, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 2, 1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 1, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 2, 1, 0, 0, 2, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, -1, -1, -2, -1, -2, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, -3, -2, -1, 0, 0, 2, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, -1, 0, -1, 1, 1, 0, 0, -1, -1, -3, -1, -2, -3, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, -2, -2, -3, -3, -3, -3, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, -2, 0, -1, -2, -3, -3, -2, -4, -3, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, 2, 1, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 2, 2, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, -1, 0, 0, 0, -2, 0, 2, -1, -1, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, 1, 0, 0, 0, 0, 1, 2, 0, 0, -1, -1, -2, -1, 1, 0, -1, -2, -1, 0, -1, -2, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 1, 0, 0, 1, 0, 2, 0, 0, -2, -2, -2, -2, 0, -1, -1, -2, 0, 0, -4, -3, -1, 0, 1, -1, -1, -2, -2, -2, -2, -3, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, -1, -1, -1, -2, -1, 0, -1, -2, 0, 0, -3, -3, -1, 0, -1, 0, -2, -1, -1, -2, -3, -3, -1, 0, 0, -1, 0, 0, 0, 2, 0, 0, 0, 0, -2, -1, 0, -1, 0, 0, 0, -1, -3, -2, 0, 0, -1, -1, -1, -1, -2, -1, -2, -2, -2, -1, -1, 0, 0, 2, 0, 2, 0, 0, -1, -2, -1, -1, 0, -1, -1, -1, 0, 0, -3, -3, -1, -1, -3, -4, -3, -2, -2, -1, 0, -1, -2, 0, 0, 0, 0, 2, 0, 3, 0, 0, -1, -1, -1, 0, 0, -2, -3, -2, 0, 0, -2, -2, -2, -2, -2, -3, -2, -3, -2, -1, 0, 0, 0, -2, -2, 0, 0, 1, 0, 2, 0, 0, 0, -2, -1, 0, 0, -3, -2, -3, -1, -2, -2, -3, -2, 0, 0, -2, -4, -2, -1, 0, 0, -1, 0, -1, -1, -1, 0, 2, -1, 3, 0, 0, 0, -2, -2, -1, 0, -1, -2, -2, -3, -4, -2, -1, -3, -1, 0, -2, -3, -3, -1, -2, 0, 0, 0, 0, 0, 0, 1, 1, -1, 4, 0, 1, 0, -2, -1, 0, -1, -1, -2, -2, -3, -3, -1, -2, -2, -2, -1, -3, -4, -3, -2, -3, -2, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, -2, -1, -1, 0, -1, -1, -2, -1, -4, -3, -1, 0, -1, -2, -2, -3, -2, -2, -3, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, -1, -1, -1, 0, 1, -1, -1, 0, -3, -3, -2, -1, -1, -1, -2, -2, -3, -2, -2, -1, 0, 1, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, -1, -1, 0, 1, 0, 0, 0, -1, 0, -1, -2, -1, -1, -1, -3, -2, -2, -2, 0, -1, 0, 2, 1, 0, 1, 1, 0, 2, 0, 1, 0, 1, -2, 0, 0, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, -1, -3, -2, -2, -1, -1, 0, -1, 0, 2, 1, 0, 0, 0, 0, 0, 3, 1, 0, -2, 0, 1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -3, -2, -1, -2, 0, -1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 2, 0, 0, -1, 1, 0, 0, 0, -1, -1, 0, 0, -1, -2, -1, 0, -2, -3, -2, -2, 0, 0, 0, -2, 0, 1, 0, 1, 2, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, -1, -2, -1, 0, -2, -3, -2, -1, -1, -1, -2, 0, 0, 0, -1, 1, 1, 0, 0, 1, 2, 0, 0, -1, 2, 0, 0, -1, -1, -1, -2, 0, -1, -3, -1, -1, -1, -2, -1, -1, -2, -2, -2, -1, 0, -1, -2, 0, 0, 0, 0, 0, 2, 1, 0, 0, 2, 0, 0, 0, -1, -2, -2, -2, 0, -1, -3, -2, -2, -3, -1, -2, -2, -2, -1, -1, 0, -1, -2, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, -2, 0, -1, -2, -1, -3, -1, -2, -1, 0, -2, -1, -1, -2, -2, -3, -2, -2, -1, -2, -2, 0, 0, 1, 0, 1, 1, 0, 0, 1, 2, -1, -1, 0, -1, 0, -1, -1, -1, -1, -1, -1, 0, -2, -2, -4, -3, -3, -2, -3, -2, -2, -1, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, -1, -1, -1, 1, -1, -1, -3, 0, 0, 0, 0, -1, -1, -2, -3, -3, -2, -1, -2, -3, -1, -2, 0, 1, 0, 0, 0, 2, 0, 0, 0, 0, 0, -2, 0, 0, -2, -2, -3, 0, 0, 0, 0, -2, -2, -2, -4, -2, -1, -2, -2, -3, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, -1, -1, 0, -2, -2, -1, -1, 0, 0, -1, -1, -2, -1, 0, -2, -2, -1, -2, -3, -2, -1, 0, 0, 0, 0, 0, 2, 0, 0, -1, 0, -1, 0, 0, 0, -1, -2, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, -2, -2, -1, -1, 0, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, -2, -2, -1, 0, -1, -1, -1, 0, 0, -2, -1, 0, 0, -1, 0, 0, -1, -1, -2, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, -1, -1, -2, 0, -1, -1, -2, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 1, 1, 1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 0, 1, 0, 0, 0, 2, 1, 1, 1, 2, 2, 1, 2, 1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 2, 2, 4, 3, 3, 2, 4, 3, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, -2, 0, -1, -1, 0, 0, 1, 1, 2, 2, 2, 2, 2, 1, 3, 3, 4, 3, 2, 3, 2, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 1, 1, 2, 2, 2, 1, 1, 0, 3, 2, 1, 2, 2, 2, 2, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 3, 2, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 3, 2, 2, 2, 2, 0, 1, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 1, 2, 3, 3, 2, 3, 3, 3, 2, 1, -1, 0, -2, -1, 0, -1, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 2, 4, 4, 4, 3, 3, 3, 3, 3, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 3, 2, 0, -1, 0, 1, 2, 3, 5, 4, 3, 3, 4, 2, 2, 0, 0, 0, 0, -2, 0, -1, 0, 1, 1, 1, 1, 1, 1, 2, 1, 0, 0, 2, 1, 0, 0, 1, 2, 3, 3, 3, 3, 5, 3, 3, 2, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, 1, 2, 3, 2, 2, 3, 4, 3, 3, 0, 0, 0, 0, 1, 1, 0, 0, -1, -2, -1, 0, 0, 0, 1, 1, 1, 0, 1, 2, 1, 2, 0, 1, 2, 4, 3, 3, 1, 1, 2, 3, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 3, 2, 0, 0, 0, 1, 2, 1, 2, 2, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 2, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 1, 0, 2, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 0, 0, 1, 2, 0, 1, 1, 1, 1, 2, 0, 0, 0, 1, 1, 1, 2, 2, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 3, 3, 3, 2, 1, 1, 2, 2, 2, 1, 2, 1, 2, 1, 0, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, 1, 2, 0, 0, 0, 1, 1, 0, 1, 1, 3, 2, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 2, 1, 2, 2, 3, 3, 1, 1, 1, 1, 2, 0, 2, 1, 1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 2, 4, 3, 0, 1, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 3, 2, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 4, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 1, 1, 1, 3, 4, 2, 1, 1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 2, 5, 3, 3, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 1, 2, 0, 2, 3, 3, 2, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 1, 0, 1, 0, 2, 1, 1, 1, 2, 2, 3, 1, 2, 1, 1, 1, 1, 0, 0, 0, 1, 2, 0, 2, 0, 2, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 2, 2, 1, 1, 1, 1, 1, 2, 0, 0, 1, 0, 1, 1, 0, 1, 1, 2, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -2, -1, 0, 0, 2, 2, 1, 2, 1, 1, 1, 1, 0, 0, 1, 1, 2, 2, 2, 1, 0, 0, -1, 0, -1, -2, -2, -2, -1, -1, -2, -3, -2, -2, -3, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 2, 0, 1, 2, 1, 0, 1, 0, 0, 2, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 2, 2, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 2, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 0, 1, 1, 1, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 2, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 2, 0, 0, 0, 1, 0, -2, -1, -1, -1, 0, 0, 0, 0, 1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -2, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 2, 1, 1, 1, 1, 2, 1, 1, 1, 0, 0, 0, 0, 1, 0, 2, 1, 0, 1, 0, 0, 2, 1, 0, 0, -1, 0, 1, 0, 1, 1, 0, 0, 1, 1, 2, 0, 0, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -2, -2, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -2, -2, -1, -2, -1, -3, -3, -3, -3, 0, 0, -2, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, -2, -2, -2, -1, -2, -2, -4, -5, -2, 0, -1, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -2, -2, -4, -3, -4, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, -1, -1, 0, 0, 0, -1, 0, -1, -2, -2, -3, -4, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -2, -2, 0, 0, -1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 1, 1, 1, 0, 0, -1, -2, -1, -2, -1, 0, 0, -2, 0, 0, 0, -1, 0, 0, 0, 1, 2, 1, 2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 1, 0, -1, -1, -1, 0, -1, -2, 0, 1, 0, 2, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, -2, 0, -1, -3, -2, -2, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, -3, -2, -2, -2, -2, -3, -2, -2, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, -1, -1, -2, -3, -3, -4, -2, -3, -3, -1, -1, 0, -1, 0, -1, -2, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, -1, -2, 0, 0, 0, -1, -1, -3, -2, -3, -4, -4, -4, -2, -1, -1, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, -2, -3, -4, -4, -4, -4, -3, -1, -2, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 0, 0, -1, -1, 0, 0, -1, 0, -1, -3, -4, -5, -5, -5, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 2, 1, 2, 2, 1, 0, 0, 0, 0, -1, 0, -2, -3, -4, -5, -6, -4, -3, -2, -1, -1, -1, 0, -1, 0, 0, 0, -1, -2, -1, 0, 1, 3, 1, 3, 2, 1, 0, 0, 1, -1, -1, -1, -2, -2, -5, -6, -5, -5, -4, -3, -1, -2, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 3, 2, 2, 2, 3, 0, 0, 0, -1, -2, -1, -2, -3, -4, -6, -5, -5, -3, -4, -2, -1, -2, 0, 0, 1, 0, -1, -1, -2, 0, 1, 2, 2, 1, 2, 1, 2, 0, -1, 0, -1, 0, 0, -2, -2, -4, -4, -4, -4, -4, -3, -1, -1, 0, 0, 0, 1, 0, -1, -1, 0, 1, 1, 2, 1, 1, 1, 1, 1, 0, -1, 1, 0, 0, 0, -1, -1, -3, -2, -3, -2, -3, -1, -1, 0, 0, 0, -1, 0, 0, -2, -1, 0, 2, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 1, -1, 0, -2, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, -1, -2, -2, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, -2, -1, 0, 0, 1, 1, 0, 0, 0, -2, -2, -2, -3, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, -2, -2, -3, -3, -3, -3, -4, -2, -1, 0, -1, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, -1, -1, -2, -1, -3, -4, -4, -5, -5, -5, -1, -1, 0, 0, -2, -2, -2, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, -2, -1, -2, -2, -2, -1, -1, -2, -2, -4, -4, -3, -3, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 1, 1, 2, 2, 3, 3, 2, 2, 2, 1, 2, 4, 3, 3, 2, 2, 0, 1, 1, 1, 0, 2, 2, 2, 1, 3, 1, 2, 1, 2, 2, 0, 1, 0, 1, 2, 3, 1, 2, 2, 1, 0, 3, 3, 2, 2, 2, 2, 1, 2, 1, 0, 0, 1, 1, 1, 2, 3, 2, 2, 2, 2, 3, 1, 0, 1, 1, 2, 1, 1, 2, 2, 1, 0, 2, 2, 2, 2, 1, 1, 2, 2, 1, 1, 0, 1, 0, 1, 2, 3, 2, 0, 2, 2, 3, 2, 0, 0, 1, 1, 0, 1, 1, 1, 1, 0, 1, 1, 0, 1, 2, 0, 1, 1, 2, 1, 1, 0, 0, 1, 2, 3, 1, 1, 0, 3, 2, 2, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 1, 1, 2, 1, 0, 0, 2, 4, 1, 1, -1, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 1, 0, 0, 0, 2, 1, 2, 1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, -1, -1, -1, 0, 0, 0, 1, 1, 2, 1, 0, -1, 0, 0, 0, 0, 1, 2, 2, 3, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -2, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 1, 1, 1, 1, 3, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, -1, -1, -1, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, -1, 0, 0, -2, -2, -1, 0, 1, 0, 1, 0, 1, 0, 0, 1, 1, 2, 4, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 1, 1, 2, 1, 0, 0, 1, 1, 4, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, 0, 0, -1, -1, 0, -1, -2, -2, -1, 1, -1, 1, 2, 3, 1, 0, -1, 0, 0, 3, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, -2, -3, 0, 0, 0, 1, 0, 3, 1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -2, -2, 0, 0, 1, 1, 2, 2, 1, 1, 1, 1, 3, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -2, -2, -2, -1, 0, 0, 0, 0, 1, 1, 2, 1, 2, 1, 0, 1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, -2, -1, 0, -1, 0, 0, 1, 1, 0, 0, 1, 1, 2, 2, 2, 0, 0, -1, 1, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, -1, -3, -1, -1, -1, -1, 0, 1, 1, 0, 0, 0, 1, 1, 1, 3, 0, 1, -1, 0, 2, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, -2, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 2, 1, 1, 2, 3, 0, 0, -2, 0, 3, 2, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 2, 1, 0, -1, 1, 2, 1, 1, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 0, 0, -1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 2, 0, 0, -2, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, -1, 0, 2, 0, 0, 0, 0, 1, 0, 0, -2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -3, -1, -1, -1, 0, 1, 1, 1, 0, 0, 0, 2, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, -1, 0, -4, -2, -3, -3, 0, 0, 1, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, -4, -2, -2, -2, 0, 2, 2, 1, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 1, 2, 0, 1, -1, 0, -3, -1, -1, -2, 0, 2, 2, 0, 1, 1, 2, 2, 0, 0, 1, 1, 1, 2, 2, 1, 1, 0, 1, 1, 1, 0, 2, 1, 2, 2, 0, 0, -2, 0, -2, -2, 1, 2, 2, 1, 2, 1, 3, 2, 0, 0, 2, 2, 2, 2, 2, 0, 0, 1, 1, 0, 1, 2, 2, 2, 3, 1, 0, 0, 0, -1, -2, -1, 0, 2, 3, 1, 2, 2, 2, 1, 1, 2, 1, 2, 2, 3, 4, 1, 1, 2, 3, 2, 2, 2, 3, 1, 3, 1, 0, 0, 0, -1, -1, -1, 0, 1, 2, 1, 1, 2, 3, 2, 2, 2, 1, 2, 2, 4, 4, 2, 2, 2, 1, 1, 2, 3, 2, 2, 4, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 2, 2, 3, 3, 2, 3, 2, 2, 2, 3, 3, 4, 3, 2, 2, 3, 3, 3, 3, 2, 2, 4, 1, 0, 0, 0, 0, 1, 0, 2, 3, 1, 1, 2, 2, 2, 2, 3, 2, 3, 2, 3, 2, 3, 3, 2, 3, 3, 2, 2, 2, 3, 4, 3, 1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 0, 0, 1, 2, 1, 1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 2, 3, 4, 4, 3, 4, 3, 2, 2, 2, 1, 1, 0, 1, 1, 2, 1, 3, 2, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 1, 2, 2, 2, 3, 5, 5, 4, 4, 3, 3, 3, 2, 2, 1, 0, 0, 0, 1, 2, 3, 2, 2, 1, 1, 0, 0, 0, -2, -1, -1, 0, 1, 1, 1, 2, 2, 3, 3, 3, 3, 4, 3, 2, 2, 1, 0, 0, 0, 1, 0, 2, 3, 3, 1, 0, 1, 2, 2, 0, -1, -2, -1, -1, 0, 1, 1, 0, 2, 1, 2, 2, 4, 3, 3, 2, 1, 1, 0, 0, 0, 0, 0, 0, 3, 2, 1, 2, 1, 2, 1, 0, 0, -2, -2, -1, 0, 1, 0, 0, 0, 1, 2, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 1, 2, 1, -1, -3, -1, -2, 0, 1, 1, 0, 2, 1, 1, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, -2, -3, -3, -2, -1, 0, 1, 1, 1, 1, 1, 0, 0, 0, -1, -3, -2, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, 1, 0, 2, 1, -1, -2, -1, -1, -1, 0, -1, 0, 0, 0, 0, -2, -3, -2, -3, -2, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 1, 2, -1, -2, -1, -2, -2, 0, -1, -1, 0, -1, -1, -3, -3, -4, -4, -3, -2, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 3, 2, 0, 0, -2, -2, -1, -1, -3, -2, -1, 0, -1, -2, -2, -2, -3, -4, -2, -3, -1, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, 0, 2, 2, 0, -1, -2, -2, -1, -3, -5, -4, -3, -2, -3, -3, -2, -2, -2, -1, -3, -2, -1, 0, 0, 0, 1, 1, 0, -1, 0, -1, 0, 0, 1, 0, -1, 0, 0, -1, -1, -4, -4, -5, -3, -3, -4, -3, -2, -1, -2, -2, -1, -2, 0, 0, 0, 2, 3, 1, 1, 0, 0, 0, -1, 0, 0, 1, 0, -1, -1, 0, -1, -2, -4, -4, -3, -3, -2, -3, -2, -2, -2, -2, 0, 0, 0, 0, 0, 2, 3, 2, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, -2, -4, -3, -3, -3, -4, -4, -2, -2, -2, -1, 0, 0, 0, 0, 0, 3, 4, 2, 1, 0, 0, 1, 1, 0, 1, 0, -1, -2, -1, 0, 0, -2, -3, -4, -3, -4, -3, -2, -2, -2, -2, -1, -1, 0, 0, 1, 1, 2, 2, 2, 1, 0, 1, 1, 1, 0, 1, 1, 0, -1, -1, 0, 0, -2, -3, -3, -4, -4, -2, -4, -2, -1, 0, -1, -1, 0, 0, 1, 1, 1, 2, 2, 0, 0, 0, 1, 3, 3, 1, 1, -1, -2, 0, 0, -1, -3, -4, -3, -3, -3, -3, -2, -2, 0, -1, 0, -1, 0, 1, 2, 1, 2, 2, 1, 0, 2, 2, 3, 4, 4, 2, 2, -2, -2, -1, 0, -2, -2, -4, -4, -2, -3, -2, -4, -1, 0, -1, -1, -1, 0, 1, 0, 1, 1, 1, 2, 1, 1, 2, 2, 4, 3, 3, 1, 0, -1, -1, 0, -1, -2, -3, -3, -3, -3, -4, -3, -1, -2, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 3, 1, 0, 0, 0, -1, -2, -1, -1, -2, -2, -2, -3, -4, -2, -3, -3, -2, -1, -2, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 1, 0, 1, 0, 0, 0, 0, -2, 0, -1, -2, 0, -1, -3, -2, -3, -3, -3, -2, -2, -2, 0, -1, -1, -1, -1, -1, -1, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, -2, -1, -1, -2, -2, -1, -2, -1, 0, 0, 0, -2, -2, -3, -2, -1, -1, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -2, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -3, -3, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, -2, -1, -2, -2, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -2, -2, -1, 0, 0, 0, 2, 2, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 1, 1, 3, 2, 2, 2, 2, 2, 2, 1, 0, 1, 0, 1, 1, 1, 2, 0, 1, 2, 1, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 1, 2, 3, 2, 3, 3, 3, 1, 2, 1, 1, 1, 1, 2, 1, 1, 1, 1, 1, 0, 2, 1, 2, 0, 0, 1, -1, 0, -2, -1, 0, 0, 1, 2, 4, 3, 3, 4, 2, 1, 1, 1, 0, 0, 2, 0, 1, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 1, 2, 2, 2, 2, 2, 3, 3, 2, 0, 1, 1, 2, 2, 2, 1, 0, 0, 1, 0, 1, 1, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 2, 0, 2, 2, 2, 0, 1, 2, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -2, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, -2, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, -1, -2, -1, 0, 0, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -1, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 2, 1, 0, 0, 0, -2, -1, 0, 0, 0, -1, -2, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -1, 0, -1, 0, 0, 0, -1, -1, 0, 1, 0, 0, 2, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, -2, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, -2, -2, -1, 0, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -2, -1, -1, -1, 0, 0, 2, 1, 1, 1, 0, 2, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -2, -1, -3, -3, -2, -1, 0, -2, -2, -1, 0, 1, 2, 1, 0, 1, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -2, -2, -2, -3, -3, -3, -3, -2, -4, -4, -2, 0, 0, 3, 1, 1, 1, 2, 0, 0, 1, 1, 1, 0, 0, 0, 2, 1, 0, -1, 0, -2, -1, -1, -2, -4, -4, -3, -3, -3, -4, -5, -2, -1, 2, 2, 1, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, -1, -1, -2, -1, -2, -1, -3, -3, -3, -2, -2, -2, -2, -3, -2, 0, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, -1, 0, 0, -1, -2, -3, -2, -2, -2, -2, -2, -2, -3, -3, -1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, -1, -2, -2, 0, -1, -1, -1, 0, 0, 0, -1, -1, -2, -1, -1, -2, -1, 0, 0, -1, -2, -1, 0, 2, 2, 2, 2, 1, 0, 0, 2, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 2, 3, 3, 2, 1, 1, 1, 3, 2, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 1, 1, 2, 1, 0, 2, 2, 4, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 1, 1, -1, 0, 0, 0, 1, 1, 1, 2, 3, 3, 3, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 3, 2, 1, 2, 1, 1, 0, -1, 0, 0, 1, 0, 1, 0, 1, 3, 4, 1, 2, 2, 1, 1, 1, 0, 0, 0, 0, -1, 0, 1, 1, 1, 3, 3, 2, 2, 2, 0, 0, 0, -1, 0, 1, 0, 0, 1, 2, 1, 2, 3, 2, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 2, 2, 4, 4, 2, 2, 1, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, -1, -1, -1, 0, 0, 0, 1, 0, 1, 1, 2, 4, 3, 3, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 2, 1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 2, 3, 3, 3, 2, 1, 1, 0, -1, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 1, 2, 2, 0, -1, 0, 0, 0, 1, 2, 1, 1, 2, 2, 3, 3, 2, 2, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, 1, 1, 0, 2, 2, 4, 3, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 2, 2, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 1, 1, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 3, 2, 3, 1, 1, 0, 1, 0, -1, 1, 1, 0, 0, -1, -2, -1, -2, 0, 0, 1, 1, 2, 1, 1, 0, 0, -1, 0, 1, 1, 2, 2, 3, 4, 2, 0, 0, 0, 0, 0, -1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 2, 2, 1, 1, 1, 3, 2, 1, 0, 0, 0, 0, 0, 2, 2, 1, 0, 1, 0, 0, 0, 0, 1, 0, 2, 1, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 2, 1, -1, 0, 0, 0, 0, 2, 2, 1, 2, 0, 1, 1, 0, 0, 1, 2, 3, 2, 1, 0, 0, -1, 1, 0, 2, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 3, 2, 1, 3, 1, 0, 0, 1, 0, 3, 3, 4, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 3, 3, 1, 1, 3, 1, 0, 2, 0, 1, 3, 2, 3, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, -1, 0, 3, 5, 1, 1, 1, 1, 0, 0, 0, 1, 2, 1, 2, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 5, 4, 3, 2, 2, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, -1, -1, 0, -1, -1, -1, -2, -2, 0, 0, 4, 5, 3, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, -1, -1, -1, -2, -2, -1, -3, -2, 0, 2, 3, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 0, 0, 0, -1, -1, -2, -1, -1, -2, 0, 0, 2, 2, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, -1, -3, -2, -1, -2, -3, -1, 0, 0, 2, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -4, -3, -2, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -1, -1, -1, -1, -2, -3, -3, -2, -2, -2, -3, -3, -2, -1, 2, 0, 1, 0, 0, 3, 2, 1, 2, 2, 1, 0, 1, 1, 2, 1, 0, 0, 2, 1, 2, 3, 2, 1, 2, 2, 4, 3, 2, 2, 2, 2, 2, 0, 1, 0, 1, 2, 1, 2, 3, 3, 2, 0, 1, 1, 3, 1, 1, 2, 2, 2, 2, 3, 2, 2, 3, 2, 2, 3, 2, 2, 3, 1, 2, 2, 2, 2, 2, 1, 0, 2, 1, 2, 1, 0, 0, 1, 1, 0, 0, 1, 1, 2, 3, 4, 1, 2, 3, 3, 3, 1, 1, 1, 3, 2, 2, 1, 3, 1, 3, 3, 2, 3, 1, 1, 2, 1, 1, 3, 0, 0, 0, 0, 0, 3, 3, 2, 1, 1, 1, 3, 2, 1, 1, 1, 1, 1, 2, 2, 2, 1, 1, 1, 2, 3, 3, 1, 1, 0, 1, 4, 3, 1, 1, 0, 0, 1, 2, 3, 3, 0, 0, 2, 2, 2, 1, 1, 2, 2, 1, 1, 2, 1, 1, 1, 1, 3, 3, 1, 0, 0, 1, 4, 4, 2, 1, 2, 1, 0, 2, 2, 1, 0, 0, 2, 2, 2, 1, 0, 2, 2, 0, 2, 2, 1, 0, 0, 1, 1, 1, 0, 1, 1, 2, 2, 2, 1, 1, 1, 1, 0, 0, 2, 0, -1, -1, 0, 1, 1, 1, 1, 2, 2, 0, 2, 1, 1, 0, 0, 0, 1, 1, 2, 2, 0, 2, 3, 2, 0, 2, 2, 0, 0, 1, 1, 1, 0, 0, 0, 1, 2, 1, 0, 1, 1, 0, 2, 4, 3, 0, 1, 2, 2, 2, 1, 2, 2, 2, 1, 3, 1, 2, 2, 0, -1, 0, 0, 2, 1, -1, 0, 1, 3, 1, 0, 1, 1, 2, 2, 2, 3, 2, 2, 0, 1, 0, 1, 1, 3, 4, 3, 2, -1, 0, 1, 0, -1, 0, 1, 1, 3, 0, 0, 2, 3, 1, 0, 1, 1, 1, 1, 3, 3, 1, 1, 0, -1, 0, -1, 0, 0, 2, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, -1, 0, 2, 1, -1, -1, 0, 1, 0, 3, 2, 0, 0, 2, 0, 0, -2, 0, 0, 2, 1, -1, -2, -1, 0, -1, 0, 0, 1, 2, 1, 0, -1, 0, 1, 0, -1, -1, 0, 1, 2, 3, 2, 0, 0, 1, 2, 0, -1, 0, -1, 0, 1, 0, -1, -1, -1, -1, -1, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 3, 3, 0, 1, 1, 2, 2, 0, 0, 1, 0, 1, 0, 1, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, -1, 1, 2, 0, 0, 0, 1, 0, 2, 3, 1, 2, 0, 2, 1, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, -1, -2, -1, 1, 1, 1, 1, 1, 1, 2, 3, 2, 2, 2, 3, 2, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -2, -3, -2, 1, 1, 0, 0, 1, 2, 5, 3, 2, 2, 2, 3, 1, 0, 0, 0, 1, 1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 1, 0, 3, 4, 3, 4, 3, 5, 2, 2, 1, 0, 2, 2, 0, -1, -2, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 2, 3, 2, 3, 3, 4, 4, 2, 1, 1, 1, 1, 0, -2, -3, 0, 0, 0, 0, 0, 1, 1, 2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 3, 1, 2, 1, 0, 1, 2, 1, 1, 0, 0, 0, -1, -4, -4, -2, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 2, 0, 0, -1, -1, 0, 0, 0, -2, -3, -2, -3, -2, -3, -2, 0, 0, 1, 0, 1, 0, 3, 2, 1, 4, 2, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -2, -2, -1, -1, -1, -2, -2, -1, 1, 0, -1, 0, 0, 2, 2, 1, 1, 3, -1, 0, 1, 1, 0, 1, 1, 2, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, 1, 2, 1, 1, 2, 2, 0, 0, 0, 1, 0, 0, 2, 2, 0, 0, -1, 1, 0, 0, -1, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 1, 1, 0, 0, 2, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 2, 1, 2, 0, 1, 2, 1, 1, 2, 2, -1, 1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, -1, 0, 1, 2, 1, 2, 3, 3, 2, 1, 1, 2, 0, 1, 0, 0, 0, 0, 1, 1, 2, 1, 1, 2, 4, 3, 2, 1, 0, 1, 0, 1, 0, 0, 1, 0, 1, 1, 2, 3, 3, 2, 1, 2, 1, 1, 0, 0, 0, 0, 1, 2, 3, 2, 1, 2, 2, 2, 4, 3, 2, 0, 0, 2, 2, 2, 1, 1, 2, 2, 4, 2, 2, 2, 2, 3, 2, 2, 2, 1, 1, 1, 1, 2, 1, 1, 0, 1, 2, 1, 2, 4, 4, 2, 2, 2, 3, 2, 2, 1, 1, 3, 4, 4, 3, 4, 4, 3, 1, 2, 1, 1, 0, 1, 1, 3, 1, 1, 0, 2, 3, 2, 3, 2, 4, 4, 4, 4, 4, 4, 4, 3, 3, 4, 4, 5, 5, 3, 3, 1, 0, 0, 0, 0, 0, 0, 0, 3, 3, 2, 1, 1, 2, 2, 2, 2, 3, 3, 3, 4, 4, 3, 4, 3, 4, 5, 5, 4, 4, 5, 3, 3, 1, 0, 1, 1, 1, 1, 0, 1, 1, 1, 1, 0, 1, 0, 0, 1, 1, 0, 1, 1, 1, 2, 2, 2, 1, 2, 2, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 2, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 0, 1, 2, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 1, 0, 0, 1, 2, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 2, 1, 2, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 2, 2, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 2, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 0, 1, 1, 1, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 2, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 2, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 2, 2, 1, 2, 1, 0, 0, 1, 2, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 0, 0, 1, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 1, 0, 2, 0, 0, 1, 1, 2, 0, 1, 1, 1, 1, 1, 1, 1, 0, 0, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 2, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 0, 1, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 1, 1, 1, 2, 2, 1, 1, 0, 0, 0, 0, -1, 0, 1, 0, 2, -1, 0, 2, 2, 1, 0, 0, 0, -1, 0, 0, -1, -2, -1, -1, 1, 2, 2, 2, 1, 1, 4, 3, 0, 0, -2, 0, 0, 0, 1, 1, 0, -2, 0, 1, 0, 0, 0, 0, 1, 0, -2, -1, -2, -3, -2, -1, 0, 0, 0, 1, 2, 2, 4, 4, 0, 2, 0, -1, 0, 0, 0, 0, 0, -2, 0, 0, -2, -3, 0, 0, 0, -1, -1, -3, -2, -2, -3, -2, -1, 0, 0, 0, 1, 1, 2, 4, 0, 1, -1, 0, 0, 0, 1, 0, -1, -2, 0, 1, -5, -5, -3, 0, 0, 0, -3, -2, -1, -2, -4, -4, -1, 0, 0, 0, 0, 1, 2, 5, 0, 0, 0, -1, 0, 0, 1, 0, -1, -2, 0, 0, -4, -4, -2, -1, -1, -2, -3, -2, -3, -4, -5, -4, -3, 0, -1, -2, -1, 0, 2, 3, 1, 0, 0, 0, -1, -2, 0, 0, -2, 0, 0, 0, -5, -4, -2, 0, -3, -4, -4, -1, -3, -5, -3, -3, -3, 0, -2, 0, 0, 2, 1, 3, 0, 0, 1, -1, -1, -2, 0, -1, -1, -1, 0, -1, -3, -5, -1, -1, -3, -5, -5, -4, -2, -2, -1, -2, -2, -1, -2, -1, 0, 3, 3, 4, 0, 1, 1, 0, -1, -1, 0, -1, -2, -1, 1, 0, -4, -5, -2, -3, -5, -6, -6, -6, -3, -1, 0, -1, -2, -1, -1, -2, 0, 2, 2, 6, 1, 1, 0, -1, -1, 0, 0, -1, -3, -2, -1, -3, -3, -4, -3, -3, -3, -6, -7, -5, -3, -2, 0, 0, -1, -1, -1, -1, -1, 1, 0, 6, 0, 0, 0, -2, -1, 0, 0, -2, -2, -4, -3, -4, -4, -3, -5, -2, -1, -4, -6, -3, -2, -2, 0, 0, 0, 0, 0, -1, 0, 1, 0, 6, 0, 2, -1, -3, -1, 0, 1, -2, -3, -3, -5, -5, -3, -3, -3, -2, -2, -4, -5, -4, -4, -3, -2, 0, 0, 0, 0, -1, 0, 2, 0, 4, 0, 2, 0, -4, 0, 0, 0, -1, -2, -2, -5, -6, -3, -2, -3, -2, -3, -5, -7, -2, -4, -4, -2, -1, 0, 0, 0, 0, 1, 2, 0, 4, 0, 1, 0, -3, -1, 1, 2, 0, -1, -1, -4, -7, -6, -3, -2, -4, -6, -5, -5, -2, -3, -3, -2, -2, -1, 0, 1, 0, 0, 2, 1, 5, 0, 1, 0, -1, 0, 1, 2, 0, -1, -1, -3, -4, -3, -4, -2, -4, -5, -6, -5, -4, -3, -3, -1, -1, 0, 0, 0, 0, 1, 2, 1, 5, 0, 1, -2, 0, 0, 1, 2, 0, -1, -2, -2, -2, -3, -3, 0, -2, -6, -5, -4, -4, -3, -3, -2, 1, 2, 0, 0, 0, 0, 1, 0, 5, 0, 0, -2, 1, 1, 0, 0, -1, 0, -1, -3, -2, -1, -1, 0, -2, -6, -6, -4, -3, -2, -2, -3, 1, 0, 0, 0, 0, 0, 0, 1, 6, 0, 0, -1, 2, 1, 0, 0, -2, -1, 0, -1, -2, -3, -1, 0, -2, -4, -5, -5, -3, -2, -2, -2, 0, 0, -2, 0, 0, -1, 0, 0, 6, 0, 0, -1, 2, 2, 0, 0, -2, 0, 0, -1, 0, -3, -3, 0, -4, -4, -4, -4, -3, -2, -3, -3, -1, 0, -2, -1, 0, -1, 0, 0, 4, 1, -1, 0, 2, 1, 0, 1, -2, -2, -4, -1, -2, -4, -4, -3, -3, -4, -1, -4, -4, -3, -2, -2, 0, -1, -4, 0, 1, 0, 0, 0, 4, 1, -1, 0, 3, 0, -2, 0, 0, -3, -4, -2, -2, -5, -6, -3, -4, -5, -4, -4, -4, -2, -3, -1, -1, -2, -4, 0, 1, 0, 0, 1, 4, 0, 0, 1, 3, -1, -2, -1, -1, -3, -5, -4, -2, -4, -5, -4, -2, -5, -5, -3, -5, -4, -4, -3, -1, -4, -3, 0, 0, -1, 0, 1, 5, 0, -1, 1, 1, -2, -4, -3, -1, -2, -3, -4, -3, -3, -3, -2, -2, -3, -4, -4, -6, -7, -4, -5, -4, -5, -3, -1, 0, 0, 0, 0, 3, 0, 0, 1, 1, -3, -5, -1, 0, -1, -3, -5, -3, -1, 0, -1, -3, -4, -6, -6, -5, -6, -5, -5, -4, -4, -3, 0, 0, 0, 0, 0, 3, 0, 0, 1, 0, -2, -3, 0, 0, -2, -3, -4, -2, 0, -1, -2, -3, -2, -6, -6, -7, -5, -4, -4, -4, -5, -2, -2, 0, 0, 0, -1, 4, 0, -1, 0, 0, -3, -3, 0, 0, -2, -4, -3, -1, 1, 0, -2, -2, -1, -3, -4, -4, -4, -4, -4, -6, -5, -2, 0, 0, 0, 1, 0, 3, 0, 1, 0, 0, -3, -3, 0, 0, -2, -2, -2, 0, 0, 0, -1, -2, -1, -1, -1, -1, -4, -4, -3, -3, -2, -1, 0, 0, 1, 2, 1, 3, 0, 1, 0, 0, -3, -4, -1, 0, -1, -2, -2, 0, 0, -1, 0, -2, -1, -1, 0, 0, -1, -2, -4, -2, -1, 0, 1, 1, 2, 2, 1, 3, 0, 0, 0, -1, -3, -4, -2, 0, -2, -4, -2, 0, 0, -1, 0, -1, -2, -2, 0, 0, 0, -1, -1, -1, 0, 1, 2, 2, 1, 2, 1, 1, 0, 0, 0, 0, -1, -2, -1, -2, -2, -3, -2, 0, 0, 0, 0, 0, -2, -1, 0, 1, -1, 0, -2, 0, -1, 1, 2, 1, 2, 1, 1, -1, 1, 0, 0, 0, -1, -1, -1, 0, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 3, 2, -2, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 2, 1, 2, 2, 1, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 2, 1, 1, 2, 3, 3, 2, 2, 1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 2, 1, 2, 1, 2, 1, 2, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 1, 0, -1, -1, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, -1, -2, 0, -1, 0, 0, 0, 1, 0, 0, 0, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -2, -1, -1, -2, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -2, -1, -1, 0, -1, -1, -2, -2, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, -1, -2, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -2, -2, -2, -2, -2, -2, -2, -1, -1, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, -1, -2, -1, -2, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -2, -2, -1, -1, -2, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, -1, 0, -2, -2, -1, -2, -3, -2, -3, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, 0, -2, -2, -2, -2, -1, -2, -1, -2, -2, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 0, -1, -1, 0, 0, -2, -1, -2, -1, -1, -2, -1, -2, -1, -1, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 1, 2, 0, 2, 0, 0, 0, -1, 0, 0, -1, -2, -3, -1, -1, -2, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 2, 1, -1, 0, 0, -1, 0, -2, -1, -2, -2, -2, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, -2, -1, -2, -2, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, -1, -1, -2, -1, -2, -1, -1, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -2, 0, 0, -1, 0, -2, -2, -1, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 2, 1, 1, 1, 1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 1, 2, 1, 1, 1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 2, 2, 1, 2, 2, 1, 1, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 2, 1, 3, 2, 2, 2, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 1, 3, 3, 3, 2, 2, 2, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 1, 1, 2, 1, 1, 1, 2, 1, 0, 0, 0, 0, 2, 1, 1, 2, 1, 1, 1, 1, 3, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 1, 2, 2, 0, -1, 0, 0, 0, 0, 2, 1, 1, 1, 1, 1, 2, 2, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 3, 2, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, -1, -1, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, -1, -1, -2, -1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, 1, 0, 1, 1, 0, 0, -1, -1, -1, -2, 0, 0, -1, 0, 0, 0, -3, -2, -2, -3, -1, -2, -2, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 2, 2, 0, -1, -1, -1, -2, 0, -1, 0, -1, 0, -2, -1, -1, -1, -3, -3, -2, -2, -3, -2, -1, 0, 0, 0, 0, -2, 0, 0, -1, 0, 1, 2, 0, 0, 0, 0, -1, -1, -1, -2, -1, -2, -1, -1, -1, -2, -3, -2, -3, -3, -3, -1, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, -2, 0, -1, -2, -1, -1, -2, -2, -1, -2, -2, -3, -1, 0, 0, 0, 1, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, -2, -2, -2, -1, -3, -3, -2, -2, -2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, -2, -3, -1, -2, -2, -2, -3, -2, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, -1, -1, -1, -1, 0, 0, -1, -1, -2, -1, -1, -1, -3, -1, -2, -3, -2, -2, -3, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, -3, -2, -2, -3, -2, -3, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, -1, 0, 0, 0, -1, -2, -1, -1, -2, -1, -2, -3, -2, -1, -2, -3, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 0, -1, -1, 0, 0, 0, -2, -2, -2, -1, -2, -2, -2, -3, -2, -1, -3, -2, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 2, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, -2, -1, -2, -2, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, -1, -1, 0, 0, 0, 0, 0, -2, -1, -1, 0, -2, -1, -2, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, -2, -1, -2, -2, -2, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, -1, -1, -2, -2, -2, -1, -2, -2, -2, 0, -2, -1, -1, -2, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, -2, -2, -1, 0, -2, -1, 0, -1, -1, -2, -2, -2, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -2, -2, -2, -1, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -2, -2, -2, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -2, -3, -3, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -2, -2, -1, -1, -1, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, -1, -2, -1, -2, -2, 0, 1, 0, 1, 1, 0, 0, 1, 0, 1, 1, 2, 2, 0, 1, 0, 1, 0, 0, 0, 2, 1, 1, 1, 1, 2, -1, 0, -1, -1, 0, -2, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 2, 1, 2, 2, 1, 0, 1, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 2, 2, 2, 2, 1, 0, 1, 0, 1, 1, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 1, 2, 1, 1, 3, 2, 2, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -2, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 2, 2, 1, 3, 1, 2, 2, 1, 0, 1, 0, 0, 0, -1, 0, 0, -1, -2, -1, -1, -1, -2, -1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 1, 2, 3, 3, 1, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 0, 2, 0, 0, 1, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 2, 1, 2, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 2, 2, 3, 3, 2, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, -2, -2, -1, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -2, -2, -1, -2, -2, -3, -1, -1, -2, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, -2, -1, -2, -1, -3, -4, -4, -2, -3, -1, -2, 0, 0, -1, -1, 0, -1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, 0, -2, -2, -4, -4, -3, -4, -3, -3, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -2, -3, -5, -4, -4, -4, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -3, -3, -5, -5, -5, -4, -4, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -5, -5, -6, -5, -3, -3, -2, -3, -2, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 2, 1, 0, 0, 2, 0, -1, 0, 0, -2, -5, -6, -5, -3, -3, -2, -3, -2, -2, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 2, 2, 2, 1, 2, 0, 0, 0, -1, -2, -3, -4, -4, -4, -4, -4, -2, -2, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 2, 2, 1, 2, 2, 2, 1, 0, 1, 0, 0, 0, -1, -2, -2, -3, -4, -3, -4, -3, -3, -1, -1, 0, 0, 0, 0, 0, -2, 0, 0, 0, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -3, -2, -3, -2, -2, -1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, -2, -2, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, -1, -2, -1, -3, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -2, -2, -1, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, 0, 0, 1, 1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 2, 1, 1, 1, 0, 2, 0, 0, 0, -1, -1, 0, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -2, -1, 0, 0, 0, 1, 2, 1, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, 0, 0, -1, 0, 1, 1, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -3, -2, -4, -3, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -2, -2, -3, -2, -4, -4, -4, -4, -2, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, -2, -3, -2, -3, -1, -3, -2, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 1, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, -2, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, 0, -2, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -2, -2, 0, 0, -2, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, 0, 0, -1, -1, -2, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, -1, -1, -1, -1, -2, 0, -1, 0, -1, -1, 0, -1, -2, -1, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -2, -2, 0, 0, 0, -1, 0, 0, -2, -1, -1, -1, 1, 0, -1, -1, -1, -1, -1, -1, -1, 0, -1, -1, -1, 0, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, 1, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, -1, 0, 0, -1, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, -1, 0, -1, 0, 0, 0, -2, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -2, 0, -1, -2, -1, -1, -1, 0, -1, 0, -2, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -2, -2, -1, -2, 0, -1, -1, 0, -1, 0, -1, -2, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -2, -1, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, -2, -1, 0, 0, -1, -1, -1, -1, -1, 0, -1, -1, -2, -1, -1, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, 0, 0, -2, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -2, 0, -1, -1, -2, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, -1, 1, 1, 0, 1, 1, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, 0, -1, -2, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -2, -1, -1, -1, -1, -1, -2, -1, -2, -1, 0, 0, 0, 0, -1, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, -1, -1, -2, -1, -2, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, 0, -1, -1, -2, -1, -1, -2, -2, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, -1, -3, -3, -1, -1, -2, 0, -2, -2, -2, -2, -2, -1, 0, 0, 0, 1, 0, 0, 2, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -1, -2, -2, -3, -1, -1, 0, -2, -2, -2, -1, -2, -1, -1, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, -3, -3, -2, -2, -2, 0, 0, -1, -3, -3, -3, -2, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -2, -3, -3, -3, -3, -1, -1, -1, -3, -3, -3, -1, -2, -1, -1, -1, -1, -1, -1, 0, 1, 3, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -3, -2, -2, -2, -1, -2, 0, -1, -2, -2, -2, -1, 0, -2, -2, -2, 0, 0, 0, 0, 1, 3, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -2, -1, -2, -3, -2, -2, -2, -2, -2, -2, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 2, 3, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, -2, -2, -2, -2, 0, -1, -2, -2, -2, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 2, 3, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -2, -2, 0, -1, -1, -2, -2, -3, -2, 0, -1, -1, -1, 0, -1, 0, 0, 1, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -1, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, -2, -1, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 1, 3, 0, 0, 1, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -2, -1, 0, 0, 0, -2, -3, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -2, -1, -1, -2, -3, -1, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 1, 2, -1, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -2, -1, -2, -1, 0, -3, -2, -1, -2, -1, 0, -2, -2, -2, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, -2, -2, -2, -3, -3, -2, -1, -1, 0, -2, -2, -2, 0, 0, 0, 0, 1, 2, 0, 0, 3, 0, -1, 0, 0, 0, -2, 0, -1, -1, -1, -1, -2, -2, -2, -2, -1, -2, -2, -2, -1, -1, -1, -2, -1, 0, 0, 0, 2, 2, 0, 0, 1, -1, 0, 0, 1, 1, -1, -1, -1, -1, -2, -1, -2, -1, -2, -1, -1, 0, -2, -3, -2, -1, -1, -1, 0, 0, 0, 0, 2, 2, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, 0, -1, -1, -1, -2, -3, -1, -2, -1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 3, 0, 0, 0, -1, 0, 0, 0, -2, -1, -1, -1, -2, -1, -1, 0, -1, -1, -2, -2, -1, 0, -2, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -2, -1, 0, 0, 0, 0, -1, -1, -1, -2, -2, 0, 0, 0, 0, 1, 2, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -2, -1, 0, -1, -2, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, -2, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 1, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, -2, -1, -2, -1, -1, 0, -1, -1, 0, 0, 0, 2, 1, 0, 1, 0, 1, 0, 2, 1, 2, 2, 1, 0, 0, 1, 1, 1, 1, 1, 0, -1, -1, -1, -1, -1, -2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 2, 1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, -1, 0, 1, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 1, 1, 0, -1, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, 0, -1, -2, -1, -1, -1, -1, -2, 0, 0, 0, 0, -1, 0, 0, 3, 1, 1, 1, 1, 0, -1, 0, 0, 0, -2, -1, 0, 0, 0, -1, -1, -2, -1, -1, -1, -1, -1, 0, -1, -2, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 1, 1, 0, 0, 0, 0, -3, -1, -1, -1, -1, -2, -2, -1, -2, -1, -1, -2, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, 2, 3, 1, 2, 1, 0, 0, 1, 2, 1, -1, -1, 0, 0, -2, -1, -2, -2, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 0, 0, 0, 2, 0, 0, -1, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 2, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, -1, -1, -1, -1, -1, 0, -2, -2, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -1, -2, -2, -2, -3, -3, -3, -1, -1, -2, -1, 0, 0, -1, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -4, -2, -3, -3, -1, -2, -3, -2, -2, -3, -2, -1, 0, 0, 0, -1, 0, 1, 1, 3, 3, 2, 0, -1, 0, 0, 1, 0, 0, 0, -1, -3, -4, -3, -4, -4, -2, -4, -2, -3, -2, -2, -2, -2, 0, -1, -1, 0, 1, 3, 2, 3, 4, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -4, -3, -3, -2, -3, -3, -3, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 3, 3, 4, 1, 0, 1, 0, 2, 3, 2, 1, 0, 0, -3, -3, -2, -1, -1, -1, -3, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 3, 3, 2, -1, 1, 1, 1, 3, 2, 0, 0, -1, -1, -1, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 2, 2, 1, 0, 1, 3, 2, 2, 2, 0, 1, 0, 0, 0, 0, -1, 0, 0, -2, -2, -1, -2, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 3, 0, 0, 1, 3, 3, 2, 0, 1, 0, 0, 0, 0, -2, -1, 0, -2, -2, -3, -2, 0, -1, -1, -2, 0, 1, 0, 1, 1, 1, 0, 1, 1, 1, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, -1, -3, -2, -1, -3, -3, -1, -3, -1, -1, -2, -1, 0, 0, 0, 2, 2, 1, 1, 1, 2, 1, 0, 4, 3, 2, 0, 0, 0, 0, 0, -1, -1, -3, -2, -1, -2, -2, -3, -3, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 2, 4, 1, 1, 0, 0, 0, 0, -1, -1, -2, -2, -2, -3, -1, -2, -3, -2, -2, -2, -1, -1, -2, -1, 0, 0, 0, -1, 1, 2, 1, 0, 4, 4, 2, 3, 2, 2, 0, 0, 0, 0, -2, -2, -2, -2, -2, -2, -4, -3, -1, -1, -2, -3, -1, -1, 0, 0, -1, 0, 1, 1, 0, 1, 5, 4, 3, 3, 3, 2, 1, 1, 0, 0, 0, 0, 0, -1, -4, -4, -3, -2, -2, -2, -1, -2, -2, -3, -1, -1, 0, 0, 0, 1, 1, 1, 4, 5, 3, 4, 5, 3, 1, 2, 0, 0, 0, 0, 0, 0, -1, -3, -2, -2, -3, -2, -2, -2, -3, -2, -1, 0, 0, 0, 1, 2, 2, 1, 4, 4, 3, 3, 3, 2, 2, 1, 1, 1, 1, 1, 0, 0, 0, -1, -1, -2, -1, -1, -3, -4, -2, -2, 0, 0, 0, 0, 0, 0, 0, 2, 4, 4, 3, 4, 4, 2, 1, 2, 1, 0, 1, 0, -1, 1, 0, -2, -1, 0, -1, -1, -2, -2, -3, -2, 0, 0, 1, 0, 0, 0, 0, 1, 5, 5, 4, 4, 4, 2, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, -2, -1, 0, 0, 0, 1, 0, 0, 2, 4, 3, 1, 3, 2, 3, 2, 1, 0, 0, 0, -2, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 2, 3, 1, 1, 2, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 2, 2, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, -1, -1, -2, -3, 0, 0, 2, 1, 0, 0, 1, 1, 2, 1, 0, 1, 2, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, -2, -2, -1, 0, 0, -1, -1, -3, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 1, 0, -1, 0, -1, -2, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -2, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, -2, -3, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, -1, -1, -2, -3, -3, -2, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 3, 1, 2, 2, 0, 1, 0, 0, 0, 0, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 2, 1, 1, 2, 2, 2, 2, 1, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 2, 2, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 2, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 2, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, -2, -1, -2, -2, -1, 0, 3, 1, 1, 1, 0, 3, 2, 1, 0, 2, 1, 0, -1, 0, 0, 1, 1, 1, 0, 1, 0, 1, 2, 2, 1, 2, 2, 2, 0, 0, 2, 0, 4, 1, 0, 0, 0, 2, 1, 1, 0, 0, -1, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 1, 0, -3, -1, 1, 2, 3, 2, 1, 0, 0, 2, 0, 0, 0, 0, 0, -2, -2, 0, 1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -5, -5, 0, 1, 4, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 5, 3, 0, -1, -1, 0, -1, 0, 0, -1, 0, 1, 0, -1, -5, -5, -1, 1, 4, 2, 0, 1, 0, -1, -1, -2, 0, -1, 0, 1, 1, 4, 4, 3, 1, 0, -2, -1, -1, -1, -1, -2, -3, 0, 0, 0, -3, -4, -1, 0, 3, 2, 0, 0, -1, -1, -2, -2, -2, -2, -1, 0, 0, 3, 3, 3, 0, 1, -1, 0, -1, -1, -1, -2, -3, -3, 0, -1, -2, -3, 0, 0, 4, 0, 0, -1, -2, -3, -2, -1, -1, -2, -3, -1, 0, 0, 1, 1, 2, 2, 0, 0, -3, -2, -1, -3, -4, -2, 0, 0, -2, -1, -1, 0, 4, 0, 0, 0, -2, -2, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 1, 0, 0, -2, -3, -1, 0, -1, -3, -2, 0, 0, 0, -2, -1, 0, 4, 1, 0, 0, 0, 0, 1, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 1, 0, -1, 0, 3, 2, -1, -1, 0, 3, 1, 1, 0, 0, 1, 2, 0, 1, 1, 0, 0, 0, 1, 1, 0, -2, -1, 0, 0, 1, 1, 3, 4, 1, 0, 0, 3, 3, 0, 0, 0, 3, 0, 1, 1, 0, 2, 3, 2, 1, 1, 1, 1, 1, 1, 0, -2, -2, -3, 0, 1, 2, 2, 5, 5, 4, 1, 2, 2, 2, 0, -2, -1, 3, 2, 1, 2, 1, 0, 4, 3, 2, 2, 1, 2, 2, 2, 2, 1, -2, -2, -1, 1, 1, 3, 5, 6, 6, 5, 3, 2, 2, -1, -1, 0, 1, 3, 2, 3, 3, 1, 3, 2, 2, 4, 3, 2, 2, 0, 1, 1, 0, -1, 0, 0, 1, 2, 5, 7, 7, 6, 3, 3, 1, 0, 0, 0, 2, 2, 2, 3, 2, 2, 3, 1, 2, 4, 5, 4, 2, 1, 0, 0, 1, 0, 0, 0, 0, 1, 3, 5, 5, 4, 3, 1, 0, 0, 0, 0, 4, 3, 3, 4, 2, 1, 1, 1, 3, 5, 4, 4, 1, -1, -1, 0, 1, 1, 2, 1, 0, 1, 3, 4, 3, 1, 1, -1, 0, 0, 0, 0, 4, 3, 3, 4, 2, 0, 0, 1, 2, 3, 4, 4, 2, 0, -2, -1, 0, 0, 2, 1, 0, 0, 3, 2, 3, 0, 0, -1, -1, 0, 0, 0, 6, 2, 2, 4, 2, 2, 1, 2, 2, 2, 2, 1, 1, 1, -2, -2, -2, -1, 0, 0, 0, 3, 3, 2, 1, 1, 0, -2, -2, 0, -1, -1, 4, 2, 0, 3, 1, 1, 0, 4, 5, 4, 3, 3, 1, 2, 0, -2, -3, -3, -2, -1, 0, 3, 4, 3, 2, 3, 1, -1, -1, -1, 0, 0, 4, 1, 0, 2, 1, 0, 0, 1, 5, 2, 2, 2, 0, 3, 0, -1, -2, -3, -1, 0, 0, 1, 4, 3, 4, 3, 1, -2, 0, 0, -1, 0, 6, 2, 0, 3, 1, 0, -1, 0, 2, 1, 0, 1, 1, 1, 0, -1, -3, -2, 0, 2, 0, 1, 1, 4, 5, 3, 1, -1, 0, 1, -1, 0, 5, 4, 1, 1, 1, 0, -1, -2, 0, 0, 1, 0, 1, 0, 0, -1, -2, -1, 0, 2, 2, 0, 0, 2, 4, 5, 1, -1, 0, 0, 0, 0, 5, 5, 1, 2, 1, 0, 0, 0, 0, 0, 1, 3, 0, 0, -1, -2, 0, 0, 0, 1, 1, 0, 0, 1, 5, 5, 1, 0, 0, 0, 0, 1, 7, 4, 0, 1, 1, 2, 0, 0, 1, 1, 3, 3, 1, 1, 0, 0, 0, 0, 1, 2, 3, 1, 0, 2, 4, 3, 0, 0, 0, 0, 0, 0, 7, 4, 0, 1, 1, 1, 0, -1, 0, 2, 4, 4, 2, 1, 0, 1, 2, 0, 0, 1, 2, 0, 0, 2, 3, 4, 1, -1, 0, 0, 1, 1, 7, 4, -1, 0, 0, 0, -1, 0, 0, 3, 4, 3, 0, 0, 1, 3, 2, 1, -2, 0, 0, 1, 0, 2, 1, 2, 0, -2, -1, 0, 1, 0, 8, 4, -1, 0, 0, -1, -3, -2, -1, 1, 2, 1, 0, 0, 1, 2, 3, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 1, 1, 1, 6, 4, -1, 0, 0, -2, -3, -3, 0, 1, 0, 0, 1, 1, 1, 1, 1, 2, 2, 4, 2, 0, 0, 1, 1, 0, 0, -1, -1, 0, 2, 1, 7, 5, 0, 0, -1, -3, -4, -2, 0, 0, 0, 0, 0, 2, 1, 0, 1, 2, 3, 6, 4, 3, 1, 1, 0, 0, 1, 2, 0, 0, 2, 1, 4, 4, 1, 0, -2, -1, -2, -2, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 4, 5, 5, 3, 3, 3, 2, 2, 2, 2, 0, 1, 2, 2, 5, 4, 0, -1, -3, -2, -3, -3, -1, 0, 0, -1, 0, 0, 0, -2, -2, -1, 0, 3, 4, 3, 2, 2, 2, 2, 3, 2, -1, 0, 4, 3, 4, 3, 0, -1, -2, -3, -2, -2, -1, 1, -1, -1, -1, -1, -1, -2, -2, -3, 0, 0, 1, 1, -1, 0, 1, 1, 2, 0, -1, -1, 1, 2, 2, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -2, 0, 0, 0, -1, -2, -1, -1, 0, -1, -1, -2, -2, 0, 2, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 3, 1, 1, 1, 1, 2, 1, 1, 0, 1, 2, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 2, 4, 3, 3, 4, 2, 2, 3, 2, 1, 3, 2, 1, 1, 2, 2, 1, 2, 2, 2, 1, 1, 1, 0, 0, -2, 0, -1, 0, 0, 1, 1, 3, 3, 5, 5, 5, 3, 2, 1, 2, 1, 1, 1, 1, 0, 0, 0, 2, 1, 1, 2, 2, 0, 1, 1, 0, -2, 0, 0, 1, 2, 2, 0, 2, 2, 4, 3, 4, 3, 2, 2, 0, 1, 0, 0, 1, 1, 2, 3, 3, 0, 1, 1, 2, 2, 1, 0, 0, 0, 0, 1, 1, 2, 1, 2, 0, 1, 3, 3, 3, 3, 2, 0, -1, -1, -2, 0, 0, 1, 2, 2, 3, 2, 1, 2, 1, 2, 2, 1, 0, -1, 0, 0, 0, 2, 1, 2, 1, 2, 3, 2, 0, 1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 3, 2, 2, 0, 1, 2, 2, 2, 1, -1, 0, 0, -1, 0, 1, 3, 3, 3, 4, 2, 0, -1, 0, 0, -2, -3, -2, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 2, 1, 2, -1, 0, 0, 0, 0, 2, 3, 4, 4, 4, 3, 1, 0, -1, -3, -4, -2, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 2, 2, -1, -2, -1, -1, 0, 0, 1, 4, 4, 2, 3, 0, -1, -2, -2, -2, -2, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 2, 4, -1, -2, -2, -1, -1, 0, 0, 0, 2, 1, 1, 0, 0, -2, -2, -2, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 2, 5, 3, -1, -3, -3, -2, -1, -2, -2, -2, -1, 0, 0, 0, -1, -3, -2, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 1, 3, 4, 4, -2, -3, -3, -2, -3, -3, -5, -4, -2, -2, -2, -1, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 2, 3, 4, -1, -2, -3, -3, -3, -5, -6, -6, -5, -3, -3, -3, -1, -1, -1, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 2, 2, 2, 0, -3, -3, -4, -2, -5, -5, -6, -6, -5, -4, -1, 0, 1, 0, 1, 2, 2, 1, 2, 2, 3, 2, 2, 0, 0, 0, 0, 1, 0, 1, 2, -2, -3, -3, -1, -2, -3, -5, -6, -4, -4, -4, -1, 0, 1, 2, 2, 3, 3, 3, 1, 3, 2, 4, 2, 1, 1, 0, 0, 0, 0, 1, 2, -1, -2, -2, -1, -2, -4, -6, -5, -5, -4, -3, -2, 0, 2, 2, 3, 3, 3, 2, 2, 2, 3, 3, 3, 2, 0, 0, 0, 0, 1, 2, 2, 0, -1, -1, -2, -3, -3, -5, -5, -4, -3, -2, 0, 0, 1, 2, 1, 2, 4, 2, 2, 2, 3, 2, 1, 1, 0, 0, 0, 2, 3, 3, 2, -1, -2, 0, -1, -4, -3, -5, -4, -3, -4, -2, 0, 1, 1, 1, 1, 0, 1, 1, 2, 2, 3, 2, 2, 2, 2, 1, 2, 3, 3, 3, 3, 0, -1, 0, -1, -4, -4, -4, -5, -3, -1, -1, -1, 1, 1, 1, 0, 0, 0, 1, 1, 1, 1, 1, 3, 3, 2, 3, 2, 3, 2, 3, 2, -1, -1, 0, -1, -2, -3, -4, -4, -2, -2, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 1, 1, 1, 1, 2, 1, -2, -1, 0, -1, -3, -4, -4, -4, -4, -2, -3, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 1, -1, 0, -1, -2, -3, -3, -3, -4, -3, -3, -2, -1, 0, 0, 1, 0, -1, -1, -2, -2, -1, -1, -1, -2, -1, 0, 0, 0, -1, -1, -1, 1, -2, 0, -1, 0, -3, -2, -1, -1, -1, -2, -1, -1, 0, 0, 0, 0, -2, -4, -2, -2, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, 0, -1, -1, 0, -1, -2, -2, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, -3, -3, -3, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 1, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, -1, -3, -5, -3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, -3, -3, -2, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 1, 3, 1, 2, 2, 2, 1, 0, 0, 0, -1, -2, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, -1, -1, 0, 0, 0, 2, 3, 3, 2, 3, 2, 2, 3, 2, 2, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 2, 2, 3, 4, 3, 3, 3, 3, 3, 3, 3, 2, 3, 2, 2, 0, 0, 1, 1, 1, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 2, 3, 2, 4, 4, 1, 3, 1, 1, 3, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, -1, 0, 1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 2, 2, 1, 2, 1, 2, 1, 1, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 3, 4, 3, 2, 2, 1, 0, 0, 2, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 2, 3, 2, 2, 2, 2, 3, 2, 1, 1, 2, 1, 1, 1, 2, 2, 2, 2, 3, 2, 2, 1, 2, 1, 0, -2, -2, 0, 1, 0, 0, 0, 1, 3, 4, 4, 3, 1, 3, 1, 1, 0, 1, 0, 0, 1, 1, 1, 1, 1, 0, 1, 2, 1, 1, 0, -1, -2, 0, 0, 1, 1, 0, 0, 0, 2, 3, 3, 3, 2, 2, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 2, 1, 1, 3, 2, 1, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 2, 2, 0, 0, -1, 0, 0, 0, 0, 1, 2, 2, 2, 0, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 2, 1, 2, 1, 0, 1, 0, 1, 1, 1, -1, 0, 0, -1, 0, 1, 2, 2, 2, 3, 1, 0, 0, -1, -1, -2, -2, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 1, 1, 2, 0, -1, -2, -1, 0, 1, 1, 3, 3, 2, 0, 0, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 1, -1, -2, -2, -2, 0, 0, 0, 0, 3, 0, 0, 0, -2, -3, -2, -2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 4, 1, -1, -1, -1, -2, -1, 0, -1, 0, 0, 1, 0, -1, -2, -1, -3, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 2, 4, 2, -1, -2, -3, -2, -2, -3, -2, -1, -1, -1, -1, 0, -2, -3, -3, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 3, 2, -2, -3, -2, -1, -2, -3, -4, -2, -2, -2, -2, 0, -1, -2, -1, -2, 0, 0, 1, 1, 0, 0, 0, 1, -1, -1, 0, 1, 0, 0, 2, 2, -2, -1, -3, -2, -2, -3, -4, -2, -3, -3, -2, 0, -1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, -1, -2, -2, -1, -2, -2, -4, -2, -2, -3, -2, -2, 0, 1, 0, 2, 1, 2, 1, 1, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 1, 0, -2, -2, 0, 0, -1, -2, -4, -2, -3, -2, -3, -2, -1, 0, 0, 1, 3, 2, 1, 2, 2, 3, 1, 1, 0, 0, -1, 0, 0, 1, 1, 1, -1, -1, -1, -1, -1, -3, -3, -4, -2, -1, -2, -2, 0, 1, 1, 2, 2, 2, 2, 1, 1, 3, 1, 1, 1, -1, -2, 0, 0, 0, 2, 2, -2, 0, 0, -1, -2, -3, -3, -2, -3, -3, -3, -1, 0, 0, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 2, 2, 3, 0, -1, -1, 0, 0, -1, -2, -2, -3, -3, -2, -2, -1, -1, 0, 1, 0, 0, 0, 1, 0, 1, 1, 2, 2, 1, 1, 0, 2, 2, 1, 2, 1, -1, 0, 0, 0, -2, -3, -2, -2, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 2, 1, 2, 1, 0, 1, 1, 0, -2, 0, 0, -1, -2, -2, -3, -3, -3, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -2, -2, -2, -2, -3, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -2, -2, -3, -3, -2, -2, -1, -2, -1, 0, 0, 0, -2, -1, -2, -1, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, -1, -3, -4, -2, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 0, -1, 0, -1, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -1, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -2, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, -2, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, -2, 0, 0, 0, 0, 1, 2, 0, 0, 2, 2, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, -1, -1, 0, -1, 1, 0, 2, 3, 2, 3, 2, 3, 1, 2, 3, 1, 2, 0, 1, 1, 0, 1, 2, 0, 0, 0, 0, 2, 0, 2, 1, 1, 0, 0, 0, 0, 1, 1, 1, 2, 3, 2, 2, 2, 2, 2, 2, 1, 2, 1, 1, 0, 1, 2, 1, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 2, 1, 1, 1, 1, 2, 1, 2, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 2, 1, 2, 1, 2, 1, 1, 2, 1, 0, 1, 1, 2, 2, 1, 2, 1, 1, 3, 3, 3, 2, 2, 2, 1, 1, 0, 2, 1, 1, 1, 2, 0, 1, 0, 0, 1, 1, 2, 1, 2, 2, 1, 1, 1, 2, 0, 0, 1, 3, 2, 2, 2, 1, 2, 3, 2, 1, 1, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 3, 2, 3, 1, 0, 0, 1, 0, 0, 2, 2, 1, 2, 3, 1, 1, 1, 2, 2, 2, 2, 1, 1, 0, 1, 1, 1, 0, 0, 1, 0, 1, 1, 1, 3, 3, 0, 0, 0, 0, 1, 1, 1, 0, 1, 2, 0, 1, 2, 2, 1, 0, 2, 2, 0, 1, 0, 0, 0, 2, 0, 0, 0, 1, 1, 0, 2, 1, 0, 0, 0, 1, 1, 2, 1, 1, 1, 1, 1, 2, 0, 0, 2, 1, 2, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 2, 1, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 2, 1, 1, 0, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, -1, 0, 1, 1, 0, 2, 2, 1, 1, 0, 0, 1, 1, 0, 1, 2, 2, 2, 0, 1, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 0, 0, 1, 2, 1, 0, 0, 2, 2, 1, 2, 3, 1, 2, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 1, 2, 2, 1, 0, 0, 1, 2, 1, 2, 1, 1, 2, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 2, 2, 1, 0, 1, 1, 1, 0, 1, 2, 1, 1, 1, 1, 0, 0, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 2, 1, 2, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, -1, -1, 0, -1, -1, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 2, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, -2, -1, -1, -1, 0, 0, 0, -1, -1, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, -1, 0, 0, 1, 1, 1, 1, 2, 2, 0, 0, 1, 1, 3, 2, 0, 1, 0, 1, 0, 0, 1, 1, -1, 0, -2, -1, -1, 0, -1, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 3, 0, 1, 3, 3, 3, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 3, 3, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 0, 2, 1, 2, 1, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 1, 1, 0, 2, 2, 1, 0, 0, 0, 0, 1, 0, 0, -2, -2, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 2, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, -2, 0, -1, 0, 0, -1, 0, 2, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 2, 2, 1, 2, 2, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 0, 2, 1, 1, 1, 1, 0, 1, 0, 1, 1, 2, 1, 2, 2, 2, 1, 1, 0, 0, 0, -1, 0, 1, 2, 0, 0, 1, 1, 2, 2, 1, 1, 1, 2, 1, 2, 2, 1, 0, 2, 2, 0, 2, 3, 1, 2, 2, 1, 1, 1, 1, 1, 0, 0, 0, 1, 2, 1, 1, 2, 1, 2, 1, 3, 2, 1, 2, 2, 2, 1, 1, 1, 2, 1, 3, 2, 3, 3, 2, 1, 0, 1, 1, 0, 0, 0, 0, 2, 1, 0, 1, 0, 2, 2, 2, 3, 3, 2, 2, 2, 3, 3, 1, 1, 2, 1, 2, 3, 4, 4, 3, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 2, 2, 2, 3, 2, 1, 2, 3, 2, 3, 2, 2, 3, 2, 3, 2, 2, 1, 0, 1, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 2, 1, 2, 0, 1, 2, 1, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 2, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 0, 2, 0, 0, 1, 1, -1, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 2, 0, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 0, 1, 1, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 2, 2, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 2, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 2, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 2, 1, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -1, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 2, 1, 1, 1, 1, 0, 0, -1, -2, -2, -1, -1, -2, 0, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 2, 1, 2, 0, 0, 2, 0, 0, 0, 1, 1, 1, 0, 0, -1, -1, -1, -1, -2, -1, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -2, -1, 0, 0, 0, -1, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, -2, -2, -2, -2, 0, -1, -1, 0, -3, -3, -1, 0, -1, 0, 0, 1, 0, 0, 1, 2, 1, 1, 0, 0, -1, 0, 1, 0, 0, 1, 1, 0, -2, -1, -2, -1, 0, 0, -1, -1, -1, -2, 0, -1, 0, 0, 0, 1, 2, 0, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, -2, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, -1, -1, -2, 0, -1, -1, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, -2, 0, 0, 0, 0, -2, 1, 1, 0, -1, -1, 0, 0, -1, -1, -1, 0, 1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 2, 1, 0, 1, 0, -1, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, -1, 1, 1, 1, 1, 2, 0, 0, 1, 1, 0, 2, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, -2, 0, 0, 0, 0, -1, 0, 0, -1, -2, -2, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 3, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -2, -1, -1, 0, -1, 0, -1, -1, -1, 0, -1, -2, -1, 0, 0, 0, 0, 1, 1, 0, 4, 1, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, -1, -3, -1, 0, -1, -1, 0, 0, 0, -1, 1, 2, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -2, -1, 0, -1, 0, -1, 0, -1, 0, 1, 1, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, -2, -1, -2, -2, -1, -1, 0, 0, 0, 0, 2, 1, 0, 3, 1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -2, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, 2, 1, 2, 2, 2, 1, 0, 2, 2, 2, 1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 2, 2, 1, 1, 1, 0, 0, -1, 0, 1, 1, 3, 2, 2, 1, 1, 1, 2, 2, 1, 2, 2, 1, 0, 1, 0, 0, 0, 0, 0, 2, 1, 1, 2, 1, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 1, 1, 0, 2, 2, 2, 1, 1, 0, 0, 0, -2, 0, 0, 0, 1, 1, 0, 1, 1, 4, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 2, 1, 1, 1, 0, -1, 0, -2, -2, -1, 0, 0, 0, 0, 1, 1, 4, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, -1, -1, 1, 1, 0, 1, -1, 1, 0, -2, -1, -1, -1, -1, -1, 0, 0, 2, 3, 0, 1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, -1, 0, 0, 0, 2, 0, 0, -2, 0, -2, -1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -2, -2, -1, -1, 0, 0, 0, -2, -3, -1, 0, 0, 0, 0, 2, 3, 0, 0, -1, -1, -1, -1, 1, 0, 0, 0, 1, 0, -2, -1, -2, -2, -1, -3, -1, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -3, -3, -1, -2, -4, -2, -1, 0, 0, 0, 0, 0, 0, -2, 0, -1, 1, 3, 0, 0, 0, 0, -1, -1, 1, 0, -2, -1, 0, 0, -1, -2, -2, -3, -1, -3, -4, -4, -3, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 2, 0, 0, 0, -1, -1, 0, 1, -1, -2, -1, 0, -1, 0, 0, -2, -2, -1, -2, -4, -3, -3, -2, 0, 0, 0, 0, 0, 0, -2, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -1, -2, -1, -2, -3, -3, -4, -3, -2, -2, 0, 1, 1, 0, -1, -2, -1, -1, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -2, -3, -2, -1, -3, -3, -5, -4, -4, -2, -2, -1, -1, 0, 1, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, -2, -2, -3, -2, -2, -3, -5, -5, -5, -5, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, -1, 0, 0, 1, 0, -1, -1, 0, -1, -3, -3, -3, -3, -5, -5, -4, -4, -4, -3, -1, -2, 0, 0, -1, 0, 0, 0, 0, 2, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -3, -2, -3, -4, -4, -3, -4, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 3, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -3, -2, -3, -1, -4, -4, -4, -3, -4, -2, -3, -2, 0, 0, -1, 0, 0, 0, 0, 2, 0, 0, -1, 0, 2, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -1, -3, -4, -3, -2, -4, -2, -2, -1, 0, -2, -2, 0, 0, 0, 0, 2, 1, 1, -1, 0, 2, 1, 2, -1, 0, 0, 0, -1, -1, -2, -2, -3, -2, -3, -2, -2, -3, -2, -2, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 0, -2, -1, -1, -2, -3, -3, -2, -3, -2, -2, -2, -1, -1, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, -1, -1, -1, -2, -3, -2, -3, -4, -2, -2, -2, -2, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -2, -2, -2, -2, -3, -2, -2, -2, -4, -3, -3, -2, -2, -1, 0, 0, -1, -1, 0, 0, 0, -1, 1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, -1, -2, 0, 0, -2, -2, -2, -2, -3, -2, -2, -1, -2, -1, -2, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -2, -2, 0, 0, 0, -2, -1, -2, 0, 0, 0, 0, -2, -3, -3, -3, -2, -2, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -3, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -3, -2, -3, -1, -1, -1, -2, -3, 0, 0, 0, 0, 0, 1, 0, 0, -2, -1, -1, -2, 0, -1, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, -1, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, -2, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 2, 0, 0, 0, 0, -1, -2, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 2, 0, 2, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 2, 1, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 2, 1, 1, 0, 1, 0, 0, -1, -1, -1, -1, -2, -2, -1, -2, -1, -1, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, -1, -2, -1, 0, 1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, -1, -2, -2, -2, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, 0, -1, -1, -2, -2, -1, 0, 0, 2, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -2, -1, -2, -2, -1, 0, -1, -1, -1, 0, 0, 2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, -1, -2, 0, 1, 1, 0, 0, -1, -1, -2, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 2, 2, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -2, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 1, 2, 2, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 2, 0, 2, 0, 0, 0, 0, 1, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 1, 2, 0, 0, 0, 0, 0, 1, 0, 2, 1, 2, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, -1, 0, 0, 0, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, -1, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 2, 1, 1, 1, 1, 1, 2, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, 1, 3, 3, 2, 2, 2, 2, 2, 1, 2, 2, 2, 1, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 3, 2, 2, 2, 2, 1, 2, 1, 2, 2, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 3, 3, 3, 2, 3, 2, 2, 1, 2, 2, 3, 3, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 4, 3, 1, 2, 1, 3, 0, 2, 1, 2, 2, 2, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 3, 3, 3, 2, 1, 1, 0, 1, 2, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, 0, 0, 2, 3, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 3, 2, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -2, -2, 0, 0, 2, 2, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -3, -2, -2, -1, 0, 2, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -2, -2, -2, -1, -1, -1, 0, -1, -1, -1, -1, -1, -2, -2, -2, -3, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -2, -1, -1, -1, 0, -2, -2, -2, -1, -1, -2, -2, -2, -3, -2, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 0, 1, 1, 1, 1, 0, 0, 1, 1, 0, 0, -2, 0, 0, -1, 0, -1, -1, -2, -1, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -2, -1, -3, -3, -3, -2, -3, -2, -1, 0, 0, 1, 1, 1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, -2, -1, -3, -3, -3, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, -1, 0, -2, -2, -2, -2, -1, -3, -2, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, -2, -2, -2, -2, -1, 0, 0, 0, 1, 0, 0, -1, -2, -2, -1, -1, -1, -2, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -2, -1, -1, 0, 0, 1, 1, 1, 0, 0, -2, -1, -1, 0, -1, -2, -2, 0, 1, 1, 0, 0, 0, 0, 0, 1, 2, 0, 0, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, -1, -2, 0, -1, -2, -2, -1, -1, -1, -2, 0, 1, 2, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, -2, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, -2, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, -1, -3, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -4, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -2, -3, -2, -1, -2, -1, 0, 0, 1, 1, 0, 0, -1, -3, -2, -3, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -2, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -3, -3, -4, -3, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 1, 1, 0, 0, -1, 0, 0, -1, -1, -2, -1, -4, -4, -3, -2, -1, 0, 1, 2, 1, 2, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, -4, -3, -2, -1, 0, 0, 3, 3, 3, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, -1, 0, 0, 1, 1, 0, -2, -3, -3, -4, -2, 0, 0, 1, 3, 2, 2, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 1, 1, 1, 0, 0, 0, 0, 2, 1, 0, 0, -2, -3, -2, -2, 0, 0, 3, 2, 1, 0, 1, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 1, 0, -2, -3, -4, -3, -3, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, 0, 0, 1, 1, 2, 2, 1, 1, 0, -1, 2, 1, -1, -1, -2, -4, -2, -2, 0, 0, 0, 1, 1, 0, -1, 0, 1, 1, 0, -1, -2, 0, 1, 1, 1, 1, 2, 2, 0, 0, 0, -1, 2, 2, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -1, -2, 0, 1, 3, 1, 0, 2, 0, -1, -1, -1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, 0, 1, 1, 0, 1, 0, -1, -1, 0, 0, 0, 2, 1, 1, 0, 0, 1, 2, 1, 1, 1, 1, 2, 2, 2, 1, 0, -2, -3, -2, 0, 0, 0, 1, 0, -1, -1, -1, -1, -2, -1, 0, -1, 1, 1, 0, 0, 1, 2, 3, 1, 1, 1, 2, 3, 4, 2, 1, 0, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 3, 2, 2, 1, 2, 4, 2, 1, 1, 1, 1, 4, 4, 3, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 2, 1, 1, 3, 4, 4, 1, 2, 2, 1, 3, 1, 0, -1, -1, -1, 1, 0, -1, -1, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 2, 3, 2, 1, 4, 4, 3, 1, 1, 1, 2, 2, 0, -2, -2, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 3, 4, 2, 3, 3, 4, 2, 2, 2, 1, 1, 0, -1, -1, -2, -2, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, -1, -1, -1, 0, -1, 0, 2, 3, 2, 2, 4, 3, 2, 2, 2, 2, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -2, -1, -1, -1, 0, 2, 2, 1, 0, 1, 3, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -2, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, -1, 0, -2, -1, 0, 0, -1, 0, 0, -2, -3, -3, -3, -3, -3, -2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, -2, 0, -1, -2, -3, -2, -3, -3, -5, -5, -4, -5, -5, -3, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, -2, -2, -2, -1, -1, -2, -2, -3, -3, -4, -3, -3, -3, -2, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -2, -2, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 1, 3, 2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 2, 3, 2, 3, 2, 3, 2, 2, 3, 2, 1, 3, 2, 2, 1, 0, 1, 2, 3, 2, 0, 0, -2, 0, 0, -1, 0, 0, -1, -2, -1, -1, 0, 1, 0, 2, 3, 3, 2, 3, 2, 3, 2, 1, 1, 1, 0, 0, 0, 2, 3, 0, 0, -1, -2, -2, -1, -2, -2, -2, -2, -2, 0, 0, 1, 1, 1, 0, 2, 3, 2, 4, 4, 2, 2, 2, 2, 0, -2, -1, 0, 1, 3, 1, 0, -1, -1, -1, -2, -2, -2, -3, -2, -2, 0, 0, 3, 1, 1, 0, 0, 2, 1, 1, 1, 2, 1, 1, 1, -1, -2, -2, -1, 0, 2, 2, 0, -1, -1, -1, -2, -2, -2, -2, -1, 0, 1, 2, 2, 1, 0, 2, 1, 1, 1, 1, 1, 1, 0, 0, 2, 0, -1, -1, -1, 1, 2, 0, 0, -1, -3, -3, -4, -2, -3, -3, -3, -1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 0, 0, 2, 1, -1, 0, 0, 1, 2, 0, -1, -2, -3, -3, -2, -3, -1, -1, -1, 0, 1, 1, 2, 1, 1, 1, 2, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 2, 0, -1, -2, -4, -4, -3, -3, -1, 0, 0, 0, 0, 3, 2, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 1, 2, 0, -1, -2, -3, -3, -3, -1, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 1, 1, 0, 0, 1, 2, 0, 0, 1, 1, 2, 0, -1, 0, 1, 0, 0, -1, -3, -1, -1, 0, 0, 1, 0, 0, 1, 3, 3, 0, 0, 0, 1, 1, 0, 1, 1, 2, 1, 2, 2, 1, 3, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, 1, 2, 0, 2, 2, 2, 2, 1, 0, 0, 1, 3, 1, 3, 3, 1, 1, 2, 2, 3, 1, 0, 0, 0, 3, 0, 0, 0, -1, -1, 0, 2, 2, 1, 2, 2, 1, 2, 2, 1, 0, 2, 2, 2, 2, 3, 2, 2, 2, 3, 3, 3, 1, -1, -1, 0, 2, 0, 0, 0, 0, -1, 0, 0, 1, 2, 3, 3, 2, 2, 1, 1, 3, 1, 1, 3, 1, 1, 1, 1, 2, 1, 2, 1, 0, 0, -1, 0, 3, 1, 1, 1, 0, 0, 0, 0, 1, 4, 5, 3, 2, 0, 0, 1, 2, 2, 1, 1, 1, 0, 0, 2, 2, 1, 0, 0, -1, -2, -2, 0, 2, 1, 1, 0, 1, 0, 0, 1, 1, 2, 3, 3, 1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, -1, -1, 0, 3, 2, 1, 1, 0, 0, 0, 1, 0, 2, 3, 2, 1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, -2, -1, -2, -1, 0, 2, 0, 1, 1, 1, -1, 0, 1, 1, 2, 3, 2, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, -2, -2, -2, -2, 1, 3, 1, 0, 0, 0, 0, 0, 1, 2, 2, 3, 2, 3, 2, 0, 0, -1, -2, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, -1, -2, -1, 1, 3, 2, 1, 1, 0, 0, 0, 1, 2, 0, 2, 1, 1, 1, 1, 0, -1, -1, -1, 0, 0, 1, 1, 2, 0, 2, 0, -2, -1, 0, -1, 0, 3, 3, 1, 1, 0, 1, 0, 1, 1, 1, 2, 0, 1, 2, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 4, 2, 1, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 2, 1, 0, -1, 0, 0, 0, 0, 4, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 3, 2, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 4, 3, 0, 0, 0, 0, 0, 1, 4, 3, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 2, 1, 2, 1, 1, 1, 1, 1, 1, 0, 2, 2, 5, 4, 1, 0, 0, 1, 1, 2, 3, 3, 0, 0, 0, 0, 0, -2, 0, 1, 2, 2, 1, 2, 1, 3, 2, 0, 0, 0, 2, 0, 1, 3, 4, 2, 1, -1, 0, 1, 1, 2, 4, 1, 0, 0, -1, 0, -3, -1, 0, 0, 1, 1, 0, 0, 0, 1, 2, 1, 0, 0, 2, 1, 2, 3, 2, 2, 0, 0, 0, 0, 0, 2, 4, 2, -1, -1, 0, -1, -4, -3, -1, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 2, 3, 2, 0, 2, 2, 0, 0, 0, 0, 0, 1, 2, 3, 1, -1, 0, -2, -3, -2, -2, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 1, 2, 4, 1, 1, 2, 0, 1, 0, 0, 0, 0, 1, 1, 3, 0, -1, -1, 0, -3, -3, -3, -1, 0, 0, 0, 1, 1, 2, 0, 1, 0, 1, 3, 3, 3, 1, 2, 1, 1, 1, 0, 0, 0, 1, 2, 3, 0, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 3, 3, 2, 3, 3, 3, 1, 2, 3, 1, 0, 0, 2, 4, 2, 2, 0, -2, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 2, 0, 1, 0, 2, 1, 2, 2, 2, 0, 0, 2, 4, 2, 2, 0, 0, -1, -1, -1, 0, -1, 0, 0, -1, -1, 0, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 1, 0, 0, 2, 4, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 1, 2, 2, 1, 1, 1, 2, 1, 2,
    -- filter=0 channel=4
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -1, -2, 0, -2, 0, -1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, -2, -1, -1, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -2, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 2, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 2, 2, 2, 2, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, 1, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 1, 2, 0, 1, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, -1, 0, 0, 2, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 1, 1, 0, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 1, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, 0, 0, -1, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 1, 0, -1, 0, -1, 0, -1, -1, -2, 0, -2, -1, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 2, 2, 2, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 2, 2, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 2, 0, 1, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 2, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 2, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, -1, -1, 0, -1, -1, 0, -1, -1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 2, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 2, 2, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, 1, 1, 2, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 1, 1, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -2, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -2, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -1, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, -3, -4, -2, -2, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -3, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -2, -3, -1, -1, -2, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 1, 1, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 3, 2, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -3, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 2, 1, 1, 1, 2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 1, 1, 2, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 1, 2, 1, 1, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -2, -2, -1, 0, 0, 0, 1, 1, 1, 1, 2, 2, 0, 1, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, -1, -1, -1, -2, -1, -1, 0, 1, 1, 1, 2, 2, 1, 2, 1, 0, 2, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -3, -2, -1, -1, 0, 0, 2, 1, 1, 1, 0, 2, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -2, -2, -2, -2, 0, -1, -2, -2, -2, -2, -1, -1, 0, 1, 0, 0, 1, 1, 1, 2, 0, 1, 0, -1, -2, -1, 0, -1, -1, 0, -2, -1, -1, -1, -1, 0, 0, -1, -1, -2, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 2, 2, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, -1, -2, 0, -1, -1, 0, -1, -1, -1, -2, 0, 0, 0, 0, -2, -1, -1, -1, -1, 0, 1, 1, 0, 0, -1, 0, -2, 0, 0, -2, 0, 0, 0, 0, -1, 0, -1, 0, 0, -2, -1, -2, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, -1, -2, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 1, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 1, 1, 1, 1, 2, 0, 0, 0, -1, -2, -2, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 2, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 0, 0, 0, 1, 1, 2, 0, 0, 0, -1, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 1, 2, 0, 0, 2, 1, 2, 1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 2, 1, 1, 2, 0, 0, 1, 2, 0, 0, 0, 0, -2, -1, 0, -2, -2, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 2, 2, 2, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -2, -2, -1, 0, -1, -2, -2, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 2, 0, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -2, -2, -2, -1, -1, -2, -2, -2, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -2, 0, 0, 0, -2, -1, -2, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -2, -2, -1, -1, -2, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, 0, 0, -1, -3, -4, -2, -4, -3, -2, 0, -1, 0, -1, 0, 0, -2, -1, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, -2, -3, -1, -1, -1, -1, -4, -3, -2, -2, -2, -3, -1, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, -1, -1, -1, -1, -1, 0, -2, -4, -2, -1, -1, -2, -1, -2, 0, 0, -1, -1, -2, -2, -2, 0, -1, 0, 0, 1, 0, 0, 1, 1, 1, 0, -1, -2, 0, -2, -1, -1, -1, -2, -2, -2, -1, -2, -1, -2, -2, -2, -1, -3, -1, -2, -3, -1, 0, 0, 1, 1, 2, 1, 1, 2, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, -2, 0, -1, -1, -1, -2, -2, -2, -2, -3, -2, -2, -3, -2, -1, -1, 0, 1, 2, 1, 1, 1, 0, 0, -1, -1, -2, -1, 0, 0, 0, -1, -1, 0, 0, 0, -2, -2, -1, -2, -1, -2, -3, -2, -2, -3, -1, -1, 0, 0, 1, 1, 2, 2, 0, 0, 0, -2, -1, 0, -1, 0, 0, -1, -1, 0, -1, -1, -1, -2, -1, -2, -2, -3, -2, -3, -3, -3, -2, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, -2, -2, -3, -4, -4, -3, -3, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, -1, 0, -1, -2, 0, 0, -1, -1, 0, 0, -1, -2, -1, -3, -1, -1, -3, -2, -5, -5, -3, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -2, -2, -1, -1, -3, -3, -3, -4, -5, -3, -1, -1, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, -1, -2, -2, 0, -1, -1, -2, -2, 0, 0, 0, -1, -2, -2, -3, -3, -4, -5, -4, -3, -2, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, -1, -1, -2, -1, -1, -1, -2, -1, -1, 0, -1, -1, -2, -2, -3, -2, -4, -5, -5, -3, -2, -1, -1, -1, -2, -1, 0, -1, 0, 0, -1, -1, -2, -3, -1, -1, -1, -3, -3, -1, 0, -1, 0, -2, -3, -2, -3, -4, -4, -5, -6, -5, -3, -2, -1, 0, -2, -1, -2, -1, 0, 0, 0, 0, -2, -2, -3, 0, -1, -3, -1, -1, -1, -1, -1, -2, -3, -2, -3, -4, -6, -7, -5, -4, -3, -3, -2, -3, -2, -1, -1, -1, 0, 0, 0, -2, -2, -1, -1, -1, -1, -3, -2, -2, -1, -2, -2, -3, -3, -3, -3, -4, -5, -5, -6, -3, -3, -2, -3, -3, -2, -2, -2, 0, 0, 0, -1, -1, -1, -2, -3, 0, 0, -2, -2, -2, -2, -2, -2, -1, -2, -2, -3, -4, -5, -5, -6, -4, -2, -2, -3, -3, -1, -2, -1, 0, 0, 0, -1, -2, -3, -3, -2, 0, -1, -1, 0, -1, 0, 0, 0, -3, -2, -3, -2, -5, -5, -6, -5, -4, -1, -2, -2, -1, -1, 0, 0, 0, -1, 0, -1, -1, -2, -2, -1, 0, -1, -2, 0, 0, -1, -1, -1, -1, -2, -2, -4, -4, -6, -5, -5, -3, -2, -2, -3, -2, -1, -1, 0, 0, 0, -1, 0, 0, -1, -2, -1, -1, -2, -2, -1, 0, -1, -1, -1, -2, -2, -3, -3, -4, -4, -5, -2, -2, -1, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, -1, -1, 0, 0, -1, -1, 0, -2, -2, -3, -3, -4, -4, -3, -4, -2, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, -3, -2, -2, -3, -2, -2, -3, -3, -2, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, -2, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, -2, -1, -2, -3, -2, -2, -3, -2, -2, -2, 0, -1, -2, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -2, -1, 0, -1, -1, -1, -1, 0, -2, -1, -2, -3, -3, -2, -4, -3, -3, -2, -2, -2, -2, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -2, -3, -2, -2, -1, -1, -2, -2, 0, -1, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, -1, -1, -1, -1, 0, 0, -1, 0, -2, -1, -3, -2, -2, -2, -3, -1, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, -1, -1, -1, -3, -1, -1, 0, 0, -2, -1, 0, -2, -1, -2, -1, -1, -1, -1, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, -2, -3, -1, 0, 0, -2, -2, -2, -1, -2, -2, -1, 0, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, -2, -1, -1, -1, -1, -1, 0, -2, -4, -2, -1, -2, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, -1, 0, -1, -1, -2, -3, -1, -1, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 2, 2, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 2, 2, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -2, -1, -2, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, -2, -3, -1, -1, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -2, -3, -2, -1, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -2, -1, -1, -2, -2, -3, -2, -2, -3, 0, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, 2, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, -2, -1, -2, -2, -2, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, -2, -3, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, -1, -1, -1, -2, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 2, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 1, 0, 1, 1, 0, 1, 1, 1, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -1, -2, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -1, 0, 0, -3, -2, -3, -2, -1, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 2, 0, 1, -1, -2, -3, -2, -1, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 0, 1, 1, 0, 1, 0, 0, -1, -2, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 1, 0, 1, 0, 0, -1, -1, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 2, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 2, 2, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 2, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 2, 2, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, -2, 0, 1, 0, 0, 2, 1, 2, 2, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, -1, 0, -1, -1, 0, -2, -1, -3, -1, 0, 0, 0, 0, 2, 2, 1, 2, 1, 0, -1, -1, -1, 0, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -4, -2, -2, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, -1, -2, -3, -4, -4, -2, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -2, -4, -4, -4, -3, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -4, -6, -6, -4, -4, -2, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -2, -2, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, -2, -3, -5, -6, -5, -5, -4, -2, -2, -2, 0, -1, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -3, -3, -3, -6, -6, -5, -6, -4, -2, -2, -2, -3, -1, 0, -1, 0, 0, 0, -1, -2, -3, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, -2, -4, -4, -7, -6, -5, -5, -4, -3, -3, -2, -2, -2, 0, -1, 0, 0, -2, -2, -2, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, -1, -4, -4, -6, -6, -6, -5, -4, -3, -3, -2, -1, -2, -1, 0, -1, 0, -2, -2, -2, -2, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, -1, -1, -2, -3, -5, -5, -4, -5, -3, -4, -2, -2, -3, 0, -1, 0, -1, -1, -1, -1, -2, -1, 0, 0, 1, 0, 0, 2, 1, 2, 0, 1, 0, -1, -2, -3, -5, -5, -4, -3, -3, -3, -3, -1, -2, -1, 0, 0, -1, -1, -2, -1, -2, 0, 0, 0, 0, 0, 2, 2, 1, 2, 3, 0, 0, -1, -2, -2, -4, -3, -4, -3, -2, -2, -1, -2, 0, -1, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 1, 1, 2, 2, 2, 1, 1, 0, 0, -1, -2, -3, -3, -3, -3, -2, -3, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 1, 1, 1, 2, 2, 3, 1, 1, 2, 0, 0, -2, -2, -4, -3, -2, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 2, 2, 2, 3, 2, 2, 0, 1, 0, 0, -2, -3, -2, -2, -2, -3, -1, -1, -2, -1, -1, -1, 0, 1, 0, 0, -1, 0, -1, 0, 1, 1, 1, 1, 2, 2, 1, 0, 1, 1, 0, -1, 0, -1, -2, -3, -2, -2, -1, 0, -1, -1, -1, 0, -1, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 2, 1, 0, 1, 1, 0, 0, 0, 0, -2, 0, -1, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, 0, 0, 0, 0, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -2, -1, -2, -1, -2, 0, 0, -1, -2, -1, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -2, -1, -2, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -3, -5, -4, -5, -4, -5, -4, -2, -1, 0, 0, -1, -2, -2, -2, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, 0, -3, -4, -7, -6, -7, -7, -7, -6, -4, -2, 0, 0, -1, -1, -1, -2, -2, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -3, -4, -7, -6, -6, -6, -7, -6, -3, -2, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 3, 2, 2, 1, 2, 0, 1, 0, -2, -2, -1, -1, -2, -3, -7, -5, -6, -4, -5, -3, -2, -1, 1, 1, 0, 0, 1, 2, 2, 1, 2, 3, 3, 4, 3, 1, 2, 1, 0, 0, 0, 0, 0, -2, -1, -3, -6, -5, -5, -4, -3, -3, -1, -1, 0, 0, 0, 0, 2, 2, 1, 2, 4, 4, 5, 4, 2, 2, 3, 2, 1, 1, 0, 0, -1, -1, -2, -4, -5, -4, -4, -3, -2, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 2, 4, 3, 3, 4, 3, 2, 2, 1, 0, 1, -1, 0, -2, -1, -4, -5, -3, -2, -2, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 2, 2, 3, 3, 2, 3, 2, 0, 1, 0, 0, 0, 0, -2, -1, -3, -3, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 1, 2, 2, 1, 2, 2, 1, 2, 0, 0, 1, 0, -1, 0, -1, -1, -2, -2, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, -1, -1, -2, -1, 0, 2, 3, 3, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 1, 2, 3, 2, 1, 2, 0, 0, 0, -1, -1, -2, -1, 0, 1, 2, 2, 4, 3, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, -2, -1, 0, 1, 3, 3, 2, 3, 2, 0, 0, 0, -2, -3, -2, -2, 0, 0, 2, 2, 3, 2, 4, 3, 2, 2, 2, 2, 3, 1, 0, 0, -1, 0, 0, 0, 1, 2, 2, 3, 1, 1, -1, -3, -3, -5, -4, -3, -2, 0, 0, 0, 2, 2, 2, 2, 2, 2, 4, 3, 3, 2, 0, -1, 0, 0, 0, 1, 0, 1, 3, 2, 1, 2, 0, -2, -3, -5, -4, -3, -2, -2, -2, -1, -1, 0, 1, 3, 4, 4, 6, 5, 5, 3, 0, -1, -1, -1, 0, 0, 1, 0, 1, 1, 3, 1, 1, -1, -2, -5, -5, -5, -5, -4, -3, -4, -4, -2, 0, 3, 4, 3, 4, 5, 4, 1, 0, 0, 0, -1, 0, 1, 1, 0, 3, 3, 3, 3, 0, -1, -3, -4, -5, -5, -6, -6, -6, -6, -7, -4, -3, 0, 3, 3, 4, 4, 2, 2, -1, -1, -1, -1, -1, 0, 0, 1, 3, 4, 3, 3, 1, 0, -2, -4, -4, -5, -6, -8, -8, -8, -7, -6, -3, 0, 2, 3, 3, 3, 2, 1, -1, 0, 0, 0, -1, 0, 1, 2, 3, 3, 3, 2, 2, 0, -2, -2, -3, -5, -6, -8, -8, -9, -9, -5, -4, 0, 1, 3, 4, 3, 3, 1, 0, -1, 0, -1, -1, 0, 1, 0, 3, 4, 5, 4, 2, 0, -1, -3, -3, -4, -4, -6, -8, -7, -6, -3, -1, 0, 1, 3, 3, 2, 1, 1, 0, -1, 0, -1, 0, 0, 0, 2, 2, 4, 4, 3, 2, 0, -1, -2, -3, -3, -4, -4, -6, -5, -4, -3, 0, 1, 2, 5, 3, 3, 2, 0, 0, -1, 0, -1, 0, 1, 0, 1, 3, 3, 4, 2, 2, 1, -1, -2, -3, -3, -2, -3, -3, -3, -1, 0, 2, 2, 3, 3, 2, 3, 1, 1, -1, -1, 0, 0, 1, 1, 2, 2, 2, 3, 3, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 3, 4, 4, 2, 3, 2, 1, 0, -1, 0, 0, 2, 2, 3, 1, 1, 1, 3, 2, 0, 1, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 3, 2, 3, 3, 2, 3, 2, 1, -1, 0, 0, -2, 1, 4, 2, 3, 0, 1, 2, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 2, 2, 4, 3, 3, 2, 0, 0, -1, 0, 2, 3, 2, 1, 0, 1, 1, 2, 1, 0, -1, 0, 0, 1, 1, 2, 1, 1, 1, 2, 2, 2, 2, 2, 2, 3, 2, 1, -1, 0, -1, -2, 0, 2, 2, 1, 1, 1, 0, 1, 1, 0, -1, -1, 0, 0, 2, 1, 3, 2, 2, 3, 3, 2, 1, 3, 2, 2, 1, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 3, 3, 3, 3, 3, 3, 4, 3, 3, 2, 1, 0, 0, -1, -1, -2, -4, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 3, 4, 2, 3, 2, 3, 3, 4, 2, 3, 0, 0, 0, -1, -1, -3, -4, -2, -2, -3, -4, -4, -2, 0, 0, 0, 0, 0, 0, 0, 1, 3, 3, 3, 4, 3, 2, 2, 1, 1, 0, 1, 1, 0, -1, 0, -2, -4, -4, -3, -4, -5, -5, -6, -5, -2, 0, 0, 0, 0, 0, 0, 2, 2, 3, 3, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -5, -7, -3, -5, -5, -5, -6, -5, -4, -3, -1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, -2, -2, -2, -1, -1, -1, -1, -3, -1, -2, -2, -3, -6, -4, -3, -3, -4, -4, -5, -3, -3, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, -3, -2, -2, -3, -3, -1, -1, -1, -1, -1, -2, -1, -2, -1, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -2, -3, -2, -2, -2, -2, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -2, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 2, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 2, 2, 1, 0, -1, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 2, 3, 2, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 3, 0, 0, 1, 4, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 2, 2, 2, 1, 1, 3, 3, 0, 0, 0, 1, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 2, 2, 1, 2, 2, 2, 0, 0, 0, 0, 2, 1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 2, 2, 2, 0, 0, 0, 0, 1, 0, 0, -2, -1, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 2, 2, 3, 2, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -2, -2, -2, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, -1, -1, -1, 0, 1, 2, 2, 2, 2, 0, 0, 0, 0, -1, 0, -2, -1, -1, -1, -3, -3, -1, -1, 0, 0, 0, 1, 3, 2, 2, 1, 1, 0, 0, 0, 0, 1, 3, 3, 3, 2, 1, 0, 0, 0, -1, -1, -1, -2, -2, -1, -2, -4, -2, -2, 0, 0, 0, 0, 2, 3, 1, 2, 1, 1, 0, 1, 1, 1, 1, 2, 4, 3, 1, 0, 1, 0, -1, -1, -2, -2, -2, -1, -1, -1, -2, -1, 0, 0, 1, 0, 2, 3, 2, 1, 1, 2, 1, 1, 2, 1, 1, 1, 3, 2, 1, 0, 1, 0, -1, 0, -1, -2, -2, 0, -2, 0, -2, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 1, 1, 2, 1, 1, 0, 1, 1, 2, 0, 1, 0, 0, 0, -1, -1, -2, -2, -1, -1, -1, -2, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -2, -2, -3, -2, -1, -1, -1, 0, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -3, -3, -2, -2, -2, -1, 0, 0, 1, 0, 1, 0, 0, -1, -1, 0, 0, -1, -2, -1, 0, 0, 2, 1, 0, -1, 0, 1, -1, -1, -1, 0, -2, -3, -1, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -2, 0, -2, -2, -1, 0, 1, 0, 0, 0, 1, 0, -1, -2, -2, -1, -1, -2, -1, 0, -1, -1, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, -2, -1, 0, 1, 2, 0, -1, 0, 0, 0, -1, -2, -1, -1, -2, -3, -4, -1, 0, 0, 0, -1, 0, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, -1, 0, 0, 0, -2, -1, -1, -1, -2, -3, -1, -1, 0, 0, 0, 0, 1, 3, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 2, 0, 0, 0, 0, 1, 0, -1, -1, -1, -1, -2, -2, -2, -1, 0, 1, 0, 0, 0, 2, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 2, 1, 0, 0, 1, 1, 0, 0, -1, -2, -1, -1, -3, -3, -2, -1, 0, 1, 2, 1, 3, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 2, 0, 0, 1, 1, 0, 0, -1, -1, -1, -2, -2, -2, -2, -1, 0, 0, 0, 2, 3, 2, 2, 0, 0, 0, 0, 1, 1, -1, 0, 0, 2, 2, 0, 0, 1, 1, 1, 0, 0, -1, -1, -1, -2, -2, -2, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 2, 2, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 1, 1, 0, 0, 1, 3, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 1, 0, 0, 0, 1, 2, 0, -1, -2, -1, 0, 2, 1, 0, 0, -1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 2, 2, 2, 1, 0, 0, 0, 0, 1, 1, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 0, -1, 0, -2, -2, -2, -1, -1, -2, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -4, -3, -2, -3, -3, -3, -2, -1, 0, 0, -1, 0, -1, -2, -1, -1, 0, 0, 1, 1, 1, 1, 0, 2, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -2, -2, -3, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 1, 2, 2, 2, 0, 0, 0, 1, 1, 1, 0, -2, -1, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 2, 2, 0, 1, 0, 1, 0, 0, -2, -1, -2, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 2, 2, 2, 1, 0, 1, 1, 2, 0, -2, 0, -2, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 1, 0, 1, 2, 2, 0, 0, 1, 0, 2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, -1, -1, -1, 0, 0, 0, 1, 2, 2, 1, 1, 0, 0, -1, 0, 0, 1, 0, -1, 0, -1, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 1, 1, 0, 0, 1, 0, 2, 1, 0, 0, -1, 0, 1, 1, 0, 0, 1, 1, 1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 2, 1, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 2, 2, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, -3, -2, -2, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -4, -1, -2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -2, -4, -2, -2, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 1, 0, -1, -2, -2, -2, -1, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 2, 1, 2, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 3, 2, 2, 0, 0, 1, 1, 2, 3, 2, 1, 0, 0, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 3, 2, 1, 1, 1, 1, 2, 1, 3, 2, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 2, 1, 2, 3, 1, 0, 0, 0, 1, 2, 2, 0, 1, 2, 1, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 1, 1, 2, 3, 2, 0, 0, 0, 1, 2, 3, 1, 2, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 3, 3, 3, 0, 2, 2, 1, 1, 3, 2, 1, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 3, 3, 3, 2, 1, 3, 2, 3, 3, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 3, 2, 3, 1, 2, 2, 2, 2, 3, 2, 0, 0, -1, 0, -1, -2, -2, 0, 0, -1, 0, -1, -2, 0, 0, 0, -1, 0, 0, 1, 0, 2, 2, 2, 1, 1, 1, 1, 1, 2, 1, 1, 0, 0, -1, -1, 0, -2, -1, 0, 0, -2, -1, -2, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 1, 2, 1, 1, 1, 1, 1, 1, 0, -1, -1, -1, -2, -1, -1, 0, -2, -1, -2, -2, -2, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, 0, 0, 0, -1, -3, -3, -2, 0, 0, -1, -1, -1, -1, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, -2, -1, -1, -1, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, -2, -2, -3, -3, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, 0, -1, 0, -2, -2, -2, -2, -3, -2, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 1, 0, -1, -1, 0, 0, 0, -1, -2, -2, -1, -1, -1, -1, -1, -2, -1, -2, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -3, -3, -3, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 2, 0, 0, -1, -1, -1, -1, 0, 1, 1, 0, -1, -3, -3, -3, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 0, -1, -1, 0, -2, 0, -1, -1, -2, -2, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, -1, 0, 0, -1, -3, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, -2, -2, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 2, 3, 1, 2, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 2, 4, 4, 4, 4, 4, 3, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, -2, -2, -1, 0, 0, 1, 2, 3, 4, 5, 5, 4, 3, 3, 1, 1, 1, 0, 0, 2, 3, 2, 0, 1, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, 2, 1, 3, 4, 6, 5, 4, 3, 2, 1, 3, 1, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 1, 2, 3, 4, 2, 2, 1, 2, 1, 2, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, -3, -4, -4, -3, -3, -2, -2, 0, 0, 1, 1, 0, 0, 2, 2, 1, 2, 1, 3, 3, 3, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -2, -3, -3, -4, -3, -2, -1, 0, 1, 1, 1, 1, 0, 0, 1, 0, 1, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, -1, -1, -3, -3, -1, -1, -1, 0, 1, 2, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, -1, -1, -3, -1, -2, -2, -1, -2, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -2, -1, -2, -2, -2, -1, -3, -2, 0, 1, -1, -1, -1, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, -2, -1, -1, -1, -3, -3, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, -2, -1, -2, -3, -1, -1, 0, -1, -2, -2, -1, -2, -1, -2, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -3, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, -3, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, -1, -1, -1, -1, 0, 0, 0, -1, -2, -2, -2, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, -2, 0, 0, -1, -1, 0, 0, 0, -2, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, -2, 0, 0, 1, 1, 0, 0, -2, -2, -2, -2, -3, -2, -3, -1, -2, -1, -2, -1, -1, -1, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, -2, -3, -2, -2, -1, -1, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -3, -2, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 2, 0, 1, 0, 0, 0, 1, 0, -1, -1, -1, -4, -2, 0, 0, -1, -2, -3, -2, -1, 0, 0, 0, 0, -1, 0, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 3, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, -2, 0, 0, 0, 2, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 2, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, -1, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 0, 0, -1, -1, 0, -2, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -2, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, 0, -1, 0, -1, 0, 0, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -2, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 2, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 2, 1, 2, 1, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, -2, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 2, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 2, 1, 0, 1, 2, 1, 2, 2, 0, 1, 1, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 2, 2, 1, 2, 1, 1, 1, 2, 1, 0, 0, 0, -2, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 1, 1, 2, 1, 1, 1, 2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 2, 0, 0, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 2, 0, 1, 0, 1, 0, 2, 1, 2, 1, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 2, 2, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 1, 2, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 2, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 3, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 2, 1, 1, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 1, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 3, 3, 2, 2, 2, 0, 0, 2, 0, 0, 1, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 2, 1, 3, 2, 3, 3, 1, 0, 0, 1, 1, 1, 1, 1, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 3, 1, 2, 1, 1, 0, 0, 0, 1, 1, 1, 1, 1, 2, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, 1, 0, 0, 1, 2, 2, 3, 2, 1, 2, 1, 0, 2, 2, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 3, 2, 2, 0, 1, 2, 2, 2, 2, 2, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 2, 1, 1, 1, 0, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 1, 0, 1, 2, 2, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, -2, -2, -2, -2, -2, -1, -2, 0, -1, 0, 0, 0, 0, -1, -2, 0, -1, 0, 1, 1, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, -1, 0, -5, -4, -4, -3, -2, -3, -2, 0, -1, 1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -3, -3, -3, -2, -2, -2, -2, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, -3, -2, -2, -1, -2, -2, -2, 0, 0, 1, 0, 0, 1, 0, 0, 0, 2, 2, 2, 2, 2, 0, 2, 1, 0, 0, 0, 0, 2, 1, 1, 0, -3, -2, -1, -2, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 1, 2, 1, 2, 1, 2, 1, 0, -1, 0, 1, 2, 0, 0, -2, -3, -3, -2, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 1, 2, 1, 3, 1, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, -2, -2, -2, -2, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 2, 2, 1, 1, 1, 1, 1, -1, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, -2, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -2, -2, -1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 2, 1, 0, -2, -2, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, -2, -2, 0, 0, 0, 1, 1, 2, 1, 2, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, -1, -2, -3, -2, 0, 0, 1, 0, 0, 1, 2, 0, 1, 0, 0, 0, 1, 1, 2, 2, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, -3, -4, -2, -1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 2, 2, 2, 1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, -3, -2, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 1, 2, 3, 1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, -1, -3, -3, -2, -3, -2, -1, 0, -1, -2, 0, -1, 0, 1, 2, 1, 2, 2, 1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 1, 2, 0, 0, -1, -3, -1, -1, -2, -2, -1, -3, -2, -2, -1, -1, 0, 1, 1, 2, 1, 1, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, 2, 2, 1, 0, -1, -2, -1, -2, -4, -4, -3, -3, -3, -2, -1, 0, 0, 0, 1, 2, 2, 1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -1, 0, -1, -2, -3, -4, -3, -2, -1, -1, 0, 0, 0, 2, 2, 2, 0, 0, 0, -2, 0, -1, -1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, -1, 0, -3, -3, -4, -2, -1, 0, -1, 0, 1, 0, 0, 1, 2, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 2, 1, 1, 0, 0, 0, -1, -1, -3, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 2, 2, 1, 0, -2, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 2, 1, 0, 0, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -2, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, -2, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 1, 0, 0, 1, 0, 0, 1, 1, 0, -1, 0, 0, 0, -2, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, -2, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 2, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -4, -2, 0, 0, -2, -3, -2, -2, -1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 2, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, -3, -3, 0, 0, -1, -3, -3, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, -1, 0, 0, -4, -3, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -2, -2, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -2, -1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 2, 2, 2, 2, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 2, 1, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 1, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 1, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 2, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 0, 0, 0, 0, -2, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 2, 1, 2, 1, 0, 0, -1, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, -1, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 2, 2, 1, 1, 1, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 2, 1, 0, -1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -2, -1, -1, -2, -2, 0, -1, 0, 0, 0, 0, 0, 1, 0, 2, 2, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 2, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 1, 2, 2, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, -1, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 1, 2, 0, 1, 1, 2, 2, 1, 0, 0, 0, -1, 0, 1, 0, 0, 1, 1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 1, 1, 1, 2, 0, 0, 1, 0, 0, 0, 0, 2, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 1, 1, 2, 2, 1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 1, 0, 0, 0, 1, 0, 2, 0, 0, -1, -1, 0, 0, 1, 1, 1, 0, -1, 0, 0, -1, 1, 2, 1, 0, 0, 0, 1, 1, 1, 2, 5, 3, 0, 0, 2, 1, 1, 0, 0, 0, -1, -1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 2, 2, 5, 3, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 3, 0, 1, 1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 1, 1, 0, 0, 0, -2, -2, 0, 1, 0, 0, -1, 1, 1, 0, -1, 2, 5, 2, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 1, 0, 0, -2, 0, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 3, 3, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, -2, -2, -1, -1, 0, -1, 0, -1, 0, -1, 0, 0, -1, 1, 3, 1, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -2, 0, -2, -1, 0, 0, -2, 0, -1, 0, -1, 0, 1, 2, 1, 1, 0, -1, -1, 0, -1, 0, 0, 1, 0, 0, 1, 1, 3, 1, 0, 0, -2, -1, -2, -2, -1, -1, -1, -3, 0, -2, 0, 0, 1, 3, 1, 0, 0, -1, -2, 0, 0, -1, 0, 1, 0, 0, 1, 2, 0, 0, -2, 0, 0, -1, -2, -3, -2, -1, -1, -1, -3, -1, -1, -2, 0, 1, 2, 0, 0, -1, -2, -1, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, -2, -2, 0, -1, -2, -3, -3, -3, -2, -3, -2, -2, -2, -1, 0, 2, 3, 0, 1, -3, -3, -2, -1, -1, -2, 0, 1, 0, 0, 2, 0, 0, 0, -2, -1, 0, -1, -3, -2, -2, -2, -3, -3, -2, -2, -1, 0, 4, 2, 0, 0, -1, -4, -3, 0, 0, -2, -2, 0, 0, 0, 1, 2, 0, 0, -1, -1, 0, -1, -1, -3, -3, -3, -4, -5, -1, -3, -1, 0, 3, 3, 0, 0, -2, -2, -2, -2, -1, -2, -2, -1, 0, 0, 1, 2, 0, 0, -2, -1, -1, -2, -2, -4, -3, -3, -3, -4, -2, -3, -1, 0, 3, 2, 0, 1, -2, -3, -2, -1, -2, -4, -3, -2, 0, 1, 1, 2, 0, 1, -1, -2, -2, -2, -4, -4, -3, -3, -4, -5, -2, -2, -1, 1, 2, 2, 0, 0, 0, -3, -3, -2, -2, -2, -3, -4, 0, 0, 0, 0, 0, 0, -1, -2, -3, -4, -4, -3, -3, -5, -4, -4, -3, -3, 0, 1, 2, 0, 0, 0, 0, -1, -2, -3, -2, -3, -5, -4, 0, 1, 1, 0, 0, 0, -1, -2, -1, -2, -3, -4, -3, -4, -4, -5, -4, -2, -1, 2, 1, 0, 0, 0, 0, -1, -3, -2, -2, -2, -3, -3, 0, 2, 2, 2, 0, 1, -1, -1, -3, -4, -2, -3, -3, -3, -3, -4, -5, -3, -1, 1, 1, 0, 0, 0, 0, 0, -3, -3, -2, -3, -4, -3, 1, 3, 3, 3, 1, 0, -1, -1, -3, -3, -2, -2, -2, -3, -5, -5, -4, -2, -1, 1, 3, -1, 0, 0, 0, -1, -2, -4, -3, 0, -2, -1, 0, 0, 4, 2, 0, 0, -1, -2, -2, -2, -2, -1, -3, -2, -4, -4, -3, -2, -1, 1, 3, 0, 0, 0, -2, 0, -3, -3, -2, -1, -1, 0, 0, 1, 4, 2, 0, 0, -2, 0, 0, -2, -2, -2, -1, -3, -2, -1, -3, -3, -3, 0, 2, 0, 0, 0, -1, -1, -2, -2, -1, 0, -1, 0, 0, 0, 4, 3, 0, 0, -1, 0, 0, -1, -2, 0, -1, -3, -2, -2, -2, -3, -1, 0, 3, 1, 0, 0, -1, -1, -2, -1, -2, 0, 0, 0, -2, 0, 5, 2, 0, 0, 0, -1, 0, 0, -1, -2, -2, -1, -1, -1, 0, -2, -2, 0, 2, 1, 0, 0, -1, -2, -2, -1, -1, 0, -1, 0, -1, 0, 3, 1, 0, 0, 0, -1, 1, 0, -1, -1, -2, -2, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -2, 0, 2, 1, 0, 0, 1, 0, -1, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, 0, -1, 0, -1, -2, -2, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, -2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, -1, -2, -2, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 3, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, -2, -1, 0, 0, -1, -1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, -1, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 3, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, 1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 3, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -2, -3, -3, -2, -2, -2, -2, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -2, -2, -3, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -3, -2, -1, -1, -2, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, -1, -3, -1, -1, -2, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -1, -2, 0, -1, -2, 0, -1, 0, -1, -2, -1, 0, -1, -1, 0, 1, 1, 1, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -3, -2, -1, -2, -1, -1, 0, 0, -1, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, -2, 0, 0, 0, 0, -1, -1, -1, -1, -2, -2, 0, 0, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, -2, -1, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, -2, -1, -1, 0, -1, 0, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, -2, -2, -1, -1, 0, -1, 0, 0, 0, 1, 2, 1, 1, 0, -1, 0, -1, 0, -1, -1, 0, -1, 0, -1, -1, -1, 0, -1, -1, -1, -2, 0, 0, -1, -3, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, -1, -1, -1, -1, -1, 0, -1, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, -1, 0, 0, 0, 0, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, -2, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -2, -1, 0, 0, 0, -1, -1, -1, -1, 0, -1, -2, 0, -1, -2, -1, -2, -2, 0, -2, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, -1, -2, -2, -1, -1, -1, -2, -1, -1, -1, -1, -1, -2, 0, 0, 0, 0, -1, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -2, -2, -1, -1, 0, 0, -1, 0, -1, -1, -3, -2, -1, 0, 0, 0, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -2, 0, -2, -1, -1, -2, 0, 0, 0, -2, -1, -1, -2, -1, 0, 0, -1, -2, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -1, 0, 0, -2, 0, 0, -1, -2, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -2, -2, 0, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -2, -1, -2, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, -1, -1, 0, 0, 0, 0, -2, -1, 0, -1, -1, -1, -2, -1, -1, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, -2, -2, -2, -1, -1, -1, -1, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, -1, -1, -1, -1, 0, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, -1, 0, -2, -1, 0, -1, -1, -2, -1, 0, 0, -1, -1, -1, -2, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -2, -2, -1, 0, -2, -2, -1, -2, -1, 0, -2, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -3, -2, 0, 0, 0, -2, -2, -1, -1, -1, 0, -2, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -2, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 0, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 1, 1, 1, 1, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 2, 2, 1, 1, 0, 1, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 0, 0, 0, 1, 1, 0, 2, 1, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 1, 1, 1, 1, 2, 2, 2, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 2, 2, 3, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 0, 2, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, -1, 0, 0, 2, 0, 1, 2, 1, 2, 1, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 2, 2, 3, 2, 1, 0, 0, -1, -1, -1, 0, 0, -1, -1, -1, 0, -1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 2, 3, 2, 2, 0, 0, 0, -2, -1, -2, -1, -1, 0, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 2, 2, 2, 2, 0, 0, -2, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 2, 2, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 3, 1, 1, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 2, 1, 2, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 2, 3, 2, 1, 0, 0, -1, 0, -1, -2, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 2, 1, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, -1, -1, -1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 2, 0, 0, 0, 1, 1, 0, -1, -1, -1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -5, -4, -5, -5, -4, -3, -2, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 2, 2, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -3, -4, -4, -3, -4, -5, -3, -2, 0, 0, 1, 0, -1, -1, 0, -1, 0, 1, 1, 2, 1, 0, 1, 1, 2, 0, 0, -1, -2, -1, 0, -1, -4, -4, -4, -3, -2, -4, -3, -2, -1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 1, 2, 1, 2, 2, 2, 1, 0, 0, -1, 0, 0, -1, -2, -3, -4, -4, -3, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 4, 3, 2, 2, 2, 1, 1, 0, 0, 0, 0, -1, -3, -4, -4, -3, -2, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 3, 4, 4, 3, 2, 1, 2, 0, 0, -1, 0, 0, 0, -1, -3, -2, -2, -2, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 3, 2, 3, 2, 2, 1, 2, 1, 0, 0, 0, 0, -2, -2, -3, -2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 2, 3, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 2, 1, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -2, -2, 0, 1, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -2, -1, 0, 1, 1, 1, 1, 3, 3, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 0, 1, 1, 0, 0, -1, -2, -1, -1, -1, 0, 0, 1, 2, 2, 3, 3, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -4, -4, -4, -2, -1, 0, 0, 0, 1, 1, 2, 1, 2, 2, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -2, -3, -3, -4, -4, -2, 0, -1, 0, 0, 0, 2, 2, 2, 4, 4, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, -5, -3, -3, -3, -2, -2, -2, -2, -1, 0, 2, 3, 3, 4, 2, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -3, -4, -3, -3, -4, -3, -3, -3, -3, -2, 0, 0, 3, 4, 3, 2, 0, 0, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -4, -3, -2, -3, -3, -5, -4, -5, -3, -1, 0, 1, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -3, -2, 0, -2, -2, -4, -5, -5, -4, -3, 0, 0, 1, 3, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -2, -2, -1, -2, -2, -4, -3, -4, -2, 0, 2, 1, 2, 1, 0, 1, 0, -2, 0, 0, -1, 0, 0, -1, 0, 2, 0, 0, 0, 0, 0, -2, -3, -2, -1, -1, -1, -1, -2, -1, 0, 1, 0, 1, 1, 2, 0, 0, -1, -1, 0, -1, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 1, 1, 2, 2, 3, 2, 2, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 3, 3, 4, 2, 2, 1, 1, 0, 0, 0, -1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 2, 1, 1, 0, 1, 1, 3, 3, 3, 1, 0, 0, 1, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 2, 1, 0, 1, 2, 2, 3, 2, 3, 2, 0, 0, 0, 0, -1, -1, -1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 3, 3, 3, 2, 1, 1, 2, 3, 3, 3, 1, 0, 0, 0, -1, 0, -1, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 2, 3, 3, 2, 3, 4, 3, 4, 2, 1, 1, -1, -1, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 4, 4, 3, 3, 3, 3, 3, 4, 3, 2, 0, 0, -2, -2, -1, -2, -2, -1, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 3, 3, 4, 2, 2, 4, 3, 2, 1, 2, 0, 0, -2, -1, -2, -2, -3, -2, -2, -3, -2, -1, -1, -1, 0, 0, 1, 0, 0, 1, 1, 3, 2, 2, 3, 3, 1, 2, 2, 0, 0, 0, 0, 0, -2, -1, 0, -3, -5, -3, -2, -2, -3, -3, -2, -2, -2, 0, 0, 0, 0, 1, 0, 1, 1, 3, 3, 1, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, -3, -5, -3, -2, -1, -3, -2, -4, -3, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -2, -4, -3, -2, -2, -1, -1, -3, -3, -2, -2, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, -2, -1, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 1, 1, 1, 1, 0, 1, 2, 2, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 2, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 1, 2, 0, 0, 0, 0, 2, 2, 2, 2, 1, 0, 0, 2, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 2, 3, 0, 1, 0, 1, 1, 0, 1, 2, 1, 1, 2, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 3, 1, 2, 2, 0, 2, 0, 2, 2, 2, 2, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 1, 1, 0, 0, 2, 2, 1, 1, 1, 1, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 2, 2, 1, 2, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 0, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 1, 2, 1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -2, -2, -1, -2, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -2, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -2, -1, -1, -2, -2, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, -1, -1, -2, -1, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 2, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -3, -2, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 2, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -2, -1, -2, -1, -2, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, -1, -1, 0, -2, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 0, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 1, 1, 2, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 0, 2, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 0, 0, 1, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 0, 1, 2, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, 2, 0, 0, 2, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -2, -2, -3, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -2, -2, -2, 0, -1, 0, -1, -3, 0, -1, -1, -2, -1, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, -2, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -2, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -2, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, -2, -1, -1, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -2, -2, -1, -3, -2, -2, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, -2, -2, -2, -2, -3, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, -3, -2, -1, -2, -2, -2, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, -1, -2, -2, -1, -1, -3, -3, -4, -2, -2, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -3, -1, 0, -1, -1, -1, -2, 0, -1, -1, -1, 0, -2, -1, -2, -3, -3, -5, -3, -2, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -2, -2, -2, -1, -1, -4, -4, -5, -4, -3, -1, 0, -1, -2, -1, 0, -1, 0, 0, -1, 0, 0, -2, -1, 0, -1, -2, -1, 0, 0, 0, -2, -2, -2, -1, -2, -3, -3, -4, -4, -3, -3, -2, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, -2, -2, -2, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, -2, -4, -4, -4, -4, -4, -3, -3, -1, -2, -1, -1, -1, -1, -1, -1, 0, -2, -2, -2, 0, 0, -1, -1, 0, 0, -1, -1, -2, -1, -2, -1, -3, -3, -3, -5, -4, -4, -3, -2, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -2, -2, -4, -4, -2, -2, -2, -1, -2, -2, -2, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -2, -2, -1, -1, -3, -3, -2, -3, -1, -1, -1, -1, -1, -2, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -3, -2, -3, -3, -1, -1, 0, -1, -2, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -3, -2, -3, -3, -3, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -2, -2, -2, -3, -2, -2, -1, 0, 0, -2, 0, 0, 0, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, -1, -2, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, -2, -2, -2, 0, -1, -1, 0, -2, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, -2, -1, 0, -2, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -2, -1, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, -1, -1, -1, -2, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, -2, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, -1, -2, -1, -2, -1, -1, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -2, -1, -1, 0, -1, 0, 0, -3, -2, -3, -4, -2, -3, -3, -2, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, -1, -2, -1, 0, -2, -1, 0, -1, -1, 0, -2, -3, -3, -4, -3, -3, -2, -2, -2, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -3, -3, -2, -3, -2, -3, -2, -2, -1, -1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 2, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -3, -2, -3, -2, -1, -2, -2, -1, -2, -1, 0, 0, 0, 2, 1, 1, 2, 1, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -1, -3, -3, -2, 0, -2, -1, -1, -1, 0, 0, 1, 2, 2, 1, 1, 1, 1, 1, 2, 1, 1, 0, 1, 0, 0, 1, 1, 0, -1, 0, -2, -1, -1, -2, -1, -1, -1, 0, -1, -1, 0, 1, 0, 0, 0, 0, 1, 2, 1, 2, 2, 2, 0, 1, 0, 1, 0, 0, 2, 1, -1, 0, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, -1, 0, -3, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 1, 1, 1, 0, 0, 0, 2, 1, 2, 0, 0, -2, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 0, 1, 1, 0, 0, 1, 2, 1, 0, 0, -2, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 1, 2, 0, 0, 2, 0, 0, 3, 2, 3, 0, 0, 0, 0, -1, 0, 1, 0, 1, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 2, 1, 0, 2, 2, 4, 3, 0, 0, -2, 0, -1, 0, 0, 1, 0, 1, 3, 1, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 4, 3, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 3, 3, 3, 1, 0, -1, 0, -1, -2, 0, -1, -1, -1, -1, 0, 1, 2, 1, 1, 1, 3, 2, 1, 0, -1, -1, -1, 0, 0, 0, 1, 2, 3, 4, 3, 1, 1, 0, -1, -2, -3, -3, -3, -3, -2, -2, -1, 0, 1, 1, 1, 1, 2, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 3, 3, 3, 2, 1, 2, 0, -1, -3, -4, -5, -4, -3, -3, -3, -2, 0, 0, 1, 1, 1, 1, 2, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 3, 2, 3, 2, 1, 0, 0, -3, -4, -3, -4, -3, -3, -2, -1, -1, 0, 0, 3, 2, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 4, 2, 3, 2, 1, 0, -1, -1, -3, -4, -3, -3, -3, -2, -1, 0, 0, 2, 2, 2, 3, 3, 0, 0, -2, 0, 0, 0, 0, 0, 1, 2, 2, 4, 3, 1, 0, 0, -1, -1, -2, -2, -2, -3, -3, -2, -1, 0, 0, 0, 1, 3, 2, 2, 0, 0, -1, -1, 0, 0, 0, 0, 2, 2, 3, 3, 2, 2, 1, 0, -1, 0, -1, -3, -1, -2, -2, -1, 0, 0, 0, 1, 2, 1, 3, 2, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 2, 2, 3, 2, 1, -1, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 1, 0, 1, 2, 2, 1, 0, -1, 0, 0, 0, 1, 1, 1, 2, 1, 2, 2, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 1, 1, 0, 1, 2, 2, 1, 0, -1, 0, 0, 0, 1, 2, 2, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 1, 0, 1, 2, 4, 3, 0, 0, -2, 0, 1, 2, 2, 2, 0, 0, 0, 0, 2, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 3, 2, 0, 0, -2, 0, 1, 1, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 1, 0, -2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 1, 1, 2, 0, 0, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, -2, 0, 0, 0, -2, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, -1, 0, 0, -2, -2, -3, -1, -1, -1, 0, 0, 1, 1, 1, 1, 2, 3, 2, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -3, 0, 0, -1, -1, -3, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 1, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, -3, -1, 0, -1, -1, -2, -3, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 3, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, -1, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, -2, -2, -1, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, -1, -1, -2, -2, 0, -2, -1, -3, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -2, -1, -2, -1, -2, -2, -1, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -2, -1, -3, -2, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -3, -2, -1, -1, -1, -2, -3, -2, -2, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, -3, -1, -2, 0, -1, -2, -4, -3, -3, -3, -3, 0, -1, -1, 0, 0, 0, 0, -1, -2, -4, -2, 0, -2, -3, -2, 0, -1, 0, 0, 0, 0, -2, -3, -2, -1, -2, -3, -3, -2, -1, -4, -1, -2, -1, 0, 1, 0, 0, 1, 0, -2, -3, -2, -2, -2, -2, -1, -2, -1, 0, 1, 0, 0, -1, -4, -3, -3, -3, -2, -3, -2, -3, -2, -1, -2, -1, -1, 1, 0, 0, 0, 0, -2, -2, -1, -2, -2, -2, -2, -1, 0, 1, 0, 0, 0, -1, -3, -2, -2, -2, -3, -2, -2, -2, -2, 0, -1, -1, 0, 2, -1, 0, 1, 0, -1, -2, -2, -3, -2, -3, -3, -1, 0, 0, 1, -1, -1, -1, -3, -2, -3, -4, -4, -2, -2, -3, -4, -2, -2, -1, 0, 2, -1, 0, 0, 0, 0, -2, -1, -1, -2, -3, -2, -2, 0, 1, 1, -1, 0, -1, -4, -2, -3, -4, -2, -3, -3, -3, -3, -3, -3, -1, 0, 2, 0, 0, 1, 0, -1, -1, -2, -3, -2, -1, -2, -2, 0, 2, 3, 0, 0, -2, -3, -2, -2, -2, -1, -3, -2, -3, -3, -2, -2, -2, 0, 2, 0, 0, 0, 0, -2, -2, -2, -4, -1, 0, -2, -2, -1, 2, 2, 0, 0, -2, -3, -1, -3, -3, -1, -2, -2, -3, -2, -2, -2, -1, -1, 2, -1, 0, 0, 0, -2, 0, -2, -2, 0, 0, -2, -1, -1, 0, 2, 0, -2, -2, -3, 0, -2, -2, -1, -1, -1, -3, -3, -1, -1, -2, -2, 1, 0, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, -2, 0, 2, 0, 0, -1, -1, 0, 0, -2, -1, 0, -2, -1, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, -1, -1, -1, -2, 0, -1, 0, 0, -2, 1, 2, 0, 0, -1, -1, 0, 0, 0, -2, -1, -1, -2, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, -2, -1, -2, -1, 0, 0, 0, 0, -1, 1, 2, 1, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, -2, 0, 1, 0, 0, -1, -1, -1, 0, -1, -1, -1, -2, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, -1, 0, -2, 0, 1, -1, 0, -1, -2, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, -1, -3, -1, -2, 0, 0, 1, 0, 0, -1, 0, 1, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -2, -2, -2, -1, 0, 0, 0, 0, -3, 0, 1, -1, 0, -1, -1, -1, -1, -1, 0, 0, -1, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 1, 1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -2, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, -1, 0, 0, -1, -2, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, -1, -1, -1, -1, -2, 0, -1, -2, 0, 0, -1, -1, -1, 0, 0, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 2, 1, 1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 1, 1, 0, 1, 1, 1, 0, 0, 1, 2, 1, 0, 0, 2, 2, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, -1, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, 1, 2, 1, 0, 0, -1, -1, -1, 0, 1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 2, 3, 2, 1, 1, 2, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 2, 3, 4, 2, 3, 2, 3, 1, 2, 1, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 2, 2, 3, 2, 3, 3, 2, 1, 2, 2, 1, 3, 2, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 2, 2, 2, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 1, 0, 1, 1, 0, 2, 3, 2, 2, 2, 1, 1, 0, -1, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 2, 3, 3, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, -2, -3, -1, -1, 0, 0, -1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 1, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -2, -1, 1, 2, 0, 0, -1, -1, -1, 0, -2, -2, 0, 0, -1, 0, 1, 2, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, -2, -2, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, -2, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 2, 1, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -2, -3, -2, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, 0, 2, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 1, 0, -1, -1, -2, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -2, -1, -2, -2, -1, 0, 0, 1, 0, 0, 0, 0, -1, -2, -1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, 0, -1, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 2, 0, -1, -2, -1, -1, 0, 1, 0, -2, 0, 0, 0, 0, 0, 2, 1, 1, 1, 1, 1, 1, 0, 1, 2, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -3, -1, -1, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 2, 1, 2, 2, 0, 1, 1, 2, 2, 3, 1, 1, 0, 0, -1, -1, 0, -1, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, -1, -2, -1, -2, -2, -2, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -2, 0, -1, 0, -1, 1, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, -2, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, -2, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, -2, -1, -2, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, -2, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, -2, -1, -1, 0, -2, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, -1, -1, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -3, -3, -3, -4, -2, -3, -3, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, -2, -4, -4, -5, -4, -3, -5, -4, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, -2, -4, -3, -5, -3, -3, -3, -2, -1, 0, 0, 1, 1, 3, 2, 2, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -4, -4, -3, -4, -4, -1, -2, 0, 0, 0, 1, 3, 2, 4, 2, 2, 3, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -3, -4, -3, -4, -2, -2, -2, -2, 0, 2, 1, 1, 3, 3, 3, 3, 3, 3, 1, 2, 2, 1, 0, 1, 1, 1, 0, 0, 0, 0, -2, -2, -3, -4, -2, -3, -3, -2, -1, -1, 0, 1, 2, 2, 1, 2, 2, 2, 1, 3, 2, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, -2, -2, -2, -3, 0, -1, -1, 0, -1, -1, 0, 1, 1, 2, 1, 2, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, -1, -1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 1, 2, 0, 1, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 2, 2, 2, 2, 0, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 1, 2, 2, 1, 1, 1, 1, 1, 2, 3, 2, 3, 2, 0, -1, 0, 0, 0, 1, 1, 1, 2, 2, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 2, 2, 2, 1, 3, 4, 5, 3, 1, -1, 0, 0, 0, 0, 0, 3, 1, 2, 2, 0, 0, 0, -1, -1, -1, -2, -3, 0, 0, 0, -1, 1, 2, 2, 1, 2, 5, 4, 4, 1, 0, 0, 0, 0, 0, 0, 1, 2, 3, 3, 4, 3, 2, 0, -1, -1, -3, -3, -3, -3, -2, -3, -2, -1, 0, 0, 2, 2, 4, 4, 5, 1, 0, -2, 0, 0, 0, 0, 0, 2, 3, 4, 4, 3, 3, 1, -1, -2, -3, -5, -6, -5, -5, -5, -4, -4, -1, 0, 1, 3, 4, 4, 4, 1, 0, 0, 0, -1, 0, 0, 1, 2, 2, 3, 6, 6, 4, 2, 0, -2, -3, -4, -7, -7, -5, -6, -5, -6, -2, -1, 0, 1, 3, 2, 3, 0, 0, -2, 0, -1, 0, 0, 1, 3, 4, 4, 5, 4, 4, 3, 1, -1, -4, -5, -7, -6, -7, -7, -7, -6, -4, -1, 0, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, 1, 1, 1, 4, 5, 6, 6, 5, 2, 1, -1, -3, -5, -7, -7, -7, -6, -7, -6, -2, -1, 0, 1, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 2, 3, 5, 4, 5, 3, 2, 0, -2, -4, -5, -6, -5, -6, -5, -4, -5, -3, -1, 0, 2, 2, 4, 2, 1, 0, -1, 0, -1, 0, 0, 0, 2, 4, 6, 6, 4, 4, 2, 0, -3, -3, -4, -3, -4, -4, -4, -2, -3, -1, 0, 1, 1, 2, 3, 3, 1, 0, 0, 0, 0, 0, 1, 1, 2, 4, 4, 6, 3, 4, 2, 0, -2, -4, -4, -3, -4, -2, -3, -2, 0, -1, 0, 2, 3, 3, 3, 3, 0, 0, 0, 0, -1, 0, 1, 2, 2, 4, 5, 3, 4, 3, 1, 1, 0, -2, -1, -1, -1, -1, -2, -1, -1, 0, 1, 0, 1, 1, 3, 4, 1, 0, -1, 0, 0, 1, 2, 2, 3, 2, 3, 3, 4, 2, 1, 0, -1, -1, 0, -1, -1, -2, -1, 0, 0, 0, 1, 0, 3, 2, 2, 3, 2, 0, 0, 0, 0, 1, 2, 3, 2, 3, 3, 3, 3, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 4, 3, 2, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 2, 2, 3, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 3, 3, 2, 2, 0, 0, 0, 0, 0, 1, 2, 2, 1, 2, 0, 2, 1, 1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 2, 1, 2, 1, 2, 2, 3, 2, 2, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 1, 1, 2, 3, 2, 1, 2, 1, 2, 3, 2, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 1, 2, 2, 1, 2, 2, 2, 1, 1, 1, 2, 1, 1, 0, 0, -2, -2, -2, -1, 0, -3, -2, -2, -1, 0, 0, 1, 1, 1, 0, 1, 1, 2, 3, 1, 3, 2, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, -2, -2, -2, -3, -2, -2, -2, -3, -3, -1, 0, 1, 2, 2, 2, 1, 3, 3, 3, 2, 2, 2, 0, -1, -1, 0, -1, 0, 0, 0, 0, -2, -1, -2, -4, -3, -3, -2, -2, -2, -2, -2, -1, 0, 1, 1, 1, 0, 1, 1, 2, 1, 2, 0, -2, -3, -2, -1, -1, -1, -1, 0, -1, -1, -2, -2, -2, -2, -2, -2, -3, -3, -2, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, -2, -2, -1, -3, -2, -1, -1, 0, -2, 0, -1, -1, 0, -1, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -2, 0, 0, 0, -1, 2, 3, 0, 1, 2, 1, 1, 1, 1, 0, 0, 0, 1, 3, 2, 2, 2, 2, 2, 0, 2, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 2, 3, 3, 2, 1, 2, 1, 3, 2, 0, 1, 2, 1, 3, 3, 2, 1, 2, 2, 1, 2, 1, 0, 1, 0, 0, -1, 0, -1, 0, 1, 0, 2, 1, 3, 1, 1, 1, 1, 2, 2, 2, 0, 1, 2, 2, 2, 1, 1, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 2, 3, 2, 2, 3, 3, 1, 2, 1, 3, 3, 1, 2, 2, 1, 2, 1, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, 1, 2, 2, 2, 2, 2, 1, 1, 1, 1, 3, 3, 3, 2, 1, 2, 2, 1, 2, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 3, 1, 1, 2, 2, 2, 2, 2, 2, 2, 0, 3, 3, 3, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 2, 2, 2, 1, 2, 1, 2, 1, 2, 2, 3, 1, 1, 0, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 2, 0, 2, 0, 1, 2, 2, 1, 2, 1, 2, 2, 1, 0, 2, 2, 2, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 2, 1, 0, 1, 0, 1, 0, 0, 0, 2, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 2, 2, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 3, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -2, -1, -2, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -2, -2, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -3, -1, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -3, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -1, -1, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 2, 2, 2, 1, 1, 1, 1, 1, 1, 0, -1, -1, 0, -1, 0, -1, -2, -3, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 2, 1, 2, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 1, 2, 2, 2, 2, 2, 1, 2, 0, 2, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 3, 2, 1, 2, 1, 1, 2, 2, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 3, 3, 3, 1, 0, 0, 2, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 2, 0, 1, 2, 1, 1, 1, 2, 1, 1, 1, 2, 2, 0, 1, 1, 0, 2, 0, -1, 0, 0, 1, 1, 1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 3, 2, 2, 3, 1, 1, 1, 2, 2, 3, 2, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 1, 1, 2, 2, 1, 2, 2, 2, 1, 3, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 3, 2, 0, 2, 2, 1, 1, 1, 2, 3, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 2, 1, 1, 2, 3, 1, 3, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 2, 2, 1, 2, 1, 1, 0, 2, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 1, 2, 1, 3, 3, 3, 2, 0, 1, 1, 0, 1, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -2, -3, -2, -2, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 2, 1, 0, 0, 0, -1, -2, 0, -1, -1, -3, -2, -2, -2, -2, 0, -1, 0, 1, 1, 0, 0, 0, 1, 0, 1, 2, 1, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -4, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 1, 1, 1, 1, 1, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, -1, -2, 0, -2, -1, -1, 0, 0, 0, 0, 1, 1, 2, 1, 3, 2, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 2, 3, 1, 1, 2, 0, 1, 0, 0, 0, 1, 1, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 2, 1, 3, 2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -2, -1, -1, 0, 0, 1, 0, 1, 2, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -3, -2, 0, 0, 0, 0, 0, 2, 1, 1, 2, 2, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -4, -3, -3, -2, 0, 0, 0, 0, 2, 2, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, -1, -2, -4, -4, -3, -3, -2, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, -2, 0, -1, 0, 0, -1, -1, -1, -1, -3, -3, -5, -3, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, -1, -3, -2, -4, -4, -5, -4, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -2, -1, 0, 0, -1, 0, 0, -1, -1, -3, -4, -5, -6, -5, -3, -3, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, -1, -1, -2, -3, -1, -4, -4, -6, -5, -5, -3, -2, -2, -2, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, -1, 0, -1, -1, -1, -2, -3, -5, -6, -6, -4, -4, -2, -3, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, -3, -5, -6, -5, -4, -2, -2, -1, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -2, -1, -3, -4, -5, -4, -3, -2, -2, -3, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, -2, -1, -4, -3, -3, -3, -3, -1, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -3, -3, -4, -3, -2, -2, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -2, -1, -2, -1, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -3, -3, -2, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, -1, -2, -1, 0, -1, -1, -1, -1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -3, -2, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, -3, -2, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, -1, -2, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -3, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -2, -2, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 1, 2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -2, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, -2, 0, 0, 2, 0, 0, 1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 1, 1, 0, 2, 1, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -2, 0, 1, 1, 0, 1, 1, 1, 2, 1, 0, 0, 0, -1, -2, 0, -1, -1, -2, -1, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 1, 2, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 2, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 1, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -1, -1, -1, -2, -1, -1, -1, 0, 0, -1, -2, -2, -2, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -3, -2, -2, -1, -1, -1, 0, -1, 0, -1, 0, 0, -1, -1, -3, -2, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, -2, -2, -1, -1, -3, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 1, 0, -1, -1, -1, -2, -1, -2, -2, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 0, 1, 1, 0, 0, 1, 0, 0, 1, 3, 3, 0, 0, -1, -2, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 1, 0, 1, 0, 0, 1, 0, 0, 2, 4, 3, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 2, 0, 2, 0, 2, 0, 2, 1, 1, 2, 3, 1, 0, 0, -2, -1, -2, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 2, 2, 1, 1, 1, 1, 1, 1, 3, 3, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 2, 3, 3, 2, 1, 1, 0, 1, 1, 0, 0, 1, 2, 1, 1, -1, -1, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 2, 1, 0, 0, 0, 0, 0, 2, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 1, 2, 3, 2, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 2, 3, 3, 1, 3, 3, 1, 0, -1, 0, 0, 0, 1, 2, 2, 2, 1, 0, -1, 0, 0, 0, 0, 0, 1, 1, -1, 0, -1, 0, 0, 1, 1, 2, 2, 2, 3, 3, 1, 0, 0, 0, 0, 1, 2, 4, 4, 2, 1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 3, 3, 3, 2, 2, 0, 0, 0, 1, 2, 1, 3, 3, 3, 3, 0, -1, 0, -2, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 2, 1, 1, 1, 0, 1, 0, 2, 1, 2, 4, 3, 4, 2, 1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 4, 3, 2, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 2, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 2, 3, 2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 2, 2, 4, 2, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 1, 3, 2, 0, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 3, 4, 2, 1, 0, 0, 1, -1, -1, -1, 0, 0, 0, 2, 3, 2, 1, 0, -1, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 1, 2, 3, 3, 4, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 2, 1, 1, 0, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, 1, 1, 0, 2, 2, 3, 3, 3, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 4, 3, 2, 0, 0, -1, 0, -1, 0, 0, 0, -2, -1, -2, 0, 0, 1, 1, 1, 3, 4, 4, 1, 1, 0, 0, 2, 1, 1, 0, 0, 0, 4, 4, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, 1, 1, 0, 2, 3, 5, 3, 2, 0, 0, 1, 3, 2, 2, 0, 0, 1, 4, 4, 1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 2, 2, 3, 2, 2, 0, 0, 1, 2, 2, 1, 2, 1, 1, 3, 3, 3, 0, 0, 0, 2, 1, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 2, 1, 2, 3, 2, 0, 0, 0, 3, 1, 1, 0, 1, 0, 3, 3, 2, 0, -1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 3, 2, 2, 2, 0, 0, 1, 2, 1, 0, 1, 0, 2, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 2, 2, 1, 2, 3, 0, 1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 2, 0, -2, 0, 0, 1, 0, -2, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 2, 2, 2, 1, 1, 1, 2, 1, 2, 2, 0, 0, 1, 2, 0, -1, 0, 0, 0, -1, -1, -3, -3, -1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 2, 0, 1, 0, 0, 0, 1, 1, 1, 2, 0, 0, 0, 0, -2, 0, 1, 0, -1, -4, -3, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, -1, 0, 2, 1, 1, 0, 1, 1, -1, -1, 0, 0, -1, -2, -3, -2, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 2, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 2, 3, 3, 1, 1, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 1, 1, 2, 1, 1, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, -2, 0, -2, 0, 0, 0, -1, -1, 0, 0, 0, -1, -2, -1, 1, 1, 0, 1, 3, 2, 2, 2, 0, 0, 0, 0, -1, 0, -2, -1, -1, -2, -2, -3, -2, -1, 0, 0, 0, -2, -1, 0, 0, 0, -2, -1, 2, 1, 0, 2, 2, 1, 0, 2, 0, 0, 0, 0, 0, -1, -2, 0, -1, -2, -3, -2, -3, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 3, 1, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, -2, -2, -3, -3, -1, 0, 0, 0, -1, 0, -1, 0, -1, -2, -2, 2, 3, 0, 1, 2, 1, 0, -1, 0, 0, 0, 0, -1, -1, -3, -1, -1, -1, -3, -3, -2, 0, 1, 1, 1, -1, 0, 0, 0, 0, -2, 0, 1, 1, 2, 1, 0, 0, 0, -1, 0, -1, -3, 0, -1, -1, -3, -2, -1, 0, -1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, -1, -1, 1, 2, 2, 0, 0, -1, -1, -1, -1, -3, -2, -2, -1, -1, -1, -1, -2, 0, -1, 0, -1, -1, 0, 0, 0, 0, -2, 0, 1, 0, -1, -1, 2, 2, 1, 0, -1, -2, -1, -1, 0, -2, -2, -1, -2, -1, 0, 0, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 3, 1, 1, -1, -2, 0, -2, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, -2, -1, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, -2, -1, 2, 1, 0, 0, -1, -2, -2, -1, -2, -2, -2, -1, -1, -1, -1, 0, 1, 0, -1, -1, -1, -2, -2, -1, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, -1, -1, -2, -2, -2, -1, -2, -4, -3, 0, 1, 0, 0, 0, 1, 2, 1, -2, -3, -3, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 2, 0, 0, -2, -4, -2, -3, -3, -2, -4, -3, 0, 2, 1, 0, 1, 3, 4, 2, 1, -1, -2, 0, 0, 0, 0, 1, 0, 1, 1, 0, -1, 1, 0, 0, -1, -3, -2, -2, -2, -2, -4, -4, -3, 0, 0, 0, 0, 3, 5, 4, 4, 3, 1, 0, 1, 1, 0, 0, 0, 1, 1, -1, 0, 2, 0, -1, -1, -2, -1, -1, -2, -2, -3, -3, -3, 0, 0, 0, 0, 2, 3, 5, 3, 3, 2, 1, 2, 1, 0, 0, 1, 2, 0, 0, 0, 1, 1, -1, -2, -2, -2, -2, -2, -1, -1, -3, -3, -1, 1, 0, 0, 1, 1, 3, 2, 3, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 2, 0, -1, 0, -3, -3, -3, -2, -2, -1, -2, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 2, 0, -1, -2, -2, -5, -4, -5, -2, -1, -1, -2, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 3, 1, 0, 0, -3, -2, -4, -4, -3, -1, -2, -3, -2, -1, 0, 0, 0, 0, -1, -1, -1, -2, 0, 0, -2, -1, -1, 0, 0, 0, -1, 0, 3, 1, 0, 0, -1, -1, -2, -3, -3, -2, -1, -2, -2, -2, 0, 0, 0, 0, 0, 0, -1, -3, -1, -1, -3, -2, -2, 0, -1, -1, 0, 0, 3, 0, 0, 0, -2, -1, -3, -2, -2, 0, -2, -1, -1, -1, 0, 1, 0, -1, -1, 0, 0, -1, -1, 0, -1, -2, 0, 0, -1, 0, -1, 0, 1, 0, -1, -2, -1, -1, -2, -2, -2, 0, -2, -1, 0, -3, -1, 1, 1, -1, -2, 0, 0, -1, -1, 0, -1, -3, -1, 0, 0, 0, 0, 0, 2, 1, -1, -1, -2, -1, -2, -2, -3, -2, -2, -1, 0, -3, -2, 0, 1, -1, -2, -2, 0, 0, 0, 0, -2, -3, -1, -1, 0, 0, 0, 0, 2, 1, -1, 0, 0, -1, -2, -1, -3, -2, -2, 0, 0, -2, -1, 0, 0, 0, -1, -2, -1, 0, 0, -1, 0, -2, -3, 0, -1, -1, -1, -1, 3, 1, 0, 0, -1, -2, -2, -2, -2, -3, -2, -1, 0, 0, -1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, -1, 3, 3, 0, 0, 0, -1, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, -2, -2, -1, -2, -1, 0, -1, -2, -2, -1, 0, 0, 0, 4, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, -1, -1, 0, -2, -2, -1, -2, -3, -3, 0, -2, -1, 0, 0, 0, 0, 0, 4, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -3, -2, 0, 0, -1, -1, -2, -1, -2, -1, -1, -2, -2, 0, -2, -2, -1, 0, 0, 0, -1, 4, 2, 0, 0, 0, 0, 1, 1, 0, 0, -2, -3, -2, 0, 0, 0, -2, -3, -2, -1, -1, -2, -4, -3, -1, 0, -2, -1, 0, -1, 0, -1, 4, 2, 0, 0, 1, 0, 0, 1, 2, 1, 0, -2, 0, 0, 0, -1, -1, 0, -1, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 2, 5, 4, 2, 1, 0, 0, 3, 4, 4, 1, 0, 0, 2, 0, 0, 1, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 1, 3, 4, 3, 1, 0, 0, 1, 2, 3, 2, 0, 0, 1, 1, 2, 3, 1, 1, 1, 1, 1, 1, 2, 3, 2, 3, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -2, -1, 0, 0, 0, -1, -3, 0, 0, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 3, 0, 1, 0, 0, 0, 0, 0, -1, -2, 0, -1, -1, -1, 0, 0, 0, -2, -2, -1, -2, -2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 4, 5, 0, 1, 0, 1, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, -3, -1, -2, -2, -2, -1, 0, -1, -2, -1, 0, 0, -1, 0, 4, 4, 0, 0, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, -3, -4, -2, -1, 0, -1, -3, -2, 0, 0, -1, 0, 3, 3, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -3, -3, -4, -3, -3, 0, 0, -1, -1, -2, -1, -2, -1, 0, 2, 2, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -2, 0, 0, 0, 0, -2, -4, -3, -3, -3, -1, 0, 0, -2, -2, 0, -1, -1, -3, 0, 1, 0, 1, -1, -2, 0, -1, -1, -2, 0, 0, 0, -2, 0, 1, 0, 0, -2, -2, -3, -3, -4, -1, -1, -2, -4, -3, -1, -1, 0, -2, 0, 1, 0, 0, -1, -2, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 1, 0, -2, -2, -3, -3, -5, -2, -2, -3, -3, -3, -1, -1, -1, -2, 0, 1, 0, 0, 0, -2, -2, -1, -1, -1, 0, 0, -1, -1, -1, 0, 0, -2, -3, -4, -1, -2, -3, -4, -4, -2, -4, -3, -3, -2, -2, 0, -1, 0, 0, 0, 0, -1, -3, -3, -1, -3, -2, 1, 0, 0, 0, 0, 0, -1, -3, -3, -1, -3, -4, -3, -3, -3, -3, -3, -3, -2, -2, -1, 0, 1, 0, 1, 0, -3, -4, -4, 0, -2, -2, 0, 0, 0, 0, 0, 0, -2, -4, -3, -2, -3, -2, -2, -4, -4, -4, -4, -2, -3, -1, 0, 0, 0, 0, 1, 0, -2, -3, -3, -1, -1, -4, -2, -1, 0, 0, 1, 0, -1, -3, -3, -4, -3, -3, -3, -4, -4, -4, -4, -3, -3, -3, -2, 0, 0, 0, 1, 0, -4, -5, -4, -2, -3, -4, -4, -1, 0, 0, 0, 1, 0, -2, -4, -4, -4, -3, -4, -3, -3, -3, -4, -4, -2, -2, -1, 0, 1, 0, 2, 0, -3, -5, -3, -3, -4, -4, -4, -2, -1, 0, 1, 0, 0, 0, -4, -2, -2, -3, -4, -3, -5, -4, -4, -3, -3, -3, -1, 1, 0, 0, 0, 0, -2, -4, -2, -4, -5, -4, -4, -4, 0, 0, 0, -1, 0, -2, -4, -4, -3, -5, -3, -3, -4, -4, -5, -3, -4, -2, 0, 1, -1, 0, 0, 0, -1, -4, -3, -4, -4, -5, -5, -2, 0, 2, 1, -1, 0, -2, -5, -3, -3, -3, -3, -3, -4, -4, -5, -5, -5, -3, 0, 2, 0, 0, 0, 0, -1, -2, -3, -4, -4, -3, -4, -3, 0, 3, 2, 0, -1, -3, -4, -3, -3, -3, -3, -3, -5, -3, -4, -5, -4, -2, 0, 1, -1, -1, 0, 0, -2, -3, -4, -6, -4, -3, -3, -3, 0, 1, 4, 1, -2, -2, -5, -3, -2, -3, -2, -4, -4, -5, -4, -5, -3, -3, 0, 3, 0, 0, 0, 0, -3, -1, -3, -5, -3, -2, -3, -3, -2, 1, 4, 1, -1, -3, -5, -1, -2, -3, -1, -3, -3, -4, -3, -3, -4, -3, 0, 2, 0, 0, 0, 0, -2, -2, -3, -5, -3, -1, -2, -1, -3, 0, 4, 0, -2, -3, -4, 0, -1, -3, -1, -1, -4, -3, -1, -2, -4, -3, -2, 1, 0, 0, 1, 0, -2, -2, -3, -3, -3, 0, -3, -1, -2, 0, 4, 0, -1, -1, -2, 0, 0, -2, -2, -1, -2, -1, 0, 0, -1, -3, -1, 0, 0, 0, 1, 0, -3, -2, -2, -2, -2, -1, -2, -2, -2, 0, 3, 1, 0, 0, -3, 0, 0, -2, -3, -2, -3, -4, -1, -1, -1, -2, -1, 0, 0, 0, 1, -2, -1, -2, -2, -2, -2, -1, -1, -1, -3, 0, 1, 1, 0, 0, -1, -1, 1, 0, -2, -1, -4, -4, -1, -1, -1, 0, 0, -1, 0, 0, 1, 0, -3, -1, -1, -3, -2, -1, -2, -1, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -4, -3, -2, -1, -2, 0, 0, 1, -1, 0, 0, -2, -3, -2, -2, -3, -3, -1, 0, -2, -1, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -3, -2, -3, -2, -1, 0, 0, 0, -2, 0, 0, -1, -2, -2, -1, -1, -2, -1, -1, -2, -2, -2, -3, -1, -1, 0, -2, -2, -1, -2, -1, 0, -2, -2, -1, 0, 0, 0, 0, 0, -2, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, -2, -1, -3, -3, -2, 0, -1, -2, -1, -2, 0, 0, -1, -1, -1, -2, 0, 0, 1, 1, -1, 0, 1, -2, -3, 0, 0, -1, 0, -2, -2, 0, -2, -1, -2, -3, -2, 0, -2, -2, -2, -2, 0, 0, -1, 0, -1, -2, -2, 0, 0, 2, 0, 0, 0, 0, -2, -1, 0, 0, 1, -1, -1, -1, -2, -1, -3, -1, -1, 0, 0, -3, -3, -2, 0, -1, -2, -1, 0, -1, 0, 0, 0, 2, 0, 0, 0, 0, -2, -2, 0, 1, 1, 0, -1, -2, -1, 0, -1, -2, -1, 0, -1, -2, -1, -1, 0, 0, 0, 0, -1, 0, -2, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -2, -2, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, -1, 0, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -2, -1, -3, -3, -2, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -3, -2, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, -2, -1, -1, -2, -3, -2, 0, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -2, -2, -2, -1, -2, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -2, -2, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 2, 2, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 2, 0, 1, 1, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 2, 2, 1, 1, 2, 2, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 2, 0, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 1, 2, 1, 2, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 2, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 2, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, -2, -1, -2, -2, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, -2, -1, -2, -2, -2, -1, -2, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -2, -2, -2, -1, -2, -1, -2, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -3, -3, -2, -2, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 1, 1, 1, 0, 1, 1, 1, -1, 0, 0, 0, 0, -1, -2, -2, -2, -3, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, -2, -2, -1, -2, -2, -2, -1, -1, -1, -1, 0, -1, -1, -1, -1, 0, -1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -2, -2, -3, -2, -1, -2, -1, -1, -1, -1, 0, -2, -2, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, -2, -1, -2, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 2, 1, 1, 1, 0, 0, 0, -1, 0, -2, -2, -1, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 2, 1, 1, 2, 1, 1, 0, 0, 0, -1, -1, -2, -2, -1, -1, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 2, 2, 2, 2, 1, 1, 1, 0, 0, 0, 0, -2, 0, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 2, 1, 2, 0, 2, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 2, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -4, -3, -3, -4, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, 0, -1, -3, -3, -3, -3, -3, -4, -2, -3, -1, 0, 0, 0, 1, 1, 3, 2, 2, 3, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, -3, -3, -1, -1, -1, -2, -1, 0, 0, 1, 1, 2, 3, 3, 2, 4, 2, 2, 2, 3, 1, 2, 1, 0, 0, 1, 0, 1, 3, 1, 0, -1, -4, -3, -2, -1, -2, -1, 0, 0, 0, 0, 0, 1, 3, 4, 2, 2, 3, 3, 3, 3, 1, 2, 1, 1, 0, 1, 0, 1, 1, 0, -1, -1, -4, -4, -3, -1, -2, 0, 0, 0, 0, 0, 1, 2, 2, 3, 3, 2, 3, 3, 2, 2, 2, 1, 2, 1, 2, 1, 1, 0, 1, 0, 0, -2, -4, -3, -1, -2, -1, -1, -1, -1, 0, 1, 1, 2, 1, 1, 2, 2, 2, 3, 3, 1, 1, 2, 2, 2, 1, 0, 0, 1, 2, 0, 0, -1, -1, -1, -1, 0, -2, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 2, 2, 2, 1, 1, 0, 1, 2, 1, 1, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 1, 2, 2, 0, 2, 2, 2, 3, 1, 3, 3, 2, 0, -1, -2, -1, 0, 2, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 2, 3, 2, 3, 2, 2, 2, 2, 3, 3, 3, 3, 3, -1, -1, -1, 0, 0, 1, 2, 2, 1, 2, 1, 0, 0, -1, 0, -1, 0, 0, 0, 2, 2, 2, 3, 4, 2, 3, 3, 3, 4, 5, 4, 1, -1, -1, -1, 0, 0, 1, 1, 2, 2, 0, 1, 0, 0, 0, -2, -1, -1, 0, 0, 1, 0, 1, 1, 2, 3, 3, 3, 3, 4, 5, 3, 2, 0, 0, -2, -1, 0, 1, 2, 1, 1, 2, 2, 0, -1, -1, -2, -3, -2, -2, -1, 0, 0, 0, 0, 1, 2, 2, 4, 3, 4, 3, 3, 0, -1, 0, -2, 0, 0, 0, 1, 2, 2, 2, 1, 0, 0, -1, -2, -3, -3, -3, -1, -1, -1, 0, 1, 2, 2, 3, 4, 3, 3, 4, 3, 1, -1, 0, 0, 0, 0, 0, 1, 2, 3, 4, 2, 2, 0, -1, -4, -4, -4, -4, -4, -4, -3, -1, -1, 0, 1, 2, 3, 2, 2, 3, 1, 0, -1, 0, -1, -1, 0, 0, 1, 3, 2, 3, 2, 1, 1, -2, -3, -4, -6, -6, -5, -6, -4, -4, -4, -1, 0, 1, 2, 2, 1, 3, 2, 0, 0, 0, 0, 0, 0, 0, 1, 2, 4, 4, 3, 3, 1, -2, -3, -4, -5, -5, -6, -4, -4, -4, -3, -2, -1, 0, 0, 1, 1, 3, 3, 0, -1, -1, 0, 0, 0, 0, 2, 3, 5, 3, 4, 2, 1, -1, -4, -4, -4, -6, -5, -4, -6, -5, -3, -1, 0, 0, 2, 2, 2, 4, 3, 0, -1, 0, -1, 0, 0, 2, 2, 4, 3, 5, 3, 2, 0, -1, -3, -4, -4, -5, -5, -5, -4, -3, -2, -1, 0, 2, 2, 3, 3, 2, 2, 0, -1, 0, -1, 0, 0, 0, 2, 4, 5, 4, 3, 1, 0, 0, -3, -5, -3, -3, -3, -3, -1, -2, -1, 0, 1, 3, 2, 2, 2, 2, 2, 2, -1, 0, -2, 0, 0, 1, 3, 3, 5, 3, 3, 2, 0, 0, -2, -4, -2, -1, 0, -1, -2, -2, 0, 0, 1, 2, 3, 2, 2, 2, 3, 2, 0, -1, 0, 0, 2, 2, 2, 3, 3, 2, 1, 0, 0, 0, -2, -3, -1, -2, -1, -1, -1, 0, 0, 1, 2, 3, 3, 3, 2, 3, 3, 1, 0, -1, 0, 0, 2, 3, 2, 4, 3, 3, 3, 1, 0, 0, -1, -2, -1, -2, -2, -1, -1, -1, 0, 0, 1, 1, 1, 2, 1, 2, 2, 0, -1, -1, -1, 0, 1, 3, 3, 2, 2, 4, 3, 1, 1, 0, -1, -1, -2, -1, -1, 0, 0, 0, 1, 0, 0, 1, 2, 2, 2, 3, 3, 1, -1, 0, -1, 0, 1, 2, 1, 2, 2, 1, 2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 3, 3, 1, 3, 3, 1, 0, 0, -1, 0, 0, 1, 2, 2, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 2, 2, 1, 0, 1, 2, 2, 3, 1, 1, 2, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 2, 2, 2, 1, 2, 3, 2, 3, 3, 2, 2, 2, 0, 0, -1, -2, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 2, 1, 2, 2, 1, 2, 3, 2, 0, 0, 0, -1, -3, -2, -2, -2, -3, -1, 0, 0, 0, 0, 1, 1, 0, 2, 3, 2, 2, 2, 3, 2, 1, 1, 1, 0, 0, 1, 2, 1, 1, 0, 0, -2, -4, -4, -2, -3, -2, -1, -2, -1, 0, 0, 2, 2, 1, 1, 2, 2, 2, 3, 3, 2, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, -1, -2, -5, -3, -2, -1, -1, -1, -2, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 2, 2, 0, 1, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, -2, -4, -3, -1, 0, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 1, 1, 1, 1, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 1, 2, 0, 1, 2, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 2, 1, 2, 2, 1, 1, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 0, 0, 0, -2, -2, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 1, 1, 1, 3, 2, 1, 1, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 2, 2, 1, 3, 2, 2, 0, 0, 0, -1, -1, -2, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 2, 1, 1, 0, 0, 0, -1, 0, -2, 0, -1, 0, 0, -1, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 1, 2, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 2, 1, 1, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, -1, -3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -2, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, -2, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, -2, -2, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, -2, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, -2, 0, 0, 0, -1, -1, -2, -1, 0, -1, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -2, -1, 0, 0, -1, -2, -2, 0, -1, -1, 0, -1, -1, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -2, -1, -1, -1, -2, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -2, -1, 0, 0, 0, 0, -1, -1, -1, 0, -2, -1, -2, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, -2, -1, -1, -1, -1, -1, 0, 1, 0, -1, -1, -1, -2, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -2, 0, -1, -2, -2, -2, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -2, -2, -1, -1, -1, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, -2, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, -1, -1, 0, 0, -1, 0, -1, -2, -2, -1, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, -2, -1, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, -2, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -2, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 2, 3, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 1, 2, 0, 1, 1, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, -1, 0, 0, 0, 1, 1, 1, 1, 2, 3, 2, 1, 2, 1, 4, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 1, 2, 2, 1, 2, 3, 2, 1, 1, 2, 3, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 2, 2, 2, 3, 3, 2, 2, 2, 2, 2, 2, 2, 3, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 2, 0, 0, 0, 0, 1, 1, 3, 4, 3, 3, 3, 3, 1, 1, 3, 3, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 1, 0, 1, 1, 0, 2, 2, 2, 2, 4, 3, 1, 2, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 1, 2, 1, 2, 2, 2, 2, 1, 2, 1, 2, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 2, 1, 2, 1, 1, 1, 1, 0, 2, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 0, 1, 0, 0, 1, 2, 2, 3, 2, 1, 0, 2, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 2, 1, 2, 1, 0, 1, 0, 0, 1, 1, 3, 1, 1, 0, 0, -1, -1, -2, 0, -1, -3, -2, 0, -1, 0, 0, 0, 1, 2, 1, 3, 2, 3, 2, 1, 1, 0, 1, 1, 1, 0, 1, 3, 2, 1, 0, 1, 0, -2, -1, -1, -2, -3, -2, -1, -1, 0, 0, 0, 0, 2, 2, 3, 2, 3, 3, 1, 2, 2, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -2, -3, -3, -2, -1, 0, 0, 1, 0, 0, 2, 1, 2, 3, 2, 1, 1, 2, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, -3, -3, -3, -2, -1, 0, 0, 0, 2, 2, 2, 2, 2, 2, 1, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, -3, -3, -4, -3, -2, 0, -1, 0, 0, 2, 4, 3, 3, 2, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -3, -3, -2, -1, 0, 1, 1, 4, 4, 4, 4, 3, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -2, -3, -3, 0, 0, 0, 1, 2, 3, 3, 4, 4, 2, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, -2, -1, -2, -2, -1, 0, 0, 1, 2, 2, 5, 5, 3, 3, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, -2, 0, 0, -2, -2, -1, -1, 1, 2, 1, 2, 4, 6, 6, 4, 2, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 1, 3, 2, 2, 4, 5, 7, 4, 2, 1, 0, 1, 3, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -2, 0, -2, -2, -1, -1, 0, 2, 2, 2, 2, 3, 4, 6, 5, 2, 1, 0, 1, 1, 2, 2, 1, 0, 0, 1, 0, -1, -1, -1, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 1, 2, 3, 4, 5, 4, 4, 4, 2, 1, 0, 1, 2, 2, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, 1, 3, 3, 3, 4, 4, 4, 3, 1, 1, 2, 2, 2, 3, 2, 2, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 2, 3, 2, 2, 2, 1, 1, 1, 2, 3, 1, 2, 2, 0, 0, -1, 0, -1, -1, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 1, 1, 3, 2, 1, 2, 1, 2, 1, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 2, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, -1, -1, -1, -1, -2, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, 0, 0, -1, -2, -3, -2, -2, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -2, -1, 0, 0, -2, -1, -3, -1, 0, -1, -1, -1, -2, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 2, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -2, 0, -1, -2, -1, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -2, -2, -1, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, -1, -1, -1, -1, -2, -2, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 2, 1, 1, 2, 1, 2, 1, 1, 1, 1, 0, -1, 0, -2, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 2, 1, 1, 2, 1, 0, 0, 0, 1, 0, 1, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 2, 2, 1, 0, 0, 1, 1, 0, 0, 1, 0, -1, 0, 0, -2, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 2, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 1, 0, 2, 1, 1, 0, 2, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 1, 1, 1, 0, 2, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, -1, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 2, 1, 1, 0, 0, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, -1, -2, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 2, 3, 2, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 1, 1, 0, 1, 0, -1, 0, -1, -2, -1, -1, -1, 0, 0, 0, 0, 1, 2, 2, 2, 1, 2, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, -2, -2, -3, -1, -2, -2, -3, -2, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -3, -1, -1, -3, -2, -2, -3, -2, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 1, 2, 0, 0, 0, -1, -2, -2, -2, -3, -3, -2, -1, -2, -1, 0, 0, 1, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 1, 0, 0, 0, -1, -3, -2, -2, -3, -3, -1, -2, 0, 0, 1, 1, 2, 2, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -2, -2, -1, -3, -2, -2, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, -1, 0, -1, -1, -1, -1, -1, -1, 0, 0, 1, 1, 2, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 1, 2, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, 1, 2, 0, 2, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 0, 2, 1, 0, 2, 1, 1, 1, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 1, 1, 1, 0, 2, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, -1, 0, -1, -1, -1, -2, -1, -1, -1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -2, 0, -2, -1, -2, -2, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -2, -2, -2, -1, -1, -2, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -3, -2, -3, -1, -1, -1, -1, -3, -3, -1, -2, -1, -1, 0, 0, 0, 0, 0, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, -2, -2, -4, -3, -3, -1, -1, 0, -1, -2, -2, -2, -1, 0, 0, 0, 2, 3, 3, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -2, 0, 1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 3, 4, 2, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 2, 2, 1, 0, 0, 0, 1, 2, 0, -1, -2, 0, 1, 0, 0, 1, 4, 6, 3, 0, 0, 0, 0, 1, 0, 1, 1, 0, -2, -2, -2, -1, 0, 1, 2, -1, -1, 0, 0, 1, 0, 0, -1, 0, 2, 1, 0, 2, 3, 6, 2, 0, -2, 0, 0, 0, 0, 0, 1, 0, -2, -3, -2, -4, -1, 0, 1, 0, -1, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 1, 3, 7, 3, -1, 0, -1, 0, 1, 0, 0, 0, 0, -1, -1, -1, -4, -3, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 2, 1, 1, 2, 3, 6, 3, 0, -1, 0, 1, 1, 1, 0, -1, -1, 0, 0, -1, -2, -2, -1, 0, 0, 1, 2, 2, 0, 1, 0, 0, 1, 0, 2, 1, 2, 3, 6, 5, 0, -1, -1, 2, 4, 3, 0, -1, -1, 0, -1, -1, -3, -2, 0, -1, 0, 1, 3, 2, 3, 1, 0, -1, 0, 0, 0, 1, 4, 5, 7, 6, 0, 0, 0, 1, 2, 3, 0, -1, 0, 0, -1, -3, -3, -2, -1, 0, 0, 1, 4, 4, 3, 1, 1, -1, -3, -2, 0, 1, 4, 6, 9, 6, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -4, -4, -3, -2, 0, 3, 2, 4, 4, 4, 2, 0, -1, -3, 0, 1, 2, 5, 8, 9, 7, 0, -1, 0, 1, 0, 0, 0, -1, 1, 1, 0, -4, -4, -3, -1, 2, 3, 5, 6, 6, 5, 4, 2, -2, -3, 1, 1, 3, 4, 7, 10, 7, 0, 0, -1, 0, -1, 0, -2, -1, 0, 0, 0, 0, -2, -2, 0, 3, 3, 4, 6, 6, 5, 5, 3, 0, 0, 1, 3, 4, 6, 7, 9, 8, 1, -1, 0, 0, -1, -2, -1, 0, 0, 1, 1, 0, 0, -1, 0, 2, 2, 3, 2, 5, 4, 4, 2, 1, 1, 2, 3, 4, 5, 6, 9, 8, 1, 0, 0, 0, -2, -3, -3, 0, 0, 2, 3, 2, 0, 1, 2, 3, 2, 0, 1, 2, 2, 3, 1, 2, 1, 1, 3, 4, 4, 6, 7, 5, 1, 0, 0, 0, -2, -2, -2, 0, 0, 0, 3, 2, 2, 3, 2, 5, 3, 0, -1, 0, 2, 1, 2, 2, 0, 0, 1, 4, 4, 4, 6, 3, 2, 0, 0, 0, 0, -2, -1, 0, 0, 0, 1, 4, 4, 5, 4, 7, 4, 0, -2, -1, 1, 0, 0, 1, -1, 0, 1, 3, 5, 4, 5, 2, 1, 0, 1, 2, 1, -1, 0, -1, -2, 0, 0, 1, 4, 3, 5, 7, 5, 2, 0, 0, 0, 1, 0, 0, -2, -1, -1, 1, 2, 4, 6, 5, 0, -1, 1, 2, 1, 0, 0, 0, -1, -2, 0, 2, 4, 4, 5, 5, 5, 4, 0, 0, 2, 0, 0, -2, -2, -2, -1, 0, 1, 2, 7, 4, 0, 0, 0, 2, 0, 0, -1, -2, -2, -2, 0, 1, 1, 1, 2, 2, 5, 4, 2, 1, 0, 0, 0, 0, -2, -2, -2, -1, 0, 4, 7, 5, 1, -1, 0, 1, 0, -1, -3, -3, -2, -2, -3, 0, 2, 1, 0, 1, 3, 5, 3, 1, -1, 0, 0, 0, 0, -2, -1, -2, 0, 5, 8, 7, 0, 0, 0, 2, 0, -1, -2, -2, -3, -3, -3, -1, 1, 1, 0, 1, 0, 3, 3, 1, 0, 0, 0, 0, -1, 0, -1, -4, -1, 4, 10, 7, 1, -1, 1, 2, 1, 1, -1, 0, -2, -4, -4, -3, 0, 1, 0, 0, 0, 1, 4, 2, -1, -2, 0, 0, 0, 0, 0, -2, 1, 5, 8, 6, 2, 0, 0, 3, 1, 1, 1, 0, -2, -4, -4, -3, -1, 0, 0, 1, 2, 1, 2, 1, 0, -2, -3, 0, 0, 1, 1, 0, 2, 4, 8, 8, 2, -1, 1, 4, 4, 3, 2, 0, -2, -4, -3, -2, -1, 0, 0, 2, 2, 2, 3, 2, 0, -1, -3, -2, 0, 1, 1, 0, 1, 3, 7, 7, 2, 0, 1, 4, 4, 3, 1, 0, -3, -3, -3, -2, -1, -3, 0, 1, 2, 0, 1, 2, 1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 5, 6, 2, 0, 1, 3, 4, 3, 1, 0, -3, -2, -1, -2, -1, -2, 0, 2, 2, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 3, 5, 1, 0, 2, 3, 3, 2, -1, -1, -2, -2, 0, 1, -1, -1, -1, 2, 3, 1, 2, 1, 1, 0, -1, 0, -1, -1, 0, 1, 2, 3, 4, 4, 2, 0, 0, 5, 4, 1, -3, -3, -3, -1, 0, 0, 0, 0, 0, 2, 2, 2, 2, 1, 0, -1, -1, 0, 0, -1, 0, 3, 3, 4, 3, 2, 1, -1, 0, 4, 4, 1, -1, -4, -4, -1, 3, 2, 1, 0, 0, 0, 3, 2, 3, 2, 1, 0, -1, -1, 0, 0, 0, 2, 5, 4, 3, 3, 0, 0, 0, 3, 4, 1, -1, -4, -4, 0, 3, 4, 1, 0, 0, 1, 2, 3, 2, 4, 4, 0, 0, 0, 0, 0, 2, 4, 5, 7, 7, 5, 2, 0, -1, 0, 2, 1, 0, -3, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, 1, 4, 5, 3, 1, 1, 1, 0, -2, -1, -2, -2, -2, -2, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, -2, -3, -3, -2, -2, -3, -2, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, -1, -1, -2, -3, 0, 0, -1, -4, -6, -6, -4, -5, -5, -3, -2, -1, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 1, 2, 1, 1, 2, 2, 1, -1, -1, -2, -1, 0, -2, -4, -5, -5, -4, -3, -4, -4, -3, -2, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 3, 3, 4, 2, 2, 2, 1, -1, -2, -1, -1, 0, 0, -3, -5, -4, -3, -3, -3, -2, -3, -2, -2, -2, -3, -2, -2, -1, 0, 0, 1, 2, 3, 3, 3, 2, 2, 0, 0, -1, -1, 0, 0, 0, 0, -3, -3, -3, -3, -2, -1, -1, -1, -3, -2, -3, -3, -3, -2, -2, -1, 0, 1, 2, 3, 4, 4, 4, 2, 1, 0, 0, -1, 0, 0, 0, -1, -1, -3, -3, -3, -2, -2, -2, -2, -2, -2, -2, -3, -1, -2, -2, -1, 0, 0, 1, 1, 3, 3, 3, 2, 2, 0, -1, -1, -1, -1, -1, 0, 0, -3, -2, -2, -2, -2, -2, -2, -2, -3, -2, -1, -1, -3, -3, -2, -1, 0, 1, 2, 3, 2, 3, 3, 0, 0, 0, -1, -2, -1, 0, 0, -2, -3, -2, -1, -2, -1, -2, -3, -2, -3, -2, -1, -3, -3, -4, -4, -1, 0, 0, 1, 3, 1, 3, 2, 0, 0, -1, -2, -2, 0, 0, 0, 0, -2, -2, -1, -1, -2, -2, -3, -2, -2, 0, -2, -2, -4, -3, -3, -2, 0, 1, 0, 2, 2, 1, 1, 0, 0, -1, -2, -1, -1, -1, 0, -1, -1, -2, 0, -1, -1, -2, -3, -2, -2, 0, -2, -2, -4, -4, -3, 0, 0, 0, 0, 1, 3, 3, 1, 0, 0, -1, -1, -2, -1, -1, -1, 0, -2, -2, -1, 0, 0, -1, -2, -1, -1, -2, -2, -5, -5, -5, -4, -1, -1, 0, 1, 0, 2, 2, 0, 1, 0, -1, -1, -1, 0, 0, 0, -1, -3, -2, -1, 0, -1, -2, -3, -3, -2, -3, -3, -4, -6, -6, -3, -2, -1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, -2, -3, -3, -1, -1, -1, -2, -3, -3, -3, -3, -4, -7, -5, -4, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, 0, 0, -2, -4, -2, -2, -2, -1, -3, -2, -2, -2, -3, -4, -4, -7, -4, -4, -1, -1, 0, -1, -2, -2, 0, 0, 1, 1, 0, -1, -1, -2, -1, 0, -1, -2, -3, -3, -3, -2, -2, -2, -2, -2, -3, -4, -5, -5, -4, -2, -1, -1, -1, -2, -2, -3, -2, 0, 0, 1, 0, -1, -1, -2, -1, 0, -1, -3, -2, -3, -2, -3, -2, -3, -3, -2, -4, -4, -6, -5, -3, -1, -2, -1, -2, -3, -3, -2, -2, 0, 0, 0, 0, 0, -1, -2, -3, 0, -1, -2, -2, -3, -2, -1, -3, -2, -2, -3, -4, -4, -6, -5, -3, -2, 0, -2, -2, -4, -2, -3, 0, 0, 0, 0, 0, 0, -2, -2, -2, -1, -1, -2, -3, -3, -2, -2, -1, -2, -2, -2, -4, -4, -4, -4, -3, -2, -1, -2, -4, -2, -1, 0, 0, 0, 0, -1, 0, -2, -1, -1, -1, 0, -2, -3, -2, -1, -2, -1, -1, -2, -2, -2, -3, -4, -5, -4, -3, 0, 0, -2, -2, -2, 0, 0, 0, 1, 0, 0, -1, -1, -2, -2, -1, -1, -2, -1, 0, 0, -2, -1, -1, -1, -2, -4, -4, -2, -4, -2, -1, -1, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, -2, -2, -2, -2, -1, 0, -1, -1, 0, 0, 0, -1, 0, -1, -2, -3, -3, -3, -2, -3, -2, -2, 0, 0, -1, 0, 0, 1, 1, 1, 2, 0, -1, -1, -1, -1, -1, 0, 0, -2, -1, 0, -2, -1, -1, -1, -1, -2, -4, -1, -3, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 1, -2, -1, -1, -1, -1, -1, -2, -1, 0, -1, -1, -1, 0, -1, -2, -2, -1, -1, -2, -2, 0, -1, 0, 0, 0, 0, -1, -1, 0, 1, 2, 0, 0, -1, -2, -1, -2, -1, -1, -3, -2, -1, -1, 0, -1, 0, -2, 0, -1, -1, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, -1, -2, -1, -1, -2, -1, 0, -1, -2, -1, -1, 0, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 3, 0, 0, -2, -2, -2, -2, -1, -3, -2, -2, -1, -1, -2, -1, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 2, 0, 0, -1, -1, -3, -1, -1, -3, -3, -2, -1, -2, -1, -2, -1, -1, -3, -2, -1, -3, -1, -2, 0, 0, 0, 1, 1, 1, 1, 0, 2, 0, 0, 0, 0, -1, -2, 0, -2, -4, -3, -3, -2, -2, -3, -3, -2, -3, -3, -3, -1, -3, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, -5, -6, -5, -3, -1, -1, -3, -3, -2, -3, -1, -1, -2, -1, -2, 0, 0, 0, 1, 2, 0, 1, 0, 0, -1, -1, -2, -2, -1, -2, 0, 0, -3, -4, -2, -1, -2, -1, -2, -3, -2, -1, -1, 0, -1, -1, -1, -1, 0, -1, 0, 1, 0, 0, 0, -1, -2, -1, -1, -1, -1, -1, -1, 0, 0, -2, -1, -2, 0, -2, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -3, -2, -2, -2, -1, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -2, -3, -2, -2, -2, -1, 0, 0, 0, -1, -1, 0, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -2, -2, -2, -1, -1, -1, -4, -3, -3, -3, -2, -1, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, -2, -1, -2, -1, 0, 0, -2, -3, -2, -2, -2, -3, -1, -1, 0, -1, -1, -2, -1, -2, -1, 0, 0, 0, 0, 1, 1, 2, 0, 0, 1, 0, 0, -2, 0, 0, 0, 0, -3, -2, -2, -2, -3, -2, 0, -1, -1, -2, -1, -1, -2, -2, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, -1, 0, -2, 0, -1, 0, -1, -3, -2, -2, -1, -1, -1, -2, -1, -2, -2, -1, -2, -3, -2, 0, 0, 0, 1, 1, 2, 2, 1, 1, 0, 0, -1, -1, -2, 0, 0, -1, 0, -1, -1, -1, -2, 0, -1, -2, -1, -2, -1, -2, -2, -2, -1, -1, -1, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, -1, -2, 0, 0, -1, -1, 0, 0, -2, -2, -2, -1, -2, -3, -1, -1, -2, -1, -2, -2, -2, -1, 0, 1, 1, 0, 0, 1, 0, 0, -1, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, -2, -1, -1, -1, -2, -3, -3, -1, 0, 0, 0, 0, 1, 2, 0, 0, 0, -2, -1, -2, -1, 0, 0, -1, 0, 0, -1, -1, -1, -2, -1, -3, -1, -1, -1, -1, -3, -3, -3, -1, 0, 0, 0, 1, 1, 1, 1, 0, -1, -1, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -2, -2, -3, -3, -1, -2, -1, 0, 0, 1, 1, 2, 1, 0, 0, -1, -2, -1, -2, 0, 0, 0, -1, -1, -2, -1, -1, -1, -1, -2, -2, -1, -3, -3, -2, -2, -1, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, -1, -2, -1, -1, -1, -2, -1, -3, -1, -2, -3, -4, -3, -3, -2, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, -1, -2, -2, -2, -1, -1, -1, -1, -3, -3, -2, -3, -3, -3, -3, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -2, -1, -2, -2, -2, -2, -2, -2, -2, -1, -2, -3, -3, -4, -2, -2, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, -2, -1, -2, -1, 0, -1, -2, -1, -3, -3, -2, -2, -2, -2, -3, -2, -3, -3, -3, -3, -2, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, -1, 0, -1, -2, -1, 0, -1, -2, -1, -2, -1, -2, -1, -3, -2, -3, -3, -4, -3, -3, -2, -1, -1, 0, -2, -2, -1, -1, 0, 0, -1, 0, -1, -2, -1, -1, -1, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2, -3, -2, -2, -5, -4, -2, -1, -1, -2, -1, -1, -2, 0, 0, -1, 0, 0, 0, -1, -1, -3, -1, -1, -2, -2, 0, -1, -1, -2, 0, -1, -2, -2, -2, -3, -4, -2, -2, -1, -1, -1, 0, -2, 0, 0, 0, 0, 0, -1, 0, -2, -1, -2, -1, 0, -1, -1, 0, 0, -1, -2, -1, -2, -2, -2, -3, -4, -2, -3, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, 0, 0, -2, -1, -1, 0, 0, 0, -1, -2, -2, -3, -2, -3, -2, -1, -2, -1, 0, 0, -1, 0, 0, 1, 1, 0, -1, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, -2, -2, -2, -3, -3, -2, -1, -2, -1, -2, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -1, 0, -1, -1, -1, -1, -1, -2, 0, -1, 0, 0, -3, -2, -3, -2, -2, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -2, -1, 0, -1, -2, -1, 0, 0, 0, -2, -1, -2, -1, -1, -1, -2, -1, -2, -2, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -2, -1, -1, 0, -1, -2, -1, -1, 0, -1, 0, -1, -1, -1, -1, 0, -1, -2, -2, -3, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, -2, -2, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -1, -3, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, -1, -2, -3, -2, -2, 0, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -3, -1, -1, -2, -2, -2, -1, -2, -2, 0, 0, 0, -2, -2, -2, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -2, -1, 0, 0, -2, -3, -2, -2, -1, -1, -2, -2, -2, 0, -1, -1, 0, -2, -2, -2, -1, -1, 0, 0, 0, 1, 0, 0, -1, -2, 0, -2, 0, -1, 0, 0, -3, -4, -2, -2, -1, -2, -1, -1, -1, -1, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, -2, 0, -1, -2, 0, -2, -1, 0, -2, -2, -2, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 2, 1, 1, 1, 2, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 2, 2, 3, 1, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, 0, 0, -1, -1, -2, 0, -2, -1, 0, 1, 1, 1, 2, 2, 1, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, 2, 2, 1, 2, 2, 2, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 1, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 2, 0, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 1, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, -1, -1, -1, -1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 1, 1, 0, -1, -1, 0, -1, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 1, 2, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, -1, -1, -2, 0, 0, 0, 0, 1, 2, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 2, 0, -1, -1, -1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 2, 3, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, -2, -1, -1, 0, 0, 0, 1, 0, 1, 2, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 2, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, -1, -2, -1, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 2, 1, 0, 0, -1, 0, -1, -1, -2, 0, -1, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -2, -1, 0, 1, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 2, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 3, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -2, 0, -1, -1, 0, 0, -1, 0, 0, 0, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, -1, -1, -1, -2, -1, 0, 0, -1, -1, -1, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 3, 3, 3, 0, 1, 2, 2, 2, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 1, 0, 0, 2, 1, 2, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 1, 0, 2, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, -1, 0, 0, -1, -2, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 1, 0, 0, 0, 1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, -2, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 1, 1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 1, 2, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -2, -2, 0, -1, 0, -1, 0, -1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -1, -2, -2, -1, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -2, -1, -1, -1, 0, -2, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -1, -1, -1, 0, -1, -1, -2, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -2, -1, -2, -1, -2, -2, 0, 0, -1, 0, 1, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -2, 0, -1, -1, 0, 0, -1, 0, 1, 1, 1, 0, -2, 0, 0, -1, 0, 0, -1, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, -2, -1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, -1, 0, 0, 1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, -1, -1, 0, 0, 0, 1, 0, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 1, 1, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, -1, -1, 0, -2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, -2, -1, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 2, 0, 1, 2, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 1, 0, 0, -1, -1, 0, -2, -2, -1, 0, 1, 0, 1, 0, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, -1, 0, -1, 0, -1, -1, -2, 0, -1, -1, 0, 0, 0, 0, 1, 0, -1, -1, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, -1, 0, -2, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, -3, -1, -2, -2, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 1, 1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, -2, -2, -2, -2, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, -1, -3, -3, -2, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -2, -1, -3, -2, -2, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, 1, 0, -1, -2, -2, -2, -1, -1, 0, 0, 0, -1, 0, -2, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -2, -1, 0, 0, -1, -1, -2, -3, -1, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, -2, -2, -2, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, -2, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, -1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -2, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, -1, -1, -1, -2, -1, -1, 0, 0, -1, -1, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 2, 3, 2, 1, 1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 2, 2, 3, 3, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, -1, 0, 0, 2, 2, 2, 3, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 4, 4, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 2, 3, 2, 1, 0, 0, -1, -1, -2, -2, 0, 0, 1, 1, 3, 3, 4, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 2, 2, 3, 1, 1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 1, 1, 3, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 2, 4, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 1, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 3, 2, 3, 4, 3, 3, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, 2, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 4, 2, 4, 4, 1, 1, 0, 1, 0, -1, -1, -1, -1, 0, 0, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 2, 3, 4, 3, 3, 2, 3, 1, 1, 2, 0, 1, 0, 0, -1, 0, 0, 1, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 2, 2, 3, 3, 2, 3, 3, 2, 1, 1, 1, 0, 0, 0, 0, 1, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 3, 3, 2, 3, 3, 2, 3, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 2, 2, 3, 1, 1, 3, 2, 2, 0, 0, 0, 0, 1, 1, 0, 0, 2, 2, 2, 1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 2, 1, 3, 4, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 3, 2, 2, 2, 1, 0, 0, 0, 0, 1, 1, 0, 1, 4, 3, 1, 0, 0, -1, 1, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 2, 3, 3, 2, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 1, 1, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 2, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, 0, 1, 0, 0, 0, -1, -3, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -2, 0, 0, 0, 1, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -4, -5, -5, -4, -4, -4, -3, -3, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -4, -5, -4, -4, -3, -4, -4, -3, -1, 0, 1, 0, 0, 0, -1, 0, 1, 0, 1, 3, 3, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -4, -4, -2, -2, -2, -3, -3, -2, 0, 1, 0, 0, 0, 0, 0, 0, 2, 2, 2, 3, 1, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -4, -4, -2, -3, -2, -3, -1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 3, 2, 3, 3, 1, 0, 1, 0, 0, 0, 0, 2, 1, 0, -1, -2, -3, -3, -1, -2, -1, -1, 0, -1, -1, -1, 0, 0, 1, 0, 2, 2, 3, 2, 4, 2, 2, 1, 1, 2, 0, 0, 0, 1, 0, 0, 0, -3, -3, -3, -2, -2, -1, -2, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 1, 3, 2, 1, 1, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, -3, -3, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, -3, -1, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -2, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, -2, -2, -1, -1, 0, 1, 1, 2, 1, 2, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, -2, 0, 1, 0, 1, 1, 1, 0, 0, 0, -1, -2, -3, -2, -1, 0, 1, 2, 2, 2, 3, 2, 0, 1, 0, 0, 0, 2, 2, 1, 0, -1, -2, 0, 0, 1, 1, 0, 1, 0, 1, -1, -2, -3, -2, -1, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 2, 3, 4, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -3, -3, -4, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 2, 2, 3, 3, 2, -1, -1, -1, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, -3, -3, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 3, 2, 4, 3, 4, 1, 0, -1, -1, 0, 0, 1, 0, 0, 1, 1, 2, 0, 0, 0, -2, -2, -3, -2, -2, -3, -4, -3, -2, -1, -1, 1, 3, 1, 2, 2, 3, 0, 0, -1, -2, 0, -1, 0, 0, 1, 1, 2, 1, 2, 0, 0, 0, -1, -2, -3, -4, -4, -3, -4, -4, -2, 0, 1, 1, 1, 1, 1, 2, 0, -1, -1, 0, 0, -1, 0, 0, 1, 2, 2, 2, 2, 0, 0, 0, 0, 0, -2, -2, -5, -4, -4, -2, -1, 0, 0, 1, 2, 1, 1, 0, 0, 0, -1, 0, -1, -1, 0, 2, 2, 3, 3, 2, 2, 0, 0, -1, 0, 0, -2, -3, -3, -4, -3, -2, -1, -1, 0, 0, 1, 2, 3, 2, 1, 0, -1, 0, -1, 0, 0, 1, 2, 1, 2, 2, 3, 0, 0, 0, 0, -1, -1, -3, -3, -3, -2, -1, 0, 0, 0, 2, 1, 1, 2, 0, 1, 0, 0, -1, 0, 1, 1, 1, 0, 0, 3, 2, 2, 1, 1, 1, 0, 0, -1, -3, -2, 0, 0, 0, 0, 1, 0, 2, 1, 1, 1, 1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 2, 2, 1, -1, -2, -1, 2, 0, 1, 2, 1, 2, 1, 2, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 1, 4, 1, 0, -2, 0, 1, 1, 0, 1, 2, 0, 0, 1, 2, 1, 1, 0, 1, 0, 0, 1, 0, -1, -1, 0, 0, 1, 1, 0, 0, 1, 2, 2, 0, 0, -1, -1, 1, 2, 1, 1, 1, 1, 0, 1, 2, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 2, 0, -2, 0, 0, 0, 2, 2, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 2, 1, 0, -1, 0, 0, 1, 2, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 1, 0, 1, 0, 2, 1, 0, -3, 0, 1, 1, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 2, 2, 1, 2, 0, 0, 0, 0, 0, -1, -3, -2, 0, 1, 0, 0, -2, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, -4, -1, 0, 0, 0, -1, -2, -3, -1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -3, -2, 0, 0, -2, -3, -3, -2, -2, 0, 0, 1, 0, 0, 1, 0, 0, 2, 2, 2, 0, 0, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, -4, -3, -1, 0, -2, -3, -4, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -2, -3, -2, -3, -2, -1, 0, -1, -1, -1, 0, -3, -2, 0, 0, 0, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, -3, -3, -3, -3, -2, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 1, 0, 1, 1, 1, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -2, -2, -1, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, -1, -1, 0, 0, 1, 3, 2, 0, 0, 1, 1, 2, 2, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 1, 0, -1, -1, -2, -1, -1, 0, 1, 1, 3, 2, 0, 0, 2, 2, 1, 2, 0, 0, 1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 1, 1, 0, 1, 1, 1, 0, 2, 1, 0, -1, -3, -2, 0, 0, 2, 1, 1, 1, 2, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 3, 4, 3, 0, 0, 1, 1, 0, 0, 0, 0, -2, -2, -3, -2, -2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 3, 2, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 3, 4, 3, 0, -1, 0, 0, 2, 2, 0, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 3, 4, 3, 1, 0, 0, 1, 1, 2, 0, 0, 0, 0, -1, -3, -2, -2, -1, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, -1, 0, 1, 1, 3, 5, 4, 1, 0, 0, 0, 1, 2, 0, 0, 0, 0, -1, -2, -3, -1, 0, 0, 0, 0, 0, 2, 0, 0, 0, -1, -2, -1, 1, 1, 3, 3, 5, 6, 1, 0, 0, 1, 0, 2, 0, 0, 1, 0, -2, -2, -3, -1, 0, 0, 2, 2, 3, 2, 1, 0, 0, -2, 0, 0, 0, 2, 3, 5, 6, 6, 2, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, -1, -1, 0, 1, 2, 2, 2, 2, 2, 1, 0, -1, -2, -1, 0, 1, 2, 3, 5, 7, 6, 2, 0, 1, 1, 1, 1, 0, 0, 1, 2, 2, 1, 0, 0, 0, 1, 3, 2, 2, 1, 1, 0, 0, -1, -1, 0, 1, 2, 4, 4, 6, 5, 1, 0, 0, 0, 0, -1, 0, 1, 2, 3, 2, 3, 1, 2, 4, 4, 2, 1, 0, 2, 0, 0, -1, 0, 0, 0, 0, 2, 3, 5, 4, 5, 1, 0, 1, 0, -1, 0, 1, 1, 1, 4, 5, 4, 4, 3, 3, 4, 3, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 3, 3, 5, 3, 1, 0, 0, 0, -2, -1, 0, 1, 3, 4, 4, 4, 4, 5, 5, 4, 4, 2, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 1, 3, 4, 3, 1, 0, 1, 1, 0, 0, 2, 2, 2, 3, 3, 4, 5, 6, 5, 6, 4, 1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 1, 3, 3, 3, 1, 0, 1, 0, 1, 1, 1, 0, 1, 1, 3, 5, 5, 4, 4, 5, 2, 2, 1, 0, 2, 0, 1, 0, -1, -2, 0, 0, 1, 3, 5, 2, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 2, 4, 6, 3, 5, 2, 2, 2, 1, 0, 2, 0, 0, -1, -2, -1, -1, 0, 0, 3, 4, 4, 1, 0, 0, 2, 0, 0, 0, -1, 0, 0, 1, 2, 3, 3, 2, 2, 2, 1, 2, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 3, 6, 4, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 3, 3, 2, 1, 1, 2, 0, 0, -1, -2, 0, 0, 0, 0, -2, -1, 0, 4, 7, 5, 2, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 1, 1, 0, 1, 0, 0, -1, -1, -1, 0, -1, 0, -1, -2, 0, 4, 6, 6, 2, 0, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, -1, -1, -1, 1, 3, 6, 5, 2, 0, 1, 2, 2, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 5, 5, 6, 3, 0, 2, 2, 3, 2, 1, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, -1, -1, -2, -2, -2, -1, 0, -1, 0, 1, 2, 3, 6, 5, 3, 0, 1, 3, 2, 2, 1, 1, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 1, 1, 3, 5, 5, 2, 0, 2, 3, 2, 2, 0, 0, 0, -2, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 2, 2, 4, 4, 4, 0, 1, 3, 4, 1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 2, 1, 2, 0, 0, 0, 0, -2, 0, 0, -2, 0, 0, 1, 2, 4, 4, 3, 1, 2, 3, 4, 2, -1, -2, -1, 0, 0, 1, 0, 0, 1, 2, 2, 2, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 3, 2, 3, 0, 1, 1, 4, 3, 2, 0, -1, -2, 0, 0, 2, 1, 1, 0, 2, 2, 1, 1, 2, 1, 0, -1, 0, 0, 0, 0, 1, 3, 4, 2, 3, 1, 1, 0, 2, 2, 2, 0, 0, -1, 0, 2, 2, 1, 0, 1, 2, 1, 2, 2, 3, 2, 0, 0, 0, 0, 0, 0, 1, 3, 4, 4, 3, 2, 0, 1, 2, 2, 1, 1, 1, 1, 1, 0, 2, 1, 1, 1, 3, 1, 1, 1, 1, 1, 0, 1, 1, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1,
    -- filter=0 channel=5
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, 0, -1, -2, -2, -2, -1, 0, 0, 1, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 1, 0, 1, 1, 2, 1, 0, 0, -1, -1, -2, -1, -2, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 2, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, -1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -2, -1, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, -2, -2, -1, 0, -1, 0, 0, 1, 1, 2, 1, 0, 0, 0, 2, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 2, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 1, 1, 0, 1, 1, 1, 0, 2, 2, 1, 2, 2, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 2, 1, 1, 2, 0, 1, 1, 2, 2, 1, 0, 1, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 2, 2, 2, 2, 2, 2, 1, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 2, 2, 2, 1, 1, 2, 2, 1, 1, 1, 2, 2, 2, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 2, 0, 1, 0, 1, 1, 0, 2, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 2, 2, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 2, 0, 3, 2, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 3, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 2, 2, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 2, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 1, 2, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 2, 1, 2, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 2, 0, 1, 2, 3, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 2, 0, 1, 1, 0, 1, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 2, 2, 0, 1, 0, 1, 2, 1, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -2, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, -2, -2, 0, -1, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -2, -1, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, -2, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -2, -2, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, 0, -1, -1, -2, -1, 0, 0, 0, 0, -2, -2, -1, 0, 0, -1, -1, -1, -2, -2, -2, -2, -1, 0, 0, -1, -1, -3, -2, -2, -3, -3, -4, -5, -5, -4, -4, -4, -3, -2, -1, 0, -3, -2, -2, -1, 0, -2, 0, -2, -1, -1, -1, -1, -1, -1, -1, -2, -3, -3, -1, -2, -2, -3, -3, -3, -3, -3, -3, -3, -1, -1, 0, 0, -2, -2, -3, -1, 0, -1, 0, -2, -1, -1, -2, -2, -3, -1, -1, -2, -1, -1, -2, -1, -2, -3, -2, -3, -3, -2, -2, -1, -1, 0, -2, 0, -2, -3, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, -2, -3, -1, 0, -1, -2, -2, 0, 0, -2, -2, -1, -2, -2, 0, 0, -1, -1, -1, 0, -2, -3, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -2, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, -2, -2, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, -2, -2, 0, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 2, 2, 2, 1, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 2, 2, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 2, 1, 2, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 2, 1, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 2, 1, 1, 0, 0, 0, 1, 1, 0, -1, 0, 0, 2, 2, 1, 4, 3, 3, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 1, 2, 2, 2, 1, 1, 0, 0, 1, 1, 1, 0, -1, 0, 0, 1, 2, 4, 4, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 2, 2, 2, 1, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 1, 3, 4, 2, 2, 1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 1, 1, 1, 1, 2, 1, 1, 0, 1, 2, 2, 0, 0, 0, 0, 2, 1, 3, 4, 3, 2, 1, 0, 0, 1, 0, 0, -2, -1, 1, 0, 0, 0, 0, 2, 3, 3, 2, 1, 1, 2, 0, 0, 0, -1, 0, 0, 1, 2, 4, 3, 3, 2, 3, 0, 0, 1, 1, 0, -1, 0, 0, 0, 1, 0, 0, 1, 2, 1, 3, 2, 2, 1, 0, 0, -1, -1, 0, 0, 1, 3, 3, 3, 4, 4, 2, 1, 0, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 3, 3, 3, 3, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 3, 2, 2, 3, 1, 3, 2, 1, 1, 0, 0, -1, -1, 0, 1, 1, 1, 0, 2, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, -2, 0, 1, 1, 2, 2, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 1, 1, 2, 0, 0, 1, 1, 1, 1, 1, 0, -2, -1, 0, 1, 0, 2, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 3, 2, 0, 2, 0, 0, 1, 0, 0, 1, 1, 0, 0, -2, -1, 0, 0, 0, 1, 1, 0, 0, 0, -2, 0, 0, 0, 0, 1, 0, 2, 0, 2, 1, 2, 2, 0, 1, 0, 1, 0, 0, 1, 0, 1, -3, -1, -1, 0, 0, 0, 1, 1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 2, 1, 1, 0, 0, 0, 1, 0, 0, 0, -2, -4, -2, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 3, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, -4, -3, -3, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -3, -3, -1, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, 0, -2, -2, -3, -1, -1, -1, -1, 0, -2, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -2, 0, -1, -1, -1, -1, -1, -2, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 1, 1, 0, 2, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, -1, -2, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, 0, -1, 0, 0, 1, 0, -2, -3, -1, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, -1, 0, 1, 1, 0, 0, -2, -3, -2, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -2, -3, -1, 0, 0, 0, -1, 1, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, 0, 0, 1, 1, 0, 0, -1, -2, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, -1, -2, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, 0, -3, -3, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 2, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 2, 2, 0, 1, -1, -3, -4, -2, -1, 0, 0, 1, 0, 1, 2, 2, 3, 4, 2, 3, 1, 1, 1, 0, 2, 1, 1, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, -2, -3, -1, 0, 0, 1, 0, 1, 1, 3, 3, 3, 3, 2, 2, 3, 2, 3, 1, 3, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -3, -2, -1, 0, 2, 1, 2, 1, 1, 3, 2, 3, 2, 2, 2, 2, 2, 4, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, 1, 1, 2, 3, 1, 1, 1, 2, 0, 1, 1, 1, 3, 2, 3, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 1, 2, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 3, 2, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -2, 0, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 3, 2, 1, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 3, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 2, 2, 2, 1, 0, 0, 0, 0, -1, 0, 0, 2, 0, 0, 0, -1, 0, 0, 1, 2, 2, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 1, 1, 0, 2, 2, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 1, 4, 3, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 2, 1, 1, 1, 1, 1, 0, 0, 0, -1, 0, -1, -2, 0, 0, 3, 3, 4, 2, 1, 1, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, 1, 1, 2, 1, 1, 3, 1, 0, 0, -1, -1, 0, 0, -1, 0, 1, 3, 5, 3, 3, 2, 2, 2, 3, 3, 3, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, -1, -2, -2, 0, -1, -2, 0, 1, 3, 3, 3, 2, 3, 3, 2, 2, 4, 3, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, -2, 0, 1, 2, 2, 3, 3, 3, 4, 3, 3, 2, 2, 1, -1, -1, -1, 0, 0, 0, 1, 1, 2, 2, 1, 0, 0, 0, -1, 0, 1, 0, -2, 0, 1, 1, 2, 2, 4, 4, 4, 2, 3, 0, 2, 0, 0, 0, 0, 1, 1, 2, 1, 2, 0, 2, 0, 0, 0, 0, 1, 1, 0, 0, -2, 0, 0, 1, 1, 1, 2, 3, 4, 2, 2, 1, 0, 1, 1, 1, 0, 2, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 0, -1, 0, 0, 0, 0, 1, 2, 3, 1, 1, 0, 1, 0, 0, 1, 2, 2, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, -1, -1, -1, -1, -1, 0, 0, 1, 2, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 2, 1, 0, 1, 2, 1, 0, -1, -2, -2, -3, -3, -2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 2, 1, 2, 0, 0, 0, 1, 1, 0, -2, -2, -3, -3, -2, -2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 2, 2, 1, 0, 0, 1, 2, 0, 0, -2, -3, -2, -1, -3, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 1, 0, 0, -2, -2, -1, -2, -3, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, -2, -1, -2, -1, -1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 1, -1, -2, -2, -1, -1, -2, -1, -1, -1, -1, -1, 0, -1, 0, 0, -1, -1, 0, -1, -1, -2, -2, -1, 0, 0, -1, -2, -1, 0, 1, 1, 0, 0, -1, -2, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, -1, -2, -1, -1, 0, -1, -2, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, -2, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, -1, -2, -1, 0, -1, -2, 0, -1, -1, -1, -2, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -2, -2, -2, -1, 0, -1, -2, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -2, -2, -2, -2, -2, -1, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -2, -2, -2, -2, -1, -1, -1, 0, -2, -1, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, -1, -1, -1, -1, -1, -1, -2, -1, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -2, -2, -1, 0, 0, -1, -1, 0, -2, -2, -1, 0, -1, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -2, -2, -1, -2, -1, -1, -1, 0, -1, -2, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -2, -1, -1, -1, 0, -1, -1, -1, -1, -1, 0, -1, -2, 0, -1, 0, -1, -1, -1, -1, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -2, -1, -1, 0, -1, -1, -1, -1, -1, -1, 0, -1, 0, -1, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -3, -2, -3, -2, -1, -2, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, -1, -1, -1, 0, -1, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -2, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, -2, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, -1, -1, 0, -1, -1, -1, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -2, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -2, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -2, -1, -2, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 1, 1, 2, 1, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 0, 0, 2, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 1, 2, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 2, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 2, 2, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 2, 3, 2, 2, 3, 2, 1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, -1, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 1, 2, 2, 1, 2, 2, 1, 1, 1, 0, 0, 0, 0, 2, 1, 1, 1, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 2, 2, 2, 0, 0, 0, 0, 2, 1, 2, 1, 1, 0, 0, -1, -2, -3, 0, -1, -1, 0, 0, 0, 0, -2, -1, -2, -2, -1, 0, -1, 0, 0, 2, 0, 1, 0, 0, 0, 1, 3, 2, 3, 1, 1, 0, -1, -4, -3, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 1, 1, 0, 0, 0, 1, 1, 2, 1, 3, 1, 0, -1, -3, -3, -2, 0, -1, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 1, 3, 1, 1, 0, -1, -2, -3, -3, -1, -1, -2, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 2, 0, 1, 3, 2, 1, 2, 2, 1, 0, -1, -1, -4, -2, -2, -1, -1, -1, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 1, 1, 1, 2, 1, 2, 3, 3, 1, 0, 0, -2, -3, -1, -1, -1, 0, 0, -1, -2, -1, 0, 0, 1, 1, 1, 0, 0, 1, 2, 2, 1, 1, 1, 1, 2, 2, 2, 1, 1, 1, 0, 0, -1, -3, -2, -2, 0, 1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 1, 2, 1, 1, 2, 1, -1, -2, -1, -1, 0, 0, 0, 1, 0, -1, -2, -1, -2, -1, 0, 0, 0, 0, 2, 2, 2, 1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -4, -3, -3, -1, -1, 0, 0, 1, 0, 1, 3, 1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, -1, -1, 0, 0, 1, 2, 1, 0, -1, -2, -3, -4, -3, -2, -1, -1, -1, 0, 1, 1, 2, 0, 1, 0, 0, 0, -1, -1, 0, 1, 1, 0, -1, -1, 0, 1, 1, 1, 2, 0, -1, -2, -4, -2, -2, -2, -1, -3, -2, 0, 1, 1, 1, 2, 0, 0, 0, 0, -1, 0, 0, 2, 0, 0, 0, 0, 0, 1, 2, 3, 3, 1, 0, -2, -3, -3, -3, -2, -3, -2, -1, -1, 0, 1, 0, 0, 1, 0, 1, 0, 0, -1, 0, 3, 1, 0, 0, 0, 0, 2, 2, 4, 2, 1, 0, -1, -1, -1, -1, -2, -3, -2, -1, -1, -1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 2, 1, 0, 0, -1, 0, 2, 3, 4, 3, 2, 0, 0, -2, -1, -1, -2, -1, -3, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 2, 0, 0, 0, 0, 0, 3, 3, 5, 2, 1, 1, 0, -1, 0, 0, 0, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 2, 4, 4, 2, 2, 0, 1, 0, 1, 1, 0, -1, -2, -2, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 4, 3, 2, 2, 2, 1, 1, 0, 0, 0, 0, -3, -2, -1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 2, 1, 2, 1, 1, 0, 0, 0, -1, -1, -1, 0, 0, 2, 1, 2, 2, 1, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, -1, 0, -1, -1, 0, 0, 1, 1, 1, 0, 2, 1, 1, 0, 1, 1, 1, 2, 3, 3, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, -1, -2, -2, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 2, 2, 2, 2, 3, 3, 3, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 2, 3, 3, 3, 2, 2, 3, 4, 3, 0, 0, -2, -1, 0, -1, 0, 0, 2, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 2, 3, 1, 3, 4, 4, 3, 3, 4, 3, 5, 2, 0, 0, -1, 0, 0, -2, 0, 0, 1, 1, 2, 1, 0, 0, 0, 2, 1, 0, 1, 0, 0, 2, 2, 2, 3, 4, 2, 3, 3, 3, 3, 2, 0, -1, -1, 0, 0, 0, -1, 1, 1, 1, 1, 1, 1, 2, 2, 3, 2, 0, 0, 0, 1, 2, 1, 2, 3, 2, 3, 1, 1, 2, 4, 2, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 2, 3, 2, 1, 1, 2, 1, 1, 0, 0, 0, 1, 0, 1, 2, 2, 0, 0, 1, 3, 3, 3, 1, 0, 0, 1, 1, 1, 0, 0, 1, 2, 2, 3, 1, 2, 1, 2, 1, 1, 0, 1, 0, 0, 0, 0, 2, 2, 1, 0, 2, 2, 2, 1, 1, 0, 0, 1, 1, 1, 0, 0, 1, 1, 2, 2, 2, 1, 1, 1, 2, 1, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 2, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -1, 0, 0, 0, -1, -2, -3, -3, -3, -4, -3, -4, -6, -5, -4, -5, -5, -5, -2, -1, 0, 0, -1, -1, 0, 0, -1, -1, -2, -2, 0, 0, -1, 0, -1, 0, -2, -2, -3, -5, -4, -4, -4, -5, -7, -7, -7, -8, -6, -6, -4, -2, 0, -2, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 1, 0, -1, -1, -2, -2, -3, -3, -3, -4, -3, -5, -5, -4, -5, -6, -5, -5, -4, -2, 0, 0, -2, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -2, -1, -2, -1, -3, -3, -3, -2, -4, -4, -4, -4, -4, -2, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, -3, -3, -2, -3, -3, -2, 0, -1, -1, -1, 0, 0, 1, 0, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, 0, 1, 0, 0, 1, 1, 0, 2, 0, 1, 1, 0, 1, 0, 1, 2, 2, 2, 3, 2, 2, 2, 2, 2, 2, 1, 0, 0, -1, -1, -1, -1, 0, 0, 1, 0, 1, 0, 2, 1, 1, 1, 1, 0, 1, 2, 2, 2, 2, 4, 3, 2, 3, 3, 3, 3, 5, 5, 2, 0, 0, 0, -1, -2, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 2, 0, 1, 0, 1, 3, 4, 5, 3, 2, 2, 3, 4, 5, 4, 4, 3, 1, 0, -1, 0, -1, 1, 2, 1, 2, 0, 2, 0, 1, 0, 2, 1, 1, 1, 2, 1, 4, 6, 4, 3, 2, 2, 4, 3, 3, 5, 4, 3, 0, -1, 0, 0, 0, 2, 3, 3, 2, 3, 2, 1, 1, 0, 1, 0, 1, 2, 2, 2, 4, 5, 5, 3, 2, 2, 3, 4, 3, 5, 4, 3, 0, 0, 0, 0, 0, 3, 3, 5, 4, 3, 2, 0, 0, 0, 0, 0, 0, 3, 4, 4, 5, 5, 5, 4, 4, 4, 4, 3, 3, 5, 4, 3, 0, 0, 1, 1, 1, 4, 5, 5, 5, 3, 2, 0, -2, -2, -1, 0, 0, 2, 2, 4, 4, 6, 4, 4, 3, 3, 3, 4, 4, 4, 3, 3, 0, -1, 1, 1, 1, 5, 7, 7, 6, 4, 1, 0, 0, -1, -1, 0, -1, 2, 3, 4, 5, 4, 4, 4, 2, 3, 3, 3, 3, 2, 3, 3, 1, 0, 0, 1, 2, 5, 8, 8, 5, 4, 3, 2, 0, 0, 0, 0, 0, 0, 2, 3, 4, 3, 4, 2, 2, 1, 2, 3, 3, 1, 2, 0, 0, -1, 0, 2, 2, 5, 7, 7, 6, 5, 3, 2, 0, 1, 0, 0, -1, 0, 1, 1, 1, 2, 1, 1, 1, 1, 2, 2, 3, 2, 1, 0, -1, -1, 0, 1, 3, 5, 7, 7, 7, 5, 3, 1, 2, 0, 1, 0, 0, 0, 0, 1, 1, 1, 2, 0, 2, 1, 2, 2, 2, 1, 0, -2, -1, -1, 1, 2, 1, 6, 7, 7, 7, 6, 4, 3, 1, 1, 1, 0, -1, 0, 1, 2, 2, 2, 1, 0, 1, 1, 2, 2, 4, 2, 0, -2, -2, -1, 0, 1, 2, 4, 6, 7, 4, 3, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 3, 2, 1, 1, 1, 1, 3, 3, 4, 2, 0, 0, -2, -2, 0, 0, 0, 3, 5, 4, 3, 2, 2, 0, 0, 0, 0, 0, -1, -1, 0, 2, 4, 4, 3, 2, 2, 2, 4, 4, 5, 3, 1, -1, -1, -2, 0, 0, -1, 1, 3, 3, 3, 2, 0, 0, 0, 0, -3, -2, -2, -1, 0, 0, 3, 4, 4, 3, 2, 3, 4, 5, 3, 2, 1, 0, -1, -1, -2, -1, -4, 0, 2, 3, 3, 2, 2, 1, 0, -1, -1, -1, -2, 0, 0, 1, 3, 5, 4, 3, 2, 2, 5, 5, 3, 2, 1, 0, 0, -1, 0, -2, -3, -2, 0, 1, 2, 1, 2, 1, 0, 0, 0, -1, 0, 0, 2, 2, 4, 4, 3, 2, 2, 4, 4, 4, 3, 1, 0, 0, 0, -1, -1, -1, -4, -2, 0, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 1, 2, 3, 2, 2, 3, 3, 3, 4, 3, 2, 2, 0, 0, 0, 0, -2, -1, -3, -6, -4, -1, -1, 0, 1, 1, 1, 0, 0, 1, 0, 1, 0, 2, 2, 3, 2, 3, 4, 3, 4, 4, 3, 1, 0, 0, 0, 0, -1, -1, -3, -6, -5, -4, -2, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 2, 2, 2, 4, 3, 2, 2, 2, 0, 0, -1, -2, 0, -1, -2, -2, -6, -4, -3, -2, 0, 1, 1, 0, 1, 0, 0, 1, 1, 1, 1, 3, 3, 3, 3, 4, 2, 3, 2, 0, 0, 0, 0, -2, -2, -1, -1, -2, -5, -3, -2, -1, 0, 1, 1, 1, 0, 0, 2, 3, 2, 1, 0, 0, 3, 2, 2, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -1, -2, -4, -2, -1, -2, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 2, 0, 2, 1, 1, 0, 0, 0, -1, -1, -1, -2, -4, -4, -1, 0, -1, -2, -2, -3, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, -1, 0, -1, -2, -3, -3, -3, -3, -3, -2, -2, 0, -1, -2, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -4, -4, -5, -4, -5, -4, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -2, -1, -2, -2, -3, -3, -3, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 2, 1, 0, 1, 0, 0, 1, 1, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 1, 1, 1, 1, 2, 1, 3, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 1, 2, 3, 2, 3, 3, 0, 0, 0, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 1, 1, 0, 1, 2, 1, 3, 2, 2, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 2, 2, 3, 1, 3, 2, 0, 0, 1, 1, 2, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 3, 2, 3, 1, 0, 0, 0, 1, 1, 2, 2, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 2, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 1, 1, 0, 2, 1, 0, 1, 1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, 2, 1, 0, 0, 1, 1, 2, 2, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, -2, -1, 0, 1, 0, -2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 2, 1, 2, 0, 0, 0, 0, -2, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 2, 2, 0, 1, 1, 0, 1, 1, 0, -1, -2, -2, -1, 0, 0, -1, 0, -2, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, -1, -2, 0, 0, 0, -1, -1, -1, -3, -1, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -1, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 2, 1, 1, 1, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, -3, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 3, 2, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 2, 0, 1, 2, 1, 1, 2, 3, 3, 2, 0, 1, 2, 2, 0, 0, 0, 0, 1, 0, -1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 3, 1, 2, 1, 3, 2, 2, 0, 1, 0, 1, 2, 0, 1, 1, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 2, 1, 0, 0, 2, 1, 1, 2, 3, 2, 0, 1, 0, 0, 1, 1, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 2, 2, 0, 1, 2, 0, 0, 1, 2, 1, 1, 0, 0, 0, 1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 3, 1, 0, 1, 2, 2, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 2, 2, 2, 2, 1, 0, 0, -1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 1, 1, 1, 2, 1, 0, 0, 1, 3, 4, 1, 1, 0, 0, -1, 0, 1, 1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, 2, 2, 2, 1, 0, -1, 0, 0, 1, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, 2, 1, 0, 0, 0, 0, 1, 2, 3, 2, 1, 0, 0, 0, 2, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 3, 2, 1, 0, 0, 0, 1, 2, 3, 0, 1, 0, 0, 2, 1, 1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 1, 2, 3, 2, 1, 2, 2, 3, 2, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -1, -1, 0, 0, 1, 1, 1, 2, 1, 1, 1, 2, 2, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, -1, -1, 0, -2, -1, -1, 0, -2, -2, -2, -2, -2, -1, -3, -3, -3, -2, -2, -3, -3, -2, -1, 0, -1, -1, -2, -2, -2, -1, 0, -2, -2, -2, -3, -2, -1, -2, -1, -1, -3, -4, -4, -3, -4, -4, -4, -4, -5, -5, -4, -5, -5, -5, -4, -1, 0, -2, -2, 0, -2, -1, -1, -1, -2, -2, -3, -2, -2, -2, -2, -2, -3, -2, -4, -2, -3, -3, -4, -3, -2, -3, -4, -4, -4, -4, -3, 0, -1, -2, -2, -2, -2, -1, 0, -1, -1, -1, -2, -1, -3, -3, -3, -1, -2, -2, -2, -3, -2, -3, -3, -3, -3, -4, -4, -4, -3, -3, -2, -1, -1, -1, -1, -2, -1, 0, 0, -1, -1, 0, -1, -1, -1, -1, -1, -2, -1, -1, -1, -2, -2, -1, -3, -2, 0, -2, -2, -3, -3, -3, -1, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, -1, 0, 0, -2, -1, 0, -1, -1, -2, -1, 0, -1, -2, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 1, 0, 0, 0, 1, 2, 1, 2, 1, 1, 0, 0, -2, -1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 0, 0, 2, 2, 1, 3, 2, 2, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 1, 2, 3, 2, 1, 2, 2, 1, 3, 4, 3, 1, 1, 0, 0, -1, 0, 0, 2, 1, 2, 3, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 1, 2, 3, 2, 1, 3, 1, 1, 3, 4, 4, 3, 2, 0, 1, 0, 0, 0, 1, 2, 3, 4, 3, 3, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 4, 3, 2, 2, 1, 1, 2, 3, 2, 3, 1, 0, 0, 0, 0, 1, 3, 3, 5, 5, 5, 2, 2, 0, 0, 0, 0, 0, 0, 1, 1, 3, 2, 2, 2, 3, 2, 3, 2, 1, 3, 2, 1, 0, 1, 0, 1, 1, 2, 4, 4, 5, 4, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 2, 2, 1, 2, 1, 3, 2, 2, 0, 0, 0, -1, 1, 1, 3, 5, 5, 4, 4, 5, 3, 2, 2, 2, 0, 0, 1, 2, 1, 2, 1, 1, 2, 2, 2, 1, 1, 2, 2, 2, 1, -1, 0, -1, 1, 2, 3, 4, 3, 4, 5, 4, 2, 2, 2, 1, 1, 0, 0, 1, 1, 1, 1, 2, 1, 2, 0, 1, 1, 2, 3, 1, 1, -1, 0, 0, 0, 2, 4, 5, 4, 5, 4, 5, 3, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 1, 2, 2, 1, 2, 1, 0, -1, 0, 0, 1, 2, 4, 3, 5, 5, 5, 4, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 2, 0, 0, -1, -1, -1, 0, 2, 2, 3, 4, 4, 5, 2, 1, 3, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, 2, 2, 2, 3, 3, 1, 0, 0, -1, 0, 0, 2, 1, 2, 2, 4, 2, 1, 2, 2, 1, 0, -1, 0, -1, 0, 1, 0, 2, 2, 0, 2, 2, 3, 2, 3, 3, 0, 0, -1, 0, -1, 0, 0, 0, 0, 2, 2, 3, 3, 2, 0, 0, 0, 0, -1, -1, 0, 1, 1, 2, 3, 1, 2, 3, 3, 2, 2, 2, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 2, 3, 3, 1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 3, 2, 2, 2, 2, 3, 2, 2, 2, 0, 0, -1, 0, -3, -2, -1, -1, -1, 0, 0, 2, 2, 1, 0, 0, 0, -1, 0, 0, 0, 1, 2, 3, 3, 1, 1, 2, 3, 1, 1, 1, 0, 0, 0, 0, -2, -2, -2, -3, -2, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 1, 2, 3, 2, 1, 1, 0, 0, 0, -1, -1, -2, -4, -3, -2, -1, -1, 0, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, 1, 1, 0, 3, 2, 2, 3, 1, 0, 0, 0, 0, -1, 0, -3, -3, -4, -4, -4, 0, 0, 0, 1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 2, 1, 1, -1, 0, -1, -1, -1, -3, -4, -3, -4, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 0, 0, -1, -1, -1, 0, -2, -3, -4, -3, -3, -3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -1, -2, -2, -2, -2, -3, -2, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -2, 0, -1, -2, -2, -3, -3, -2, -3, -1, -1, -2, -1, -1, -1, 0, -1, 0, 0, -2, -2, -1, -2, -1, -1, 0, -1, -3, -1, -3, -2, -3, -4, 0, 0, -1, -1, -2, -2, -2, -2, -2, -1, -1, -2, -2, -2, 0, -1, 0, 0, 0, -2, 0, -2, -2, -1, -2, -3, -3, -2, -4, -4, -4, -3, 0, -1, 0, -1, -2, -2, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, -2, -1, -1, -2, -1, -3, -2, -3, -3, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -1, -2, -2, -2, -2, -3, -3, -2, -3, -2, -1, -1, -2, -3, 0, 0, 0, 2, 3, 2, 2, 2, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, -1, -2, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 3, 2, 2, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 2, 1, 2, 0, 1, 0, 0, 0, 1, 2, 1, 1, 1, 0, -2, -2, -1, -2, -2, -2, -1, -2, -1, -1, -1, 0, -1, 0, 0, 1, 2, 3, 3, 3, 2, 1, 2, 0, 0, 1, 2, 1, 1, 0, 1, 0, 0, -1, -1, -1, -1, -1, -1, 0, -1, -1, -2, 0, -1, -1, 0, 2, 2, 3, 3, 2, 1, 1, 1, 2, 1, 1, 2, 1, 1, 2, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 2, 3, 4, 3, 2, 3, 3, 2, 3, 4, 3, 1, 1, 2, 1, 2, 2, 3, 3, 4, 3, 2, 2, 4, 1, 1, -1, 0, 2, 3, 2, 2, 2, 3, 4, 3, 4, 4, 4, 2, 3, 3, 2, 2, 2, 0, 2, 2, 4, 5, 6, 5, 4, 4, 5, 5, 2, 1, 0, 0, 1, 1, 2, 0, 2, 2, 4, 5, 6, 4, 5, 2, 1, 0, 0, 2, 0, 0, 1, 4, 3, 4, 4, 4, 4, 4, 5, 2, 0, 1, 0, 0, 0, 0, 1, 1, 2, 4, 5, 5, 6, 5, 4, 4, 1, 0, 1, 0, 3, 3, 4, 3, 3, 2, 0, 2, 3, 4, 2, 1, 0, 0, 0, 0, 2, 1, 0, 2, 5, 5, 4, 4, 4, 4, 4, 4, 3, 3, 3, 3, 3, 2, 4, 4, 4, 3, 0, 1, 3, 1, 1, 2, 1, 0, 0, 0, 0, 0, 1, 3, 5, 4, 6, 4, 4, 4, 4, 4, 5, 3, 3, 1, 2, 2, 2, 2, 3, 4, 2, 3, 3, 1, 1, 2, 0, 0, 0, 0, 1, 1, 1, 3, 4, 4, 5, 5, 4, 3, 2, 3, 4, 4, 2, 1, 0, 0, 2, 0, 1, 2, 3, 3, 1, 1, 2, 1, 0, 0, 0, -1, -1, 0, 1, 2, 3, 4, 4, 5, 5, 6, 4, 3, 3, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 3, 2, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 4, 4, 4, 5, 4, 3, 3, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 3, 4, 4, 3, 1, 0, 0, 0, 0, 0, 0, 1, 3, 3, 2, 3, 3, 2, 0, 0, 1, 0, 0, 1, 1, 3, 2, 3, 1, 2, 2, 2, 3, 2, 3, 1, 1, 0, -1, 0, 1, 2, 3, 4, 4, 4, 4, 4, 4, 4, 1, 3, 2, 1, 1, 0, 2, 3, 2, 3, 3, 4, 3, 2, 2, 2, 2, 0, 0, 0, 0, 2, 2, 3, 5, 5, 5, 5, 5, 6, 7, 6, 5, 4, 4, 4, 2, 1, 1, 2, 2, 3, 3, 2, 3, 3, 3, 4, 5, 0, -1, 0, 2, 3, 3, 4, 4, 3, 4, 4, 4, 5, 8, 6, 6, 4, 5, 4, 2, 1, 1, 1, 0, 1, 1, 2, 2, 3, 3, 3, 3, 0, 0, 0, 2, 3, 4, 2, 2, 2, 4, 4, 5, 3, 4, 4, 4, 3, 3, 4, 2, 4, 3, 3, 1, 1, 2, 3, 2, 1, 3, 2, 2, 0, 0, 0, 0, 2, 0, 0, 2, 4, 3, 5, 4, 4, 3, 1, 2, 0, 0, 2, 2, 4, 4, 3, 2, 1, 2, 1, 1, 2, 3, 4, 2, 1, 1, 0, 0, 1, 0, 0, 0, 2, 2, 4, 2, 2, 3, 3, 1, 1, 1, 3, 4, 4, 5, 4, 1, 2, 1, 1, 3, 2, 3, 4, 4, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 3, 2, 2, 1, 2, 1, 0, 0, 1, 1, 3, 2, 3, 2, 3, 2, 2, 4, 6, 5, 5, 2, 0, 0, 0, -1, 1, 2, 2, 1, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 1, 3, 4, 3, 3, 2, 2, 2, 2, 0, 0, 0, -1, 0, 0, 2, 1, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 1, 2, 3, 1, 1, 1, 0, 1, 0, 0, 0, -4, -2, -2, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 2, 2, 2, 1, 2, 1, 0, 0, 1, 2, 0, -1, 0, 0, -1, -1, -1, -3, -1, -1, 0, 0, 0, 1, 1, 3, 2, 1, 0, 0, 2, 0, 1, 2, 1, 2, 3, 1, 1, 2, 1, 2, 2, 2, 0, 0, -1, -2, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 2, 2, 2, 0, 2, 1, 0, -1, 0, 1, 2, 1, 1, 3, 3, 4, 2, 1, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, -2, -1, -2, 0, 0, 1, 2, 2, 3, 2, 2, 2, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 1, 1, 1, 2, 0, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 1, 2, 0, 1, 1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 2, 2, 2, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 2, 0, 0, 2, 2, 2, 1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 2, 1, 2, 2, 0, 1, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 2, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 1, 1, 1, 1, 2, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 0, 1, 1, 1, 1, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 2, 2, 0, 0, 0, 1, 1, 1, 1, 3, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 1, 0, 1, 3, 2, 2, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 2, 1, 1, 1, 2, 0, 1, 1, 2, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 2, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -2, -1, -1, -1, -2, -2, -1, -1, -2, -2, -2, -1, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 2, 1, 1, 1, 1, 0, 0, 0, 1, 1, 0, -1, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 1, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 2, 2, 3, 2, 1, 1, 0, -1, 0, 1, 1, 1, 0, 1, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 2, 3, 2, 1, 0, 0, 0, 0, 0, 1, 2, 0, 2, 2, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 2, 1, 2, 1, 0, 0, 1, 0, 0, 1, 2, 2, 2, 1, 2, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 2, 1, 1, 2, 2, 3, 2, 0, 0, 0, 0, 0, 1, 2, 3, 2, 2, 1, 2, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 2, 1, 1, 2, 2, 0, 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 0, 0, 0, -1, 0, 2, 1, 1, 1, 2, 0, 2, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 2, 0, 0, -1, 0, 2, 1, 2, 1, 0, 2, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 1, 2, 1, 0, 1, 0, 0, -1, 0, 1, 0, 0, 2, 1, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 2, 2, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 2, 1, 1, 1, 0, -1, 0, 0, -1, -1, 0, 1, 2, 1, 2, 0, 1, 1, 1, 1, 1, 1, 1, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 2, 2, 0, 1, 1, 1, 1, 1, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 2, 1, 0, 2, 1, 0, 1, 0, 0, 0, -1, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 2, 0, 0, 0, -1, -1, 0, 0, 0, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, -2, -2, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -2, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, -2, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -2, -1, -1, -2, 0, -2, -1, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, -1, -1, -2, -1, 0, -2, -2, -1, -1, -3, -1, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -3, -3, -2, -2, -2, -1, 0, 0, -1, 0, -1, 0, 0, 2, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -4, -3, -3, -2, -4, -3, -2, -2, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -2, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 2, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 2, 0, 0, 0, 0, 1, 1, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -2, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, -2, -2, -1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 1, 2, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, -1, -1, 0, 0, 1, 0, -1, -2, 0, 0, 0, 2, 3, 2, 1, 2, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, -2, -1, 0, 0, 1, -1, -1, -1, 0, 0, 1, 2, 3, 2, 2, 1, 0, -1, -2, -2, -1, 0, 0, 0, 0, 2, 2, 3, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, -1, 0, 0, 0, 2, 3, 3, 4, 2, 1, 0, -1, -3, -3, -2, 0, -1, 0, 1, 1, 2, 2, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, -1, 0, 0, 0, 2, 3, 4, 4, 2, 0, -1, 0, -2, -2, -3, -2, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 3, 3, 4, 3, 1, 1, 0, 0, -1, -1, -2, -2, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 2, 3, 4, 2, 1, 1, 0, 0, -2, 0, -2, -1, -1, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, -1, 0, -2, -1, -1, 0, 0, 2, 3, 3, 3, 2, 1, 1, -1, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, -2, -2, -1, 1, 0, 2, 5, 3, 1, 2, 0, 0, -1, 0, -1, -2, -2, -1, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, -1, -1, 0, -1, -1, -2, 0, 0, 0, 2, 2, 2, 0, 0, 1, 0, 0, 0, -1, -3, -2, -1, -2, 0, 0, 2, 2, 1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -2, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -3, -2, -3, -2, -1, 0, 2, 1, 2, 2, 1, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, -1, 0, 2, 1, 0, 1, 1, 1, 0, -2, -3, -2, -3, -3, -1, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -2, 0, 0, 1, 0, 0, 1, 1, 0, -1, -2, -1, -1, -1, 0, 0, 0, 2, 1, 1, 1, 1, 0, 1, 0, -1, 0, 0, 0, -1, -1, 0, -3, -1, 0, 1, 2, 1, 2, 1, 0, -2, -2, -1, 0, -1, 0, 1, 1, 0, 1, 0, 1, 0, 1, 1, 0, -1, 0, 0, 0, -1, 0, 0, -3, -2, 0, 0, 1, 2, 1, 1, 0, -1, -1, -1, 0, 1, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -4, -3, -1, 0, 0, 2, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 1, 2, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -4, -2, -1, 0, 0, 1, 0, 2, 0, 0, -1, 1, 1, 2, 1, 1, 1, 0, 2, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, 2, 1, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -2, -1, 0, 0, 0, 2, 2, 0, 1, 1, 0, 1, 2, 0, 1, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, -1, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -2, -1, 0, -1, 0, -2, -1, -1, -2, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, -1, -1, -2, -1, -2, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, -1, 0, -1, -2, -2, -1, -1, -1, -1, -2, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, -2, 0, 0, -2, -1, 0, -1, -1, 0, -1, -1, 0, 0, -2, -1, -1, -1, -2, -1, -2, -1, -1, 0, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, -1, -2, -2, -1, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, -2, -1, -3, -1, -2, -2, -2, -1, -1, -1, 0, 0, -1, 1, 0, 0, 0, -1, -2, -2, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, -1, -2, -2, -1, -2, -1, -1, 0, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -2, -2, -3, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, 0, 0, -1, -1, -1, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, -2, -1, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 2, 0, 1, 0, -1, 0, 0, -1, -1, -2, -2, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -2, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, -2, -2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -2, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -2, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -2, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, 0, 1, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 1, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, -2, -1, -1, -2, 0, -2, -1, 0, 0, 0, -2, -1, 0, 0, -1, -1, -1, -1, -2, 0, -1, -3, -1, 0, -2, -2, -1, -2, -2, -1, 0, -2, -2, -1, -3, -3, -3, -2, -2, -1, 0, -1, -2, -1, 0, -1, -2, -1, -2, -2, -3, -3, -4, -4, -1, 0, -2, -2, -1, -1, -2, 0, 0, -1, -2, -2, -3, -4, -2, -3, -3, -2, -1, -1, -1, -2, -2, -3, -2, -1, -1, -2, -2, -2, -5, -4, -1, -1, -2, -1, -1, -1, -3, -2, 0, -2, -2, -2, -4, -4, -2, -4, -3, -2, -2, -1, -1, -2, -2, -2, -1, -2, -2, -2, -2, -3, -4, -3, -2, 0, 0, 0, 0, 0, -1, -2, 0, -2, -2, -4, -3, -4, -3, -4, -2, -3, -4, -3, -2, -1, -2, -2, -1, 0, -2, -3, -3, -3, -3, -2, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, -4, -3, -4, -3, -3, -4, -2, -3, -4, -2, -1, -2, -2, -1, 0, -4, -3, -3, -3, -3, -1, -2, 0, 1, 0, 0, 0, 0, -1, 0, -2, -2, -3, -1, -2, -4, -4, -3, -1, -2, -4, -4, -3, -2, -1, -2, -1, -2, -4, -5, -3, -4, 0, 0, 0, 1, 1, 1, 1, 0, 0, -1, -1, -2, -2, -1, -2, -2, -4, -4, -2, -2, -4, -5, -2, -1, -2, -3, -1, -3, -3, -5, -3, -3, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, -2, -2, -1, -1, -1, -2, -3, -3, -3, -2, -3, -4, -3, -2, -2, -2, -1, -2, -4, -4, -4, -3, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, -2, -3, -4, -3, -2, -2, -2, -1, -3, -3, -2, -3, -3, -2, -3, -2, 0, 0, 0, 0, 2, 1, 1, 0, 0, 3, 2, 0, 0, 0, 1, 0, -1, -2, -3, -4, -2, -1, 0, -2, -2, -3, -1, -3, -3, -1, -3, -2, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 3, 1, 1, 0, 0, 0, 0, -1, -2, -4, -4, -2, -1, -2, -3, -2, -2, -2, -3, -1, -4, -2, 0, -1, 0, 0, 1, 3, 3, 3, 2, 3, 3, 2, 1, 1, 1, 0, 0, 0, -1, -2, -4, -3, 0, -1, -2, -1, -2, -3, -2, -2, -3, -1, 0, -1, 0, 2, 3, 1, 2, 3, 3, 4, 4, 2, 0, 2, 2, 0, 0, 0, 0, -1, -3, -2, -2, -2, -1, -2, -2, -2, -3, -2, -3, 0, 0, -1, 0, 1, 2, 1, 3, 3, 1, 3, 2, 3, 0, 2, 2, 0, 1, 0, -1, -2, -1, -2, -1, -2, -1, 0, -2, -3, -2, -1, 0, -1, 0, -1, 0, 2, 2, 1, 3, 3, 1, 1, 2, 3, 1, 1, 1, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, -3, -2, -3, -3, 0, -1, 0, -1, 0, 2, 2, 1, 3, 3, 2, 1, 3, 3, 0, 3, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, -3, -3, -2, -2, 0, 0, 0, -2, 0, 1, 0, 2, 1, 2, 2, 2, 3, 4, 1, 2, 1, 0, 1, 1, 0, -1, -2, -3, -2, -1, 0, -3, -3, -1, -2, 0, 0, 1, 0, -2, 0, 1, 0, 1, 0, 0, 2, 3, 2, 3, 3, 1, 1, 0, 0, 1, 0, 0, -1, -1, -2, -1, -2, -3, -3, -3, -1, 0, 0, 0, 0, -1, 0, 0, 2, 1, 0, 0, 1, 4, 3, 3, 3, 1, 0, 0, 0, 0, 0, -2, -2, -2, 0, -1, -3, -3, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 2, 2, 2, 3, 3, 0, -1, 0, 0, 0, -2, -4, -2, -1, 0, -2, -3, -2, -2, -1, -3, -1, 0, -1, -1, 0, 0, 1, 2, 1, 0, 0, 1, 1, 1, 3, 3, 0, 0, -1, 0, 0, -2, -3, -1, 0, 0, -1, -2, -3, -1, -3, -3, -1, -2, -2, -2, -1, 0, 0, 0, 2, 0, 1, 0, 0, 1, 2, 2, 0, -2, -2, 0, 0, -3, -3, -2, 0, 0, 0, -1, -3, -3, -3, -2, 0, -1, -3, -2, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 2, 1, -1, -4, -1, -2, -1, -3, -4, -2, 0, 0, -2, -1, -1, 0, -2, -3, -2, -1, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, -3, -4, -2, 0, -2, -3, -3, -3, -1, -2, -3, -2, 0, 0, 0, -2, -1, -2, 0, 0, -2, 0, -1, -1, 1, 0, -2, 0, 0, 1, 0, -2, -3, -3, -4, -1, -3, -2, -4, -3, -2, -2, -3, -2, 0, 1, 0, -1, -2, -2, -1, 0, -2, 0, -1, 0, 0, 0, -2, 0, 0, 0, 0, -3, -3, -3, -3, -1, -1, -3, -3, -3, -2, -2, -2, -3, 0, 0, 0, 0, -1, -3, 0, -1, -2, 0, -1, 0, 1, -1, -3, -2, 0, 0, 0, -1, -3, -2, -2, -2, 0, -3, -2, -3, -3, -3, -3, -2, 0, 0, 0, -1, -1, -2, 0, 0, -1, 0, -1, -1, 0, 0, -1, -2, 0, 0, 0, -2, -3, -2, -3, -1, -1, -1, -3, -1, -3, -2, -3, -3, 0, -1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -3, -3, -1, -2, -2, 0, -2, -3, -2, -3, -3, -2, -2, -1, 1, -1, -1, 0, -2, -1, 0, 0, 0, -1, -1, 0, 0, 0, -2, 0, -1, -1, -1, -1, -1, -2, -2, 0, -1, -2, -1, -2, -1, -2, -2, 0, 0, 0, 0, -1, -1, -1, 0, -2, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, -1, -1, -3, -2, -2, -1, -1, -2, 0, -1, 0, -1, -3, -4, -2, -4, -5, -4, -6, -5, -5, -5, -5, -5, -3, -2, 0, -2, -2, -1, 0, 0, 0, -2, -1, -1, -2, -1, -1, 0, -1, 0, -1, 0, -2, -2, -3, -2, -4, -4, -3, -4, -5, -4, -3, -3, -2, -2, 0, -1, -2, -2, -1, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, -1, -1, -2, -1, -1, -2, -1, -3, -2, -2, -3, -2, -3, -2, -1, -3, -1, 0, -2, -3, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, -2, -1, 0, -1, 0, -1, -1, -2, -1, -3, -2, -2, -2, -3, -2, -2, -3, -1, -2, 0, -2, -3, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, -2, 0, -1, 0, -1, -2, -1, -2, 0, -1, 0, -2, -2, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 2, 2, 1, 0, 1, 1, 2, 2, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 1, 1, 1, 3, 3, 2, 3, 2, 2, 2, 0, 1, 1, 1, 1, 0, 0, 2, 1, 1, 2, 1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 1, 1, 2, 2, 1, 1, 1, 1, 0, 1, 1, 0, 1, 1, 2, 0, 0, 0, -1, -1, -1, 0, 1, 0, 2, 2, 2, 2, 2, 2, 2, 3, 2, 2, 2, 2, 4, 2, 2, 0, 1, 2, 0, 1, 1, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 3, 3, 2, 2, 2, 3, 1, 1, 2, 3, 3, 2, 3, 2, 1, 1, 0, 1, 1, 1, 1, 3, 1, 0, 0, 0, -1, 0, 1, 1, 2, 3, 3, 3, 2, 1, 0, 0, 1, 2, 2, 2, 3, 4, 4, 3, 1, 1, 1, 2, 0, 1, 0, 2, 0, 0, 0, 0, 0, 1, 1, 2, 2, 3, 3, 3, 3, 2, 1, 0, 0, 2, 3, 1, 2, 3, 3, 2, 1, 2, 2, 2, 2, 2, 0, 1, 0, 0, -1, 0, -1, 1, 3, 3, 3, 2, 2, 3, 3, 3, 3, 0, 1, 0, 2, 2, 2, 3, 3, 1, 1, 1, 1, 1, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 1, 3, 2, 3, 2, 2, 2, 3, 3, 3, 3, 1, 1, 2, 3, 2, 2, 1, 1, 1, 1, 1, 0, 1, 2, 2, 1, 0, 0, 0, 0, 0, 1, 3, 2, 2, 1, 3, 3, 3, 2, 2, 2, 2, 1, 2, 1, 2, 2, 2, 1, 1, 1, 0, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 2, 2, 3, 4, 2, 3, 2, 2, 3, 2, 1, 1, 2, 2, 1, 2, 1, 2, 2, 2, 2, 1, 2, 1, 0, 0, -1, -1, -1, 0, 0, 0, 2, 4, 3, 4, 5, 5, 4, 2, 5, 2, 2, 2, 1, 2, 2, 2, 1, 1, 1, 2, 2, 1, 2, 1, 0, 0, -1, -1, 0, 0, 0, 0, 2, 3, 3, 3, 3, 3, 2, 3, 3, 4, 3, 2, 2, 0, 2, 2, 2, 1, 0, 0, 0, 2, 1, 1, 0, -1, -1, -1, 0, 0, 0, 0, 2, 3, 4, 3, 2, 4, 3, 3, 3, 2, 1, 1, 0, 0, 1, 2, 2, 1, 1, 1, 2, 2, 1, 0, 0, 1, 0, 0, -1, -1, -1, 0, 1, 1, 3, 4, 3, 4, 2, 2, 2, 2, 2, 0, 0, 0, 1, 3, 2, 2, 2, 1, 2, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 3, 4, 4, 2, 1, 1, 2, 1, 1, 1, 2, 3, 3, 1, 2, 2, 1, 2, 2, 1, 2, 0, 0, 1, 0, 0, 0, -1, 0, 1, 1, 2, 3, 4, 2, 1, 1, 1, 1, 2, 1, 2, 3, 3, 2, 2, 2, 0, 1, 1, 1, 1, 1, 0, 1, 0, 0, -1, -2, 0, -1, 0, 0, 1, 2, 2, 2, 1, 1, 0, 0, 1, 1, 2, 2, 1, 2, 2, 1, 2, 1, 1, 0, 1, 0, 1, 1, 0, -1, 0, -2, -2, -1, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 2, 1, 3, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -2, -2, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 2, 3, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 2, 0, 1, 2, 1, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, -1, -2, -1, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -2, -1, -2, -1, 0, 0, -2, -1, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -2, -1, -2, -1, -2, -2, -1, -1, -1, -1, -1, -2, 0, -1, -1, -1, -1, -1, 0, 0, -1, 0, -2, -1, 0, 0, -2, -1, -1, -1, -1, -1, -1, 0, 0, -1, -2, -2, -1, 0, -1, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, 0, -2, -2, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 1, 1, 2, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 1, 1, 2, 1, 1, 2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 2, 2, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -2, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -2, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 2, 1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 1, 0, 0, 1, 0, 1, 1, 1, 1, 0, 1, 0, 0, 2, 1, 2, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 1, 0, 1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 2, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, 2, 1, 1, 1, 1, 0, 0, 1, 0, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 1, 2, 1, 1, 0, 1, 0, 1, 0, 1, 0, 1, 2, 1, 2, 1, 0, 0, 1, 1, 1, 1, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, 2, 1, 1, 2, 1, 1, 1, 1, 1, 0, 1, 0, 1, 0, 1, 2, 0, 1, 1, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 0, 0, 1, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, -2, -1, -1, -2, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, -2, -2, -1, -1, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, -2, 0, 0, 0, -1, 0, -1, -2, -2, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -2, 0, -1, -2, -1, 0, -1, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -2, -1, -2, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -1, -2, -1, 0, -2, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 2, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -2, -1, -1, -2, -2, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -3, -2, -2, -1, -2, -1, 0, -1, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, -1, -1, -2, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, -1, 0, -1, -1, -1, 0, -1, 0, -1, -1, -1, 0, -2, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 2, 2, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 2, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 1, 2, 1, 0, 1, 2, 1, 0, 0, 1, 1, 1, 1, 2, 0, 2, 1, 1, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 1, 1, 2, 0, 1, 1, 1, 1, 2, 2, 2, 1, 1, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 1, 0, 1, 1, 2, 1, 2, 0, 2, 0, 2, 1, 2, 0, 1, 2, 1, 1, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 1, 1, 0, -1, -1, -1, -1, 0, -1, 0, -2, -2, -3, -2, -2, -2, -2, -1, -2, -2, -3, -3, -5, -5, -5, -6, -6, -6, -7, -7, -8, -6, -4, -3, 0, 0, -2, -3, -2, -1, -2, 0, -2, -1, -1, -2, -1, -2, -1, -1, -2, -2, -3, -4, -5, -4, -4, -6, -6, -6, -6, -7, -7, -5, -4, -3, 0, -2, -3, -4, -3, -3, -2, -2, -3, -2, -2, -2, -1, -3, -2, -3, -2, -4, -4, -3, -3, -4, -4, -6, -6, -5, -5, -6, -6, -5, -5, -4, -1, 0, -3, -4, -4, -2, -2, -1, -1, -2, 0, -2, -1, -2, -2, -3, -3, -3, -2, -3, -2, -4, -3, -4, -5, -4, -4, -5, -6, -6, -4, -4, -2, -2, -3, -4, -2, 0, -1, 0, -1, 0, -1, -1, -2, 0, -2, -3, -2, -1, -1, -3, -2, -2, -2, -4, -4, -3, -2, -4, -3, -3, -3, -3, -2, -1, -2, -3, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -3, -3, -1, -1, -1, 0, -2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 2, 2, 1, 0, 1, 1, 0, -1, -1, -3, -2, 0, 0, -1, 0, -1, 0, 1, 1, 2, 2, 1, 0, 2, 0, 1, 1, 2, 3, 1, 1, 0, 1, 3, 3, 2, 4, 1, 0, 0, -1, -2, -2, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 2, 0, 2, 2, 3, 3, 2, 1, 1, 1, 3, 2, 4, 3, 3, 1, 0, -1, -1, -2, -1, 0, 1, 1, 1, 1, 1, 2, 2, 0, 1, 1, 0, 0, 1, 2, 4, 4, 5, 3, 3, 1, 2, 2, 4, 5, 4, 2, 0, -1, 0, -1, 0, 1, 2, 3, 2, 1, 1, 1, 1, 0, 0, 1, 1, 0, 1, 3, 4, 6, 5, 4, 3, 3, 3, 2, 3, 4, 3, 1, 1, -1, 0, 0, 1, 2, 3, 3, 4, 4, 1, 0, 0, 0, 0, 0, 1, 2, 2, 3, 4, 4, 5, 3, 4, 3, 4, 2, 4, 4, 4, 2, 0, 0, 0, 0, 1, 4, 5, 5, 5, 5, 3, 1, 0, 0, 0, 0, 0, 0, 2, 4, 3, 5, 5, 4, 3, 2, 3, 2, 2, 3, 2, 2, 0, -1, 1, 0, 2, 4, 7, 7, 7, 4, 3, 4, 1, 1, 1, 0, 0, 0, 2, 3, 2, 4, 3, 2, 3, 2, 2, 1, 2, 2, 3, 2, 0, 0, 0, 0, 2, 5, 6, 7, 5, 4, 4, 2, 2, 2, 1, 0, 1, 1, 2, 3, 3, 3, 2, 3, 2, 2, 1, 2, 2, 2, 1, 1, 0, 0, 0, 1, 1, 3, 6, 6, 6, 5, 3, 3, 1, 2, 1, 1, 1, 0, 1, 0, 1, 2, 2, 2, 2, 2, 3, 2, 2, 2, 0, 0, 0, -1, 0, 0, 1, 4, 7, 6, 6, 6, 5, 3, 2, 1, 1, 0, 0, 1, 0, 1, 0, 1, 2, 3, 2, 2, 2, 4, 3, 1, 0, 0, -2, -1, 0, 0, 2, 4, 5, 7, 7, 5, 4, 5, 2, 2, 3, 0, -1, 0, 1, 1, 1, 2, 1, 0, 3, 3, 3, 2, 2, 2, 0, -1, -1, -2, 0, 0, 1, 3, 5, 5, 5, 4, 3, 2, 2, 2, 1, 1, -1, 0, 0, 0, 1, 2, 1, 1, 2, 2, 3, 4, 3, 3, 1, -2, -1, -1, 0, -1, 1, 3, 3, 4, 3, 3, 2, 2, 1, 2, 0, -1, -1, 0, 0, 1, 3, 4, 2, 2, 3, 4, 4, 5, 4, 3, 0, 0, -1, 0, 0, -2, 0, 1, 3, 4, 4, 3, 5, 2, 0, 0, 0, -2, 0, -2, 0, 2, 3, 4, 4, 4, 2, 2, 5, 3, 2, 3, 0, 0, 0, 0, -1, -3, -2, -1, 0, 2, 2, 4, 4, 2, 2, 0, 0, 0, 0, 0, 0, 3, 3, 4, 5, 3, 2, 3, 4, 3, 3, 3, 1, 0, 0, 0, 0, -3, -3, -2, 0, 0, 2, 3, 3, 3, 0, 0, 0, 0, 0, 1, 2, 3, 3, 3, 4, 4, 1, 2, 4, 2, 1, 1, 1, 0, 0, 0, -2, -4, -5, -2, -1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 2, 1, 1, 3, 3, 3, 3, 5, 5, 4, 3, 2, 1, 1, 0, -1, 0, -2, -4, -5, -3, -2, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 1, 3, 3, 3, 3, 5, 2, 1, 0, 0, -1, -1, 0, -1, -2, -5, -6, -5, -4, -3, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 1, 1, 2, 2, 3, 1, 2, 1, 1, 0, -2, -1, 0, 0, -1, -5, -6, -4, -4, -3, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 1, 1, 1, 1, 2, 2, 0, 0, 0, 0, -2, -1, -1, -2, -1, -3, -4, -4, -4, -3, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -2, -1, -1, -2, -2, -3, -4, -4, -3, -4, -2, -1, -1, -1, -1, -2, -1, -1, -1, -2, -1, -1, -2, -1, 0, -1, -1, -1, 0, -2, -2, -3, -2, -2, -2, -2, -1, -4, -3, -4, -4, -3, -3, -2, -2, -1, -1, -1, -1, -2, -1, 0, -1, -1, -1, -2, -3, -2, -4, -2, -3, -4, -6, -5, -4, -4, -4, -3, -1, -2, -4, -3, -3, -1, -3, -1, -1, -1, -2, -1, -1, -1, -1, -2, -1, -2, 0, -1, -2, -3, -5, -4, -3, -5, -4, -5, -5, -3, -2, -2, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 2, 1, 2, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, -2, -1, -1, 0, -1, -2, 0, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -2, -1, -2, -2, -1, -1, 0, 0, -1, -2, 0, -1, -1, -2, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, -2, -2, -2, -3, -1, -2, 0, 0, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -1, -2, -2, -2, -2, 0, -1, -1, -1, -1, -1, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -2, -3, -2, -1, -1, -2, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -2, 0, -1, 0, -2, -2, 0, -1, -3, -2, -1, -1, 0, 0, -1, 0, -1, -2, -1, -1, -2, -2, -1, -2, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -2, -2, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, -2, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -2, 0, 0, -2, -1, 0, -1, -1, 0, 0, 0, -1, -1, -1, -1, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, -2, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -2, -2, -1, -2, 0, -1, -1, -2, -1, -1, -1, -1, 0, -1, -1, -1, -2, -1, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, -1, -1, -2, -1, -1, -2, -2, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, -1, -2, 0, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, -1, -2, -2, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -2, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -2, -1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, -2, -3, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, -1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, -2, -3, -1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 1, 1, 2, 2, 0, 0, 2, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, -1, -2, -2, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -2, 0, 0, -1, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 0, -1, -2, -2, -2, -1, -2, -2, -1, -2, 0, -1, -1, -2, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 1, 0, 1, 0, -2, -3, -2, -2, -2, -2, -1, -2, 0, -1, -1, -1, -2, -2, -1, -1, -2, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -2, -3, -2, -2, -2, -1, -1, -1, 0, 0, -1, -2, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 1, 0, 0, -3, -3, -2, -1, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 2, 1, 1, 1, 1, 1, 0, -2, -2, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 2, 2, 1, 0, 1, 0, -2, -3, -2, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, -2, -2, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 1, 0, 0, 0, 2, 2, 1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, -2, -2, -1, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, -1, -2, -1, -1, -2, -1, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -3, -1, -2, -2, -1, -2, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, -1, 0, 0, 2, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, -1, -2, -2, -1, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 0, -1, 0, 0, 1, 2, 0, 0, -1, 1, 1, 2, 1, 1, 0, 0, 0, -2, -1, 0, -1, -2, 0, 0, 0, -1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 1, 1, 3, 1, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 3, 2, 3, 1, 1, 1, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 3, 1, 2, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 2, 2, 3, 3, 2, 0, 1, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 2, 1, -1, 0, 0, 0, 1, 0, 2, 2, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 2, 1, -1, -1, -1, 0, 0, 0, 0, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 2, 1, 2, 1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 1, 2, 1, 1, 0, 3, 3, 1, 0, -2, -1, 0, -1, -1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 0, 1, 1, 1, 2, 1, 0, 0, 0, -1, -2, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, -1, -1, 0, 0, 0, 1, 2, 2, 2, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, -1, -1, -1, 0, -1, -1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 1, 1, 2, 0, 0, 1, 0, 0, 0, 1, 1, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 0, 1, 1, 1, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 1, 2, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, -2, -1, -1, -1, -1, -1, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, -1, -2, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, -1, -2, -2, -1, -2, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, -1, -3, -4, -3, -2, -2, -2, -1, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, -1, -4, -3, -3, -2, -2, -2, 0, 1, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 2, 3, 2, 1, 0, 0, -2, -3, -5, -5, -3, -2, -3, -1, 0, 1, 2, 0, 1, 2, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 3, 3, 1, 2, 0, 0, -3, -3, -4, -2, -3, -2, -1, 0, 0, 1, 1, 2, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 2, 3, 2, 2, 1, 0, -1, -1, -4, -3, -4, -2, -2, -2, 0, 0, 0, 1, 1, 1, 1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 3, 2, 1, 2, 2, 0, 0, -1, -3, -3, -4, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 3, 1, 2, 2, 0, 0, -1, -2, -3, -2, -3, -1, 0, 0, 0, 1, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 3, 2, 1, 1, 0, -1, -1, -3, -3, -3, -2, -1, -1, 0, 1, 1, 2, 0, 1, 0, -1, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 2, 2, 1, 2, 2, 1, -1, -2, -3, -3, -3, -3, -2, -2, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -3, -4, -2, -3, -3, -2, -1, -1, 1, 1, 2, 1, 0, -1, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, -2, 1, 0, 0, 1, 1, 0, 0, -2, -1, -2, -3, -2, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 2, 0, 0, -1, -2, -2, -1, 0, -1, -1, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, -3, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, -4, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 1, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 2, 1, 1, 0, 1, 2, 2, 0, 1, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -3, -1, 0, 0, 1, 2, 2, 1, 1, 2, 1, 1, 1, 1, 2, 1, 2, 2, 2, 2, 2, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -2, -1, 0, 1, 0, 2, 3, 1, 1, 2, 2, 2, 1, 3, 2, 3, 2, 1, 3, 3, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 2, 1, 2, 2, 2, 2, 3, 1, 3, 3, 2, 3, 2, 3, 2, 2, 2, 2, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 2, 2, 3, 2, 1, 1, 2, 1, 1, 2, 2, 2, 3, 2, 2, 2, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 2, 0, 1, 1, 0, 1, 1, 1, 1, 2, 0, 2, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, -2, -1, -1, 0, 0, -1, -1, -2, -3, -2, -1, -2, -2, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, -1, -2, -2, -1, 0, -1, -2, -1, -1, -2, -2, 0, 0, 0, -2, -1, -1, -2, -1, -2, -1, -1, 0, 0, 0, 0, -1, -1, -2, 0, -1, -2, -2, -2, -3, -3, 0, 0, -2, 0, 0, -2, -1, 0, 0, 0, -1, -2, -3, -3, -1, -3, -1, -2, -1, -1, 0, 0, -1, -2, -1, -1, -1, -2, -1, -2, -3, -1, 0, -1, 0, -1, -1, -1, -1, -1, 0, 0, -1, -1, -2, -2, -2, -4, -2, -3, -2, -1, -1, -1, -1, -2, 0, -1, 0, 0, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, -2, -2, -2, -3, -4, -1, -1, -3, -1, -1, -2, -1, 0, -1, 0, -1, 0, -1, -1, -3, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -3, -1, -3, -2, -3, -1, 0, -2, -2, -2, -1, 0, 0, 0, 0, 0, -2, -2, -2, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, -2, -1, -2, -2, -1, -1, -2, -3, -1, -1, -3, -3, -3, -1, -1, 0, 0, 0, -1, -2, -4, -2, 0, 1, 0, 1, 0, 1, 2, 0, 0, 0, 0, -1, -2, -1, 0, 0, -2, -1, -1, -2, -2, -3, -3, -2, -1, 0, -2, -1, -1, -1, -3, -3, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, -2, -2, -3, -2, -2, -3, -3, -2, -3, 0, -1, -1, -2, -2, -2, -1, 0, 0, 0, 1, 1, 2, 0, -1, 0, 2, 0, -1, 0, 0, 0, 0, -1, -1, -3, -2, -2, -2, -1, -1, -3, -2, -2, -1, -1, -1, -3, -1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 2, 2, 0, -1, 0, 0, 0, -1, -1, -1, -3, -3, -2, -1, -1, -2, -2, -1, -3, -1, -1, -2, -1, -1, 0, 0, 2, 1, 0, 2, 2, 2, 3, 2, 0, 0, 1, 0, 0, -1, -1, -2, -3, -3, 0, -1, -1, -1, -1, -1, -3, -1, -2, -2, 0, 0, 0, 0, 2, 1, 3, 3, 3, 2, 3, 2, 0, 0, 0, 0, -1, 0, -2, -1, -2, -2, -2, -1, -1, 0, 0, -1, -1, -1, -1, -2, 0, 0, 0, 0, 2, 0, 1, 2, 3, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -2, -2, -1, -1, -1, 0, -1, -2, -2, -2, -2, -1, 1, 0, 0, 0, 2, 2, 2, 2, 2, 0, 0, 2, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, -2, -1, 0, 0, 0, -2, -1, -1, -2, 0, 2, 0, 0, 0, 2, 0, 1, 3, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, -1, 0, -1, -1, -2, -2, 0, 0, -1, -3, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 1, 0, 2, 1, 0, 1, 0, -1, 0, 0, -1, -1, -1, -2, -1, -1, 0, -2, -3, 0, 0, 0, 0, 1, -2, 0, 0, 0, 0, 1, 1, 1, 1, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -1, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 2, 2, 0, 2, 2, 1, 0, 2, 1, 0, -1, -1, 0, -1, -1, -2, -1, -1, -1, -2, -2, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 1, 2, 1, 0, 0, 1, 2, 1, 2, 2, 0, 0, 0, 0, 0, -2, -3, 0, 0, 0, -1, -3, -1, 0, -2, -2, 0, -2, -3, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 2, 2, 1, 0, -1, 0, 0, -1, -3, -3, 0, 0, 0, -2, -3, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 2, 2, 1, -1, -1, -1, 0, -1, -3, -3, -1, 0, 0, -1, -2, -2, -2, -1, -3, 0, 0, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 0, -2, -1, -3, 0, -1, -2, -2, -1, -1, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 2, 0, -1, 0, 0, 2, 1, -1, -2, -2, -3, -2, -3, -2, -3, -2, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 1, 1, 0, 0, -2, 0, 0, -1, 0, 0, 0, 2, 0, -1, -2, -4, -1, -1, -1, -1, -3, -2, -1, -1, -2, -1, 0, 0, 0, -1, -1, -2, 1, 0, 0, -1, -1, 1, 1, -1, -2, 0, 0, 0, 0, -1, -3, -2, -2, 0, -2, -2, -2, -3, -2, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, -1, 0, 1, -1, -2, 0, 0, 0, -1, -2, -1, -2, -2, 0, -1, -1, -2, -2, -2, -1, -1, -1, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, -1, -1, -2, -1, -1, 0, 0, -2, -2, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -2, -1, 0, 0, -1, -2, 0, -1, -1, -3, -1, -2, -2, -1, -1, -2, -2, -2, -3, -2, -2, -2, 0, 1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -2, 0, -2, -1, -1, -1, 0, -1, -1, -1, 0, -2, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 1, 2, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -2, -1, -1, -2, -1, 0, -1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, -2, -2, -2, -3, -2, -2, -2, -2, -2, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -1, -1, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -2, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -2, -2, -2, -3, -3, -2, -2, -1, -1, 0, -1, 0, 0, -1, 0, 0, 2, 1, 0, 2, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -2, -3, -3, -2, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 2, 0, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 0, 0, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 2, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 2, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, 1, 1, 1, 4, 2, 1, 0, 1, 2, 0, 0, 0, 1, 0, 0, -1, -2, 0, 0, 1, 2, 2, 1, 0, -1, 0, 0, 1, 1, 0, 1, 1, 1, 0, 1, 3, 4, 2, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 2, 3, 2, 2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 2, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 3, 1, 1, 2, 0, 1, 2, 0, 1, 2, 2, 1, 1, 0, 1, 2, 1, 0, -1, 0, 0, 0, 2, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 3, 1, 1, 1, 0, 1, 2, 2, 2, 2, 2, 1, 3, 1, 1, 0, 0, 0, 0, 2, 0, 1, 1, 2, 1, 1, 1, 1, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 2, 1, 3, 2, 1, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 1, 2, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 1, 1, 1, 2, 2, 1, 1, 2, 0, 1, 0, 0, -1, 0, -1, 1, 0, 2, 2, 2, 1, 0, 0, 2, 1, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 1, 2, 1, 0, 0, 0, 1, 3, 2, 0, 1, 0, 0, 2, 0, 1, 0, 0, 0, 0, 1, 1, 1, 3, 2, 3, 3, 2, 1, 1, 0, 1, 0, 2, 2, 2, 0, 0, 0, 0, 3, 3, 3, 1, 0, 0, 2, 1, 1, 0, 1, 0, 1, 1, 1, 4, 3, 4, 4, 1, 2, 3, 3, 2, 2, 2, 1, 2, 1, 0, -1, 0, 1, 1, 1, 1, 2, 0, 1, 2, 0, 0, 1, 0, 2, 4, 3, 4, 3, 4, 2, 2, 1, 1, 2, 3, 1, 2, 2, 4, 3, 1, 0, -1, 0, 0, 1, 1, 2, 1, 1, 0, 1, 1, 0, 0, 2, 3, 4, 3, 3, 3, 2, 3, 1, 1, 0, 1, 1, 1, 1, 1, 2, 1, 0, 1, 1, 1, 1, 0, 1, 2, 1, 0, 0, 0, 0, -1, 0, 1, 2, 2, 3, 3, 4, 3, 2, 1, 1, 1, 2, 1, 1, 1, 2, 3, 3, 2, 1, 1, 2, 0, 1, 0, 1, 1, 2, 0, 0, -1, 1, 1, 1, 0, 2, 1, 4, 3, 2, 2, 2, 2, 2, 1, 2, 1, 3, 2, 2, 2, 1, 0, 2, 0, 2, 2, 3, 1, 0, 1, 0, 0, 1, 2, 1, 1, 0, 1, 1, 1, 1, 0, 0, 1, 2, 0, 0, 0, 2, 3, 3, 2, 1, 2, 1, 1, 1, 3, 3, 2, 0, 1, 0, -2, 0, 2, 3, 4, 4, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 2, 3, 3, 2, 0, 0, 1, 2, 2, 0, 1, -3, -1, 0, 1, 2, 4, 2, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 2, 1, 2, 3, 3, 2, 2, 0, 0, 0, 0, 1, 0, 1, -4, -3, -2, -1, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 1, 2, 2, 1, 1, 1, -1, 0, 0, 0, 0, -2, -3, -2, 0, 0, 2, 1, 2, 2, 1, 2, 0, 0, 1, 1, 1, 1, 0, 2, 2, 2, 1, 1, 2, 3, 2, 1, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, -2, 0, 1, 0, 0, 1, 0, 1, 2, 3, 3, 2, 0, 1, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -2, -2, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -1, -2, -1, -1, -1, -2, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, -1, -1, -2, 0, -1, 0, -2, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, -2, -1, -2, -2, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -2, -2, -1, -2, -3, -2, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 2, 0, 2, 0, 1, 0, 1, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 2, 1, 2, 1, 1, 2, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 2, 3, 2, 3, 2, 2, 2, 1, 1, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 1, 1, 0, 1, 2, 1, 2, 2, 1, 2, 0, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 1, 0, 1, 1, 2, 1, 1, 1, 1, 2, 1, 1, 1, 1, 0, 1, 2, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 2, 0, 2, 0, 2, 1, 2, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 1, 2, 1, 0, 0, 1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 1, 1, 1, 1, 2, 1, 1, 1, 0, 1, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 1, 1, 0, 1, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 2, 1, 1, 2, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 1, 0, 0, 1, 2, 2, 1, 2, 1, 2, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 2, 1, 2, 1, 2, 1, 1, 1, 1, 1, 0, 1, 0, 1, 1, 2, 0, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 3, 2, 1, 0, 1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 3, 2, 0, 0, 2, 1, 0, 2, 1, 1, 2, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 1, 1, 1, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, 1, 1, 1, 2, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -2, -2, -1, 0, -2, -3, -3, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, -1, -1, -1, -3, -3, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -2, -2, -2, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 2, 2, 1, 2, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 1, 1, 0, 1, 2, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, -1, -1, -1, 0, 0, 1, 1, 1, 1, 1, 2, 1, 1, 2, 3, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 1, 1, 1, 2, 2, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 1, 0, 1, 1, 2, 2, 2, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, -2, -1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 3, 1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, -1, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 0, 2, 4, 2, 0, 0, 0, 0, 0, 1, 2, 1, 1, -1, -1, -2, -3, -3, -2, -2, 0, 0, 1, 1, 2, 1, 1, 1, 1, 0, 1, 2, 2, 1, 2, 3, 1, 0, 1, 1, 1, 1, 2, 3, 2, 0, -1, -3, -2, -4, -4, -3, -2, 0, 0, 1, 2, 1, 1, 0, 2, 0, 1, 2, 1, 2, 2, 1, 0, 0, 2, 2, 0, 1, 3, 2, 1, 0, 0, -1, -2, -2, -3, -3, -2, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 2, 1, 2, 1, 1, 0, 2, 2, 1, 3, 3, 2, 1, 0, 0, 0, -1, -1, -1, -4, -3, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 2, 2, 1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 3, 1, 0, -1, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 2, 3, 1, 0, 0, 0, -1, -1, -2, -1, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 0, 0, 1, 0, 0, 1, 0, 0, 2, 2, 1, 2, 1, 0, 0, -2, -2, -2, -3, -2, -1, 0, 0, 1, 0, 0, -1, 0, 0, 1, 2, 3, 2, 0, 1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, -2, -3, -3, -2, -2, -2, 0, 1, 0, 1, 0, 0, 0, 0, 1, 2, 1, 1, 2, 1, 0, 0, 0, -1, -2, 0, 0, 0, 0, -1, 0, -2, -2, -2, -2, -1, -1, -2, 0, 0, 0, 0, 0, 1, 0, 1, 1, 4, 3, 2, 1, 1, 1, 0, 0, 0, -2, 0, 0, 0, 0, -1, 0, -1, -1, -2, -2, -3, -1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 2, 1, 2, 2, 1, 1, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 3, 1, 0, 1, 1, 1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, 1, 0, -1, 0, -3, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 1, 0, -1, -2, -2, -2, -1, -1, 0, 1, 1, 1, 0, 1, 1, 1, 2, 1, 1, 1, 0, 1, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -3, -2, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 3, 2, 1, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, 1, 0, 0, 1, 0, 1, 2, 2, 2, 2, 2, 2, 1, 2, 0, 2, 0, 2, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 1, 1, 2, 3, 2, 2, 1, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 1, 1, 2, 3, 2, 2, 1, 0, 0, 1, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 1, 1, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, -1, -2, -1, -2, -1, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -3, -1, -2, -2, -1, -1, -1, -1, -2, -1, -2, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -2, -3, -2, -3, -3, -3, -3, -1, -2, -2, -1, -2, -2, -3, -3, -1, -1, 0, -1, 0, 0, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -4, -3, -4, -4, -3, -2, -1, -2, -2, -1, -2, -2, -2, -2, -1, -2, 0, 0, -1, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, -3, -3, -3, -4, -3, -2, -2, -2, -3, -3, -1, -2, -3, -3, -2, -1, -1, -2, 0, -1, -1, -1, -2, 0, 1, 0, 0, -1, -1, 0, -3, -3, -2, -3, -3, -4, -1, -2, -1, -3, -2, -3, -3, -2, -1, -3, -3, -2, -3, -2, -2, -1, -2, -3, -1, 0, 0, 0, -1, 0, 0, 0, -2, -1, 0, -1, -3, -3, -1, -2, -1, -1, -2, -1, -2, -3, -2, -1, -3, -3, -2, -3, -2, -1, -3, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -2, -1, -1, -2, -1, -3, -2, -2, -1, -2, -2, 0, -3, -2, -2, -3, -3, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -1, -1, -3, -2, -3, -2, -2, -1, -2, -2, -2, -2, -3, -3, -1, -1, -3, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -2, -3, -1, -1, 0, -2, -2, -1, 0, -2, -2, 0, -1, -1, -1, -3, -4, 0, -2, -2, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, -2, -3, -2, -2, -2, -1, -2, -2, -1, 0, -1, 0, 0, 0, -2, -1, -3, -1, -2, -3, 0, 0, -1, 1, 0, 0, 0, 0, 0, -1, -1, -2, -3, -2, -1, -2, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -2, 0, -2, -2, -2, -1, 0, 0, 0, 0, -1, 0, -1, -2, -3, -2, -1, -2, -1, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, -2, -1, 0, -1, -1, 0, -2, -1, -1, -2, 0, -1, -2, -1, -2, 0, -3, -2, -2, -2, -2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, -1, -1, -1, -1, -1, 0, -1, -1, 0, -2, -1, -1, -2, -1, -1, -1, -2, -3, -3, -2, -1, -1, -2, 0, -1, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -2, -2, -3, -1, -2, -2, -1, -2, 0, 0, 0, 1, 1, 1, 2, 0, -1, -1, -1, 0, -2, 0, -1, -1, -2, -1, -1, -2, -1, -2, -1, -1, -2, -2, -2, -3, -2, -1, -1, -2, -1, 0, 0, 0, 2, 2, 2, 0, 0, -1, -2, -1, 0, 0, -1, -1, -1, -2, -2, -3, -2, -2, -1, 0, -2, -3, -3, -2, -2, -1, 0, -1, 0, 0, 0, 1, 3, 2, 2, 1, 0, 0, -1, -1, 0, -1, -2, -3, -1, -1, -2, -2, -1, -1, 0, -1, -1, -1, -1, -2, -1, 0, 0, -1, -1, 0, 1, 2, 1, 1, 2, 0, 0, 0, -2, 0, 0, -1, -1, -2, -2, -1, -2, -3, -1, -2, -1, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 1, 0, 1, 1, 2, 3, 2, 1, -1, -1, 0, 0, -1, -1, -3, -3, -1, -2, -1, -2, -1, -2, 0, -2, -1, 0, -1, 0, -1, -1, 0, 1, 1, 0, 0, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, -2, -2, -3, -1, -2, 0, -1, -1, -2, -2, -1, -3, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 2, 1, -1, -1, -1, -1, 0, 0, -1, -2, -2, 0, -1, -2, -1, -1, -1, 0, -1, -3, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 1, 0, 0, 0, -1, 0, 0, -2, 0, -1, 0, 0, 0, -1, -2, -2, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 0, -1, 0, -1, -1, -1, -1, -1, -1, 0, -1, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 2, 2, 2, 2, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, -2, -4, -1, -1, -1, -1, 0, -1, 0, -1, -2, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, -3, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, -1, -1, -2, -4, -1, -1, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, -2, -4, -3, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 2, 0, 0, 1, 0, 1, 1, 1, 2, 0, 1, -2, -3, -4, -3, -1, 0, -1, -2, -2, -1, 0, 1, 2, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 2, 2, 1, 0, -1, -2, -2, -2, 0, -1, 0, 0, 0, -1, 0, 2, 1, 2, 1, 2, 0, 1, 2, 2, 0, 1, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, 0, -2, -4, -2, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 1, 0, 2, 1, 1, 2, 1, 1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, -2, -1, 0, 1, 1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, -2, -1, 0, 0, 1, 1, 1, 0, -1, -2, -2, 0, -2, 0, -1, 0, 1, 0, 3, 3, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, -1, -3, -3, -1, -1, 0, -1, -1, 0, 0, 0, 2, 1, 1, 0, 0, 0, -1, 0, -1, 0, 2, 1, 1, 0, 0, -1, 0, 0, 1, 1, 0, -1, -2, -2, -2, -1, 0, 0, -2, -1, 0, 0, 2, 2, 0, 1, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, -1, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, -1, 0, 0, 2, 0, 0, 0, -1, -2, 0, 0, 2, 2, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 2, 0, 1, 0, 0, 0, 1, 1, -1, 0, -1, 0, 1, 2, 2, 2, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 2, 1, 2, 1, 0, 1, 0, 1, 0, 0, 0, -1, -1, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 2, 1, 1, 1, 0, 1, 1, 1, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 1, 1, 0, 1, 0, 2, 2, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 0, 0, -1, 0, -1, -1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 1, 2, 1, 1, 0, 0, -2, -1, -1, 0, 0, 1, 2, 1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 2, 2, 1, 2, 0, -1, -1, -2, -1, -1, -1, -1, 0, 0, 2, 0, -1, -1, -1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 1, 1, 1, 2, 1, 2, 3, 1, 0, 0, -1, -1, -1, -1, -1, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 3, 2, 2, 2, 0, 1, 2, 3, 0, 0, 0, -2, -2, -2, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 1, 2, 3, 0, 0, -1, -1, -1, -2, -2, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -2, -1, -2, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 2, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 2, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, -2, -1, -1, -1, -1, -1, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -3, -1, -1, -2, 0, 0, -2, 0, 0, 0, -1, 0, 2, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, -1, -3, -2, -2, -2, -2, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -1, -2, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, -2, -2, -1, -1, 0, 1, -1, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -2, -1, -1, -2, -2, -2, 0, 0, -1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, -2, -1, -2, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 2, 2, 1, 1, 1, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 3, 2, 1, 0, 0, 0, 0, 0, 1, 3, 2, 1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 1, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 1, 3, 1, 0, 0, 0, 0, 0, 0, 3, 2, 1, 1, 0, 0, 0, 1, 1, 2, 1, 1, 2, 1, -1, -2, -1, -2, 0, 0, 0, 0, 0, 1, 2, 2, 2, 0, 0, 1, 0, 0, 1, 3, 1, 0, 0, 0, 0, 2, 2, 2, 2, 2, 1, 0, 0, -3, -3, -3, -2, 0, 0, 0, 0, 0, 2, 2, 2, 2, 2, 1, 0, 0, 0, 1, 2, 0, 0, -1, 1, 2, 4, 2, 3, 2, 3, 0, 0, -2, -3, -5, -3, -2, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 1, 0, 0, 1, 1, 2, 4, 4, 3, 2, 2, 1, 0, -3, -3, -4, -2, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, -1, 0, 0, 2, 3, 3, 3, 2, 3, 2, 0, -1, -2, -2, -2, -3, -1, -1, -1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 3, 2, 3, 2, 2, 2, 1, 0, -1, -1, -2, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 3, 3, 1, 0, 1, 2, 0, -1, -1, -2, -2, -2, -3, -1, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 2, 3, 4, 2, 1, 2, 1, 0, 0, -2, -3, -2, -3, -4, -2, 0, 0, 1, 0, 0, 2, 2, 0, 2, 0, 1, 1, 0, 0, 0, 0, 1, 1, 2, 2, 0, 1, 2, 1, 1, -1, -2, -1, -4, -4, -3, -2, -1, 2, 2, 1, 1, 0, 1, 1, 2, 1, 2, 1, 1, 0, 0, 0, 1, 0, 2, 1, 2, 1, 2, 2, 1, -1, -3, -2, -2, -3, -2, -1, 0, 2, 3, 3, 2, 0, 1, 1, 2, 1, 1, 1, 1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 2, 0, 1, -1, -2, -3, -2, -1, -1, -1, 0, 1, 2, 4, 2, 2, 1, 2, 1, 2, 1, 2, 1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, -1, -2, -3, -2, -2, -1, 0, 0, 2, 4, 3, 3, 3, 1, 2, 2, 2, 0, 0, 0, 0, -1, -1, 1, -3, -2, -1, -1, 0, 0, 1, 1, -2, -1, -2, 0, 0, 0, 0, 1, 2, 3, 3, 2, 2, 2, 1, 2, 1, 2, 0, 0, -1, -1, 0, 0, -2, -1, 0, 0, 0, 1, 0, 0, -1, -2, 0, 0, 0, 1, 1, 1, 1, 2, 2, 3, 2, 2, 2, 1, 1, 1, 1, 1, 0, -1, 0, 1, -3, -2, -1, 0, 1, 2, 0, 0, 0, -1, -1, 1, 1, 1, 0, 1, 1, 2, 3, 2, 1, 2, 2, 2, 1, 1, 0, 0, 0, -1, 0, 2, -2, -2, 0, 0, 0, 1, 2, 0, 0, -1, 0, 1, 2, 0, 1, 0, 1, 1, 2, 2, 1, 2, 3, 1, 1, 1, 0, 0, -1, 0, 0, 0, -2, -2, -2, -1, 0, 2, 1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 1, 2, 2, 0, 2, 2, 2, 1, 0, 0, -1, 0, 0, 1, -2, -1, -1, 0, 0, 2, 1, 2, 1, 1, 2, 2, 3, 0, 1, 0, 0, 0, 1, 2, 0, 2, 1, 2, 2, 1, 0, 0, 0, -1, 0, 1, -2, -1, -1, 0, 0, 0, 1, 1, 0, 0, 1, 2, 1, 1, 1, 0, 0, 0, 2, 0, 0, 2, 1, 1, 0, 1, 1, 0, 0, 0, 1, 2, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 2, 1, 3, 2, 2, 2, 2, 2, 1, 2, 2, 2, 3, 2, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 2, 0, 0, 0, 2, 0, 0, 1, 1, 3, 3, 3, 2, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 2, 0, 0, 1, 0, 0, 2, 2, 3, 1, 3, 1, 1, 0, 0, -1, 1, 2, 2, 0, 0, 1, 0, 1, 0, 1, 1, 1, 2, 1, 0, 2, 2, 1, 1, 0, 0, 0, 1, 3, 3, 1, 2, 1, 1, 0, 0, 0, 1, 3, 3, 1, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 3, 2, 1, 0, 0, 0, 0, 0, 0, 1, 3, 1, 1, 1, 3, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 2, 1, 2, 1, 1, 2, 0, 0, 0, 0, 1, 2, 0, 0, -1, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -2, 0, 0, 1, 1, 1, 2, 1, 2, 0, 1, 2, 3, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 1, 0, 0, 1, 0, 0, -1, 0, 1, 2, 1, 0, 0, 1, 1, 0, 2, 3, 4, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 1, -2, -1, 0, 0, 0, 3, 1, 1, 3, 3, 1, 1, 1, 3, 4, 2, 2, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 1, -1, 1, -1, -1, 0, 0, 0, 0, 3, 2, 2, 4, 3, 3, 2, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, 1, 0, 0, 0, 1, 0, 0, 1, 2, 2, 2, 4, 1, 1, 1, 2, 0, -1, 0, 1, 0, 1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 3, 0, 0, 1, 2, 0, 1, 0, 0, 0, 2, 2, 0, 1, 2, 1, 0, 0, 0, 1, 2, 2, 0, 0, 0, 1, 0, -1, -2, 0, 0, -1, 1, 0, 0, 2, 1, 0, 0, 1, 1, 0, 0, 2, 0, 0, 2, 2, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 0, -1, -2, 0, 2, 2, 0, 0, 0, 1, 1, 1, 1, 2, 2, 1, -1, 0, 0, 0, 1, 2, 1, 0, 0, -1, -2, -3, -1, 0, 0, 0, 0, -2, -3, -2, 0, 1, 0, 0, 0, 1, 3, 2, 2, 3, 3, 1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, -2, -2, -2, -2, 0, -1, 0, -2, -3, -2, 0, 1, 1, 0, 2, 3, 3, 3, 3, 4, 4, 2, 0, 1, 0, 2, 1, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, -1, 2, 0, -2, 0, 0, 1, 0, 0, 2, 1, 2, 1, 2, 2, 3, 1, 0, 0, 0, 1, 3, 0, 1, 0, 0, -1, -1, -1, -2, -2, 0, 0, 0, 0, -2, 0, 1, 3, 4, 3, 2, 1, 3, 3, 2, 4, 3, 4, 1, 0, -1, 0, 2, 2, 1, 0, -1, -1, -1, 0, 0, -1, 0, -1, 1, 0, 0, 1, 2, 4, 3, 3, 2, 3, 5, 4, 4, 4, 5, 3, 2, 1, 0, -1, 0, 2, 0, 0, 0, -1, -2, -2, 0, 1, 1, 0, 2, 2, 0, 1, 3, 3, 4, 2, 1, 2, 2, 5, 6, 5, 4, 5, 3, 2, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, 1, 0, 1, 1, 1, 1, 2, 3, 4, 3, 2, 3, 2, 3, 3, 3, 4, 3, 3, 2, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 2, 3, 3, 2, 2, 3, 4, 3, 1, 2, 3, 1, 2, 1, 0, 0, -1, 0, -1, -3, -2, -2, -1, -1, 1, 1, 1, 0, 1, 2, 3, 2, 0, 2, 1, 1, 1, 0, 2, 3, 1, 1, 0, 0, 2, 2, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 2, 0, 0, 3, 4, 3, 2, 0, 1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 2, 3, 3, 4, 3, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 1, 2, 3, 3, 2, 1, 0, -1, -2, 0, 1, 0, -1, 0, -1, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 1, 2, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, -3, -1, -2, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, 1, 0, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, -1, -1, -2, 0, 0, -1, 2, 2, 1, 1, 0, 1, 2, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, -2, -4, -4, -3, -2, -2, -2, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, -1, -1, -1, -1, -1, -1, -2, 0, -1, 0, -1, 0, -2, -3, -3, -3, -3, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 2, 0, 0, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 1, 0, -2, 0, -2, -2, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, -2, 1, -1, -3, -3, -2, -2, -3, 0, 0, -2, -2, -2, -4, -2, -1, -2, -1, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, 0, -2, -3, -4, -4, 0, 0, -3, 0, -2, -2, -3, 0, 0, 0, -3, -2, -5, -4, -4, -3, -2, -3, -1, -1, 0, 0, 0, -3, -2, -2, 0, -1, -2, -3, -5, -3, 0, 0, -1, 0, 0, -1, -3, -2, -1, -1, -1, -3, -4, -3, -3, -3, -3, -3, -4, -1, 0, 0, -1, -3, -2, 0, 0, 0, -2, -2, -4, -2, 0, 0, 0, 0, 0, -1, -2, -2, -2, -2, -4, -4, -2, -3, -4, -4, -3, -4, -4, -3, -1, -2, -3, -1, 0, -1, -2, -1, -2, -2, -2, -3, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -4, -3, -2, -3, -4, -4, -2, -2, -4, -5, -3, -3, -2, -2, 0, 0, -2, -3, -3, -1, -2, 0, 0, 0, 1, 1, 0, 0, 0, -2, -2, -2, -2, -3, -2, -3, -5, -4, -2, -2, -3, -4, -4, -3, -1, -1, -1, 0, 0, -3, -3, -3, -1, 0, 0, 0, 1, 2, 2, 0, 0, 0, -1, -3, -4, -3, -3, -1, -4, -5, -4, -2, -2, -4, -5, -3, -1, -3, -2, -1, -2, -2, -4, -4, -2, 0, 0, 0, 0, 0, 2, 0, -1, 0, -1, -4, -4, -3, -2, -2, -3, -5, -4, -2, -4, -3, -4, -4, -2, -3, -2, -2, -3, -2, -4, -6, -2, 1, 0, 0, 0, 1, 2, 0, -3, 0, 1, -2, -4, -2, -1, 0, -1, -3, -4, -4, -3, -3, -2, -2, -3, -4, -1, -4, -3, -1, -2, -6, -2, 0, 0, 0, 2, 1, 2, 1, 0, 0, 3, 2, -2, 0, -1, 0, -2, -2, -4, -4, -6, -4, 0, 0, -3, -4, -3, -3, -5, -1, -2, -4, -1, -1, 0, 0, 3, 3, 1, 2, 2, 3, 4, 2, 1, 0, 0, 0, -1, -1, -3, -3, -6, -5, -1, 0, -2, -3, -1, -1, -4, -1, -3, -4, -1, -1, 0, 0, 3, 3, 3, 3, 5, 5, 4, 4, 1, 1, 2, 0, 0, -1, -2, -3, -5, -5, -3, -2, -2, -2, -2, -3, -2, 0, -1, -4, 0, 0, 0, 0, 4, 2, 1, 3, 4, 4, 4, 3, 0, 0, 4, 1, 0, 0, -1, -1, -4, -3, -2, -3, -1, 0, -1, -3, -2, -2, -1, -3, 1, 0, 0, 1, 3, 2, 3, 3, 4, 2, 2, 2, 0, 0, 2, 3, 0, 0, -1, -1, -1, -1, -3, -2, 0, 0, -1, -4, -3, -2, -2, -2, 1, -1, 0, 0, 4, 3, 2, 4, 4, 1, 0, 3, 0, 0, 2, 0, 0, 0, -2, 0, 0, -2, -2, -1, 0, 0, -2, -3, -1, -2, 0, 0, 2, -2, 0, 1, 3, 2, 4, 4, 4, 2, 2, 4, 2, 1, 3, 0, 0, -2, -1, -1, 0, -1, -2, -3, -1, 0, -4, -4, -1, -1, -1, 0, 3, -2, 0, 0, 2, 3, 3, 3, 3, 3, 2, 3, 4, 2, 3, 0, -1, -1, -2, -1, -1, -2, -3, -1, -1, -2, -5, -4, -1, 0, 0, 0, 1, 0, 0, 0, 2, 4, 2, 1, 4, 3, 3, 3, 2, 3, 3, 0, -1, 0, 0, -3, -2, -3, -1, -2, -2, -3, -3, -2, -3, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 0, 3, 4, 4, 2, 3, 3, 2, 0, -2, 0, 0, -3, -4, -2, -1, -1, -3, -4, -3, -1, -3, -2, 0, 0, -1, 0, 0, 1, 3, 4, 3, 0, 2, 4, 3, 4, 4, 4, 1, 0, -2, -1, -2, -4, -4, -2, 0, 0, -3, -4, -4, -2, -2, -1, -1, -2, -2, -1, 0, 0, 2, 2, 2, 1, 2, 3, 3, 5, 6, 2, -1, -2, -2, -1, -2, -4, -4, -1, 0, 1, 0, -3, -3, -2, -2, -2, 0, 0, -2, 0, 0, 0, 1, 3, 2, 1, 1, 1, 2, 4, 5, 2, -1, -2, -2, -2, -4, -5, -5, -3, 0, 2, -1, -1, -3, -1, -2, -1, 0, 0, -1, 0, 0, 1, 1, 1, 2, 2, 0, 1, 0, 3, 3, 0, -3, -4, -2, -2, -3, -4, -5, -2, 0, 0, -2, -1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, -1, 0, 1, 2, 1, -1, -5, -5, -3, -3, -3, -4, -4, -2, -1, -2, -3, -1, 0, 1, 0, -1, -1, 0, 3, 0, 0, 0, 0, 2, 2, 0, -1, 0, 1, 2, 1, -1, -4, -4, -3, -1, -3, -2, -3, -2, 0, -2, -3, -2, 1, 1, 0, 0, -2, 0, 1, 0, 0, 0, 0, 1, 1, -1, -2, 0, 2, 1, 0, -1, -2, -3, -4, 0, -2, -1, -2, -3, -1, 0, -3, -2, -1, 1, 0, 0, -1, -2, 0, 1, 0, 0, 0, 1, 3, -1, -3, 0, 0, 2, 1, -1, -2, -2, -2, 0, 0, -1, -3, -3, -2, -1, -2, -1, 0, 0, 1, 1, -1, -1, 1, 1, 0, 0, -2, 0, 0, 0, -3, -2, 0, 1, 0, -1, -2, -1, -3, 0, -1, -1, -3, -2, -2, -2, -3, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, 0, 0, 0, -2, -2, -1, -1, -2, 0, -1, -1, -2, -1, 0, -2, -1, 0, -1, -2, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -2, -2, 0, 0, -2, -2, 0, -1, 0, 0, -3, -2, -1, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, -2, -2, -1, -1, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -2, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, -2, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, -2, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 1, 2, 1, 0, 0, -1, -1, -2, -1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 1, 1, 1, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 2, 1, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, 0, 1, 2, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 3, 2, 1, 2, 1, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, 2, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 1, 2, 2, 2, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 2, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, 1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 1, 1, 2, 1, 3, 3, 3, 2, 3, 1, 1, 0, 0, 1, 1, 1, 2, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, -1, 0, 0, 1, 0, 0, 1, 1, 2, 2, 1, 1, 1, 0, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 1, 1, 0, 1, 1, 0, 2, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 2, 1, 0, 1, 1, 2, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 1, 1, 1, 1, 2, 1, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, -1, -2, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, -3, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 2, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -3, -2, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, -2, -1, -3, -2, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -2, -1, 0, -1, 0, -1, -1, -2, -2, -3, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, -1, -1, -1, -3, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, -2, -1, -1, -2, -1, 0, -2, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, -2, -3, -2, 0, -1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 2, 0, 1, 0, 0, 1, 1, 0, 1, 0, -1, -1, -1, -2, -2, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, -1, -1, -1, -2, -1, -2, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 2, 2, 1, 1, 0, 0, -1, 0, 0, -1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, 2, 2, 1, 2, 0, 1, 0, 0, -1, 0, -1, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 1, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 1, 2, 1, 0, 1, 1, 2, 2, 1, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 1, 2, 2, 0, 1, 0, 2, 2, 1, 2, 1, 1, 1, 1, 0, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 2, 2, 3, 2, 3, 2, 1, 1, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 2, 2, 3, 3, 1, 3, 1, 0, 0, 0, 2, 0, 1, 1, 1, 1, 2, 1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 2, 3, 2, 2, 4, 1, 1, 0, 1, 2, 1, 1, 1, 0, 1, 1, 1, 1, 0, 2, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 2, 1, 1, 2, 2, 3, 2, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 1, 1, 1, 2, 1, 2, 2, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 2, 1, 3, 2, 2, 1, 1, 1, 2, 1, 2, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 1, 1, 1, 1, 2, 2, 1, 2, 1, 1, 0, 1, 1, 2, 1, 1, 0, 0, 1, 1, 2, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, -1, 0, 0, -2, -2, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 2, 1, 1, 0, 1, 0, 0, 0, -1, -1, -1, -1, 0, -2, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 1, 1, 2, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 1, 1, 1, 1, 1, 0, 0, 1, 1, 1, 0, 2, 2, 2, 2, 2, 2, 2, 1, 2, 2, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 1, 1, 0, 1, 0, 0, -1, 0, 0, 1, 1, 3, 3, 1, 2, 1, 1, 3, 2, 3, 3, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, 1, 0, 1, 0, -1, -1, 0, 0, 0, 1, 1, 1, 2, 1, 1, 3, 2, 2, 3, 2, 2, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 1, 2, 3, 3, 2, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 1, 2, 2, 2, 3, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 1, 2, 4, 3, 3, 0, 1, 0, -1, 1, 0, 1, 0, 0, 0, -2, -2, -3, -4, -2, -2, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 1, 2, 3, 2, 2, 1, 1, 0, 0, 1, 1, 2, 1, 0, 0, -1, -1, -3, -3, -2, -1, 0, 0, 0, 2, 0, 1, 1, 0, 1, 0, 0, 1, 2, 2, 3, 1, 1, 0, 0, -1, 0, 1, 2, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 2, 2, 2, 1, 2, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 1, 0, 1, 3, 2, 1, 0, 0, 0, 1, 1, 3, 1, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 2, 0, 1, 0, 0, 2, 2, 2, 2, 0, 0, 1, 1, 0, 2, 2, 3, 2, 2, 1, 0, -1, -1, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 2, 0, 0, 0, 0, 2, 2, 3, 2, 1, 0, 0, -1, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 2, 1, 1, 0, 0, 1, 0, 0, 1, 1, 1, 2, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 2, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 2, 2, 2, 3, 3, 1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 3, 1, 3, 3, 2, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 2, 1, 3, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 3, 2, 2, 3, 4, 2, 1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 3, 3, 2, 4, 2, 3, 2, 3, 1, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 1, 2, 2, 3, 2, 3, 2, 1, 2, 2, 1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 2, 1, 0, 1, 1, 1, 1, 2, 1, 1, 1, 2, 1, 3, 2, 3, 3, 2, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 2, 2, 2, 2, 2, 0, 1, 0, 1, 0, 0, 2, 1, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 2, 2, 2, 0, 1, 1, 0, 1, 1, 2, 3, 1, 1, 0, 2, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -2, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -2, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -1, -2, -1, -1, 0, -2, -1, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, -1, -1, -2, -1, -1, -2, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, -2, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, -2, -2, -1, -1, 0, -1, 0, -1, 0, -1, -1, 0, -1, -1, 0, -1, -1, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -2, -2, -2, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -2, -1, -1, -1, 0, -1, 0, -1, -1, -1, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, -2, -2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -2, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 1, 1, 2, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, 1, 1, 0, 1, 2, 1, 2, 1, 1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 2, 1, 2, 1, 1, 0, 1, 2, 1, 0, 0, 1, 1, 1, 2, 1, 1, 0, 1, 0, 1, 2, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 2, 1, 2, 0, 0, 1, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 1, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 1, 2, 0, 1, 0, 0, 0, -1, 0, 0, -1, -2, -1, 0, -1, -1, -1, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, -2, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -2, -1, -2, -1, 0, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, 0, -1, -2, -2, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -2, -1, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -3, -2, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 0, 0, 1, 0, 0, 0, 2, 2, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 2, 1, 0, 2, 0, 1, 1, 0, -1, 0, 0, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, 1, 1, 1, 2, 1, 0, 3, 2, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, -2, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 2, 0, 0, 0, 1, 0, -1, -2, -2, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 2, 2, 0, -1, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, 1, 0, 2, 1, 0, 1, 0, 1, 1, 1, 0, -1, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 1, 0, 1, 2, 2, 2, 1, 1, 0, -1, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 1, 3, 3, 2, 2, 3, 1, -1, -1, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 2, 1, 1, 2, 1, 1, 3, 1, 2, 1, 1, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 2, 2, 0, 0, 1, 1, 1, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 2, 2, 2, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, -1, 1, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 2, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, -2, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, -1, -1, -1, -1, 0, -1, -1, -1, 0, -1, -1, -1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -2, 0, 0, -2, -2, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, -1, -1, -2, -1, -2, -1, 0, -2, -1, -1, -1, -1, -2, -1, -1, 0, 0, -2, -1, -1, -2, -1, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, -1, -1, -1, -1, -1, -2, -2, 0, -1, 0, -1, -1, 0, -2, -1, 0, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -2, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 2, 3, 4, 1, 0, 0, 2, 1, 1, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 2, 2, 0, 1, 0, 1, 3, 2, 2, 3, 3, 2, 0, 0, 2, 1, 2, 1, 1, 3, 2, 0, 0, 0, 0, -2, -2, -1, -1, 0, 0, 1, 1, 2, 1, 0, 1, 2, 4, 3, 3, 3, 3, 2, 0, 1, 2, 3, 1, 2, 2, 4, 3, 2, 0, 0, 0, -2, -2, -2, 0, 0, 1, 1, 3, 2, 0, 1, 0, 2, 2, 3, 2, 2, 3, 1, 0, 0, 2, 2, 3, 4, 4, 4, 4, 1, 1, 0, 0, -1, 0, -2, -1, -1, 1, 2, 2, 2, 2, 1, 1, 2, 2, 2, 1, 2, 2, 0, 0, 1, 3, 3, 4, 4, 4, 4, 3, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 2, 3, 3, 1, 2, 2, 0, 0, 1, 1, 4, 3, 4, 5, 4, 3, 2, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 1, 1, 2, 2, 1, 2, 1, 2, 2, 2, 1, 1, 0, 1, 2, 2, 4, 3, 4, 5, 4, 2, 1, 0, -1, -1, -2, -2, -2, -2, -2, -1, 0, 1, 1, 2, 1, 1, 1, 1, 2, 2, 0, 0, 0, 0, 0, 2, 3, 2, 3, 4, 3, 2, 2, 0, 0, -1, -1, -2, -2, -1, -2, -1, 0, 0, 1, 1, 1, 1, 2, 3, 4, 3, 1, 1, 0, 0, 2, 2, 2, 3, 2, 4, 3, 1, 1, 0, -2, -2, -3, -2, -2, -3, -2, 0, 0, 1, 1, 0, 0, 1, 2, 2, 4, 2, 1, 0, 0, 1, 2, 2, 2, 2, 4, 3, 2, 1, 0, 0, -1, -2, -2, -2, -2, -2, -2, -1, 0, 0, 0, 1, 2, 1, 2, 2, 3, 2, 0, 1, 0, 0, 1, 2, 1, 1, 3, 3, 3, 2, 2, 1, 0, -2, -3, -1, -3, -3, -2, -1, 0, 1, 0, 1, 0, 1, 2, 3, 3, 3, 1, 0, 0, 0, 1, 2, 1, 1, 3, 3, 3, 2, 1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 1, 0, 1, 1, 0, 2, 3, 4, 2, 0, 1, 0, 1, 1, 1, 1, 1, 2, 3, 3, 2, 2, 0, 0, -1, -1, -2, -2, 0, 0, 1, 1, 0, 1, 2, 1, 0, 2, 2, 3, 3, 0, 1, 0, 0, -1, 0, 0, 0, 0, 2, 1, 2, 0, 0, -1, 0, 0, -1, -1, 0, 1, 2, 2, 0, 1, 0, 1, 1, 1, 3, 3, 1, 0, 0, 0, -1, 0, -2, -1, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 3, 1, 0, 0, 1, 0, 2, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, -2, -2, 0, 1, 0, 0, -1, -1, -2, 0, 0, -2, 0, -1, 1, 2, 2, 1, 2, 1, 1, 1, 2, 2, 1, 0, 0, 0, -1, -2, 0, 0, -2, 0, -1, -1, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, -1, 0, 0, 1, 1, 3, 2, 1, 0, 2, 1, 0, -1, 0, -1, -2, -1, -1, -2, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, -2, -1, 0, -1, 0, 0, 2, 2, 0, 1, 1, 1, 0, 0, 0, -2, -2, -2, -1, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, -2, -2, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, -1, -3, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -3, -2, -1, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, -2, 0, -1, -2, -1, 0, 0, 0, -2, -1, 0, 0, -1, 0, 1, 0, 0, -1, -2, -1, -2, -1, -1, 0, 0, 1, 0, 1, 0, 1, 1, 0, -2, 0, 0, -2, -2, -1, -1, -1, -1, -2, -2, -1, -1, 0, 0, -1, -1, -2, -2, -3, -3, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -2, -3, -2, -1, -2, 0, 0, -1, 0, -1, -1, -1, -3, -3, -3, -3, -2, -2, -1, 0, 0, -2, -2, -2, -2, -2, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 1, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 2, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 2, 2, 1, 2, 1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 2, 2, 1, 0, 1, 0, 1, 0, 0, 1, 2, 1, 2, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 2, 2, 0, 0, 0, 0, 1, 1, 1, 2, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 2, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 2, 1, 2, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 1, 0, 1, 1, 0, 1, 0, 1, 0, 1, 1, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -3, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 1, 0, 0, 2, 2, 2, 2, 1, 0, 0, 2, 3, 3, 1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 2, 1, 1, 3, 1, 1, 1, 1, 2, 1, 2, 3, 2, 2, 2, 3, 1, 1, 3, 3, 2, 0, 0, 0, 2, 0, 0, 1, 0, 0, 3, 3, 3, 2, 2, 3, 4, 3, 4, 4, 3, 2, 0, 3, 2, 1, 2, 3, 2, 2, 4, 3, 2, 1, 1, 2, 2, 1, 2, 1, -1, 0, 2, 3, 3, 2, 2, 3, 5, 5, 5, 4, 2, 1, 1, 1, 1, 0, 0, 2, 1, 2, 2, 3, 1, 1, 3, 2, 3, 1, 1, 2, 0, 0, 1, 2, 1, 2, 2, 2, 1, 4, 3, 3, 2, 0, 0, 0, 1, 0, 0, 1, 1, 1, 3, 3, 2, 3, 2, 2, 3, 2, 4, 2, 1, 0, 0, 0, 0, 1, 0, -1, 1, 2, 2, 0, 0, 0, 0, -2, -1, 0, 0, 1, 1, 2, 3, 4, 1, 3, 4, 3, 3, 2, 4, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, -1, -3, -4, -3, 0, 0, 0, 1, 2, 2, 0, 0, 2, 2, 2, 3, 3, 4, 2, 2, 1, 2, 2, 2, 1, 0, -1, -1, -1, 0, 0, -1, -3, -4, -4, -4, -1, 0, 0, 1, 2, 0, 0, 0, 1, 3, 2, 2, 3, 3, 3, 3, 2, 2, 4, 2, 3, 0, -1, -3, -2, -2, -2, -2, -2, -3, -4, -5, -2, -1, 0, 3, 2, 2, 0, 0, 1, 0, 1, 0, 0, 3, 3, 2, 2, 1, 5, 5, 3, 1, -1, -3, -4, -5, -5, -3, -1, -2, -5, -7, -4, 0, 0, 3, 4, 2, 0, 2, 1, 0, 0, -1, 0, 2, 2, 1, 1, 0, 3, 3, 2, 0, -2, -2, -5, -7, -6, -5, 0, 0, -3, -6, -3, 0, 0, 2, 4, 2, 1, 2, 1, -1, -3, -4, -5, 0, 0, 0, 0, 0, 0, 0, 1, -1, -2, -1, -3, -6, -6, -4, -1, 0, -3, -6, -3, 0, 0, 4, 5, 5, 2, 1, 0, -1, -5, -6, -6, -5, -2, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, -2, -4, -5, -1, 0, -3, -4, -2, 0, 0, 4, 4, 4, 4, 2, 0, -2, -4, -7, -9, -8, -5, -4, -1, -1, -1, -1, -1, -3, -3, 0, 0, -1, -4, -4, -3, -1, -1, -3, -2, 0, 0, 2, 4, 4, 2, 1, 0, -1, -3, -6, -8, -9, -6, -4, -3, -1, -2, -4, -4, -5, -4, 0, 1, -1, -3, -4, -3, -2, -3, -4, -2, 0, 0, 2, 4, 2, 1, 0, 0, 0, -4, -6, -7, -8, -5, -3, -2, -1, -3, -3, -6, -5, -3, 0, -1, -3, -3, -4, -2, -3, -6, -5, -1, -1, 0, 2, 3, 1, -1, -2, 0, 0, -5, -5, -7, -8, -5, -2, -2, 0, 0, -3, -2, -3, -2, -1, -2, -3, -3, -4, -1, -3, -4, -3, -2, 0, 0, 2, 4, 1, -2, -1, -1, -1, -4, -5, -5, -5, -5, -4, -1, 0, 0, -2, -1, -1, -1, 0, -2, -3, -3, -3, -2, -3, -3, -4, -2, -1, 0, 2, 3, 0, -1, -1, 1, 0, -3, -5, -4, -5, -4, -4, -2, 0, 1, 0, 0, -1, -2, 0, 0, -2, -1, -3, -2, -2, -1, -2, -2, -1, 0, 3, 3, 1, 0, 1, 1, 2, 0, -2, -5, -5, -3, -4, -3, 0, 1, 3, 2, -1, -3, -1, 0, 0, -1, -1, 0, -1, -2, -2, -1, 0, 0, 2, 3, 1, 1, 1, 3, 3, 1, -2, -4, -6, -2, -3, -1, 0, 4, 5, 3, 0, -2, -2, -1, 0, -1, -1, -1, -2, -1, -3, -1, 0, 0, 0, 1, 2, 1, 1, 2, 2, 1, -1, -4, -5, -2, 0, 0, 1, 3, 4, 3, 0, -1, -2, -2, 0, -1, -2, -2, -2, -1, -2, -2, 1, 0, -2, 0, 1, 2, 3, 2, 2, 1, -1, -3, -2, -1, 0, 0, 1, 3, 2, 2, 2, -1, -1, -1, 0, -1, -4, -3, -1, -1, -2, -1, 1, 0, -3, -2, 1, 3, 2, 3, 2, 1, 0, 0, -2, 0, 2, 0, 1, 1, 2, 2, 0, 0, 0, -1, -2, -2, -2, -2, -1, 0, -2, -1, 1, 0, -2, -1, 1, 5, 4, 2, 3, 2, 0, 0, 0, 2, 2, 0, 1, 1, 1, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -2, -1, 1, 1, -3, -1, 4, 6, 5, 4, 3, 1, 0, 0, 1, 3, 3, 1, 0, 0, 0, 1, 0, -1, 0, 2, 3, 0, 0, -1, -1, 0, -1, 0, 1, 0, -3, -1, 3, 6, 7, 6, 5, 3, 0, 0, 2, 3, 3, 0, 0, 0, 0, 0, -1, -2, -1, 1, 1, 1, 0, 0, -2, -1, -1, 0, 1, 1, -3, -3, 2, 4, 7, 5, 5, 4, 2, 1, 2, 2, 2, 0, -1, 0, -1, 0, -1, -3, 0, 0, 0, 2, 3, 0, -2, -1, -1, 1, 3, 1, -2, -1, 3, 4, 6, 7, 4, 4, 2, 1, 2, 3, 3, 1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 4, 3, 0, 0, 0, 3, 5, 2, -1, -1, 1, 2, 3, 6, 4, 4, 3, 1, 2, 1, 2, 1, 0, -1, -1, 0, 1, 1, 0, 1, 1, 3, 2, 2, 2, 2, 2, 2, 4, 3, -1, -2, -1, 0, 0, 2, 0, 2, 0, 0, 2, 1, 1, 0, 0, -1, -2, 0, -1, -1, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 3, 2, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, 0, -1, -1, -1, 0, 0, -1, -2, -1, -1, -1, -2, 0, 0, 0, 0, -1, -1, -1, -3, -2, -3, -4, -4, -3, -5, -4, -3, -3, -2, -2, -1, -1, -3, -3, -2, -1, -1, -1, -3, -3, -2, -1, -1, -1, 0, 0, 0, 0, 0, -1, -2, -3, -3, -4, -4, -4, -4, -4, -4, -3, -3, -1, -1, -2, -4, -5, -3, -1, -2, -3, -4, -4, -4, -3, -3, -3, -2, 0, -1, -2, -2, -2, -3, -3, -3, -5, -7, -7, -6, -5, -7, -5, -3, -3, -1, -1, -4, -5, -3, -2, -2, -3, -2, -3, -1, -1, -2, -3, -2, -2, -2, -3, -2, -2, -3, -3, -3, -5, -4, -4, -4, -5, -4, -5, -3, -2, -2, -1, -4, -6, -4, -2, -2, -1, -1, 0, 0, 0, -1, -1, -3, -2, -2, -2, -1, -2, -2, -2, -3, -3, -4, -4, -4, -3, -2, -2, -2, -2, -1, -1, -4, -5, -4, -2, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -2, -1, -1, -2, -1, -1, -2, -2, -3, -1, 0, -1, 0, 0, -1, -1, -1, -1, -5, -4, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -5, -3, -2, -1, 0, 0, 0, 0, 1, 1, 0, 2, 2, 0, 1, 0, 1, 0, 0, 2, 0, 1, 1, 0, 1, 3, 3, 1, 0, 1, 0, -2, -3, -2, -1, 0, 0, 0, 0, 1, 2, 3, 3, 2, 3, 2, 2, 2, 1, 2, 2, 1, 1, 1, 0, 0, 2, 3, 2, 2, 1, 0, -1, 0, -3, -2, 0, 0, 0, 1, 1, 2, 3, 3, 4, 4, 3, 1, 2, 1, 2, 3, 3, 2, 1, 1, 1, 0, 1, 2, 2, 2, 0, 0, 0, 0, -3, -3, 0, 0, 1, 2, 1, 1, 1, 2, 3, 3, 2, 1, 1, 2, 4, 5, 4, 3, 2, 0, 1, 1, 1, 1, 2, 2, 1, 0, 0, 0, -2, 0, 0, 2, 2, 4, 4, 3, 2, 2, 1, 2, 1, 2, 1, 2, 4, 4, 6, 4, 3, 2, 0, 2, 1, 1, 2, 1, 1, 0, -1, -1, -2, 1, 1, 3, 4, 4, 5, 4, 2, 1, 1, 0, 0, 1, 2, 2, 4, 4, 4, 4, 3, 1, 2, 2, 0, 2, 2, 2, 2, 0, -1, 0, 0, 1, 2, 4, 5, 6, 4, 4, 2, 1, 0, 0, 0, 0, 0, 1, 3, 4, 4, 3, 2, 1, 2, 1, 0, 0, 1, 2, 2, 0, -1, 0, -1, 0, 3, 4, 5, 5, 3, 2, 2, 2, 2, 1, 0, 1, 2, 2, 4, 4, 3, 4, 2, 1, 2, 1, 1, 1, 2, 2, 3, 1, 0, 0, -1, 1, 2, 4, 5, 5, 4, 4, 2, 1, 3, 2, 2, 0, 0, 2, 3, 4, 3, 3, 4, 3, 2, 2, 1, 2, 2, 2, 2, 0, -2, 0, -1, 1, 3, 6, 6, 6, 5, 4, 3, 3, 2, 2, 2, 0, 1, 2, 2, 3, 2, 2, 4, 4, 3, 3, 3, 1, 1, 1, 0, 0, -2, -1, -1, 0, 2, 7, 7, 7, 5, 5, 5, 3, 4, 3, 1, 0, 0, 3, 2, 1, 2, 2, 3, 3, 3, 3, 2, 3, 1, -1, -2, -2, -1, -1, -1, 0, 4, 6, 6, 7, 5, 5, 5, 5, 3, 4, 1, 0, 0, 1, 2, 2, 3, 1, 1, 1, 2, 3, 2, 1, 1, 0, -3, -2, -2, -1, -2, 0, 4, 6, 6, 6, 5, 5, 5, 5, 4, 3, 1, 0, 0, 0, 0, 1, 1, 2, 2, 2, 1, 3, 2, 2, 2, 1, -1, -3, -1, -1, 0, 0, 2, 3, 6, 5, 5, 5, 5, 4, 4, 3, 0, -1, -2, -1, 0, 2, 2, 2, 2, 2, 2, 3, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 3, 4, 4, 6, 5, 6, 3, 3, 1, 2, 0, -1, 0, 1, 3, 3, 4, 3, 1, 3, 2, 3, 2, 1, 1, 1, 0, 1, 0, -1, -1, 0, 1, 2, 3, 5, 6, 5, 3, 1, 0, 1, 1, 1, 1, 2, 4, 3, 2, 3, 2, 2, 2, 2, 1, 2, 2, 0, 1, 0, -1, -1, -2, 0, 0, 1, 2, 5, 4, 4, 1, 0, 0, 0, 0, 1, 3, 3, 2, 3, 3, 2, 2, 2, 2, 1, 1, 0, 1, 2, 1, 0, -1, -3, -3, -3, -1, 0, 3, 2, 3, 2, 1, -1, -1, 0, 0, 2, 2, 1, 1, 2, 2, 2, 4, 4, 3, 2, 1, 0, 0, 0, 1, 0, -1, -4, -6, -4, -4, -1, 1, 1, 1, 0, 0, -1, 0, 0, 1, 0, 1, 1, 1, 1, 3, 4, 4, 4, 4, 2, 2, 0, 0, 1, 0, 0, -1, -3, -6, -6, -5, -3, -1, 0, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 2, 3, 3, 2, 2, 0, 0, 0, 0, 0, 0, -1, -4, -5, -6, -4, -3, -2, -1, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -4, -4, -5, -3, -3, -2, -2, -1, -2, -1, -1, 0, 0, -1, -2, -2, -1, -2, -1, 0, 0, 0, 0, -1, -1, -2, 0, -1, 0, -1, -1, -1, -4, -4, -4, -4, -5, -4, -2, -3, -2, -2, -1, -2, -1, -1, -2, -2, -2, -2, -2, -1, -1, 0, 0, -1, -3, -2, -2, 0, -1, -2, -1, -1, -3, -4, -3, -4, -3, -2, -1, -1, -2, -1, -1, -1, 0, -2, 0, -1, -2, 0, -1, -2, -2, -2, 0, -2, -2, -3, -3, -1, -1, -1, -1, 0, -1, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -2, -2, 0, 0, -1, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -1, 0, -1, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, -1, -1, -2, -2, -2, -3, -3, -3, -4, -4, -3, -3, -2, -2, 0, 0, -2, -2, -1, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -2, -2, -3, -3, -2, -3, -1, 0, -1, 0, 0, -3, -4, -2, -2, -2, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, -1, -2, -1, 0, 0, -3, -3, -4, -3, -3, -2, -3, -2, -1, 0, 0, -1, -3, -4, -3, -1, -1, 0, -1, 0, 0, 0, -1, 0, -2, -1, -2, 0, -1, 0, 0, -1, -1, -1, -3, -1, -1, -2, -1, -1, 0, 0, 0, -1, -3, -3, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, -1, 0, 0, -1, -3, -3, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -4, -2, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 2, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 0, -2, -3, -2, 0, 0, -1, 0, 0, 0, 1, 2, 1, 3, 1, 3, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 2, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 1, 2, 2, 4, 3, 2, 3, 1, 2, 1, 1, 2, 1, 1, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 2, 2, 1, 4, 4, 4, 3, 2, 1, 1, 2, 2, 2, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, -1, -2, 0, 1, 0, 2, 2, 1, 1, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 0, 0, 1, 1, 0, 0, 1, 0, 2, 0, 0, 0, 0, -1, -1, 0, 1, 1, 2, 2, 1, 1, 1, 0, 0, 0, 2, 2, 2, 3, 2, 3, 2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 3, 1, 1, 1, 0, 0, 0, 0, 2, 2, 2, 4, 4, 3, 2, 1, 1, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 1, 1, 1, 3, 3, 1, 1, 1, 1, 2, 0, 1, 0, 0, 0, 2, 3, 3, 2, 1, 0, 1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 2, 2, 3, 0, 1, 1, 2, 3, 2, 1, 1, 0, 1, 1, 3, 2, 2, 2, 2, 1, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 2, 4, 4, 2, 1, 1, 1, 2, 1, 1, 0, 1, 2, 2, 1, 2, 1, 2, 2, 3, 2, 2, 2, 0, 1, 1, 1, 0, 0, -1, 0, 0, 2, 3, 4, 3, 3, 2, 2, 2, 3, 1, 1, 2, 1, 2, 1, 2, 1, 1, 3, 3, 3, 3, 2, 2, 1, 1, 0, -2, 0, 0, -1, 0, 2, 5, 5, 4, 4, 4, 3, 2, 3, 3, 1, 2, 0, 1, 2, 2, 1, 1, 0, 1, 1, 2, 1, 2, 1, 0, 0, -2, 0, 0, 0, 0, 2, 5, 5, 3, 4, 3, 2, 2, 3, 2, 1, 2, 0, 1, 1, 1, 0, 1, 1, 1, 1, 0, 2, 0, 0, 0, -1, -1, -1, 0, 0, 0, 2, 4, 4, 3, 4, 3, 4, 4, 2, 2, 1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 2, 5, 3, 4, 3, 3, 1, 1, 1, 0, 0, -1, 0, 1, 2, 2, 0, 1, 1, 2, 1, 1, 2, 0, 1, 1, 1, 0, 0, 0, 1, 1, 3, 3, 3, 4, 4, 2, 1, 2, 1, 1, 0, 0, 1, 2, 2, 2, 2, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 3, 4, 4, 3, 1, 1, 0, 1, 1, 0, 1, 2, 1, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 1, 1, 3, 2, 2, 0, 1, 1, 0, 1, 1, 2, 1, 0, 2, 1, 0, 0, 1, 1, 0, 0, 0, 0, 2, 0, 1, -1, -2, -3, -2, -1, 0, 1, 2, 2, 1, 0, 0, -1, 0, 0, 1, 1, 1, 1, 1, 2, 1, 2, 2, 3, 1, 0, 0, 1, 0, 1, 0, 0, -3, -2, -3, -3, -1, 0, 1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, 2, 2, 3, 3, 1, 1, 0, 1, 0, 0, 0, 0, -1, -2, -2, -3, -3, -2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, -1, -1, -1, -2, -2, -2, -2, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, -3, -3, -2, -3, -2, -1, 0, -1, -1, -1, 0, 0, 0, -2, -3, -2, -1, -2, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, -3, -3, -2, -2, -1, -2, -1, -1, 0, 0, -1, 0, -1, -2, -1, -1, -1, -1, -2, -2, -1, -2, -1, 0, -2, -2, -2, 0, 0, -1, -1, -1, -1, -2, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -2, -2, -1, 0, 0, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 2, 0, 1, 0, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 2, 2, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 2, 2, 2, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, -2, -2, -1, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 2, 0, 3, 3, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 2, 2, 1, 2, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 2, 2, 1, 1, 1, 2, 1, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 1, 1, 1, 2, 1, 1, 1, 1, 0, 1, 1, 0, -1, -1, 0, 1, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 1, 0, 1, 1, 1, 2, 0, 2, 2, 2, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -2, -2, -2, -1, 0, 0, 1, -1, -1, 0, 1, 1, 1, 0, 1, 2, 1, 3, 1, 1, 2, 1, 0, 0, 0, 1, 0, 1, 0, -1, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 2, 2, 1, 2, 2, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -2, -2, -1, -1, -1, 0, 0, -1, 0, 1, 1, 1, 1, 1, 1, 2, 3, 2, 1, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, -2, -1, -1, -1, 0, -1, 0, 0, 0, 0, 2, 3, 2, 3, 1, 1, 1, 3, 3, 2, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, -3, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 3, 2, 2, 1, 1, 2, 3, 2, 1, 1, 2, 0, 0, -1, 0, -1, 1, 0, 0, 0, -2, 0, 0, 0, 1, 1, 0, 0, 1, 2, 1, 2, 2, 3, 3, 1, 2, 3, 2, 2, 2, 1, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 1, 1, 2, 2, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -2, -2, -2, -2, 0, -1, 0, 0, 0, 0, 1, 1, 2, 1, 2, 1, 2, 0, 1, 1, 2, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 1, 2, 3, 2, 2, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, -2, 0, 0, 2, 0, 1, 1, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, -2, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, -1, -1, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, -1, 0, -1, 0, -1, -2, -1, -1, -1, -1, -1, -2, -1, -1, -1, -1, -1, 0, -1, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, -2, 0, -1, -1, -1, 0, -1, 0, -1, 0, -2, -2, -1, -1, 0, -1, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, -1, 0, -1, -2, -1, -2, -2, -2, 0, -2, 0, 0, 0, -2, -1, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, -1, -1, 0, -1, -2, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 2, 1, 2, 2, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 2, 3, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 2, 1, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 1, 2, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 2, 2, 3, 2, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 1, 1, 3, 1, 2, 1, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 2, 2, 2, 2, 0, 1, 0, 0, 0, 0, 0, -2, -1, 0, 1, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 2, 1, 2, 1, 2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 2, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -2, -2, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -2, -2, -2, -1, -2, -1, -2, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, -2, -1, -1, 0, 0, -1, -1, -1, -2, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, -1, -2, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, -2, -1, -1, -1, -2, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, -2, 0, -1, -1, 0, 0, 0, 0, -2, -2, 0, -1, -1, -2, -2, -2, -3, -2, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -2, -2, -1, -1, -1, -1, -1, 0, -2, -2, -2, -1, -1, -1, -2, -1, -2, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, -2, 0, -1, -1, -1, 0, -2, -2, -1, -2, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, -1, 0, -1, -1, -2, -1, 0, 0, 0, -2, -2, -2, 0, -1, 0, -1, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, -1, -1, 0, -1, -2, -1, 0, -2, 0, -1, -1, 0, 0, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -2, 0, 0, 0, -1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -2, 0, -1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 2, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, -2, 0, 0, 0, 1, 3, 3, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, -2, 0, 0, 0, 2, 1, 1, 3, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 1, 2, 3, 1, 1, 2, 1, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 2, 1, 2, 0, 0, 1, 0, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 2, 2, 1, 2, 2, 2, 2, 0, 1, 1, 0, -1, -1, 0, 1, 1, 0, 0, -2, 0, 2, 1, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 2, 1, 2, 2, 2, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 2, 2, 1, 2, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 0, 2, 2, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 1, 1, 2, 1, 2, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 2, 2, 1, 2, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 1, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 2, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -3, -1, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, -1, 0, 0, 0, -2, -2, 0, -1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 2, 2, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 1, 0, 1, 0, 3, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 1, 2, 0, 2, 1, 2, 1, 3, 2, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, -2, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -2, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, -1, 0, -2, -2, -2, -2, -1, -2, -1, -1, -1, 0, -1, -2, -2, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, -3, -3, -3, -2, -1, -1, 0, 0, -2, -2, 0, 0, -1, -1, -1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -3, -2, -3, -3, -2, -2, -1, 0, -1, -1, -1, -1, -1, -1, -2, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -3, -2, -2, -3, -3, -3, -1, -2, -1, -2, -2, -2, -2, -1, 0, -2, -2, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -2, -1, 0, -2, -1, -2, -2, -2, -1, 0, -1, -1, -3, -2, -3, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, -1, -1, -2, -2, -3, -1, 0, 0, -3, -3, -2, -1, -1, 0, -1, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, -2, -1, -2, -1, -2, -2, -1, -1, -1, -1, -2, -1, -2, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -3, 0, 0, 0, -1, 0, -1, -2, -2, -1, 0, -1, -2, -1, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, -2, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 2, 2, 0, -1, 1, 0, 0, 1, 1, 0, 0, -1, -1, -2, -2, -1, -2, -1, -1, 0, 0, 0, -1, -1, 0, -1, -2, -1, 0, -1, 0, 1, 3, 2, 0, 0, 1, 0, 2, 0, 1, 0, 0, 0, -1, -1, 0, -1, -1, -2, -1, -1, -1, 0, 0, -1, 0, -1, -2, -1, 0, -1, -1, 0, 2, 0, 0, -1, 1, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, -1, -2, -1, -2, -1, -1, -1, -1, 0, -1, -1, -1, -1, -1, 0, 0, 2, 1, 0, 0, 1, 2, 2, 0, 1, 0, 0, 0, 0, -1, -1, -1, -2, -1, -2, -2, -1, -1, -1, -1, -1, -1, -2, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 3, 1, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, -2, -1, -2, -2, 0, 0, 0, -1, -1, -2, -2, -1, -1, 0, 0, 0, 2, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, -1, -1, -2, -1, -2, -3, -1, 0, -1, 1, -1, -1, -1, -1, -1, -1, 0, 1, 0, 1, 0, 0, 0, 2, 2, 0, 0, 0, 0, 1, 1, 0, -1, -2, -1, -1, 0, -1, -2, -2, -1, 0, 0, 0, -2, -2, 0, 0, 0, 0, 2, 3, 0, 1, 1, 1, 2, 1, 1, 1, 0, 0, 1, 0, 0, -2, -3, -2, -2, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 3, 0, 2, 3, 2, 2, 0, 0, 0, 1, 1, 0, 0, -1, -2, -1, -2, -2, 0, -2, -1, 0, 0, -1, -2, -1, 0, 1, 1, 1, 0, 2, 3, 0, 1, 1, 2, 2, 1, 0, 0, 1, 1, 1, 0, 0, -2, -1, 0, -1, 0, -2, -1, 0, 0, 0, 0, -1, 0, 1, 1, 1, 1, 1, 3, 0, 0, 0, 2, 2, 2, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 3, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 2, 4, 0, 0, 1, 2, 1, 1, 1, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 1, 1, 2, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 1, 1, 2, 1, 1, 2, 1, 1, 3, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 2, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, 0, -2, -2, -2, -1, -3, -1, -1, -2, -1, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, -1, -1, -1, -1, -1, 0, -1, 0, -1, -1, 0, -2, 0, 0, -1, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 1, 0, 2, 1, 1, 2, 1, 1, 1, 1, 1, 0, 0, 0, 0, 2, 1, 1, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 2, 0, 2, 1, 1, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, 0, 1, 1, 1, 0, 1, 2, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 2, 1, 2, 2, 1, 1, 1, 1, 1, 0, 0, 1, 0, 1, 2, 1, 2, 3, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 2, 1, 1, 2, 2, 1, 1, 0, 1, 2, 0, 1, 0, 1, 1, 2, 2, 2, 1, 2, 1, 1, 1, 1, 1, 0, 1, 1, 2, 1, 0, 1, 0, 1, 2, 2, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 2, 1, 0, 0, 1, 1, 0, 0, 2, 1, 0, 1, 0, 1, 1, 0, 1, 3, 1, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 2, 3, 2, 2, 1, 1, 1, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 3, 3, 2, 3, 3, 1, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 3, 1, 1, 2, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 1, 2, 2, 3, 1, 0, 0, -1, -1, -1, -2, 0, -1, -1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 2, 2, 1, 1, 2, 1, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 2, 2, 1, 1, 0, -1, -1, -2, -2, 0, -2, -1, -2, -1, -2, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 1, 1, 0, 0, 0, -1, -2, -2, -2, -1, -2, -2, -1, -3, -2, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -2, -2, -3, -2, -2, -2, -1, -2, -2, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -2, -2, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, 0, -1, -1, -2, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -2, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -2, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, -2, -1, -2, -2, -2, -4, -3, -3, -3, -4, -5, -4, -3, -3, -1, 0, -2, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, -2, -3, -2, -4, -3, -2, -3, -3, -3, -3, -2, -1, -1, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 2, 2, 0, 1, 0, 2, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, 1, 2, 0, 1, 1, 0, 1, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 2, 1, 0, 0, 0, -1, 0, 0, -1, 0, 2, 3, 1, 1, 2, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 2, 1, 1, 0, 0, -2, 0, 1, 2, 1, 0, 0, 0, 0, 2, 1, 1, 2, 1, 1, 1, 0, 0, 2, 2, 1, 0, 2, 2, 1, 2, 2, 1, 2, 0, 0, 0, -2, -1, 1, 1, 1, 1, 0, 0, 1, 2, 2, 2, 0, 0, 0, 1, 1, 0, 1, 2, 2, 0, 0, 0, 1, 2, 1, 2, 1, 1, 0, 0, -1, 0, 1, 2, 1, 1, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 2, 1, 1, 0, -1, -1, -1, 0, 2, 1, 3, 1, 0, 0, 0, 0, 0, 2, 1, 2, 2, 2, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 2, 2, 2, 0, 0, 0, -1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 3, 2, 0, 1, 0, 0, -1, 0, 1, 0, 0, 1, 2, 1, 2, 0, 2, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 2, 1, 3, 3, 2, 1, 0, -1, -2, 0, 0, 0, 1, 1, 2, 3, 3, 2, 2, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 3, 2, 4, 3, 2, 0, -1, -2, -1, -3, -2, 0, 0, 2, 4, 4, 2, 1, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 1, 3, 4, 4, 4, 1, 0, 0, -2, -2, -1, -2, 0, 0, 1, 3, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, -1, 0, 0, 1, 2, 3, 3, 3, 1, 0, -1, -2, -1, 0, 0, 0, 0, 1, 3, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 2, 4, 2, 2, 1, 1, 0, 0, -1, -1, -1, -2, 0, 0, 2, 2, 0, 0, 0, 1, 0, 0, 0, 0, -1, 1, 0, -1, -1, -1, 0, 0, 2, 3, 4, 2, 1, 2, 0, -1, -2, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, -2, 0, 0, 0, 0, -2, -2, 0, 0, 0, 2, 4, 3, 1, 1, 0, 1, -1, -1, -1, 0, -2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 2, 2, 2, 0, 0, 0, 0, -3, -3, -2, -2, -1, -1, -1, 0, 2, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, 1, 1, 0, 0, 0, -1, -1, -2, -3, -4, -3, -3, -2, -1, 0, 2, 3, 3, 2, 1, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -2, -2, -3, -4, -2, -2, -1, 0, 2, 2, 4, 1, 1, 0, 1, 2, 0, 2, 1, 1, 0, -1, -1, 0, -2, -2, 0, 0, -1, 0, 0, 0, -1, -2, -3, -3, -2, -1, 0, 1, 3, 2, 3, 1, 2, 0, 1, 0, 0, 1, 0, 1, 0, -1, 0, 0, -2, -2, -1, -2, 0, 0, 0, 0, -1, -2, -2, -3, -1, 0, 0, 1, 2, 2, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -3, -3, -2, 0, 0, 0, 0, 0, -1, -3, -1, 0, 0, 0, 0, 2, 2, 1, 1, 1, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -3, -4, -1, -1, -1, 0, 0, 0, -1, -2, -2, 0, 0, 0, 2, 2, 1, 2, 1, 2, 2, 2, 2, 1, 1, 0, 0, 0, 0, -1, 0, 0, -5, -3, -2, -2, -1, 0, 0, 0, 0, -1, 0, 0, 2, 2, 2, 2, 1, 1, 1, 2, 2, 2, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -4, -2, -1, -1, -1, 1, 0, 1, 0, 0, 0, 2, 2, 3, 3, 2, 0, 1, 1, 3, 1, 0, 1, 0, 0, -1, 0, 0, 0, -2, -1, 0, -2, -2, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 3, 2, 1, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, 1, -2, -1, 0, 0, 0, 1, 2, 1, 0, 1, 1, 0, 1, 2, 1, 0, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 3, 2, 1, 0, 0, 0, 0, -2, -1, -2, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 2, 0, 1, 1, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 2, 1, 0, 1, 0, 0, 1, 1, 3, 3, 2, 2, 2, 2, 1, 1, 1, 1, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 2, 1, 0, 2, 2, 1, 2, 2, 1, 3, 3, 4, 5, 4, 4, 4, 3, 2, 1, 2, 2, 1, 2, 2, 2, 0, 1, 1, 0, 1, 1, 1, 1, 0, 1, 1, 2, 2, 2, 3, 1, 3, 2, 3, 5, 3, 3, 3, 2, 2, 3, 2, 1, 1, 1, 2, 2, 0, 0, 1, 2, 2, 1, 2, 2, 2, 2, 2, 1, 1, 0, 1, 1, 1, 2, 2, 3, 2, 2, 1, 2, 3, 1, 1, 2, 1, 2, 3, 3, 1, 2, 2, 1, 2, 1, 2, 3, 2, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 2, 1, 0, 0, 0, 1, 0, 1, 0, 0, 2, 1, 0, 2, 2, 3, 3, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 3, 1, 0, 1, 1, 3, 3, 2, 2, 2, 2, 1, 0, 0, 1, 0, 0, -1, -1, -2, -2, -1, -2, -2, -2, -3, -2, -1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 2, 1, 2, 1, 2, 2, 1, 0, 1, 0, 1, 0, 0, -2, -4, -2, -3, -3, -2, -3, -2, -3, -3, -2, 0, -1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 1, 2, 1, 1, 2, 1, -1, -3, -3, -4, -6, -6, -5, -3, -2, -4, -4, -3, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 0, -1, -2, -3, -5, -7, -6, -5, -4, -3, -5, -5, -4, -1, 0, 1, 2, 0, 0, 1, 0, -1, -1, -2, -2, -1, 0, 0, 0, 1, 1, 1, -1, -1, -3, -3, -4, -6, -5, -4, -3, -2, -4, -5, -1, -1, -1, 0, 2, 2, 0, 0, 0, -3, -4, -5, -6, -4, -1, 0, 0, 0, 0, 0, -1, -2, -3, -3, -3, -5, -5, -5, -4, -2, -2, -3, -1, 0, -1, 0, 2, 1, 0, 0, -1, -2, -3, -5, -5, -6, -4, -3, -2, 0, -2, -1, -2, -3, -3, -4, -4, -4, -4, -5, -4, -2, -3, -1, -1, 0, -1, 1, 1, 1, 0, -2, -2, -2, -3, -5, -5, -6, -4, -2, -1, -2, -3, -2, -2, -2, -3, -2, -2, -3, -4, -5, -3, -4, -3, -1, 0, 1, -1, 1, 2, 0, -2, -2, -2, -3, -3, -6, -5, -6, -4, -2, -1, -1, -2, -2, -2, -3, -3, -3, -2, -3, -4, -4, -3, -4, -4, -3, 0, 0, -1, 2, 2, 0, -2, -4, -3, -2, -5, -5, -5, -6, -4, -2, 0, 0, -1, -3, -3, -3, -2, -2, -3, -5, -4, -3, -2, -2, -3, -2, -2, 0, -1, 1, 2, -1, -3, -3, -1, -3, -5, -4, -5, -4, -5, -2, 0, 0, 0, 0, 0, -1, -3, -2, -4, -5, -3, -3, -2, -3, -2, -2, -2, -1, -1, 0, 1, 0, -3, -2, 0, -3, -4, -3, -4, -5, -2, -2, 0, 0, 1, 0, 0, -1, -1, -2, -3, -3, -2, -4, -2, -1, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, -2, -3, -5, -4, -2, -1, 0, 0, 0, 2, 0, -1, -2, -2, -1, -1, -3, -1, -3, -1, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -2, -4, -3, -3, -2, 0, 1, 1, 1, 1, -1, -2, -3, -1, -1, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -4, -4, -3, -1, 0, 1, 2, 0, 0, 0, -2, -2, -2, -3, -2, -4, -2, -1, 0, -2, 0, 1, 1, -1, 0, 0, 1, 1, 0, 1, 0, -1, -1, -2, -2, 0, 0, 2, 2, 0, 0, -1, -1, -2, -2, -2, -2, -4, -2, -2, -2, -1, -1, 1, 0, -1, 0, 0, 1, 1, 1, 1, 1, 0, -2, -1, 1, 1, 0, 1, 1, 0, 0, 0, -2, -2, -2, -2, -3, -4, -3, -2, -2, -1, -1, 0, 0, -1, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, -1, -2, -1, -2, -1, -2, -3, -3, -2, -1, -1, 0, 0, 0, -2, 0, 1, 3, 2, 2, 1, 0, 0, 0, 2, 3, 2, 2, 0, 1, 0, 0, -1, -1, -2, 0, 0, -1, -2, -3, -2, -1, -2, -1, 1, 1, 0, 0, 1, 2, 2, 2, 2, 0, 0, 1, 1, 3, 3, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, -1, -2, 0, 0, 1, 0, -1, 0, 1, 2, 3, 3, 2, 1, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 1, 2, 3, 3, 2, 3, 1, 2, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 1, 3, 3, 2, -1, 0, 1, 1, 0, 2, 2, 2, 0, 1, 0, 0, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 2, 3, 2, 1, 1, -1, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, -1, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    -- filter=0 channel=6
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -2, -2, -1, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, -1, -1, 0, -1, -2, -2, -1, -2, -3, -2, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 2, 0, 0, 0, -1, -1, -1, 0, 0, 0, -2, -1, -1, -1, -1, -1, -2, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, -1, -2, -2, -1, -2, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -2, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -2, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 1, 2, 2, 2, 1, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 3, 2, 2, 4, 3, 3, 2, 2, 2, 0, 0, 0, 0, -1, -2, -2, -1, -1, -1, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 2, 2, 3, 3, 4, 3, 3, 3, 3, 2, 0, 0, 0, -1, -1, -1, -2, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 3, 3, 4, 3, 4, 4, 4, 4, 3, 2, 2, 0, 1, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, 0, 0, 1, 0, -1, 0, 1, 2, 1, 1, 3, 3, 4, 3, 3, 2, 3, 3, 2, 2, 1, 1, 0, 0, -1, 0, -1, 0, -2, -1, -1, -1, 0, 0, 0, 0, -1, 0, 1, 2, 1, 3, 4, 4, 4, 2, 2, 3, 3, 2, 3, 3, 1, 1, 0, -1, -1, -1, -1, -1, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 1, 1, 1, 2, 3, 4, 4, 2, 2, 2, 2, 1, 2, 2, 2, 0, 0, 0, -1, 0, 0, -1, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 2, 3, 3, 3, 3, 2, 1, 4, 2, 2, 2, 3, 0, 0, 0, 0, -1, -1, 0, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 3, 2, 3, 1, 3, 3, 3, 3, 2, 1, 0, 0, -1, -1, -1, -2, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 2, 1, 0, 1, 1, 0, 2, 1, 1, 1, 2, 0, 0, 0, 0, -2, -1, 0, 0, 0, -1, -1, -1, -1, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, -2, -2, -2, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, -2, -1, 0, -1, -1, -1, 0, -1, 0, -1, 0, -1, 0, -2, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, -2, -1, -2, -2, -3, -3, -1, -2, -1, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -2, -2, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -2, -3, -1, -2, -2, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -2, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, -2, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, -1, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 2, 2, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, -1, 0, 0, -1, -1, -2, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -2, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -2, 0, -1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -2, -2, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, -1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -2, -2, -2, 0, 0, 0, 1, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -2, -3, -2, -2, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -1, -1, -3, -2, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -2, -1, -2, 0, 0, -1, -2, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, -2, -2, -1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, 0, 0, -2, -1, -2, -1, -1, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, -2, 0, -1, -1, 0, -1, -2, -1, -2, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, -1, -1, -1, 0, -2, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 1, 1, 2, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 3, 3, 3, 3, 2, 3, 3, 3, 3, 2, 2, 2, 1, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 2, 1, 1, 2, 2, 1, 1, 1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 0, 1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, -1, -2, -1, -1, 0, -1, -1, -1, -1, 0, -1, 0, 0, 1, 1, 2, 0, 1, 0, 0, 0, 0, -1, 0, 0, -2, -1, -1, -1, -1, -3, -2, -2, -3, -1, -1, -1, -1, -1, -2, 0, -1, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -3, -3, -2, -2, -3, -3, -2, -3, -2, -1, -1, -2, -2, -1, 0, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -2, -3, -3, -4, -2, -2, -4, -3, -2, -3, -3, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -3, -3, -3, -3, -3, -3, -3, -3, -2, -2, -2, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, -1, -1, -3, -3, -4, -2, -3, -2, -1, -3, -2, -2, -2, -3, -1, -1, -1, 0, 0, 1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -3, -1, -2, -2, -3, -3, -3, -1, -2, -3, -2, -1, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, -2, -1, -2, -1, -3, -3, -2, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -2, -2, -2, -1, -3, -2, -2, -1, -1, 0, -1, -1, -2, 0, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -2, -2, -2, -1, -1, -1, -2, -2, -1, -1, -1, -1, -2, -1, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -2, -2, -2, -2, -3, -1, -1, -1, -1, 0, -2, -2, -1, -2, -2, -1, -2, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -3, -2, -2, -2, -1, -1, -1, 0, -1, -1, -1, -1, -2, -2, -2, -2, -2, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, -2, -2, -1, -2, -1, -2, -1, 0, 0, 0, 0, -2, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -1, -2, -1, -2, -1, -1, 0, -1, -1, 0, -1, -2, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, -1, -2, -1, -1, -2, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -2, 0, 0, -1, 0, -1, -1, -1, 0, -1, -2, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, -2, -2, -2, -1, -2, -2, -3, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, -1, -1, -1, -1, -2, -2, -2, -2, -2, -3, -2, -3, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, -1, -1, -1, -1, -2, -3, -3, -2, -2, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -3, -2, -1, -1, -2, -2, -2, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, -1, 0, -2, -2, -1, -2, -2, -2, -2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 2, 2, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 2, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 1, 1, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 2, 1, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 2, 0, 1, 1, 1, 0, 1, 0, 0, 2, 2, 2, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 2, 1, 2, 0, -1, -2, -3, -1, -1, 0, 0, 0, 0, -2, -1, 0, 0, -1, 0, 2, 1, 2, 2, 2, 1, 2, 2, 1, 1, 1, 2, 2, 2, 2, 1, 0, -2, -3, -2, -2, 0, 0, 0, 0, -2, -1, -1, -1, -1, -1, 0, 0, 1, 1, 0, 2, 0, 1, 0, 2, 0, 1, 1, 1, 3, 2, 3, 2, -2, -1, -2, 0, 0, 0, 1, 0, 0, -1, -1, -2, -1, -2, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 3, 3, 4, 2, 1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, -2, -1, -3, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 3, 2, 2, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, -2, -2, -2, -2, -2, -3, -2, -2, -1, -1, 0, 0, 0, -2, -2, -1, 0, 1, 1, 2, 1, 1, 0, -1, 0, 0, -1, 0, 0, 0, -1, -2, -1, -1, -2, -2, -3, -4, -3, -3, -1, -2, -1, 0, 0, -1, -2, 0, -1, 0, 0, 1, 2, 1, 0, -1, -1, 0, -1, 0, -2, -2, -2, -2, -1, -1, -3, -4, -2, -3, -3, -3, -2, -3, -1, -2, -2, 0, -1, -1, 0, 0, 0, 2, 1, 1, -1, -2, 0, 0, 0, 0, -1, -1, -1, -1, -2, -1, -2, -2, -2, -3, -3, -4, -4, -4, -3, -3, -3, -2, -2, -1, -1, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -2, -1, -2, 0, -1, -1, -2, -2, -1, -1, -3, -2, -3, -3, -4, -4, -3, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -2, -1, -2, -1, -1, -1, -2, 0, -3, -4, -4, -4, -4, -4, -3, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, -1, -1, -2, -2, -2, -2, -1, -1, -1, -1, -2, -4, -4, -3, -4, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, -1, 0, -1, -3, -2, -1, -1, -1, 0, 0, -2, -3, -4, -3, -3, -3, -3, -1, 0, 1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, -2, -1, -2, -2, -2, -2, 0, 0, -2, -2, -4, -3, -2, -3, -3, -1, 0, 0, 0, 0, -1, 0, 0, -1, -2, 0, 0, 1, 0, 0, 0, -1, -1, -2, -2, -2, -1, -1, -1, -1, -2, -2, -2, -2, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, -1, -1, -1, -2, -2, -2, -3, -1, -1, 0, -1, -3, -3, -2, -2, -2, -2, -2, -2, -1, 0, 0, -2, 0, 0, 0, -1, 0, 2, 0, 1, 0, 0, 0, -2, -2, -2, -2, -2, -1, 0, 0, -2, -1, -2, -1, -2, -2, -2, -3, -2, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, -2, -2, -2, -2, -2, -2, -1, -1, -1, -2, -1, -1, -1, -2, -3, -4, -3, -2, 0, -1, 0, 0, 1, 0, -1, 1, 1, 0, 0, 0, 0, -2, -3, -2, -3, -3, -1, 0, -1, 0, -2, 0, 0, -1, -1, -1, -3, -4, -1, -3, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, -3, -2, -2, -1, 0, 0, -1, -2, -1, 0, -1, -1, -2, -2, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -4, -2, -2, -1, 0, -1, -1, -2, -2, -1, -2, -1, -2, -2, 0, 0, 0, 0, 0, 0, 1, -1, -1, -1, -1, 0, 0, 1, -1, -2, -3, -3, -2, -2, -1, -2, -2, -2, -2, -1, -2, -3, -1, 0, 0, -2, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 1, -1, -2, -3, -2, -1, -2, -1, -2, -2, -2, -2, -3, -3, -2, -2, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, -2, -2, -3, -1, -1, -2, -2, -3, -3, -3, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 0, -1, -1, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, -3, -2, -2, -3, -1, -2, -1, -1, 0, -1, 0, 0, 0, 0, 1, 2, 2, 2, 0, 0, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 3, 4, 2, 0, 0, -2, -2, 0, 0, 0, 0, -1, 0, -1, 0, 0, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 3, 3, 3, 2, 0, -2, -1, -1, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 3, 4, 3, 1, 0, -1, -3, -2, -1, 0, 0, -1, -1, -2, -1, -2, -2, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 4, 3, 2, 2, 0, 0, -2, -4, -3, -3, -2, -2, -1, -3, -2, -2, -1, -1, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 2, 2, 2, 1, 1, -1, -3, -3, -4, -1, -2, -1, -2, -2, -2, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 2, 0, 1, 1, 2, 3, 1, 2, 0, 0, -2, -3, -3, -2, -1, -2, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 2, 0, 1, 1, 2, 2, 1, 1, 3, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 1, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, -2, -1, -2, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, -2, -2, -1, -2, -1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -2, -2, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -2, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, -2, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -2, -1, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -2, -2, -2, -1, -1, 0, -1, 0, 0, 0, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, -1, -1, -2, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -2, -1, -1, -1, -2, -1, -1, -1, 0, 0, -1, -1, -2, -1, -1, -1, 0, -1, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, -2, -1, -2, -1, -1, -2, 0, 0, -1, 0, -1, 0, -1, 0, 0, -2, -1, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -2, -2, -2, -3, -1, -1, -2, -1, -2, 0, 1, 0, 0, -1, -2, -2, -1, -1, -1, -1, -1, -2, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, -2, -1, -3, -1, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, -2, -1, 0, -2, 0, -1, 0, 0, -1, -1, -1, 0, -1, -2, -2, 0, -1, -1, -2, 0, -1, 0, 0, -1, -1, -1, -1, 0, -1, -2, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -2, -3, -2, -1, -2, -1, 0, -2, 1, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, -2, -2, -1, 0, 0, -1, 0, -2, -1, -1, -1, -2, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, -2, 0, -1, -1, 0, 0, 0, 0, 0, -1, -2, -2, -1, 0, -1, 0, -1, -2, 0, 0, -1, -1, -2, -2, -2, -1, -1, -1, 0, 1, 0, -1, 0, -2, -2, -1, 0, -1, 0, -1, -1, -2, -2, -1, 0, 0, 0, -2, -1, -1, -1, -1, -1, -2, 0, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, -2, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, -2, 0, -1, -1, 0, -1, -2, -1, -1, -1, 0, 0, 0, 1, 0, -1, 0, -1, -1, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, -2, -2, -1, -2, -1, 0, -1, 1, 1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -2, -1, -1, 0, -1, 0, -2, 0, -2, -1, -2, -2, -1, -1, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -2, -1, 0, -1, 0, -2, -2, -1, -1, -1, -1, -1, -1, 0, 0, 0, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, -2, 0, -1, -1, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, -2, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -2, -1, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, -1, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -4, -5, -3, -2, 0, 0, 0, -1, -2, -2, -1, -2, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, -1, -4, -4, -2, -1, 0, 0, 0, 0, -1, -1, -1, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, -2, -3, -4, -2, -1, 0, 0, 0, 0, 0, -1, -1, -2, -3, -1, -2, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, -1, -2, -1, 0, 0, 0, -1, 0, 0, -1, -2, -2, -2, -3, -4, -4, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, -1, -3, -1, 0, -1, 0, -1, -1, -1, -1, -1, -3, -4, -4, -4, -4, -4, -3, -2, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -2, -1, -1, -1, -1, -1, -1, -2, -2, -2, -3, -2, -2, -2, -2, -3, -4, -2, -3, -1, -2, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, -3, -2, 0, -1, -2, -1, -1, -2, -3, -2, -2, -2, -2, -2, -3, -3, -4, -4, -3, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, -2, -3, -1, -1, -2, -1, -1, -2, -1, -1, -1, -1, -2, -2, -3, -1, -3, -3, -2, -2, -4, -3, -2, -2, -1, -1, -1, -2, -1, 0, 0, 0, -1, -2, -2, -1, -2, -2, -2, -3, -2, -2, -1, -2, -1, -2, -2, -1, -1, -3, -4, -4, -3, -2, -3, -2, -2, -2, -2, -1, -2, 0, 0, -1, -1, -1, -2, 0, -1, -2, -2, -1, -1, -1, -2, -3, -3, -2, 0, 0, -1, -1, -2, -3, -3, -3, -3, -3, -2, -2, -1, -1, 0, -1, -1, -1, 0, -2, -2, 0, 0, -1, -2, -3, -2, -2, -3, -2, -2, -2, -1, 0, -1, -1, -1, -3, -4, -4, -3, -5, -2, 0, 0, -1, -1, -2, -2, 0, -1, -1, -1, -2, -1, -1, -1, -2, -2, -1, -3, -2, -1, -2, 0, -1, 0, -1, -1, -2, -3, -4, -4, -3, -3, -2, 0, 0, -1, -1, -1, -2, -1, -2, -2, 0, 0, 0, 0, -2, -1, -1, -1, -3, -2, -1, 0, 0, 0, 0, -1, -1, -2, -2, -4, -5, -3, -2, -1, -2, -2, -3, -1, -1, 0, -2, -1, 0, 0, 0, 0, 0, -1, -3, -3, -2, -2, -1, -1, 0, 0, -1, 0, -2, -2, -3, -3, -4, -5, -3, -3, -1, -3, -2, -3, -1, 0, 0, 0, -1, 0, 0, 0, -2, -1, -2, -2, -1, -2, -1, 0, 0, 0, 0, -1, 0, -2, -3, -2, -4, -4, -4, -3, -2, -3, -4, -4, -1, -1, -1, -1, -1, 0, 0, 0, -2, -3, -3, -3, -2, -1, -1, 0, 0, -1, 0, 0, -2, -1, -3, -2, -4, -4, -4, -4, -2, -3, -2, -3, -1, 0, -2, -1, 0, -1, -1, -1, -2, -2, -4, -3, -1, -1, -2, -1, -2, 0, 0, -2, -1, -1, -2, -2, -4, -4, -5, -4, -2, -3, -3, -2, 0, -1, -2, 0, -1, -1, -2, -1, -2, -2, -3, -3, -2, -2, -2, -1, -1, -1, 0, -2, -1, -1, -2, -2, -5, -4, -4, -2, -2, -2, -2, -2, -1, -1, -2, -1, 0, -2, -2, -2, -1, -3, -3, -3, -2, -4, -3, -1, -1, 0, -2, -1, -2, -1, -2, -4, -5, -5, -4, -2, -3, -3, -1, -2, 0, -1, -2, -2, 0, 0, -1, -1, -1, -3, -4, -5, -4, -4, -2, -1, -1, -2, -3, -1, -2, -2, -3, -2, -4, -4, -3, -4, -2, -2, -2, -2, 0, -2, -2, -2, -2, 0, 0, 0, 0, -2, -3, -3, -3, -3, -3, -2, -3, -3, -3, -3, -2, -4, -2, -3, -3, -2, -3, -4, -1, -2, -2, -2, 0, -1, -2, -3, 0, -1, 0, 0, -1, -3, -2, -4, -2, -2, -2, -3, -4, -3, -3, -4, -3, -3, -2, -1, -1, -2, -2, -2, -2, -1, -2, -1, 0, 0, -2, -2, -1, -1, 0, 0, 0, -1, -3, -3, -2, -3, -3, -4, -3, -4, -4, -4, -2, -2, -1, 0, -1, -1, -1, -2, -1, 0, -2, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, -2, -1, -1, -3, -4, -3, -3, -4, -3, -3, -2, 0, 0, -1, -1, 0, -1, 0, -2, 0, 0, 0, 1, -2, -2, -1, 0, 0, 0, 0, -1, -1, 0, 0, -2, -1, -3, -3, -4, -4, -2, -1, -1, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -2, -1, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, -2, -3, -2, -3, -2, -2, -2, -2, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, -2, -2, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 2, 2, 2, 1, -1, -4, -4, -2, -2, 0, 0, 0, -1, -1, -1, -1, -2, -1, 0, 0, 0, 0, -1, 0, -1, -2, 0, -1, -1, -1, 0, 1, 0, 1, 2, 1, -1, -4, -4, -4, -3, -2, 0, -1, 0, -2, -1, 0, -1, -1, 0, 0, 1, 0, -1, 0, -1, -1, 0, 0, -1, -1, 0, 2, 1, 1, 1, 0, -1, -3, -5, -4, -2, -1, -1, 0, -2, -1, -1, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 3, 2, 0, 1, 0, 0, -3, -2, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 2, 2, 0, 0, 0, 1, 0, 2, 1, 0, 1, 1, 1, 2, 1, 0, 2, 2, 1, 2, 1, 3, 1, 2, 2, 3, 3, 3, 1, 2, 2, 3, 2, 1, 1, 0, 2, 2, 3, 1, 2, 1, 1, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 2, 3, 2, 3, 3, 4, 5, 4, 2, 1, 0, 1, 3, 2, 0, 1, 0, 0, 1, 0, 0, -1, -2, -1, -3, -4, -3, -2, -1, 0, 0, 0, 1, 1, 2, 3, 3, 3, 4, 4, 3, 3, 0, 1, 2, 2, 2, 1, 0, 0, 0, 0, -1, -2, -2, -3, -3, -4, -4, -3, -2, -1, 0, 0, 0, 0, 0, 1, 1, 3, 5, 5, 3, 1, 1, 1, 2, 2, 0, 1, 0, -1, 0, 0, -1, -1, -3, -4, -4, -6, -5, -3, -2, 0, 0, 0, 0, -1, 0, 0, 0, 2, 3, 3, 3, 1, 1, 0, 1, 0, 1, 0, 0, -1, 0, -1, -3, -4, -3, -4, -7, -6, -6, -4, -3, 0, 0, 0, 0, -2, -2, 0, 0, 2, 2, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -4, -6, -5, -5, -6, -6, -8, -5, -4, -2, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -2, -2, -1, -3, -6, -5, -6, -6, -7, -7, -7, -7, -5, -4, -4, -3, -2, -2, -2, 0, -1, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, -2, -1, -1, -1, -4, -5, -6, -7, -7, -7, -7, -6, -5, -5, -3, -4, -2, -3, -1, -1, 0, 0, 0, -1, -1, -1, 0, -1, 1, 0, 0, 0, 0, -1, 0, -2, -4, -4, -4, -5, -7, -6, -5, -4, -2, -3, -3, -3, -2, -2, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 1, 1, 1, 0, 0, 0, -1, 0, -2, -3, -3, -2, -3, -2, -1, -1, 0, 0, -2, -2, -2, -2, -2, -2, -1, 0, 0, -1, -1, -2, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 3, 2, 0, 0, -1, 0, -3, -3, -2, -2, -1, -1, -1, -2, -3, -1, -1, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 2, 2, 3, 5, 4, 5, 4, 3, 1, 0, 0, -2, -2, -3, -3, -2, -2, -3, -2, -2, -2, -1, 1, 0, 0, -1, -1, -2, 0, 0, 0, 1, 2, 2, 3, 5, 6, 6, 6, 3, 3, 1, 0, 0, -1, -2, -4, -3, -3, -4, -3, -3, -3, -1, 1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 3, 2, 3, 5, 6, 6, 5, 4, 3, 4, 2, 2, -1, -4, -5, -4, -4, -5, -2, -3, -2, -1, 0, 0, -1, -1, -1, 0, 1, 0, 2, 2, 2, 4, 3, 4, 4, 4, 5, 4, 5, 6, 5, 2, 0, -3, -4, -5, -4, -4, -3, -3, -1, 0, 0, 0, -1, -1, -1, -1, 1, 0, 1, 2, 2, 3, 4, 4, 5, 4, 4, 6, 7, 5, 3, 3, 0, -2, -3, -3, -4, -4, -2, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 4, 4, 3, 3, 4, 6, 6, 6, 7, 6, 4, 1, -1, -3, -6, -4, -4, -3, -3, -2, -1, -1, 0, -1, -2, -2, -1, 0, 0, 0, 0, 2, 2, 2, 3, 3, 6, 5, 6, 6, 7, 6, 3, 0, -2, -6, -5, -5, -5, -3, -3, 0, -1, -1, 0, -1, -1, -2, -1, 0, -1, 1, 1, 2, 1, 4, 3, 4, 4, 6, 5, 6, 6, 2, 0, -2, -4, -5, -6, -3, -4, -4, -2, -2, -2, 0, -1, -1, -2, -2, -2, -1, 0, 0, 1, 0, 1, 2, 3, 2, 4, 4, 3, 1, 1, 0, -2, -5, -5, -4, -4, -4, -2, -2, -1, -2, 0, 0, -1, 0, -1, -2, -2, -1, 0, 0, 0, -1, -1, 0, 1, 0, 0, 1, 1, 0, 0, -2, -4, -4, -3, -3, -3, -3, -2, -3, -1, -2, -1, 0, 0, 0, -1, -1, -2, -1, -1, -2, 0, -3, -2, -1, -2, -2, -1, -3, -2, -1, -1, -3, -4, -3, -2, -2, -1, -2, -1, -1, -3, -3, 0, -1, 1, 0, -1, 0, -2, -2, -1, -2, -1, -2, -2, -3, -3, -6, -6, -6, -5, -3, -2, -4, -3, 0, -2, 0, 0, 0, -1, -1, -2, -2, 0, 0, 1, 1, 0, 0, -1, -2, -1, -1, -1, -1, -2, -4, -6, -6, -7, -6, -6, -6, -4, -3, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 0, 0, 0, -2, 0, -1, -1, -3, -4, -4, -5, -6, -6, -6, -4, -3, -3, -1, 1, 2, 2, 2, 2, 1, 1, 1, 1, 2, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, -3, -3, -3, -5, -6, -5, -4, -3, -3, -1, -1, 1, 3, 2, 2, 2, 2, 3, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -4, -4, -3, -2, -2, -2, -1, 0, 0, 2, 3, 2, 4, 3, 2, 2, 3, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, -1, -1, 0, -1, 1, 0, 2, 3, 3, 4, 4, 3, 3, 2, 1, 0, 1, 0, 0, 2, 1, 1, 2, 2, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 5, 5, 4, 4, 2, 1, 2, 1, 0, 1, 0, 0, 1, 1, 1, 2, 1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 2, 4, 4, 4, 4, 5, 2, 2, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 2, 3, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -2, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -3, -1, -2, 0, -1, 0, 0, 0, 0, -2, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -2, 0, -2, -1, -2, -2, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -2, -2, -2, -3, -2, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 2, 2, 3, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 2, 2, 4, 4, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, -2, 0, 0, 0, 1, 0, 1, 1, 1, 2, 2, 3, 4, 4, 4, 4, 3, 1, 0, 0, 0, 0, -2, -1, -2, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 2, 2, 2, 3, 5, 5, 6, 6, 3, 3, 2, 1, 0, -1, -1, -3, -1, -1, 0, 0, 1, 1, 1, 1, 0, -1, -1, 0, 1, 0, 0, 2, 2, 1, 3, 3, 3, 3, 4, 6, 3, 2, 1, 0, 0, -1, 0, -2, -2, 0, 0, 0, 1, 1, 2, 2, 1, -1, 0, 0, -1, 0, 0, 0, 2, 2, 3, 3, 4, 3, 4, 4, 3, 0, 1, 0, 0, -2, 0, -1, -2, -1, 0, 1, 1, 0, 1, 3, 1, 0, 0, 0, -2, -1, 0, 1, 2, 2, 3, 3, 4, 3, 2, 4, 3, 1, 0, -1, -1, -1, -1, -1, -2, 0, 0, 3, 3, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 2, 2, 3, 3, 4, 3, 3, 2, 1, 0, 0, 0, -1, 0, 0, 1, 1, 2, 2, 2, 4, 2, 1, 2, 0, 0, 0, 0, -1, 0, 2, 1, 1, 3, 3, 4, 2, 3, 1, 1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 2, 3, 2, 2, 2, 1, 1, 0, 1, 0, 0, 0, 0, 2, 2, 3, 2, 3, 4, 4, 1, 2, 2, 2, 0, -1, 0, -1, 0, 0, 0, 1, 2, 2, 1, 1, 2, 0, 0, 0, 1, 0, 1, 0, 1, 3, 3, 2, 2, 2, 4, 3, 2, 0, 1, 2, 1, -1, -1, -1, -1, 0, 1, 2, 2, 3, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 2, 2, 2, 1, 2, 3, 1, 0, 0, 1, 0, -1, -3, -2, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 2, 1, 0, 0, -1, -1, -2, -2, -1, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, -2, -1, -3, -3, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 2, 1, 1, 0, 0, -2, -1, -2, -3, -3, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -2, -2, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 2, 0, 0, -1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 1, 2, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -2, -1, 1, 2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 2, 0, 0, 1, 1, 2, 3, 2, 2, 2, 1, 0, 1, 2, 1, 2, 1, 1, 0, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 1, 0, 1, 0, 1, 2, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 2, 1, 0, 2, 2, 1, 0, 1, 1, -1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 1, -1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -2, -2, -2, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, -1, 0, -1, 0, -1, -2, -2, -2, -2, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -2, -2, -2, -2, -1, -3, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, -2, 0, -2, -2, -1, -3, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, -1, -1, -1, -1, -2, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -2, -1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 0, 0, 0, -1, 0, -1, -1, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 2, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, -2, -1, -1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 1, 2, 1, 1, 1, 1, 2, 0, 1, 1, 2, 0, 0, -1, 0, 0, -1, -2, -2, 0, -2, -1, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 2, 2, 2, 2, 1, 1, 2, 2, 1, 0, 0, 0, 0, -2, -1, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 2, 2, 0, 0, 0, 1, 3, 3, 2, 1, 0, -1, -1, -1, -1, -1, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 1, 0, 1, 0, 2, 1, 4, 3, 1, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 2, 2, 1, 1, 1, 1, 2, 1, 3, 2, 2, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 2, 0, 2, 2, 0, 2, 2, 2, 3, 1, 0, -2, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 1, 1, 0, 1, 2, 1, 2, 0, 1, 1, 1, 2, 2, 1, 1, 0, -1, -2, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 2, 1, 2, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 1, 1, -1, -1, 0, 0, 0, -1, 0, -1, 0, -2, -2, -2, 0, 0, -1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -2, -1, -2, -2, -2, -1, -1, 0, 0, 0, 1, 1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, -1, -3, -3, -3, -1, -1, -2, -3, -1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -2, -2, -2, -2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -1, -2, -1, -1, -1, -1, 0, 1, 0, 1, 1, 0, 1, 2, 1, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 2, 2, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 2, 2, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, -1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 1, 1, 2, 1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 1, 0, 1, 1, 1, 0, 1, 1, 0, 1, 1, 2, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 1, 2, 2, 2, 2, 1, 2, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -1, -1, -1, 0, 1, 2, 1, 3, 4, 4, 5, 5, 4, 2, 3, 3, 4, 5, 5, 5, 3, 2, 0, 0, 1, 1, 0, 0, -1, -1, -1, -2, 0, -1, -1, -1, -1, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 3, 3, 4, 3, 4, 2, 2, 0, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 3, 4, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 1, 0, 1, 2, 3, 4, 3, 2, 2, 0, 1, 1, 1, 2, 2, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, -1, -3, -3, -3, 0, 0, 1, 1, 2, 1, 2, 2, 1, 2, 3, 1, 2, 2, 2, 1, 1, 1, 1, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 1, 2, 0, 0, 0, 0, 1, 2, 2, 2, 0, 1, 1, 0, 0, 0, 0, -2, -2, 0, 0, -2, -1, -2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 2, 0, 1, 1, 0, -1, -2, -2, -3, -1, -2, -1, -3, -2, -2, 0, -2, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, -1, -1, -2, -1, -1, -2, -2, -2, -3, -2, -3, -3, -3, -3, -2, -2, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, -2, -3, -3, -3, -5, -4, -4, -5, -5, -5, -4, -2, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, -1, 0, -2, -2, -3, -5, -4, -4, -5, -5, -5, -6, -5, -6, -5, -3, -3, 0, 0, 1, 2, 2, 1, 2, 1, 1, 1, 1, 0, 0, 1, 0, 0, -2, -2, -2, -3, -4, -3, -3, -4, -3, -3, -5, -5, -5, -3, -5, -2, -2, 0, 1, 2, 2, 2, 3, 2, 1, 0, 0, 0, 0, 1, 1, 1, -2, -3, -3, -3, -2, -3, -1, -3, -2, -4, -4, -3, -4, -5, -4, -3, 0, 0, 2, 3, 2, 2, 4, 2, 1, 0, 0, 0, 0, 0, -1, -1, -2, -2, -3, -2, -4, -4, -4, -3, -3, -3, -3, -3, -5, -5, -3, -2, 0, 0, 2, 4, 2, 0, 1, 0, 0, -1, 0, -1, 0, 0, -2, 0, 0, -1, -1, -2, -3, -3, -4, -3, -4, -2, -4, -3, -5, -4, -3, 0, 0, 2, 2, 1, 0, 0, -2, -1, -1, -2, 0, -1, -1, 0, -1, -1, 0, -1, -2, -3, -3, -4, -4, -2, -1, -2, -3, -4, -3, -4, -2, -1, 1, 3, 2, 2, 3, 3, 1, 0, 0, 0, -1, 0, -1, 0, -2, -2, -3, -3, -2, -3, -3, -2, -3, -2, -2, -3, -4, -3, -3, -1, 0, 1, 4, 5, 3, 2, 3, 4, 3, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -4, -2, -1, -2, -2, -3, -2, -2, -1, -2, -1, 0, 0, 0, 3, 3, 2, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -2, -2, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 2, 2, 2, 2, 2, 2, 1, 0, 1, 1, 1, 1, 1, 1, 0, 0, -2, -1, 0, 0, 1, 1, 1, 0, 0, 2, 1, 0, 0, 2, 0, 1, 1, 1, 1, 3, 2, 3, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 2, 2, 2, 3, 2, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 3, 2, 2, 2, 2, 2, 0, 0, -1, 0, 1, 0, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 1, 3, 2, 1, 1, 2, 1, 1, 1, 1, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, 0, -2, -1, 0, 0, 3, 2, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 4, 2, 2, 2, 1, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 2, 4, 4, 4, 2, 2, 2, 1, 0, 0, 2, 1, 0, 2, 2, 2, 0, 1, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 2, 3, 3, 2, 2, 3, 0, 2, 1, 2, 2, 2, 2, 0, 2, 1, 0, 0, 1, 1, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 2, 4, 5, 5, 1, 1, 2, 3, 2, 1, 1, 3, 3, 2, 1, 0, 1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 1, 1, 1, 1, 0, 0, 0, 1, 2, 2, 1, 1, 1, 1, 1, 0, 1, 2, 2, 2, 1, 1, 1, 1, 0, 0, 0, 0, -1, -2, -1, -2, -2, -1, 0, 0, 0, 0, -1, -2, -2, -1, -2, -3, -3, -4, -2, 0, -1, 0, 0, 3, 1, -1, -1, -1, -1, -1, -1, -1, -2, -1, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -2, -1, 0, 2, 1, 0, -1, 0, 1, -1, 0, 1, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 2, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 1, 1, 1, 2, 1, 0, -1, -1, 0, -1, 0, -2, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 2, 1, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, -1, -2, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 2, 1, 1, 0, 1, 0, 0, 0, -1, -1, -1, -1, -1, -2, -2, -2, -2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -1, -2, 0, -1, -1, -1, 0, 1, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 2, 1, 1, 2, 1, 1, 0, -1, -1, 0, -2, -1, -1, -1, -1, 0, -2, -1, -1, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 0, 0, 0, 0, 0, -1, -2, 0, 0, -2, -1, -2, -2, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 2, 1, 0, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 1, 2, 0, 1, 1, 0, 0, 0, 1, 1, 2, 2, 0, 1, 1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -2, -1, 0, 1, 1, 1, 1, 2, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 1, 1, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 2, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 2, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, -1, -1, -1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 0, 1, 2, 1, 2, 1, 1, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 4, 4, 3, 3, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 3, 3, 2, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 3, 3, 3, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 2, 2, 2, 3, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 2, 2, 3, 2, 3, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 2, 2, 1, 1, 2, 3, 1, 1, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 2, 2, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -3, -3, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -2, -2, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -2, -2, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 2, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, -1, -1, -2, -1, -3, -3, -3, -2, -2, -2, -1, 0, -1, -2, -1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -2, -1, -2, -3, -3, -4, -4, -4, -2, -1, -1, -2, 0, -1, -2, -1, 0, 2, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -2, -2, -3, -3, -3, -2, -2, -2, -1, -2, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -2, -1, 0, -2, -3, -4, -3, -2, 0, 0, 0, 0, -2, -2, -2, -1, -2, -1, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -2, -3, -3, -3, -1, 0, -1, 0, -1, 0, -1, -2, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -3, -2, -2, -2, -4, -3, -3, -1, -1, -1, -1, -1, 0, -1, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, -2, -1, -2, -2, -3, -1, -1, -3, -1, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, -2, -2, -2, 0, 1, 0, 0, -1, 0, 1, 0, -2, -2, -2, -2, -1, -1, -1, -1, -2, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, -2, -3, -2, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -2, 0, -1, 0, 0, 0, -1, 0, 0, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, -1, -2, -2, -1, 0, 0, 0, 0, 0, -2, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 2, 1, 3, 3, 3, 3, 1, 0, 0, 1, 0, -1, -2, -1, 0, -1, -2, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 1, 2, 3, 4, 3, 3, 2, 1, 2, 2, 1, 0, -2, -1, 0, -1, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 4, 5, 3, 2, 2, 2, 2, 1, 0, 0, -1, -1, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 3, 2, 4, 4, 3, 2, 2, 2, 3, 4, 2, 0, -2, -3, -2, -1, -2, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 4, 3, 2, 4, 4, 3, 2, 4, 5, 3, 4, 0, -1, -3, -1, -1, 0, -1, 0, 0, 0, 1, 0, -1, -2, 0, 0, 0, 0, 0, 2, 2, 3, 2, 3, 4, 3, 2, 3, 4, 4, 3, 3, 0, -1, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 2, 3, 3, 3, 4, 3, 3, 4, 3, 4, 2, 1, 0, -2, -4, -2, -2, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 2, 2, 3, 3, 4, 4, 2, 3, 3, 2, 0, -1, -2, -3, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, -1, 0, 3, 2, 2, 1, 2, 3, 2, 2, 1, 0, -1, -2, -2, -1, -1, 0, -1, 0, 0, 0, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 1, 1, 0, -2, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 1, 0, -1, -2, -2, -2, -1, -1, -1, -1, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, -1, -2, -3, -4, -3, -4, -3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -2, -2, -1, 0, 0, 0, -2, -2, -1, -3, -4, -3, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -2, -2, -3, -3, -2, -2, -1, -1, 0, 0, 0, 0, 0, 1, 0, 2, 2, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, -2, -2, -2, -3, -1, 0, 0, 0, 0, 1, 1, 2, 2, 2, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -2, -2, -1, -2, -2, 0, -1, 0, 0, 1, 1, 1, 3, 2, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, -2, 0, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 3, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 1, -1, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, -1, 0, 1, 0, 1, 0, 0, 2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 1, 2, 2, 3, 1, 3, 2, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 1, 2, 2, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 2, 2, 2, 2, 1, 1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, -1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 2, 1, 2, 3, 3, 1, 0, 1, 0, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, -1, 0, 1, 1, 0, 1, 0, 1, 1, 2, 3, 2, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 1, 1, 2, 2, 2, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 2, 2, 1, 1, 2, 2, 2, 0, 0, 1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 0, 1, 2, 2, 2, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 2, 1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 2, 1, 0, 1, 2, 1, 0, 0, 0, 1, 0, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 1, 2, 2, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -2, -2, -1, 0, 0, 0, 0, -1, 0, -2, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, -2, 0, 0, -1, -2, 0, -1, 0, 0, 0, 1, 0, 0, -2, 0, 0, -2, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -2, -1, -1, -1, -2, 1, 0, -1, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 2, 1, 2, 1, 0, 1, 0, -1, -1, -1, -1, -1, 0, 1, 2, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 3, 2, 2, 0, 1, 0, 0, -1, -1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 2, 2, 2, 2, 1, 2, 1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 1, 0, 0, 2, 0, 0, 0, -1, 0, 1, 0, 0, 3, 3, 2, 1, 1, 2, 3, 1, 1, 0, 1, 0, 0, 2, 2, 1, 2, 1, 0, 2, 1, 1, 2, 1, 0, -1, 0, 0, 1, 0, -1, 0, 3, 3, 3, 0, 2, 1, 0, 2, 2, 1, 1, 0, 1, 3, 2, 1, 1, 1, 1, 2, 2, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 3, 1, 1, 1, 1, 0, 1, 2, 1, 1, 1, 1, 3, 2, 1, 1, 2, 2, 4, 2, 2, 2, 0, -2, -1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, 1, 1, 0, 0, 1, 2, 0, 1, 2, 0, 2, 2, 2, 2, 1, 2, -1, -1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 1, 2, 0, -1, 0, 0, 1, 1, 1, 1, 3, 1, 0, 1, 2, 1, 2, 2, 1, 1, 1, -1, -2, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, -1, -1, -2, -2, 0, 0, 0, 1, 2, 2, 1, 1, 2, 2, 2, 2, 0, 1, 2, 0, -1, 0, -1, 0, 1, 3, 0, 0, 0, 0, 0, 0, -2, -1, -3, -2, -1, 0, 0, 1, 2, 2, 0, 0, 1, 1, 2, 1, 0, 0, 1, -1, -2, 0, -2, 0, 0, 2, 0, 0, 0, 0, 1, 0, -2, 0, -2, -1, -2, -2, 0, 0, 1, 3, 1, 1, 2, 1, 3, 0, 1, 0, 1, 0, -1, 0, -1, -2, -1, 0, 0, 0, 0, 1, 1, 0, -2, -2, 0, 0, -2, -2, 0, 0, 1, 1, 1, 0, 0, 1, 3, 1, 2, 0, 0, 0, -1, 0, -1, -3, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -1, 0, -3, -2, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 3, 1, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, 3, 2, 2, 1, 3, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, -2, 0, 1, 0, 0, 0, 1, 0, 1, 2, 1, 0, 1, 2, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, -1, -2, -1, -1, 0, 0, 0, 1, 1, 2, 0, 0, 3, 1, 0, 1, 3, 3, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 4, 2, 1, 3, 3, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 2, 5, 2, 0, 3, 2, 2, 0, -1, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 3, 3, 0, 0, 2, 1, 0, 0, 0, 2, 1, 1, 1, 1, 2, 2, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 2, 2, 2, 1, 2, 2, 0, 1, 1, 0, 1, 0, 0, 2, 1, 2, 1, 0, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 2, 2, 2, 2, 3, 2, 1, 2, 1, 0, 0, 0, 0, 0, 2, 1, 1, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 3, 1, 1, 3, 1, 2, 3, 2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 1, 3, 2, 3, 2, 2, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 1, 2, 2, 1, 0, 0, 0, 0, 1, 1, -1, 0, 0, -2, -1, -1, 0, -1, 0, 1, 0, 0, -1, 1, 0, 0, 2, 0, 0, 1, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -3, -1, 0, -1, 0, 0, 0, 0, -1, 1, 1, 0, 1, 2, 0, 0, 1, 3, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, -1, -2, -3, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, -2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, -2, -1, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 3, 2, 4, 2, 3, 1, 2, 2, 2, 2, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 3, 1, 1, 1, 1, 1, 1, 2, 1, 2, 1, 2, 0, 2, 0, 0, -1, -2, 0, -1, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 1, 2, 2, 1, 2, 3, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 1, 1, 2, 2, 2, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -2, -2, -1, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, -1, 0, 0, 0, -1, 0, -2, -2, -3, -1, -3, -2, -2, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -3, -2, -2, -3, -3, -2, -3, -2, -3, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, -2, -1, -3, -3, -3, -1, -3, -3, -3, -1, -2, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -2, -1, 0, -1, -2, -2, -2, -1, -1, 0, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -2, -3, -3, -1, -1, -1, -1, -1, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, -2, -1, 0, 0, -2, -1, -2, -2, -3, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, -1, -1, -1, -2, -2, 0, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, -1, 0, -1, -1, -2, -2, -3, -1, -1, 0, -2, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 2, 1, 0, 0, -1, 0, -2, -1, -2, -3, -2, -3, -1, -2, -3, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -3, -2, -4, -3, -2, -2, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, -2, -1, -3, -2, -3, -3, -1, -2, -1, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -2, -1, -2, -2, -2, -3, -2, -2, -2, -2, -2, -1, 0, 0, 0, 1, 0, -1, -1, -2, -1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, -1, 0, -1, -2, -1, -2, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -2, -2, -1, -2, -1, 0, -1, 0, 0, 0, -1, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -2, -2, -2, -2, -1, -1, -2, 0, -1, -2, -2, -2, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, -1, -1, -1, -2, -1, -2, 0, -2, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, -2, 0, -1, -2, -2, -1, -2, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 2, 1, 1, 0, 1, 2, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 2, 3, 2, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, -2, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 1, 2, 2, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 1, 0, 1, 2, 2, 1, 2, 0, 1, 2, 1, 1, 0, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, -2, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 1, 0, 1, 0, -1, 0, -1, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -3, -2, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 2, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -2, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 2, 1, 2, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -2, 0, -2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 1, 0, 1, 2, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 2, 2, 2, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, -1, 0, -1, -1, -1, 0, 0, 1, 1, 2, 3, 2, 3, 3, 2, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, -2, 0, 0, 0, 1, 2, 1, 2, 3, 3, 4, 3, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 1, 0, 2, 3, 1, 3, 2, 3, 2, 3, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 1, 0, -1, 0, -1, -1, 0, 0, 0, 2, 2, 2, 2, 2, 3, 2, 1, 1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 2, 2, 3, 2, 2, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 2, 2, 3, 2, 1, 0, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, 0, 0, 1, 0, 0, 2, 2, 2, 1, 2, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 2, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 1, 2, 0, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 2, 0, 1, 0, 0, 0, 1, 1, 0, 1, 2, 2, 2, 0, 1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 2, 0, 0, 1, 1, 2, 1, 2, 1, 3, 4, 2, 2, 1, 2, 1, 1, 2, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 2, 1, 3, 2, 3, 3, 4, 3, 2, 1, 1, 0, 0, 1, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 3, 4, 3, 3, 3, 1, 0, 1, 0, 1, 0, 1, 0, 2, 2, 1, 1, 0, -1, 0, -2, -1, -1, -2, 0, 0, 1, 2, 1, 0, 1, 0, 2, 2, 2, 2, 3, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -2, -1, -4, -2, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 2, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -2, -2, -2, -2, -3, -4, -4, -2, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 2, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -4, -3, -4, -4, -5, -5, -5, -4, -3, -2, -1, 0, 0, -1, -1, 0, 1, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, -1, -1, -1, -3, -4, -4, -4, -4, -5, -4, -4, -4, -3, -3, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -2, -1, 0, -2, -2, -4, -5, -5, -4, -4, -4, -4, -4, -4, -3, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 2, 1, -1, 0, -1, -1, -1, -3, -4, -5, -3, -2, -2, -2, -3, -3, -3, -1, -1, -2, -1, -2, 0, 1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, -3, -3, 0, -1, 0, -1, -1, -1, -2, -2, -3, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, -2, -2, -2, -2, -2, -2, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 2, 1, 1, 3, 2, 1, 2, 3, 2, 1, 1, 0, -1, 0, -1, -2, -3, -3, 0, -1, -1, -3, 0, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 2, 1, 2, 3, 2, 0, 1, 1, 0, -1, -1, -2, -2, -2, -3, -2, -3, -2, -2, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 1, 1, 1, 2, 1, 2, 1, 2, 0, 0, 0, -2, -3, -3, -4, -3, -3, -3, -2, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 0, 1, 1, 1, 2, 1, 1, 1, 2, 1, 1, 1, 0, -1, -2, -3, -2, -3, -3, -1, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 1, 3, 4, 3, 3, 0, -2, -2, -2, -3, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 2, 3, 4, 2, 1, 2, 0, -2, -3, -3, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 0, 1, 0, 3, 2, 3, 3, 4, 2, 0, -1, -3, -4, -4, -3, -2, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 3, 3, 2, 2, 1, 0, -1, -2, -3, -4, -2, -2, 0, 0, -1, 0, 1, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -3, -2, -3, -3, -2, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -2, -2, -1, -1, -1, 0, -1, -1, -2, -1, -3, -4, -3, -3, -1, -3, -1, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -3, -2, -3, -3, -2, -2, -3, -2, -3, -2, 0, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -4, -3, -4, -4, -5, -4, -5, -4, -5, -3, -2, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, -2, -3, -3, -3, -6, -5, -5, -5, -4, -5, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, -1, -3, -3, -3, -5, -5, -4, -3, -4, -2, -2, -1, 0, 0, 0, 1, 1, 1, 2, 3, 2, 3, 0, 1, 2, 1, 1, 2, 1, 0, -1, 0, -1, -2, -3, -3, -3, -3, -3, -2, -2, -2, -1, 0, 0, 1, 0, 0, 1, 2, 2, 3, 2, 2, 1, 0, 1, 0, 1, 1, 0, -1, 0, 0, -1, -1, -1, -1, -1, -1, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 1, 1, 3, 2, 1, 2, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, -1, -2, -1, -1, -1, -1, 1, 1, 1, 3, 3, 3, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 2, 2, 3, 3, 3, 3, 3, 2, 1, 1, 0, -1, -1, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 1, 2, 1, 1, 2, 2, 1, 2, 1, 2, 4, 4, 2, 4, 4, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 1, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, -1, -1, -1, -2, -2, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -2, -2, -2, -2, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, -1, -2, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -2, -1, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, -2, -1, 0, -1, 0, -1, -1, 0, -1, 0, -1, -2, -2, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, -1, -2, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, -1, -1, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, -1, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, 0, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, -1, 0, 1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, -1, -1, -1, -2, -2, -1, -2, -1, -1, 0, 1, -1, -1, -1, 0, -1, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, -2, -2, -3, -2, -1, 0, 0, 0, 1, -1, 0, -1, -1, 0, -1, 0, -1, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, -2, -3, -2, -2, -2, 0, -1, 0, 1, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -3, -2, -3, -1, -2, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -2, -2, -2, -1, -1, -2, -2, 0, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, -1, -1, -1, -2, -1, 0, 0, -1, -1, -2, -2, 0, -1, -2, 0, -2, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, -2, -2, -1, -2, -2, -1, -1, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, -2, -2, -1, -1, 0, -1, -1, 0, -1, 0, 0, -1, -2, -2, -2, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, -2, -1, -1, -2, -2, -1, -2, -1, -2, -2, 0, -1, 0, 0, -1, 0, -1, -1, -2, -1, -1, -1, -1, 0, -2, 0, 0, 0, -1, -1, 0, -2, -1, 0, -1, -3, -2, -2, -2, -2, -1, -1, 0, -1, 0, 0, -1, 0, -2, -2, 0, -1, -2, -2, -2, -2, -1, -2, -2, -1, -1, -1, 0, -2, -1, -1, -2, -2, -1, -1, -3, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -2, 0, -2, 0, -1, -1, -2, -1, -1, -2, 0, -1, 0, 0, 0, -2, -2, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, -1, -1, -1, -2, -2, -1, 0, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, -1, -1, 0, -1, -2, -2, 0, -1, -1, -1, -1, 0, -1, -1, 0, -2, -1, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -1, -1, -2, -1, 0, 0, -1, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, 0, -1, -1, -1, -1, 0, -1, 0, -1, -1, -2, -2, -1, -1, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, -1, -2, -1, -2, -1, 0, -2, 0, -2, -2, -2, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, -2, -1, 0, 0, -1, -2, -1, -1, -1, -1, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -2, -1, -1, -2, -1, -2, -2, -1, -1, -1, 0, -1, 1, 1, 0, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, -1, -1, -1, -2, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -2, -2, 0, 0, 0, 1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 2, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 1, 2, 1, 0, -2, -3, -2, -1, -1, 0, 1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, -1, -2, -2, -1, 0, 1, 1, 1, 0, 0, -1, 0, -1, -2, -2, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -2, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 1, 3, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -2, -3, -1, -3, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -2, -2, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, -2, -1, -2, -2, -2, -2, -2, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -2, -2, -1, -2, -2, -2, -1, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -2, -1, -1, 0, -1, -1, -1, -1, -1, -2, -2, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -2, 0, -1, -1, 0, -1, 0, -1, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, -2, -1, -2, -3, -2, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, -1, 0, -2, -2, -3, -2, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -2, -3, -3, -2, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, -1, 0, -2, -1, -1, 0, 0, 0, 0, -1, -1, -2, 0, -2, -2, -2, -2, -2, 0, -1, -2, -2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, -1, -2, -2, 0, -1, 0, -1, -1, -2, -2, -2, -1, -3, -2, -3, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, 0, -1, 0, 0, -2, 0, -1, -1, -1, -2, -3, -3, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, -1, 0, 0, -1, -1, -1, -1, -3, -2, -3, -3, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -2, -1, -1, -1, -1, -1, -1, -1, 0, -1, -2, 0, 0, 0, -2, -3, -2, -2, -3, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -2, -2, -1, 0, 0, 0, -1, -2, 0, -1, 0, -2, -2, -1, -2, -2, -1, -1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -3, -2, 0, -1, 0, -1, -1, -2, -1, -2, -2, -3, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -2, -1, -1, -1, -2, -2, 0, 0, -2, 0, -2, -1, -2, -2, -2, -2, -2, 0, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, -2, -2, -1, -3, -3, -1, -1, -2, -2, 0, 0, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, -2, -3, -2, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -2, -2, -2, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 0, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 2, 1, 1, 1, 2, 0, -2, -2, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 0, 0, 1, 0, -3, -2, -1, -1, 0, -1, -2, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 3, 1, 0, 1, 0, 0, -1, -2, -2, -1, 0, -1, -1, 0, 0, 0, 1, 0, 1, 1, 2, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 2, 1, 1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 2, 1, 1, 0, 1, 1, 0, 0, 0, -1, -1, -1, -2, -2, -1, -1, -1, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 2, 3, 2, 1, 0, 1, 0, 0, 0, -1, -2, -1, -2, -2, -3, -2, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 2, 2, 2, 1, 0, 0, -1, 0, 0, -1, -2, -3, -2, -2, -3, -2, -2, -1, -1, -1, 0, 0, 0, -1, 0, 1, 1, 2, 1, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -3, -3, -3, -3, -2, -2, 0, 0, 0, -2, -2, -2, 0, 1, 2, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -3, -2, -3, -2, -1, -1, 0, 0, -2, -1, -2, -1, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, -1, -2, 0, -1, -2, -2, -3, -2, -2, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -2, -2, -3, -3, -3, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, -2, -1, -1, -2, -2, -1, -2, -2, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, -1, -2, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -2, -2, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 2, 3, 2, 1, 1, 1, 0, -2, -1, -1, -1, 0, 0, -1, -2, -2, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 2, 1, 3, 3, 3, 5, 5, 3, 4, 3, 1, 0, 0, -1, -2, -2, -1, -2, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 4, 3, 4, 4, 5, 5, 5, 5, 5, 2, 1, 0, -2, -2, -2, -2, -2, -2, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 3, 4, 4, 6, 5, 6, 5, 5, 4, 4, 2, 0, 0, -1, -3, -3, -1, -2, -1, -1, 0, 0, 0, -1, 1, 0, 0, 0, 1, 2, 1, 2, 4, 3, 4, 6, 4, 6, 6, 5, 6, 4, 3, 0, -1, -2, -2, -3, -1, -1, -1, 0, -1, 0, 0, -1, 1, 0, 0, 0, 1, 0, 1, 3, 3, 5, 6, 4, 5, 5, 6, 7, 6, 6, 3, 1, -2, -3, -3, -3, -2, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 3, 2, 3, 5, 5, 4, 5, 5, 5, 6, 6, 5, 3, 0, 0, -3, -3, -1, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 3, 4, 5, 4, 4, 5, 5, 5, 6, 5, 4, 3, 1, -1, -4, -3, -3, -3, -2, -2, -1, -2, 0, 0, 0, 0, -2, 0, 0, 0, 1, 1, 2, 4, 4, 3, 5, 4, 5, 4, 5, 4, 3, 1, 0, -1, -3, -3, -2, -2, -2, -1, 0, -1, 0, 0, 0, -1, -2, -1, 0, 0, 0, 1, 2, 2, 3, 3, 4, 4, 3, 4, 3, 3, 2, 0, -1, -1, -3, -3, -3, -2, -2, -1, -1, -1, 0, 0, 0, -1, -1, -2, 0, 0, 0, 1, 0, 1, 3, 0, 2, 2, 1, 2, 2, 3, 0, 0, -2, -3, -3, -3, -2, -2, -1, 0, 0, -2, 0, 0, 0, 0, -2, -1, 0, 0, -1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -3, -2, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, -1, -3, -2, -2, -2, 0, 0, 0, -1, 0, -2, -1, 0, 0, 0, 0, -2, -1, -2, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -3, -4, -4, -4, -3, -4, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -3, -3, -5, -5, -3, -2, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -4, -5, -5, -3, -2, -1, -1, -1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -3, -4, -4, -3, -2, -1, -2, -1, 0, 0, 1, 2, 1, 1, 2, 1, 0, 0, -1, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -3, -3, -4, -2, -1, -1, -2, 0, 1, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, 1, 1, 2, 1, 1, 2, 1, 0, 0, 0, 0, -1, -3, -2, -3, -2, -1, -2, -1, -2, -1, 0, 0, 1, 1, 2, 1, 0, 0, -1, 0, 0, 2, 1, 0, 0, 1, 2, 2, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -2, -2, -1, 0, 0, 1, 2, 2, 1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -2, -1, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -3, -1, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, -1, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 2, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 1, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, 0, -1, 0, 1, 2, 1, 0, 0, 1, 2, 1, 2, 0, 0, 0, -1, 0, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 1, 2, 0, 1, 0, 1, 2, 2, 1, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 1, 0, 2, 1, 0, 0, 0, 1, 3, 1, 0, 1, 0, 1, 2, 1, 1, -1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 1, 1, 0, 0, 1, 0, 0, 1, 2, 3, 1, 1, 0, 0, 1, 2, 1, 0, 0, 0, -2, 0, 0, 0, 0, 1, 0, 1, 0, -1, 1, 3, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 1, 2, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -2, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 2, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, -2, -1, 0, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, -2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, 0, 0, -1, -1, 0, 0, 1, 1, 1, 2, 1, 0, -1, 0, -1, -2, -2, 0, 1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, -1, 0, 0, 0, -2, -3, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 1, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 1, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, -1, 1, 2, 2, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 1, 1, 1, -1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 2, 2, 1, 1, 2, 1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 1, 3, 1, 1, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 2, 2, 1, 1, 2, 2, 1, 1, 1, 1, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 2, 0, 2, 2, 2, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -2, -3, -2, 1, 1, 0, -1, 0, 0, 0, -2, 0, 0, 0, 0, 1, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 1, 1, 1, 2, 1, 2, 2, 1, 1, 1, 2, 2, 0, 0, 0, 2, 2, 1, 1, 0, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 3, 2, 2, 0, 1, 2, 2, 3, 3, 3, 1, 1, 0, 1, 0, 0, 0, 0, -1, -2, -1, -1, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 1, 2, 3, 3, 4, 3, 2, 1, 0, 0, 1, 1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 3, 2, 2, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 2, 2, 1, 1, 1, 1, 2, 2, 1, 2, 1, 1, 1, 2, 1, 1, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 2, 1, 2, 0, 1, 2, 2, 2, 2, 1, 2, 1, 0, 2, 2, 3, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 1, 0, 0, 0, 1, 1, 2, 3, 1, 2, 1, 0, 0, 1, 1, 2, 1, 1, 1, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -3, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 1, 1, 1, 1, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, -2, -2, 0, 0, -1, -2, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 1, 0, 1, 1, 2, 1, -1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 1, 2, 2, 2, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 2, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 0, 0, 0, 0, -1, 0, 1, 2, 0, 0, 1, 1, 0, -1, 0, -2, -1, -1, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 1, 1, 1, 1, 1, 2, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 4, 4, 2, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, -1, 0, 0, 1, 2, 1, 0, 1, 1, 0, 0, 0, 1, 2, 2, 3, 1, 1, 1, 2, 3, 2, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 3, 1, 1, 0, 1, 2, 0, 0, 0, 2, 2, 2, 3, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 3, 3, 1, 0, 1, 2, 1, 1, 1, 2, 1, 3, 1, 2, 2, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 3, 3, 2, 1, 1, 2, 1, 2, 0, 0, 2, 0, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 2, 1, 0, 0, 0, 1, 0, -1, 0, -2, -1, 0, 1, 2, 0, 1, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 1, 2, 1, 0, 0, 0, -2, -2, -3, -2, -3, -2, 0, 1, 1, 1, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 2, 2, 2, 0, 0, 0, -1, 0, -2, -2, -1, -1, 0, 0, 0, 2, 3, 2, 0, 0, 1, 1, 0, 0, 0, 0, 1, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -2, -1, -1, -2, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, -1, -3, -1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, 0, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -2, -3, -3, -1, 0, -1, 0, -1, -4, -3, -2, -2, -2, -1, -2, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 1, 0, 2, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 2, 2, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -2, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -2, -2, -2, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -1, -2, -1, -2, -1, -1, -1, -1, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, -1, -1, -1, -2, -2, -2, -1, -1, -1, 0, -2, -1, -1, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, -2, -2, -1, -2, -1, -2, -1, -2, -2, -1, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, -2, -2, 0, -1, -1, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -2, -1, 0, -1, -1, 0, -1, -1, -2, -1, 0, -2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, -2, -1, -1, 0, -1, 0, -1, -1, -1, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -2, -2, -2, -2, -1, -1, 0, -2, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -2, -3, -3, -2, -2, -1, -2, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -2, -2, -1, -3, -2, -1, -2, -2, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -2, -1, -1, -1, -2, -1, -2, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, 0, -1, -1, -2, -1, -2, -1, -2, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, -2, -2, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -2, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -2, -1, -2, -1, 0, 0, -1, -1, -2, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -2, -2, -2, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -2, 0, 0, -2, -1, 0, -1, 0, 0, -1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, -2, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 2, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 2, 1, 2, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 2, 1, 0, 1, 1, 0, 2, 4, 3, 2, 2, 0, 0, 0, 0, 0, 0, 0, -2, -1, -3, -4, -2, -2, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 1, 2, 1, 0, 2, 3, 1, 1, 0, 1, 0, 0, 0, -1, -2, -1, -2, -2, -4, -4, -4, -2, -2, -1, 0, -1, 0, 0, 1, 2, 3, 2, 2, 3, 1, 0, 2, 3, 2, 2, 1, 0, 0, -1, -1, -1, -2, -2, -3, -5, -5, -4, -3, -2, -3, 0, 0, 0, -1, 0, 0, 1, 1, 4, 2, 4, 3, 0, 2, 2, 2, 0, 0, 0, 0, 0, 0, -2, -1, -2, -3, -4, -4, -4, -3, -2, -1, 0, -1, -1, -1, 0, 0, 1, 2, 3, 1, 3, 3, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, -2, -2, -3, -3, -4, -3, -2, -2, -1, 0, 0, -1, -2, 0, 0, 0, 1, 2, 2, 2, 2, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -3, -2, -3, -4, -2, -3, -2, -2, -1, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -3, -2, -4, -3, -4, -3, -2, -2, -2, 0, -1, -2, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, -2, -1, -3, -3, -3, -3, -1, -2, -2, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, -1, -1, -2, -1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 1, 1, 0, -1, -1, -1, 0, -1, 0, 1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 1, 0, 2, 3, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 2, 2, 3, 3, 4, 4, 3, 2, 1, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, -1, 1, 0, 0, 0, -2, -2, -1, 0, 0, 2, 2, 2, 4, 5, 6, 6, 6, 5, 3, 2, 1, -1, -1, -2, -2, -1, -2, -1, -2, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 2, 1, 2, 4, 5, 6, 6, 7, 8, 6, 4, 3, 0, 0, -2, -1, -3, -3, -3, -1, -2, -2, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 4, 4, 4, 7, 7, 9, 8, 7, 5, 4, 2, 0, 0, -3, -2, -2, -1, -2, -2, -1, -1, 0, 1, 1, 0, -1, -1, -1, 0, 1, 2, 3, 3, 4, 5, 6, 7, 8, 8, 6, 7, 5, 2, 1, -1, -3, -3, -2, -1, -1, -1, 0, 0, 0, 1, 1, -1, 0, -1, -1, 0, 1, 0, 3, 3, 5, 5, 5, 6, 7, 6, 8, 7, 5, 3, 2, 0, -3, -3, -2, -2, -2, -1, 0, 0, -1, 1, 0, -1, -2, -2, 0, 0, 0, 1, 3, 5, 5, 4, 5, 7, 8, 6, 8, 6, 5, 2, 1, 0, -4, -3, -3, -3, -2, -1, 0, 0, 0, 1, 0, -2, -2, -1, -1, 0, 1, 0, 2, 3, 5, 4, 4, 6, 8, 6, 6, 6, 3, 2, 0, -1, -2, -4, -3, -3, -1, -1, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, 1, 1, 1, 2, 4, 4, 5, 6, 8, 6, 5, 4, 2, 1, -1, -2, -4, -5, -3, -4, -2, -1, 0, 0, 0, 1, -1, -1, -1, -2, -1, 0, 0, 0, 0, 1, 3, 4, 4, 5, 6, 4, 4, 1, 0, -1, -2, -3, -4, -4, -4, -3, -2, -1, -1, 0, 0, 1, 0, -2, -2, -2, -2, -2, 0, 0, 0, 1, 2, 1, 2, 2, 1, 1, 1, 1, 0, -1, -2, -3, -4, -3, -2, -1, -1, -3, 0, 0, 0, 0, 0, -1, -3, -3, -3, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -2, -2, -4, -4, -2, -2, -2, -2, -1, 0, 0, 0, 0, -1, -2, -2, -2, 0, 0, 0, 0, -1, -1, -1, -2, -3, -3, -3, -1, -1, -2, -2, -2, -1, -1, 0, -1, -2, 0, -1, -1, 0, 0, 1, 1, -1, -1, -1, -2, -1, -1, 0, -1, -2, -2, -3, -3, -4, -4, -3, -2, -2, -2, -3, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -3, -4, -5, -4, -2, -1, -2, -1, -1, 0, 0, 1, 2, 0, 0, 0, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -3, -2, -4, -4, -3, -1, -2, -1, 0, 1, 1, 2, 1, 3, 1, 1, 0, 1, 0, 0, 1, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -3, -4, -4, -2, 0, -2, -1, -1, 0, 1, 3, 2, 3, 3, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, -1, -3, -4, -3, -2, 0, -1, -2, -1, 0, 1, 1, 2, 3, 2, 2, 1, 0, 1, 0, 2, 2, 1, 1, 1, 2, 2, 2, 2, 1, 0, -1, -1, -2, -1, -1, -1, 0, -1, 0, 0, 0, 1, 3, 4, 4, 3, 3, 1, 0, 0, 1, 2, 2, 1, 2, 1, 1, 2, 2, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 2, 2, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 2, 1, 1, 1, 0, 1, -1, -2, -1, -2, -2, 0, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -2, -3, -2, -2, -1, 0, -1, -1, -1, -1, -2, 0, -1, -1, -1, 0, -1, -1, -2, -1, -2, -2, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, -2, -1, -2, -1, -1, 0, 0, -1, -1, -2, -1, 0, 0, -1, -1, -1, -1, -2, -1, -3, -2, -2, -2, -1, -2, -1, 0, 0, -1, 0, 0, 0, -2, -2, 0, 0, -1, 0, 0, 0, 0, -2, -2, -1, -1, -1, 0, -1, -1, -2, -1, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -2, -2, -1, -1, -1, 0, -2, 0, 0, -1, -1, -1, 0, -1, -2, -1, -3, -1, -1, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, 0, -1, -2, -2, -1, -1, 0, -1, 0, 0, -1, -2, -2, -2, -2, 0, -1, -1, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, -2, -3, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, -2, 0, -2, 0, -1, 0, 0, -1, 0, -1, 0, 0, 1, -1, -1, 0, -1, -1, -2, -2, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, -2, -2, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, -2, 0, -1, 0, 0, 0, 1, 1, 0, -1, -1, -1, -1, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, -1, -2, 0, -2, 0, 1, 1, 0, -1, -1, 0, -1, -2, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, 0, 0, -1, -1, -2, 0, -2, -1, 1, 1, 0, 0, 0, 0, -2, -2, -2, -1, -1, -1, 0, 0, 1, 0, -1, 0, 0, 0, -2, 0, -1, 0, 0, -1, -1, -2, -1, -1, -1, 0, 1, 1, 1, 0, 0, -1, -2, -2, -2, -2, 0, -1, 0, 0, 1, -1, -2, -1, -1, -1, 0, -2, -2, 0, -1, -1, -1, -1, -2, -3, -2, -1, 0, 0, 0, -1, 0, 0, -2, -3, -2, -1, -2, -2, 0, 0, 0, 0, -2, 0, 0, -1, 0, -2, -1, -2, -2, -2, -2, -2, -2, -3, -2, 0, 0, 0, -1, -1, 0, 0, -3, -3, -3, -3, -1, -2, -1, 0, 1, 0, -2, -1, 0, -1, -1, -1, -1, -2, -2, -1, -1, -2, -1, -1, -2, -1, 0, -1, 0, -2, -1, -3, -3, -2, -2, -2, -2, -1, -2, 0, 0, 0, -1, -1, -2, -2, -2, -1, -2, -1, -2, -2, -2, -2, -1, -1, -2, -1, 0, 0, -2, -2, -2, -2, -2, 0, -2, -2, -1, -2, -2, 0, 1, 0, 0, -1, -2, -1, -2, -1, -2, -2, -3, -2, -1, -1, -1, -2, -2, -2, 0, 0, 0, -2, -1, -1, -1, 0, -2, -2, -1, -2, -2, 0, 1, 0, 0, 0, -3, -2, -2, -1, -1, -2, -2, -2, -1, -2, -1, -1, -2, -1, 0, -2, -1, -1, 0, -2, -2, 0, -2, -3, -2, -1, -1, 0, 0, 0, -1, -1, -2, -1, -2, -1, -3, -3, -1, -2, -2, -3, -1, -1, -2, -2, -1, -1, -2, -1, 0, -2, -2, 0, -1, -2, 0, -2, -2, 0, 0, 0, 0, 0, -2, -2, -1, -1, -2, -1, -1, -2, -2, -3, -3, -1, -1, 0, -2, -1, -2, -1, 0, -2, -1, -2, -3, -2, -2, -1, -2, 1, 0, 0, -1, -1, -1, -2, -1, -2, -2, -1, -2, -1, -2, -2, -2, -1, 0, 0, -1, -2, -1, -1, -1, -3, -1, -1, -1, -1, -2, -2, -2, 1, 0, 0, 1, -1, -1, -1, -1, 0, -2, -1, -2, -1, -1, -2, -3, -1, -1, 0, -1, -1, 0, -1, 0, -2, -2, -1, -1, -1, -1, -2, -2, 1, 0, 0, 1, 0, -3, -1, -1, 0, -1, -1, -1, -1, 0, -2, -3, -2, 0, 0, -1, -2, 0, -1, -2, -1, -1, -1, -2, -2, -1, -1, -1, 2, 0, 0, 0, 0, -2, -2, -1, -1, -2, -1, 0, 0, 0, 0, -1, -1, -2, 0, -1, -1, -1, -1, -1, -2, -4, -2, -3, -1, -2, -2, -1, 1, 0, 0, 0, -1, -1, -1, 0, 0, -2, -2, 0, 0, -1, 0, -1, -1, -1, -2, -2, -3, -2, -1, -2, -2, -4, -3, -2, -3, -2, -3, -1, 2, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, -1, -1, 0, -1, -1, -2, -3, -3, -1, -1, -3, -2, -4, -4, -3, -3, -3, -2, -1, 2, 0, 0, 0, 0, -2, 0, 0, -1, -1, 0, -1, -1, -1, -2, 0, -1, -1, -2, -3, -2, -1, 0, -2, -3, -4, -4, -4, -2, -3, -3, -1, 1, 0, 0, -1, 0, -1, -1, 0, -1, -2, 0, 0, 0, 0, -1, -1, -1, -2, -2, -1, -3, -1, -2, -2, -2, -2, -3, -2, -2, -2, -1, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, -2, -2, 0, 0, 0, 0, -2, -1, -1, -1, -2, -2, -2, -3, -2, -2, -3, -2, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, -1, 0, -1, -2, -2, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -2, -2, -1, -2, -1, -1, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 1, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -3, -1, -1, -1, 0, 0, -1, -2, 0, -2, -1, -1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 2, 1, 0, 1, 0, 2, 1, 1, -1, -3, -2, -2, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 2, 3, 2, 1, -2, -2, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 2, 3, 2, 0, -1, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, -1, -2, -3, -2, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 2, 2, 1, -1, -2, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -3, -2, -2, -3, -2, -2, -1, -2, 0, 0, -1, 0, -1, -1, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, -2, -2, -3, -3, -3, -4, -4, -3, -3, -3, -2, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -2, -2, -3, -3, -3, -3, -3, -3, -2, 0, 0, 0, -1, -1, -1, 1, 1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, -1, -1, -1, -2, -1, -3, -3, -3, -3, -3, -2, -2, -1, 0, 0, -1, 0, 1, 1, 0, -1, -2, 0, 0, -1, -1, 0, -1, -1, 0, -1, -1, -1, -1, -1, -2, 0, -2, -2, -4, -3, -3, -3, -3, -2, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -2, -1, -1, -1, 0, 0, -1, -3, -3, -3, -2, -3, -2, -1, -1, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, 0, 0, 0, 0, -1, 0, -3, -4, -4, -3, -3, -3, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, -3, -3, -4, -3, -3, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -3, -4, -4, -3, -2, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, -2, -1, -2, -3, -3, -3, -2, -1, -1, -1, 0, -1, 0, -1, -2, 0, 0, 0, 0, 1, 0, 0, -1, -2, -1, -2, 0, 0, 0, -1, 0, -1, -2, -1, -1, -2, -3, -2, -2, 0, 0, -1, -2, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, -2, -2, -3, -4, -2, -2, -1, -1, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, -1, -1, 0, 0, 0, -1, 0, -2, -1, -3, -4, -4, -3, -1, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -2, -1, -1, -1, 0, -1, -1, 0, 0, -1, -3, -4, -3, -3, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, -3, -1, -2, -2, -1, -2, 0, -1, -1, 0, 0, -1, -3, -3, -3, -2, -1, -2, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -3, -2, -3, -2, -1, 0, -1, -1, -1, -1, 0, -1, -2, -3, -2, -1, -2, -2, -1, -1, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -2, -1, -2, -3, -1, -1, -1, -1, -2, -3, -1, -3, -2, -1, -1, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, -1, -2, -2, -2, -2, -3, -2, -3, -2, -3, -3, -3, -2, -2, 0, -2, -1, -1, -1, -1, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, -1, -2, -1, -2, -1, -3, -3, -3, -2, -3, -2, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 1, 1, 0, 0, -1, 0, -1, -1, -3, -2, -3, -3, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, -2, -1, -2, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 2, 2, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 3, 3, 2, 3, -2, -1, -1, -2, -1, 0, 1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 3, 2, 3, -2, -3, -3, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 2, 1, -1, -3, -3, -2, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 1, 3, 0, 0, -1, -2, -2, -2, 0, -2, -1, -2, -1, -1, 0, 1, 0, 1, 1, 2, 1, 0, 0, 1, 0, 0, 1, 1, 0, 1, 3, 3, 2, 2, 2, 0, 0, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 2, 2, 1, 2, 1, 0, 2, 2, 2, 0, 0, 0, 0, -1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -2, -2, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, -1, -2, -2, -1, 0, 0, 0, 1, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 1, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, -1, -2, -2, 0, -1, -2, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -2, -1, -1, -2, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 1, 2, 1, 2, 1, 1, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 5, 2, 3, 2, 2, 2, 2, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -2, -1, -1, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 2, 4, 2, 1, 2, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -3, -2, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, -3, -3, -3, -4, -3, -2, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, -1, -1, 0, 0, 0, 0, -1, -1, -2, -3, -4, -3, -2, -1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, -1, 1, 1, 0, 0, 0, 0, -2, -3, -2, -1, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 1, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 2, 1, 0, 1, 3, 0, -1, -2, -1, -1, -1, 0, -2, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 0, -1, -1, -2, -1, -2, -1, 0, -1, -1, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, -2, 0, 1, 1, 0, -1, -1, 0, 0, 0, -2, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, -1, -3, -3, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, -1, -1, -1, -1, 0, 0, 0, -1, -2, -2, -2, -2, 0, 2, 0, 0, 0, 1, 0, 0, 1, 2, 3, 3, 2, 3, 3, 3, 2, 0, 1, 0, -1, -1, -1, -1, 0, -1, -1, -2, -2, -1, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 6, 6, 5, 5, 5, 3, 2, 2, 2, 1, 0, -1, -1, -1, -2, -2, -3, -2, -1, -2, -3, -1, 0, 1, 0, 0, 0, 0, 0, 2, 3, 6, 7, 9, 8, 8, 7, 6, 4, 3, 2, 2, 1, 0, -1, -2, -1, -3, -1, -1, -2, -2, -3, -1, 0, 0, 1, 0, 0, 0, 0, 2, 3, 6, 7, 8, 10, 9, 8, 6, 6, 5, 4, 4, 3, 0, -1, -1, -2, -3, -2, -1, -1, -1, -2, -1, 0, 0, 0, 0, 1, 0, 1, 3, 5, 6, 7, 7, 8, 8, 6, 6, 4, 5, 6, 5, 4, 0, -2, -2, -1, -3, -1, -2, -2, -1, -2, 0, 0, -1, 0, 0, 0, 1, 2, 4, 5, 8, 8, 8, 9, 8, 6, 5, 4, 5, 6, 5, 2, 0, -3, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 3, 5, 7, 8, 7, 9, 8, 5, 5, 4, 5, 4, 4, 3, 0, -2, -1, -1, 0, 1, 0, -1, 0, -1, 0, 1, -1, -1, 0, -1, 1, 2, 3, 6, 6, 8, 7, 7, 6, 4, 4, 5, 4, 3, 4, 2, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 2, 4, 5, 7, 7, 8, 6, 6, 5, 4, 5, 4, 3, 3, 2, 0, -1, 0, -1, 0, 0, 0, 1, -1, -1, 0, 0, 0, -1, -1, 0, 1, 2, 3, 3, 5, 6, 7, 6, 5, 5, 3, 3, 3, 0, 1, 1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 2, 1, 2, 2, 2, 6, 4, 3, 3, 3, 2, 2, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, -2, -1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 2, 2, 3, 0, 0, 0, 0, 0, -2, -2, -2, -1, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, -1, -1, -2, -2, -2, -4, -4, -2, 0, 0, 0, -1, 0, -1, -2, -1, -1, -2, -2, -3, -2, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -2, -2, -2, -3, -4, -4, -4, -3, -2, 0, 0, -1, -1, 0, 0, -1, -2, -1, 0, -1, -1, -2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -4, -4, -5, -5, -6, -4, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 1, 1, 2, 0, 0, 1, 0, 1, 0, 0, 0, -1, -3, -4, -5, -6, -6, -4, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -2, -2, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, -1, -2, -4, -3, -4, -5, -3, -2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 1, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -4, -3, -4, -3, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, -3, -2, -4, -3, -2, -2, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 2, 3, 2, 0, 0, 0, 0, 0, 0, 0, -2, -2, -3, -2, -1, -1, -1, -2, -3, -2, -2, -1, -1, -1, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, -1, -2, -1, -1, -1, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, -1, -1, 0, 0, 0, -2, 0, -1, 0, -1, -1, 0, -1, -1, -1, 0, 0, 1, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, -1, -1, 1, 0, 0, 3, 1, 1, 1, 1, 0, 2, 1, 1, 1, 1, 0, 0, 0, 0, 2, 2, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, 2, 0, 0, 0, 0, 0, 0, -1, -1, 1, 2, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -2, -1, -2, -1, 0, 0, -1, -1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 2, 0, 0, 0, 1, 0, 0, 2, -1, -1, -1, -1, 0, 0, 0, -2, -2, 0, 0, -1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 2, 0, -1, 0, 0, 0, 0, -2, -1, 0, 0, -1, 0, 0, 2, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 2, 0, 0, 0, 1, 1, 0, -2, -2, 0, 0, 0, -1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 1, 1, 0, 0, 2, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, -1, -2, -2, -1, -2, -3, -2, -1, 0, 0, 0, 0, 2, 3, 0, -1, -2, 0, 0, 0, 2, 2, 1, 2, 3, 3, 2, 2, 2, 1, 0, -1, -3, -3, -2, -3, -4, -4, -3, -3, -1, 0, 1, 1, 2, 4, 1, 0, -1, 0, 0, 0, 2, 0, 1, 2, 3, 2, 3, 3, 1, 2, 1, 0, -3, -5, -3, -4, -6, -6, -5, -5, -2, -2, 0, 1, 3, 2, 3, 0, 0, 0, 0, 0, 1, 3, 3, 4, 3, 2, 3, 3, 2, 3, 2, 0, -2, -2, -4, -5, -6, -6, -6, -4, -4, -2, 0, 1, 1, 2, 4, 3, 0, -1, 0, 0, 1, 2, 3, 4, 3, 2, 3, 2, 3, 1, 0, 0, -1, -2, -3, -3, -4, -5, -6, -4, -4, -1, 0, 0, 1, 3, 5, 5, 2, 0, 0, -1, 0, 0, 2, 2, 4, 3, 3, 1, 2, 1, 0, -1, -2, -3, -5, -5, -3, -4, -4, -4, -3, -1, 1, 1, 1, 2, 3, 3, 1, 0, -1, -1, 0, 0, 1, 3, 4, 3, 2, 0, 1, 0, 0, 0, -2, -3, -3, -4, -4, -5, -5, -2, -1, 0, 2, 3, 1, 2, 2, 2, 1, 0, 0, 0, 0, 1, 2, 3, 3, 2, 1, 0, 0, -1, 0, 0, 0, -2, -3, -5, -4, -4, -3, -1, 0, 0, 2, 2, 1, 3, 3, 3, 1, 2, 0, 0, 0, 0, 1, 2, 3, 2, 1, 0, 0, 0, -1, 0, -1, -2, -2, -4, -4, -3, 0, 1, 1, 1, 3, 3, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 2, 3, 3, 2, 0, 1, 0, 1, -1, -1, -1, 0, -2, -3, -2, -1, 1, 0, 2, 2, 2, 3, 2, 0, 0, 1, 0, 1, 0, 0, 2, 1, 2, 3, 4, 2, 0, 0, 2, 0, 0, -1, -1, 0, 0, -2, -4, 0, 1, 1, 2, 4, 2, 3, 1, 0, -1, 1, 1, 1, 0, 0, 3, 3, 4, 4, 4, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, -2, -2, 0, 2, 3, 0, 3, 2, 3, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -2, 0, 2, 2, 1, 2, 2, 1, -1, -1, -1, 0, 0, 0, -1, -1, 1, 0, 0, 1, 3, 4, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 2, 2, 0, 1, 0, 0, -2, -3, -2, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, 4, 2, 0, 1, 0, 1, 2, 2, 0, -2, -1, 0, 2, 3, 1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 2, 2, 3, 2, 1, 0, 0, 0, 0, 0, -1, 0, 1, 3, 2, 1, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 2, 2, 2, 2, 1, 2, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 3, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 3, 1, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, 2, 0, 0, 1, 1, 1, 1, 2, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, -3, -2, -1, 0, 1, 1, 1, 0, 0, 0, 2, 2, 1, 0, 0, 0, 0, 0, -1, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, -2, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, -2, 0, 0, -1, -2, -1, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, -2, -1, -2, -1, -2, -2, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, -3, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -3, -1, -2, -3, 0, 0, -1, -3, -1, 0, -1, 0, -2, 0, 0, -3, -3, -2, 0, 0, 0, 1, 0, 1, 1, 1, 0, -1, 1, 0, -1, -1, -2, -2, -2, -1, 2, 0, 0, -2, -2, 0, -1, 0, -2, 0, -2, -1, -1, -2, 0, 0, 0, 0, 1, 1, 1, 2, 1, -1, 1, 0, 0, -1, 0, -2, -1, -1, 2, 1, -1, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, -2, 0, 0, 0, 0, 1, 4, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, -1, 0, 0, -2, 0, -1, 0, -1, 1, 2, 0, 0, 3, 5, 3, 0, 2, 1, 0, -1, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 3, -1, 0, 0, -1, 0, -1, 0, 0, 3, 1, 1, 0, 1, 3, 3, 3, 4, 3, 3, 0, 3, 3, 1, 1, 0, 1, 1, 1, 2, 0, 0, 3, -1, -1, 0, -1, 0, -1, -1, 0, 1, 1, 0, 1, 1, 2, 2, 2, 2, 3, 3, 2, 3, 4, 0, 1, 1, 1, 1, 2, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 3, 2, 0, 0, 3, 3, 1, 2, 2, 4, 4, 2, 0, 2, 0, 0, 3, 2, 0, 0, 1, -2, 0, 1, 0, 1, 0, -1, -1, 0, -1, 0, 3, 2, 0, 0, 1, 1, 1, 2, 4, 3, 3, 1, 0, 2, 0, 0, 3, 1, 0, 0, 2, -2, 0, 0, 1, 2, 0, 0, 0, 0, -1, 1, 3, 1, 0, 0, -1, 0, 1, 1, 3, 3, 2, 2, 1, 1, 1, 1, 1, 2, 1, 1, 2, -1, 0, 0, 0, 0, 2, 2, -1, -1, -1, 0, 1, 0, -1, -1, -3, -1, 0, 0, 3, 3, 3, 3, 1, 0, 0, 1, 0, 2, 0, 0, 3, -1, 0, 0, -1, 0, 1, 2, 0, 0, 0, 0, 1, 0, -2, -1, -3, -3, -2, 0, 0, 3, 2, 4, 1, 0, 1, 1, 0, 1, 1, -1, 0, -1, 1, -1, -3, -1, 0, 0, 0, 0, 0, 1, 0, 0, -2, 0, -1, -4, -2, -1, 0, 0, 0, 1, 0, 0, 0, 2, 0, 1, 0, -1, -1, -1, 0, 0, -3, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -3, -1, -1, -3, 0, 0, -2, 0, 2, 1, 0, 2, 3, 1, 0, 1, 0, -1, -1, 0, 0, -1, -3, -1, -1, 0, 0, -1, 0, 0, -1, -2, -3, -1, -1, -2, 0, 0, 0, 0, 1, 0, -1, 2, 3, 2, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 1, 0, 0, 0, -2, 0, -1, -3, 0, 0, 0, 0, 0, 2, 0, 1, 3, 1, 0, 2, 0, 0, 0, 0, 0, 0, 1, -2, 0, -1, -1, 0, 0, 0, 1, 0, -4, -2, 0, -2, 0, 0, 0, -1, 2, 0, 0, 2, 5, 0, 0, 2, 0, 2, 2, 0, 0, 0, 1, -1, -3, -2, -1, 0, 2, 0, 2, 1, -2, -1, 0, -2, 0, 0, 0, 0, 1, 1, 0, 2, 4, 0, 0, 3, 0, 3, 0, 0, 0, 1, 0, -1, -2, 0, 0, 0, 1, 1, 2, 1, -1, -2, 0, 1, 0, -1, 0, 0, 1, 0, -1, 2, 4, -1, 0, 2, 1, 2, 0, 0, 0, 1, 1, -1, 0, 1, 2, 3, 1, 2, 2, 1, -2, -1, 0, 0, 0, -1, -1, 1, 1, 0, 0, 3, 4, -1, 0, 1, 1, 2, -1, 0, 1, 0, 0, -1, -1, 2, 4, 2, 2, 2, 3, 2, -1, -1, 0, 0, 0, 0, 0, 2, 0, 1, 1, 3, 3, 0, 0, 0, -1, 0, 0, 0, 1, 1, -1, -2, 0, 0, 4, 3, 2, 3, 3, 2, 1, 0, 0, 0, 0, 0, 0, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, 1, 3, 1, 1, 2, 2, 3, 2, 1, 2, 0, 0, 0, 0, 3, 1, 0, 0, -1, 0, 0, -1, 0, -1, 1, 2, 0, 0, 0, 0, 0, 0, 1, 4, 1, 1, 1, 3, 1, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, 1, 0, 0, 1, 1, 2, 2, 0, 1, 1, 0, 1, 1, 1, 0, 0, -1, 0, 1, 0, 0, -1, -1, -1, -2, -2, -3, -3, 1, 2, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 1, 0, -2, -1, -2, -3, -3, -2, -1, -2, 2, 1, 0, -1, -1, 2, 0, 0, 1, 0, 1, 0, 1, 1, 0, -1, -1, 0, 0, 1, -2, 0, 0, -2, -1, 0, -2, -3, -2, -1, 0, -2, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -2, -3, -2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -1, 0, -1, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 1, 1, 0, 0, -1, -1, -2, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 2, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, -2, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 2, 1, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, -2, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, -1, 0, -1, -2, -2, -2, -2, -2, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -1, 0, 0, 0, -1, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -2, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, 0, -1, -1, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, -1, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -2, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, -2, -1, -2, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -1, 0, -1, 0, 0, -1, 0, -2, -1, -1, -2, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, -1, 0, -1, -2, -2, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -2, 0, 0, -1, -2, -2, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 2, 0, -2, -2, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 1, 1, 1, 1, 1, 1, 2, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -3, -2, -2, -2, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, -2, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, -1, -2, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -2, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -2, -2, -1, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 1, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, -2, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, -2, -2, -1, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, -1, -2, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -3, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, -2, -2, -2, -2, -2, 0, -2, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, -1, -2, -1, 0, -1, 0, -1, 0, -1, 0, -1, -1, -2, -3, -1, -1, -1, -2, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, -2, -1, -2, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, -2, -2, -1, -1, -2, -3, -2, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -2, -1, -1, -2, -1, -1, 0, -2, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, -2, -1, -1, -2, 0, 0, 0, 0, -1, -2, -1, 0, -2, -2, -2, -1, -2, -1, -1, -1, -1, -2, 0, 0, -1, -1, 0, -1, -1, -1, -2, -1, -2, -1, -2, -1, 0, 0, -1, 0, -1, -1, -2, -2, -1, -2, -1, -1, -2, -1, 0, -1, -1, -2, -1, 0, -1, 0, -1, -1, -3, -3, -1, -2, -1, -1, 0, 0, 0, 0, -1, -1, -2, 0, -1, -2, -1, -1, -1, -2, -1, 0, -2, -1, -1, -1, -2, 0, -2, 0, -1, -2, -2, -1, 0, -2, -1, -2, -2, -2, 0, 0, 0, 0, 0, -2, -1, -2, -1, -1, -1, -2, -1, -1, -2, 0, -2, -1, -1, -1, -2, -1, -1, -1, -1, -3, -3, -1, -3, -1, -1, -1, 0, 0, -1, -1, 0, -1, 0, -1, -1, -2, -1, -2, -1, -1, -2, -1, -2, -1, -1, -1, -2, -2, -1, 0, -1, -1, -1, -2, -3, -2, -2, -2, 0, 0, -2, 0, 0, -1, -1, 0, -1, -1, -1, -2, -1, -1, -1, -3, -1, 0, 0, -2, -2, -2, -2, 0, -1, -1, -2, -3, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -2, -2, -3, -2, -2, -1, -1, -1, -1, -1, 0, 0, -2, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, -2, -1, -2, -2, -1, -1, 0, -1, 0, -1, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, -2, -1, -1, -1, -1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, -1, 0, -1, -1, -1, -2, -2, -2, 0, 0, -1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -2, 0, -1, -1, 0, 0, -2, 0, -2, -1, -1, -1, -2, -2, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, -2, -1, -1, -1, -1, 0, -1, 0, 0, -2, -1, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, -1, -1, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 2, 2, 2, 2, 0, 2, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -2, -2, -2, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 3, 3, 3, 2, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -2, -3, -1, -1, 0, 0, 0, 1, 1, 1, 2, 3, 3, 4, 4, 3, 1, 1, 1, 1, 2, 2, 0, 1, 0, 0, 0, 0, -1, -1, -1, -2, -3, -2, -1, -2, -2, 0, 0, 0, 0, 0, 1, 2, 2, 3, 3, 2, 1, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, -1, -1, -2, -3, -3, -3, -3, -2, -1, -2, 0, -1, 0, 0, 1, 1, 2, 3, 4, 3, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, -1, -2, -3, -4, -4, -4, -4, -4, -3, -3, -1, -2, 0, -1, 0, 1, 1, 2, 2, 2, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -3, -4, -5, -5, -4, -5, -5, -4, -4, -2, -2, 0, 0, 0, 1, 1, 2, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -3, -4, -3, -3, -5, -4, -4, -4, -4, -3, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -2, -3, -3, -4, -3, -3, -2, -2, -3, -3, -3, -2, -2, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, -1, -2, -2, -2, -2, -3, -1, -1, 0, -1, -2, -2, -2, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, -2, -3, -1, -2, -1, -1, 0, 1, 0, 0, 1, -1, 1, 0, 0, 0, -1, -1, -1, -1, 0, -2, 0, 0, 0, 0, 1, 2, 3, 2, 0, -1, -1, -1, -2, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 2, 2, 4, 3, 1, 0, 0, -1, -1, -1, -3, -3, -1, -1, 0, 0, 0, 0, 2, 1, -1, 0, -1, -1, -1, -1, -2, -2, 0, -1, 0, 1, 2, 3, 3, 4, 1, 2, 0, 0, -2, -3, -3, -2, -2, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, -2, 0, 0, 1, 2, 2, 4, 5, 3, 2, 3, 1, 1, -1, -2, -3, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, -2, -1, -1, -1, -2, -1, 0, 1, 0, 2, 1, 3, 3, 3, 2, 3, 3, 1, 1, 0, -2, -3, -2, -1, 0, 0, 0, 0, 0, 1, 0, -2, -1, -1, -1, -3, -2, -1, -1, 0, 0, 2, 3, 2, 3, 4, 3, 3, 1, 2, 0, 0, -2, -2, -2, -1, 0, 0, 0, 0, 1, 1, 0, 0, -2, -2, -1, -3, -3, -2, 0, 0, 1, 0, 3, 3, 4, 4, 5, 4, 3, 1, 0, 0, -3, -4, -2, -3, -1, 0, 1, 1, 1, 1, 0, 0, -1, -1, -1, -2, -1, -2, -2, 0, 0, 1, 2, 3, 3, 4, 4, 4, 3, 1, 0, -2, -3, -4, -3, -2, -2, 0, 1, 0, 0, 1, 0, 0, -2, 0, -1, -1, -1, -3, -1, 0, 0, 1, 2, 2, 3, 2, 2, 1, 0, 0, -1, -1, -3, -3, -2, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -2, -2, 0, 0, -1, -2, -2, 0, 0, 1, 1, 2, 0, 0, 0, -1, 0, -1, -1, -2, -3, -2, -1, 0, -1, -1, -1, 0, 1, 0, -2, -1, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, -1, 0, -1, -2, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, -1, -2, -1, -1, -2, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, -2, -2, -4, -3, -2, -2, -1, -1, 0, 0, 1, 0, 1, 0, 0, 1, 2, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -2, -2, -2, -1, -1, -1, 0, 0, 1, 0, 2, 2, 0, 1, 1, 2, 2, 2, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -2, -2, -2, -1, -2, 0, 0, 1, 1, 1, 2, 1, 1, 1, 1, 2, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -2, 0, 0, -2, 0, 0, 0, 1, 2, 1, 2, 2, 2, 1, 2, 1, 2, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 1, 3, 2, 3, 3, 4, 3, 1, 2, 2, 0, 0, 0, 0, 2, 0, 3, 1, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 4, 4, 4, 4, 4, 3, 3, 1, 2, 1, 0, 1, 2, 1, 3, 2, 2, 2, 3, 3, 1, 2, 1, 1, 0, 0, 2, 2, 1, 2, 1, 1, 2, 3, 4, 3, 5, 3, 3, 2, 2, 0, 1, 0, 1, 0, 2, 2, 2, 2, 0, 1, 0, 1, 1, 0, 0, 1, 1, 1, 1, 1, 0, 2, 1, 2, 2, 0, 1, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 2, 2, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 1, 2, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 2, 3, 2, 2, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 2, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 2, 2, 1, 3, 3, 4, 2, 0, 0, 1, -1, 0, 0, 1, 0, 1, 2, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 3, 2, 2, 3, 3, 3, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 2, 1, 0, 0, 0, 1, 0, 1, 1, 2, 1, 2, 2, 3, 3, 2, 2, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 2, 2, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 0, 1, 2, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 2, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 1, 1, 2, 1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 2, 1, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 1, 1, 1, 0, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -2, 0, 1, 1, 0, 0, 1, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, -1, 0, -1, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, -2, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, -1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, -2, -1, -2, -1, 0, -1, -1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -2, -2, -1, 0, -2, -1, -2, -2, 0, 0, 0, -1, 0, 0, 2, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -2, -2, -2, -2, -2, 0, 0, -1, -1, 0, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, 0, -1, -2, -1, 0, 0, -1, -2, 0, 0, 0, 0, 2, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, 0, -2, -2, 0, -1, -1, 0, 0, 0, 3, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 1, 0, 0, -3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, -1, 0, -1, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 2, 1, 1, 2, 2, 2, 1, 2, 2, 1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 1, 0, 1, 0, 1, 1, 2, 1, 2, 1, 2, 2, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 1, 0, 1, 0, 1, 0, 2, 1, 1, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, 0, -1, 0, 0, -1, -1, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -3, -2, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 2, 0, -1, 0, 0, 2, 1, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, -1, -1, -2, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -2, -3, -3, -1, 0, -2, 0, -1, -1, 0, 2, 1, 0, 1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -2, -3, -3, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 1, 3, 1, 1, 0, 0, 0, -1, 0, 1, 0, 1, 1, 0, -1, -2, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 1, 2, 3, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -2, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 1, 2, 1, 2, 2, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, -1, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, 0, 0, 2, 1, 1, 1, 1, 1, 0, 0, 2, 2, 3, 2, 1, 0, 0, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -2, 1, 2, 1, 1, 0, 0, 0, 0, 2, 2, 2, 4, 3, 0, 0, 0, -2, -3, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 1, 0, -1, 0, 1, 1, 1, 2, 2, 1, 0, 0, -1, -2, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 1, 0, -1, -2, -4, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, -4, -3, -2, -1, -1, 1, 0, 0, 0, 2, 1, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 2, 1, 2, 1, 0, 0, -2, -3, -2, -2, 0, -1, 1, 0, 0, 0, 1, 2, 1, 2, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 0, -1, -2, -1, -2, -1, 0, 1, 0, 0, 0, 1, 1, 1, 0, 2, 0, 0, 0, 1, 0, 2, 1, 2, 2, 2, 1, 1, 1, 1, 1, 0, 0, 0, -2, -1, -1, -1, -1, -1, 0, 0, 2, 2, 2, 2, 1, 2, 0, 0, 0, 0, 2, 3, 2, 2, 3, 2, 1, 1, 0, 0, 1, 0, 0, -1, -2, -3, -1, -1, -2, -1, -1, 0, 3, 3, 2, 2, 1, 1, 2, 0, 0, 0, 2, 2, 2, 1, 3, 2, 0, 1, 0, 0, 0, -1, -1, -2, -1, -3, -2, -3, -2, -1, 0, 0, 2, 2, 2, 2, 1, 1, 1, 0, 0, 0, 0, 2, 2, 2, 1, 2, 1, 0, 0, -1, -1, -2, -2, -2, -2, -3, -4, -3, -3, 0, 0, 1, 1, 1, 2, 0, 1, 0, 1, 0, 0, 0, 0, 1, 2, 1, 2, 3, 1, 0, 0, 1, 0, -1, -2, -2, -2, -2, -2, -2, -2, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 2, 1, 2, 3, 2, 0, 0, -1, -1, -1, -2, -2, -2, -3, -3, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 2, 1, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 2, 2, 1, 0, 1, 2, 3, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 3, 2, 2, 2, 0, 1, 3, 2, 3, 1, 1, 0, 1, 1, 1, 0, 1, 1, 0, 0, -1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 2, 1, 3, 2, 2, 0, 1, 3, 2, 1, 0, 0, 2, 0, 0, 0, 2, 0, 2, 1, 0, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 2, 2, 3, 2, 2, 0, 1, 2, 3, 1, 1, 1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 1, 0, 0, 0, 2, 2, 2, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 2, 1, 1, 1, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -2, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -2, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -2, -1, -2, -2, -2, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -2, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -1, -1, -2, -1, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, -1, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 3, 2, 3, 2, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 2, 2, 3, 2, 3, 1, 2, 1, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 2, 1, 1, 2, 2, 2, 1, 2, 1, 0, 0, -1, -1, 0, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 2, 2, 1, 2, 3, 1, 2, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 2, 2, 1, 2, 1, 2, 2, 1, 2, 1, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 2, 3, 2, 3, 2, 3, 2, 1, -1, -1, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 2, 2, 3, 2, 2, 1, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 2, 1, 2, 1, 2, 1, 0, 1, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, -1, 0, 1, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 2, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 2, 2, 2, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 2, 2, 1, 1, 2, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 2, 2, 2, 1, 1, 0, 0, 0, 1, 0, 5, 5, 2, 3, 2, 2, 3, 2, 0, -1, 0, 0, -2, -2, -4, -5, -3, -3, -3, -3, -3, -2, -1, -2, -3, -2, 0, -1, 0, 0, 0, 1, 7, 6, 4, 3, 2, 1, 2, 2, 1, 0, -1, -3, -3, -5, -7, -8, -7, -6, -6, -6, -4, -3, -3, -3, -2, -1, -2, -2, -1, 1, 0, 0, 4, 5, 4, 2, 0, 0, 0, 0, 0, -2, -3, -4, -5, -7, -10, -8, -6, -5, -5, -5, -4, -2, -3, -2, -1, 0, 0, 0, 0, 1, 2, 1, 3, 3, 2, 0, -1, -3, -2, 0, -1, -1, -4, -5, -6, -9, -9, -8, -3, -2, -1, -2, -2, -1, -2, -1, -1, 0, 1, 1, 1, 2, 2, 2, 2, 3, 0, -1, -2, -3, -1, 0, -2, -1, -2, -5, -5, -6, -6, -4, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 2, 2, 2, 3, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -4, -3, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 1, 1, 1, 2, 3, 3, 1, 2, 4, 3, 1, -1, -2, 0, 0, 1, -1, 0, 2, 2, 4, 3, 1, 1, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 1, 3, 1, 0, 0, 4, 4, 2, 0, -1, 0, 1, 2, 1, 0, 3, 2, 3, 3, 2, 2, 0, 0, 0, 2, 1, 0, -1, -1, -1, 0, 2, 2, 2, 0, -1, 0, 3, 3, 0, 0, -2, 1, 1, 2, 4, 5, 3, 4, 2, 3, 2, 0, 0, -1, 0, 2, 2, 0, -2, -4, -2, 0, 1, 2, 1, -1, -4, -2, 0, 1, 0, -1, 1, 2, 2, 4, 7, 7, 5, 4, 4, 4, 1, 1, 0, -1, 0, 0, 1, 0, -3, -4, -5, -1, 1, 1, 0, -1, -1, -1, 1, 0, 0, 1, 4, 5, 6, 6, 7, 6, 5, 5, 4, 2, 2, 0, 0, 0, 1, 0, 0, -2, -2, -4, -4, -3, 0, 0, 0, -1, 0, 0, 0, 0, 1, 3, 7, 10, 9, 9, 9, 9, 6, 4, 4, 3, 2, -1, -2, -1, 0, 0, -2, 0, 0, -2, -4, -2, 0, 0, 1, 1, 0, 0, 0, 2, 3, 7, 11, 12, 12, 12, 11, 10, 7, 5, 5, 5, 3, 0, -1, -1, -2, -3, -2, -1, 0, 0, -2, -3, -1, 0, 0, 0, 2, 0, 1, 3, 6, 10, 13, 14, 16, 15, 14, 12, 8, 7, 8, 8, 5, 2, 0, -1, -3, -4, -1, 0, 2, 1, -2, -2, 0, 0, 0, 0, 2, 2, 2, 4, 6, 10, 13, 13, 15, 17, 16, 14, 11, 10, 11, 10, 7, 1, 0, -2, -2, -1, -1, 0, 4, 4, 1, -2, 0, 1, 0, 1, 1, 3, 4, 5, 7, 11, 14, 14, 14, 15, 16, 12, 9, 9, 12, 10, 6, 1, -1, -4, -3, 0, 0, 2, 2, 4, 2, 0, 1, 0, -1, 0, 0, 3, 4, 6, 8, 12, 15, 14, 13, 13, 14, 10, 8, 10, 12, 10, 5, 1, -2, -4, -2, 1, 3, 1, 2, 3, 2, 2, 1, 1, -2, -3, 0, 2, 2, 5, 8, 12, 14, 14, 12, 13, 12, 9, 9, 9, 9, 8, 4, 2, 0, -2, -2, 1, 4, 2, 1, 3, 2, 3, 3, 0, -3, -4, 0, 0, 3, 6, 7, 11, 13, 13, 13, 11, 10, 9, 8, 8, 8, 6, 4, 3, 1, 0, 0, 1, 4, 3, 2, 2, 0, 0, 1, 1, -2, -4, -1, 2, 3, 5, 5, 9, 11, 12, 12, 10, 7, 9, 7, 7, 6, 6, 4, 4, 2, 1, 2, 2, 1, 1, 1, 2, 0, -1, 0, 0, -1, -2, 0, 3, 5, 4, 3, 6, 9, 12, 12, 7, 5, 6, 8, 5, 4, 2, 5, 3, 1, 3, 4, 1, 0, 0, 0, 0, 0, -2, 0, 1, 0, -1, 0, 2, 3, 3, 1, 3, 8, 10, 9, 6, 3, 3, 4, 4, 0, 0, 1, 2, 0, 2, 4, 2, 0, -1, 0, 0, -3, -3, -1, 0, 0, 0, 0, 0, 2, 2, 0, 1, 4, 8, 6, 3, 0, 1, 2, 1, -2, -1, 1, 2, 0, 1, 3, 2, 0, 0, -1, -3, -1, -2, -3, 0, 0, 1, 0, -1, 1, 0, 0, 1, 3, 4, 2, 0, -1, -1, -1, -2, -3, -3, 1, 3, 1, 1, 0, 0, -2, -3, -2, -1, -2, -3, -2, 0, 0, 1, 0, -1, -1, 1, 2, 0, 0, 0, 0, -1, -2, -4, -6, -6, -7, -3, 0, 3, 1, 0, 0, 0, -2, -1, -2, 0, -1, -4, -3, -1, 2, 0, -1, -1, 0, 1, 3, 1, 0, 0, 0, -3, -5, -7, -7, -7, -7, -2, 1, 1, 1, 0, 0, 0, 0, 2, 1, 1, -2, -4, -2, -1, 2, 1, 0, -1, -1, 2, 3, 2, 0, 0, 0, -4, -6, -7, -8, -8, -6, -3, 0, 1, 0, 1, 1, 2, 2, 4, 2, 2, -1, -2, -3, 0, 3, 2, 0, -2, 0, 1, 3, 1, 0, 0, -1, -5, -6, -7, -9, -7, -6, -2, 0, 0, 0, 0, 1, 2, 2, 2, 1, 1, 0, -1, -2, -1, 4, 3, 0, -1, -1, 0, 0, 0, 0, -1, -2, -6, -8, -8, -7, -7, -5, -2, -1, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, -2, -3, -1, 4, 3, 0, 0, 0, 0, -1, 0, -1, -2, -4, -7, -8, -7, -7, -6, -6, -4, -3, -2, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -2, -1, 4, 4, 2, 1, 1, 0, 0, 0, -1, -3, -4, -5, -8, -7, -6, -6, -5, -4, -4, -3, -1, -1, 0, 0, 0, 1, -2, -3, 0, 2, 0, 0, 2, 2, 3, 1, 1, 0, 0, 0, 0, -2, -2, -3, -4, -4, -3, -3, -2, -3, -3, -2, 0, 0, 0, 0, 0, 1, 0, -2, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 2, 2, 2, 3, 2, 3, 3, 3, 3, 1, 3, 1, 2, 0, 1, 1, 2, 1, 1, 0, -2, -2, 0, 0, -1, 0, 0, -2, -1, -1, -1, 0, 0, 2, 2, 2, 2, 3, 2, 2, 1, 3, 3, 3, 2, 1, 3, 3, 3, 3, 1, -1, -3, -3, 0, 0, 1, 2, 1, 0, 0, 0, 0, -1, 0, 2, 4, 2, 2, 2, 3, 3, 2, 2, 2, 3, 2, 3, 3, 4, 4, 2, 2, -1, -2, 0, 0, 0, 2, 2, 2, 1, 1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 1, 0, 1, 1, 2, 4, 5, 3, 2, 1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -2, -1, -2, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 3, 2, 0, -1, -1, 0, 1, 0, 0, 0, -1, -1, -1, -2, -3, -3, -3, -3, -3, -2, -1, 0, 0, 0, 0, -1, -2, 0, -1, 0, 1, 2, 2, 2, 0, -1, 0, 0, 0, 0, -1, 0, -2, -2, -3, -2, -4, -5, -4, -5, -5, -3, -3, -3, -1, -2, -1, -2, -1, -1, -1, 0, 0, 2, 1, 0, 0, -1, -1, 0, 0, -1, -1, 0, -3, -3, -4, -2, -3, -4, -5, -4, -5, -4, -4, -4, -4, -2, -2, -1, -2, -1, -1, -1, 1, 0, 1, 1, 0, 0, -2, 0, 0, -1, -1, 0, -1, -3, -4, -5, -5, -4, -5, -6, -5, -4, -5, -4, -4, -2, -3, -2, -2, -2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, -2, -4, -5, -6, -6, -4, -3, -5, -5, -3, -5, -4, -4, -4, -2, -3, -2, 0, 0, 0, 1, 1, -1, -1, 0, 0, 1, 0, -1, -1, 0, 0, -1, -2, -3, -5, -5, -3, -3, -3, -3, -4, -5, -5, -4, -3, -3, -2, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -2, -4, -4, -3, -1, -2, -2, -2, -3, -3, -4, -3, -3, -2, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, -1, -3, -2, -2, -1, 0, 0, -2, -2, -3, -3, -3, -3, -3, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 1, 0, 1, 0, -1, -1, -2, -2, -3, -2, -2, -1, 0, -1, -3, -3, -4, -2, -4, -3, -3, -1, 0, 0, 0, -1, -2, -2, -1, 1, 1, 2, 1, 2, 1, 0, 0, 0, -3, -3, -3, -2, -2, -2, -2, -3, -3, -3, -2, -1, -2, -2, -2, -1, -2, -1, -2, -2, -2, -2, -1, 1, 0, 2, 1, 1, 1, 0, 0, -1, -3, -2, -3, -2, -2, -1, -1, -2, -2, -2, -2, -1, 0, -2, -2, -4, -3, -1, -2, -3, -3, -1, -1, 0, 0, 1, 1, 2, 0, 0, -1, -2, -2, -4, -3, -3, -2, -1, -3, -1, -2, -2, -1, -1, -1, -2, -3, -4, -3, -2, 0, 0, -2, 0, 0, 0, 0, 2, 2, 1, 0, 0, -2, -3, -2, -3, -2, -4, -2, -2, -3, -2, -1, 0, -1, 0, 1, -2, -4, -4, -4, -3, -2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -2, -3, -4, -3, -4, -4, -1, -1, -1, -1, -1, 0, 0, 0, -1, -2, -4, -3, -2, -1, -2, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, -1, -2, -3, -4, -3, -4, 0, 0, 0, 0, 0, 0, 0, -1, -2, -4, -4, -2, -1, -1, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -3, -3, -3, -4, -4, -2, -1, -1, -1, 0, 0, -2, -2, -3, -3, -4, -2, -1, -2, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, -2, -3, -4, -4, -4, -3, -3, -2, -3, -3, -1, -2, -3, -3, -2, -3, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, -1, -4, -3, -4, -3, -3, -4, -4, -3, -3, -2, -3, -3, -3, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, -1, -3, -3, -3, -3, -4, -3, -3, -4, -4, -4, -3, -2, -2, -1, 0, -1, -1, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 2, 1, -1, -1, -2, -2, -2, -2, -4, -3, -4, -3, -3, -2, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 0, 1, 1, 0, 1, 1, 1, 0, 0, -1, -2, -1, -1, -4, -3, -2, -3, -3, -1, -1, -1, 0, 0, 0, 0, 0, 1, 2, 3, 3, 3, 2, 0, 0, 2, 1, 2, 2, 1, 0, 0, 0, 0, -1, 0, -2, -2, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 3, 4, 4, 1, 0, 0, 0, 2, 1, 0, 1, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 2, 2, 5, 4, 4, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 1, 1, 0, 0, 0, -1, -2, 0, 0, 0, 1, 2, 3, 3, 2, 2, 3, 2, 0, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 2, 2, 2, 2, 1, 0, 0, 0, 0, 0, 1, 2, 4, 5, 2, 2, 2, 1, -2, -2, -3, -1, -1, 0, 0, -1, 0, 0, 1, 1, 2, 2, 2, 2, 3, 2, 1, 3, 2, 1, 2, 1, 1, 3, 4, 5, 3, 2, 1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 1, 1, 2, 2, 2, 1, 0, 1, 3, 3, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 3, 4, 3, 2, 3, 1, 2, 3, 2, 1, 3, 2, 1, 1, 0, 1, 1, 0, 0, -2, -2, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 2, 1, 1, 1, 2, 1, 2, 1, 3, 2, 3, 2, 2, 2, 2, 2, 1, -2, 0, -1, 0, 0, 1, 1, 2, 0, 0, 0, -1, -1, 0, 0, 2, 2, 0, 2, 1, 2, 1, 1, 2, 2, 1, 2, 3, 4, 3, 2, 1, 0, -1, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 0, 1, 0, 2, 2, 3, 4, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 2, 2, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -2, -1, -2, -2, -3, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 2, 0, -1, 0, 0, 0, 0, -1, 0, -1, -2, -1, -2, -2, -2, -3, -3, -3, -3, -2, -2, -1, -1, -1, 0, 0, 0, -1, 0, 1, 2, 2, 1, 0, -1, 0, 0, 0, 0, 0, -1, -2, -2, -2, -1, -3, -2, -4, -4, -3, -4, -3, -2, -2, -1, -2, -1, -1, 0, -1, -1, 0, 1, 1, 1, 0, -1, -1, 0, 0, -1, 0, -1, -1, -2, -2, -2, -3, -2, -2, -3, -3, -3, -2, -3, -3, -3, -1, -1, -2, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -3, -3, -2, -1, -1, -1, -1, -3, -3, -3, -3, -3, -2, -3, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -3, -2, -2, -1, -1, -2, -1, -3, -4, -4, -2, -4, -2, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -2, -2, -3, -2, -2, -1, -1, -2, -3, -4, -4, -4, -4, -2, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, -2, -1, -2, -2, -1, -1, -2, -2, -2, -2, -3, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, -1, -2, -2, -2, -1, -2, 0, -1, -3, -2, -3, -2, -1, -2, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 2, 0, 0, 0, -1, -2, -2, -3, -2, -3, -1, -2, -3, -2, -2, -1, -1, -2, -2, -1, -2, 0, -1, -1, -1, -1, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, -2, -1, -3, -3, -3, -2, -1, -2, -2, -2, -2, -1, -1, 0, -1, -2, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -2, -2, -3, -3, -3, -2, -2, -1, -3, -3, -1, 0, 0, -1, -3, -3, -3, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, -2, -1, -3, -2, -3, -2, -1, -3, -2, -1, -2, -1, 0, 0, -1, -2, -3, -4, -3, 0, -1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -2, -3, -3, -3, -3, -2, -1, -1, 0, -1, -2, 0, -1, 0, -1, -3, -2, -2, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, -1, -1, -3, -2, -2, -2, -2, -1, 0, 0, -1, -1, 0, -1, -1, -2, -2, -2, -2, -1, 0, 1, 2, 2, 0, 0, 0, 1, 0, 0, 1, 0, -1, -1, -2, -4, -4, -3, -1, -1, -2, 0, -1, -1, -1, -1, -1, -2, -1, -1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -3, -3, -3, -3, -2, -1, -3, -2, -1, -2, -3, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -3, -2, -2, -2, -1, -2, -3, -1, -2, -2, -1, -2, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -3, -2, -3, -3, -3, -1, -2, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, -2, -1, -3, -2, -2, -1, -2, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 3, 1, 0, 0, 1, 0, 0, 2, 1, 1, 0, -1, 0, 0, 0, -1, -2, -1, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 3, 4, 1, 1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 3, 3, 1, 1, 0, -1, 0, 0, 1, 1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 3, 3, 2, 0, 0, -1, 0, 0, -1, 0, -1, -1, -2, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 2, 2, 2, 2, 0, 2, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 1, 2, 1, 0, 1, 0, 1, 0, 0, 2, 3, 2, 2, 1, 1, 0, 0, -1, -3, -2, -1, -2, 0, -1, 0, 0, 1, 0, 0, 0, 1, 2, 1, 1, 0, 2, 2, 1, 2, 2, 0, 1, 1, 3, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, -1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -2, -1, 0, 0, -1, 1, 1, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, 1, 1, 0, -1, -1, 0, -1, -2, -2, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, 2, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, 0, -2, -1, 1, 1, 0, 0, 0, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -2, -1, 0, -1, -2, -1, -1, -1, -2, 0, 1, 1, 0, 1, 0, 1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, 0, -1, -2, -2, -2, -2, -2, -2, 0, 1, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, -1, 0, -2, -3, -3, -2, -3, -2, -2, -2, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, -1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -3, -3, -3, -4, -2, -2, -2, -1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, -2, -2, -1, -3, -3, -3, -2, -3, -2, -1, -1, 0, 1, 1, 0, 3, 3, 0, 0, 0, -1, 0, 0, 2, 1, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, -3, -2, -3, -3, -2, -2, -2, 0, 0, 0, 1, 0, 2, 2, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -2, 0, -1, -2, -1, -2, -2, -2, -3, -3, -1, -2, -1, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -2, -1, -1, 0, -2, 0, 0, -1, -2, -3, -3, -2, 0, 0, 1, 2, 1, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -2, -2, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -3, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 1, 1, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -2, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, 1, 0, 0, 1, 2, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 2, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -2, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, -2, -2, -2, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -2, -1, -2, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, -1, 0, -1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, -2, -1, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, -2, -1, -1, -1, -1, -2, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 2, 1, 2, 2, 1, 0, 1, 1, 0, -1, 0, -1, 0, 0, 0, -1, -2, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 1, 0, 1, 1, 2, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 2, 2, 2, 2, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, -2, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 2, 2, 0, 0, 1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, 1, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 2, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 2, 1, 2, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -2, -2, -1, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, 0, -1, -2, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -2, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, -2, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, -1, -3, -3, -3, -1, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, -1, -2, -2, -1, -1, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, -2, -3, -2, -1, -1, 0, 0, -1, -1, 0, 0, -1, -2, -1, 0, 0, -2, -2, -2, -2, 0, -1, -1, -1, -1, -2, -1, -1, 0, 0, 0, 0, -2, -2, -3, -1, -1, -1, 0, 0, 0, -2, 0, 0, 0, 0, -1, -1, 0, -1, -1, -2, 0, 0, 0, 0, -2, -1, 0, 0, -1, 0, -1, 0, -2, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -2, 0, -1, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -2, -2, -1, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -3, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, -1, 0, -2, 0, 0, 1, 0, 0, 0, 0, -1, -1, -2, -1, 0, -2, -2, -1, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, -1, -2, -1, -2, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -2, -1, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, 2, 2, 1, -1, -1, 0, -1, -2, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -2, -1, 0, 0, -1, 0, 1, 1, 0, 0, 0, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, -2, 0, 0, 2, 0, 0, 1, -1, -1, -3, -3, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -2, -1, -1, 0, 0, 1, 1, 0, -1, 0, -2, -2, -1, -1, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, -1, -2, -1, -1, -2, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, -2, -1, -2, 0, -2, -1, -2, 0, 0, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, -1, -1, -1, -2, 0, 0, -1, -2, -2, -2, -2, -2, -1, -1, 0, 0, -1, -1, -2, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, -1, -1, -2, 0, 0, -2, -1, 0, 0, -2, -1, -3, -3, -1, 0, 0, -1, 0, -1, -2, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, 0, -1, -2, 0, -1, 0, -1, -1, -1, -2, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -2, 0, 0, 0, -1, -1, -2, -1, -1, -2, -1, -1, -2, 0, -3, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -1, 0, 0, -2, -1, -1, -2, -2, -1, -1, 0, -1, -2, -1, -1, 0, -1, -2, -1, -2, -2, -1, -2, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -2, -1, 0, -2, -1, -1, 0, 0, -2, -1, -2, -2, 0, 0, -2, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -1, -1, -1, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -2, -2, -2, -1, 0, 0, 0, -1, -1, -2, -1, -1, -1, -2, -2, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, 0, 0, -1, 0, -2, -1, -1, -1, -2, -3, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -2, -1, 0, -1, -1, -3, -3, -3, -3, -3, -2, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -2, -2, -2, -1, -3, -2, -3, -2, -3, -3, -1, -3, -2, 0, 0, 0, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -2, -1, 0, -2, -1, -2, -2, -3, -3, -3, -1, -2, -2, 0, 0, 0, -2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -2, -2, -1, -2, -2, -2, 0, -1, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 2, 2, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 2, 3, 1, 1, 0, 1, 2, 1, 0, 0, 0, -1, -1, -3, -3, -4, -4, -3, -2, -3, -1, -1, -1, -2, 0, -1, 0, -2, 0, -1, 0, 1, 2, 3, 0, 0, 0, 0, 0, 0, -1, -1, -1, -3, -4, -4, -5, -5, -3, -3, -2, -2, -2, -1, -1, -2, -1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -4, -4, -5, -5, -2, -2, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -3, -3, -4, -2, -2, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, -3, -3, -3, -2, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, -1, 0, 0, -1, -1, -2, 0, -1, -1, -2, 0, 0, 1, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 2, 2, 0, 0, 0, 1, 0, 1, 0, 2, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, -1, -1, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 2, 1, 3, 2, 1, 0, 1, 0, 0, 1, 2, 1, 0, 0, -1, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 2, 3, 4, 5, 4, 4, 3, 3, 3, 3, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 1, 4, 5, 7, 6, 6, 6, 5, 4, 2, 2, 1, 0, 1, 0, 0, 0, 0, -2, -1, -2, -2, -2, -3, 0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 6, 6, 6, 5, 5, 5, 4, 5, 4, 3, 1, 2, 0, 0, 0, -1, -1, 0, -1, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 5, 5, 5, 5, 6, 5, 4, 4, 3, 4, 4, 3, 1, 0, 0, 0, 0, -1, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 2, 3, 5, 6, 7, 7, 5, 6, 3, 3, 3, 3, 2, 2, 2, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 4, 6, 7, 6, 6, 6, 3, 3, 3, 4, 3, 2, 1, 1, 0, 0, 2, 1, 0, 1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 1, 2, 2, 5, 6, 7, 6, 5, 3, 3, 3, 4, 4, 4, 2, 1, 1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, -1, -1, -1, 0, 0, 2, 2, 3, 6, 6, 7, 6, 5, 4, 5, 3, 3, 4, 3, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 2, 2, 4, 5, 5, 6, 5, 4, 4, 4, 3, 2, 2, 2, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 2, 3, 3, 3, 4, 5, 3, 2, 4, 3, 2, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 2, 1, 3, 3, 5, 3, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 3, 2, 1, 0, 0, -1, 0, -1, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, -2, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, -1, -1, -2, -3, -4, -3, -3, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -3, -1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -2, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -3, -3, -1, -1, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 1, 2, 0, 1, -1, -1, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -2, -2, -2, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 2, 1, 2, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -2, -2, -3, -2, -1, -1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -2, -2, -2, -4, -4, -5, -6, -4, -3, -2, -1, 0, 0, -1, -1, 0, 0, 2, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, -1, -1, -2, -2, -2, -2, -2, -4, -5, -4, -4, -4, -1, -1, 0, -1, 0, -2, -2, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -2, -2, -4, -4, -4, -2, -1, -1, -1, -2, -2, -2, -3, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, -1, -1, -2, -3, -4, -4, -4, -2, 0, -1, 0, -2, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -3, -4, -4, -4, -3, -3, -2, -2, -2, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -3, -1, -1, -2, -4, -3, -4, -3, -2, -3, -1, -2, -1, -1, -1, -1, 0, -1, 0, -1, -2, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, -2, -3, -2, -1, -2, -2, -2, -1, -2, -1, -2, 0, -2, -1, -1, 0, 0, 0, 0, 0, -1, -2, -2, -1, 0, 1, 1, 0, 0, 1, 2, 0, -1, -2, -1, -2, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, -2, -1, -3, -1, 0, 0, 0, 0, 0, 1, 2, 0, -1, 0, -1, -1, 0, 2, 1, 2, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, -1, -2, -1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 2, 4, 3, 5, 4, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -3, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 4, 5, 5, 6, 6, 3, 2, 2, 2, 1, -1, -1, -1, -1, -1, -2, -3, -2, -2, -3, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 2, 4, 3, 5, 6, 4, 4, 2, 3, 3, 3, 1, 0, 0, -1, -3, -3, -2, -3, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 3, 3, 4, 4, 5, 4, 3, 4, 3, 4, 3, 2, 0, -2, -3, -2, -1, -2, -2, -2, -3, 0, 1, 0, -1, 0, 0, 0, 1, 0, 1, 2, 3, 2, 4, 6, 6, 4, 4, 4, 5, 5, 4, 1, 0, -3, -2, -2, -1, 0, -2, -2, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 3, 3, 5, 4, 6, 4, 4, 4, 5, 5, 6, 4, 3, 0, -2, -2, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 3, 4, 4, 5, 5, 5, 5, 5, 5, 7, 6, 4, 1, -1, -4, -3, -3, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 4, 3, 4, 5, 5, 5, 7, 6, 7, 4, 3, 0, -3, -5, -4, -1, -2, -3, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 2, 3, 5, 4, 6, 6, 4, 5, 3, 3, 0, -1, -3, -2, -3, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 3, 4, 3, 3, 4, 2, 3, 3, 1, 0, -2, -1, -2, -1, -2, -2, -1, 0, 0, -1, -2, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, -1, -1, -1, -2, -1, -1, -1, 0, 0, 0, -2, -2, 0, 0, -1, 0, 0, -1, 0, 0, -2, -3, 0, 0, 0, 0, -2, -1, -2, -1, 0, 0, 0, -1, 0, 0, -1, 0, -2, -1, 0, -2, -2, -2, 0, 0, -1, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, -2, -2, -2, -2, -3, -1, -1, -1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, 1, 1, 1, 1, 0, 0, -2, -2, -2, -2, 0, 0, -1, -3, -2, -3, -4, -4, -3, -3, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, -2, -1, -2, -1, 0, -1, -1, -1, -2, -3, -3, -2, -2, -2, -1, 0, 0, 0, 1, 1, 0, 1, 2, 1, 1, 0, 1, 0, 2, 0, 0, 0, -2, 0, -1, -1, -1, -1, -1, 0, -1, -1, -2, -2, -2, -2, 0, 0, 0, 0, 0, 2, 1, 2, 3, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, -2, -2, -2, -2, -1, 0, 0, 0, 0, 1, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, -1, -1, -1, -1, -2, 0, -2, 0, 0, 0, 0, 1, 2, 3, 3, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 1, 1, 1, 4, 4, 3, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 2, 1, 1, 1, 1, 0, -1, 0, -1, -1, 0, 0, 1, 0, 1, 2, 2, 2, 2, 4, 2, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 4, 4, 2, 2, 0, 1, 0, 0, 0, 0, -1, -1, -1, -3, -4, -3, -3, -3, -2, -2, -2, -1, 0, -2, 0, -2, 0, 0, 0, 1, 2, 0, 5, 4, 3, 2, 1, 0, 0, 0, 0, -1, -1, -2, -3, -6, -7, -6, -5, -5, -4, -4, -2, -3, 0, -1, -1, 0, 0, 0, 0, 1, 1, 2, 4, 4, 3, 2, 1, 0, 0, 0, 0, -2, -2, -3, -5, -7, -7, -6, -5, -5, -2, -4, -4, -2, -3, -3, -1, -1, 1, 1, 0, 1, 1, 0, 2, 3, 3, 0, 0, 0, -1, 0, 0, -1, -1, -3, -3, -6, -6, -6, -3, -1, -1, -2, 0, -1, -2, -2, -1, 0, 1, 2, 2, 3, 2, 2, 3, 4, 2, 1, 0, 0, -1, -1, 0, 0, 0, -3, -3, -2, -3, -2, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 1, 3, 2, 3, 2, 2, 1, 3, 1, 1, 1, 2, 0, 0, 0, 1, 0, -2, -2, -3, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 3, 2, 1, 1, 2, 2, 0, 0, 2, 3, 2, 0, -1, 0, 2, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 3, 1, 2, 0, 0, 0, 3, 4, 4, 2, 0, 2, 2, 1, 1, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 2, 2, 1, 0, 0, 0, 3, 3, 3, 0, 0, 3, 2, 2, 2, 3, 2, 1, 2, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, -1, -1, 0, 0, 2, 0, 0, -1, 0, 1, 1, 1, 1, 1, 3, 2, 2, 5, 3, 4, 3, 3, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 4, 4, 4, 4, 6, 4, 5, 5, 4, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 3, 6, 6, 7, 5, 6, 7, 5, 6, 3, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 4, 6, 7, 7, 8, 9, 8, 7, 6, 5, 5, 4, 1, 1, 1, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 1, 2, 0, 1, 1, 2, 3, 6, 6, 7, 8, 9, 8, 9, 7, 7, 7, 6, 4, 0, 0, -1, 0, 0, 1, 3, 1, 1, 0, 0, 1, 1, 1, 2, 1, 1, 2, 2, 4, 5, 7, 7, 9, 10, 9, 8, 8, 8, 7, 7, 3, 0, 0, 0, 0, 1, 3, 4, 2, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 3, 4, 7, 7, 7, 9, 9, 7, 6, 8, 9, 8, 5, 3, 0, -1, 0, 1, 2, 3, 4, 4, 2, 2, 1, 1, 0, 1, 1, 1, 2, 1, 4, 5, 8, 8, 8, 9, 8, 7, 7, 8, 9, 7, 4, 1, 0, -1, 0, 1, 3, 2, 3, 3, 2, 3, 3, 1, 0, 0, 1, 2, 2, 2, 4, 5, 7, 6, 7, 7, 6, 7, 7, 8, 9, 6, 4, 2, 1, 0, 0, 0, 1, 1, 2, 3, 2, 3, 1, 2, 0, -1, 1, 1, 2, 2, 3, 4, 7, 8, 6, 7, 7, 6, 6, 7, 7, 5, 4, 4, 2, 0, 0, 0, 0, 1, 2, 3, 2, 0, 2, 1, 0, 0, 0, 0, 2, 3, 3, 3, 5, 6, 7, 6, 5, 6, 6, 6, 5, 5, 4, 4, 2, 2, 0, 2, 1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 1, 2, 1, 1, 2, 5, 7, 6, 4, 4, 5, 5, 6, 5, 3, 4, 4, 3, 2, 2, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 1, 4, 6, 4, 2, 3, 2, 3, 3, 2, 2, 4, 4, 3, 2, 1, 1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 2, 3, 3, 1, 0, 1, 1, 2, 1, 2, 3, 3, 1, 0, 2, 1, -1, -2, -1, 0, 0, -1, -1, -1, 0, 0, -1, -2, -1, -1, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 2, 1, 1, 1, -1, -1, -1, -1, 0, 0, -1, -1, 1, 1, 0, -2, -2, 0, 1, 0, 0, 1, 0, 0, 0, 0, -2, -2, -1, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -2, 2, 2, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -2, -2, -3, 0, 2, 2, 0, 0, 1, 0, 1, 2, 3, 2, 1, -1, -2, -2, 1, 1, 0, -1, -1, 0, 1, 1, 0, 0, 0, -1, -3, -3, -3, -3, -2, 0, 0, 2, 0, 0, 1, 2, 3, 3, 3, 3, 1, -1, -2, 0, 1, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, -1, -3, -3, -5, -4, -1, 0, 0, 0, 0, 0, 1, 2, 3, 3, 2, 0, 1, -1, -2, -1, 3, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, -3, -5, -5, -4, -3, -2, 0, 0, -1, 0, 1, 1, 2, 2, 1, 0, 0, 0, 0, -1, -2, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -4, -6, -4, -4, -3, -2, -2, -2, -1, 0, 1, 2, 2, 1, 1, 1, 0, 0, 0, -1, -1, 3, 3, 2, 0, 1, 0, 0, 0, 0, -1, -2, -2, -3, -4, -4, -2, -2, -1, -1, -1, 0, 1, 1, 2, 1, 1, 0, -1, 0, 1, 1, 0, 2, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -2, -3, -2, -1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0,
    -- filter=0 channel=7
    0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 2, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 2, 2, 1, 1, 2, 2, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 2, 1, 1, 1, 1, 1, 1, 0, 1, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 2, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 2, 2, 1, 2, 1, 2, 2, 0, 1, 1, 1, 1, 3, 0, 1, 0, -1, -1, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 2, 1, 2, 1, 2, 1, 0, 0, 2, 2, 1, 2, 1, 1, 2, 3, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 1, -1, -2, -2, 0, -1, -1, 0, -1, -1, -1, -2, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -2, -2, 0, -1, 0, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, -2, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, -2, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -2, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -2, -1, -2, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -2, -3, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, -1, -3, -3, -3, -2, -2, 0, 1, 0, 0, 0, -1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -2, -3, -2, -2, -1, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -2, -2, 0, 0, 2, 2, 3, 1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, -2, -1, -1, 0, 1, 2, 3, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, -2, -2, -2, -1, -1, 0, 1, 3, 1, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -2, -3, -3, -2, -1, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -2, -3, -4, -4, -3, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -2, -2, -1, -2, -2, -3, -2, -3, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, -2, -2, -2, -2, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, 0, -2, 0, 0, 0, -1, 0, -1, 0, -2, -2, -3, -3, -2, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 1, 0, -1, -1, -1, -2, -1, 0, -1, -1, -2, -1, -2, 0, -2, -2, -1, -2, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, -1, -2, 0, -1, -2, -2, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -2, -2, -2, -2, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, -1, -1, 0, -1, 0, 0, -1, -1, -3, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -2, -1, -1, 0, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 2, 0, 1, 0, -1, -1, -1, -1, 0, -1, -1, -2, -1, -1, 0, -1, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 1, -1, -1, -1, 0, -1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 2, 0, 2, 1, 1, 1, 0, 0, 0, 1, 1, 1, 1, 2, 2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 0, 1, 1, 0, 1, 2, 1, 2, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, -1, 0, -1, -1, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -2, -1, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, -1, -2, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 0, -1, -1, 0, -1, -2, -2, -1, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 2, 2, 0, 2, 1, 2, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, -2, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 2, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 2, 1, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -2, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 2, 2, 1, 1, 1, 2, 0, 1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 1, 1, 1, 1, 2, 3, 2, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 3, 2, 2, 2, 1, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 2, 1, 2, 1, 3, 2, 2, 2, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 2, 3, 2, 2, 1, 1, 0, 1, 0, -1, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 3, 3, 2, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 3, 3, 2, 2, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 2, 2, 3, 1, 2, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 2, 2, 2, 1, 2, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 2, 2, 2, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 1, 1, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 1, 1, 2, 3, 2, 1, 2, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, -1, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 1, 2, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 2, 1, 1, 1, 1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 3, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 3, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 1, 0, 2, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, -1, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 1, 0, 1, 1, 1, 3, 2, 1, 1, 1, 0, 0, -1, -2, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 3, 3, 2, 3, 3, 3, 1, 2, 0, -1, -2, -2, -1, -1, -1, -2, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 2, 3, 3, 3, 3, 3, 1, 0, -2, -2, -3, -3, -1, 0, -1, -2, -2, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, 1, 1, 1, 3, 3, 2, 3, 1, 3, 0, 0, -2, -3, -2, -3, 0, 0, -1, 0, -2, -1, -1, -1, -1, -1, -1, 0, 0, -1, 0, -1, -1, 0, 1, 2, 2, 3, 1, 2, 2, 2, 1, 0, -1, -3, -2, -1, -1, 0, 1, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -2, 0, 0, 0, 0, 2, 2, 1, 0, 1, 2, 1, 0, 0, -1, -2, -2, -2, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 2, 1, 2, 2, 1, 0, 2, 0, 0, -2, -3, -2, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 2, 1, 2, 2, 1, 1, 1, 1, 0, -2, -3, -2, -1, -1, 1, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 1, 1, 2, 2, 1, 2, 1, 0, 1, 0, -1, -3, -2, -2, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 2, 2, 0, 0, 0, 0, -2, -3, -1, -2, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 2, 2, 2, 0, 1, 0, 0, -2, -2, -2, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 2, 3, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 2, 2, 1, 2, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 2, 1, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 1, 1, 0, 0, 2, 1, 2, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 2, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 2, 4, 2, 1, 1, 0, 1, 0, 0, -2, -2, -2, -1, 0, 1, 2, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, -1, 0, 2, 3, 4, 2, 2, 1, 0, 0, -2, -2, -2, -3, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, -2, -2, -3, -2, 0, 0, -2, -2, -3, -1, 2, 4, 3, 1, 0, 0, -1, -1, 0, -1, -1, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -2, -2, -2, 0, 2, 2, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -2, -1, -2, 0, 0, 0, -2, -2, -2, -1, 2, 3, 2, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, -1, -1, 0, -1, -1, 0, 0, -2, -1, -2, -1, 1, 2, 1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 3, 1, 0, -1, 0, 0, 0, 0, -2, 0, 0, 1, 1, 0, 0, 1, 2, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, -1, 0, 1, 3, 1, 2, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 2, 3, 2, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 3, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 3, 3, 2, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 3, 2, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 3, 4, 3, 1, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, -1, 0, -1, -1, -1, 1, 1, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 3, 2, 2, 2, 0, -1, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 2, 1, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 2, 3, 4, 3, 2, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, -2, -2, -2, 0, 0, 0, 0, 0, -1, 1, 2, 3, 2, 2, 0, -1, -2, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 1, 1, 0, -2, -3, -3, -2, 0, 0, 0, 0, 0, 2, 3, 3, 3, 3, 2, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 1, 0, -2, -2, -1, 0, 0, 1, 2, 0, 0, 1, 5, 5, 4, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -1, 1, 2, 1, 0, 0, 0, 0, 2, 1, 1, 1, 2, 3, 3, 5, 4, 2, 2, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -1, 2, 3, 0, 0, 0, 0, 1, 2, 1, 1, 3, 3, 4, 5, 5, 4, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, -2, 2, 4, 2, 1, 0, 0, 1, 2, 2, 2, 2, 3, 4, 4, 3, 2, 2, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 3, 3, 2, 1, 1, 1, 1, 0, 1, 3, 3, 2, 2, 2, 2, 2, 2, 0, 1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, -1, -2, 0, 3, 3, 1, 2, 0, 1, 0, 2, 3, 3, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, -1, -1, 0, 3, 4, 1, 1, 0, 0, 0, 2, 1, 3, 2, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 3, 3, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, -3, -2, 3, 2, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -3, -1, -2, 3, 4, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, -1, -2, -2, 3, 3, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, -1, -2, -2, -2, 3, 5, 3, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, -1, -1, -1, -1, -1, -2, -3, -3, -2, 4, 4, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, -2, -2, -2, -2, 2, 5, 4, 3, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, -1, 0, -1, 0, -1, -1, -2, -2, 0, 1, 2, 2, 3, 2, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, 1, 0, 2, 1, 1, 1, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -3, -1, 0, 0, 0, 1, 1, 1, 0, 1, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -2, -4, -2, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -2, -3, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, 0, 0, -1, -1, 0, -1, -1, -1, 0, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -2, -1, -1, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -3, -2, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -3, -1, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -2, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 1, -1, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -2, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 1, -1, 0, 0, 0, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, -2, 0, -1, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, -1, 0, 0, -2, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -2, -1, -1, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -2, -2, -1, -2, -1, 0, 0, -1, -2, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -1, -1, -2, -1, -1, -1, -2, -2, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, -2, -1, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, -3, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, -3, -2, 0, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -3, -2, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -3, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, -1, 0, -1, 0, -1, -4, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -3, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 1, 1, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 2, 3, 2, 1, 2, 2, 1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, 2, 0, 0, 0, -2, -2, -1, -1, -1, -1, -3, -2, 0, 3, 3, 1, 2, 3, 1, 2, 1, 0, -1, -1, 0, 0, 1, 0, 0, 1, 2, 0, 2, 0, 0, 0, -2, -2, -1, -3, -2, -2, -4, -3, 0, 2, 2, 1, 2, 1, 1, 1, 1, -1, -1, -1, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, -1, 0, -2, -1, 0, -2, -1, -2, -3, -3, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, -1, 0, -2, -1, -1, -1, -3, -3, 0, 1, 2, 0, -1, 0, 0, -1, -2, -1, -1, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -2, -1, -1, -2, -3, 0, 1, 0, 0, -1, -1, -2, -1, -3, -3, -2, -1, -2, -1, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, -1, -2, -1, -1, -1, -2, -3, -3, -3, -3, -3, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 2, 1, 0, 0, 0, 0, 0, -1, -2, -3, -3, -4, -2, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -1, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -3, -3, -4, -2, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, 0, 2, 2, 1, 1, 0, 0, 0, 0, -3, -2, -2, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 3, 2, 1, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, -1, 0, 2, 2, 1, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, -2, 0, -1, 0, 2, 1, 0, 0, 0, 2, 0, 0, -2, -1, -1, -1, 1, 1, 0, 0, 0, -2, -3, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, -2, -2, 0, 0, 1, -1, 0, 0, 0, 1, 0, -1, -2, 0, 0, 1, 1, 2, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, 0, 2, 1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 1, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 2, 1, 0, 0, -1, -2, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, -1, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -2, 0, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 1, 2, 1, 0, 0, 0, 0, 0, -2, -2, -1, -1, 0, 1, 0, 0, -1, -2, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, 1, 3, 1, 1, 0, -1, -1, -2, -1, -1, -1, -1, 0, 1, 0, 0, -1, -1, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, 1, 3, 2, 1, 0, -1, -2, -1, -2, -2, 0, 0, -1, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 3, 2, 1, 0, 0, 0, -2, -2, -2, -1, -1, -1, -2, -1, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, 1, 3, 2, 1, 0, 0, -1, -1, -2, -1, -1, -2, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -3, 0, 3, 3, 0, 0, -1, -1, -1, -2, -3, -2, -2, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 1, 2, 0, 0, 0, 0, -1, -2, -3, -2, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, 0, 2, 1, 0, 0, -1, -1, -1, -1, -2, -1, -2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, -2, -3, 1, 2, 3, 0, 0, -1, 0, 0, 0, -1, -2, 0, -1, 0, 1, 0, 0, -1, 0, 0, 2, 2, 1, 0, 0, 0, -1, 0, 0, 0, -3, -3, 0, 3, 4, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 2, 2, 1, 1, 1, 0, 0, -1, 0, -1, -1, -3, -4, 0, 2, 3, 3, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, -1, -4, -3, 1, 2, 4, 3, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, -1, -1, -2, -1, -3, 0, 2, 2, 2, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 3, 3, 3, 3, 2, 2, 1, 2, 2, 1, 1, 2, 3, 2, 3, 2, 1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 2, 3, 5, 6, 7, 7, 4, 4, 2, 2, 2, 2, 1, 1, 2, 1, 3, 4, 4, 1, -1, -2, -2, -3, -2, 0, 0, -1, -1, -2, -1, 0, 1, 2, 4, 5, 5, 6, 5, 3, 1, 1, 1, 2, 0, 0, 1, 0, 1, 3, 1, 1, -2, -2, -3, -2, -2, -1, -1, -1, -2, -2, -2, -1, 0, 1, 3, 3, 3, 3, 4, 2, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, -1, -2, -3, -2, -1, -2, -2, -4, -4, -4, -2, -1, 1, 1, 2, 2, 3, 4, 3, 2, 1, 1, 1, 0, 1, 0, 1, 2, 0, 0, 0, 0, -2, -1, -4, -2, -2, -2, -3, -4, -4, -3, -2, -1, 0, 1, 1, 3, 3, 3, 2, 0, 1, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 1, -1, -2, -3, -2, -3, -2, -1, -2, -5, -4, -3, 0, 2, 0, 1, 1, 1, 3, 2, 1, 2, 0, 2, 1, 0, -1, -1, 0, 1, 0, 1, 1, 0, -2, -3, -4, -3, -2, -1, -2, -2, -3, -3, -2, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 2, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -3, -2, -2, -2, -1, 0, -2, -2, -2, -2, -1, 0, -1, -1, 0, 0, 2, 1, 2, 1, 1, 2, 0, 0, 1, 1, 1, 2, 0, 0, -1, -1, -2, -2, -2, -1, -1, 0, 0, -2, -1, 0, 0, -2, -1, 0, -1, 0, 0, 0, 2, 3, 3, 4, 2, 1, 0, 1, 2, 2, 1, 0, -1, 0, -1, -1, -1, 0, -1, -2, -1, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, 0, 2, 3, 3, 4, 3, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -3, -3, -5, -5, -4, 0, 1, 3, 1, 2, 1, 0, 0, 1, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -3, -5, -7, -8, -4, -2, 0, 3, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -4, -7, -7, -5, -3, 0, 5, 6, 5, 3, 2, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -3, -6, -6, -4, -2, 2, 7, 9, 7, 5, 2, 2, 1, 1, 0, 0, 0, -1, 0, -3, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, -3, -7, -7, -4, 0, 3, 7, 9, 8, 6, 2, 0, 0, 1, 1, 1, 0, -1, 0, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -4, -6, -7, -5, -1, 1, 6, 7, 7, 5, 2, 0, -1, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -4, -7, -7, -5, -3, 1, 4, 7, 7, 3, 1, 0, -1, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -3, -5, -7, -8, -7, -2, 0, 4, 4, 5, 3, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 1, 0, -1, -1, -3, -4, -5, -7, -6, -3, 0, 3, 4, 3, 2, 0, -1, 0, 1, 0, 0, 1, 0, -1, -1, 0, -1, -2, 0, 0, 0, 0, 1, 0, -3, -3, -3, -5, -5, -5, -5, -1, 0, 3, 3, 5, 4, 1, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, -1, -1, 0, 0, 1, 0, 0, -1, -3, -4, -4, -3, -5, -3, -1, 0, 2, 3, 5, 5, 4, 0, 1, 0, 1, 2, 0, 0, -1, 0, -1, -2, -2, -1, -1, 0, 0, 0, 0, -2, -5, -5, -3, -3, -3, -2, -1, 2, 3, 4, 4, 4, 3, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, -1, -3, -2, -2, -1, -1, -3, -3, -4, -4, -4, -3, -2, -1, -2, 0, 1, 2, 3, 3, 3, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -3, -1, -3, -2, -4, -3, -4, -3, -3, -2, -3, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -1, -2, -3, -3, -3, -4, -5, -4, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 1, -2, -3, -3, -3, -1, -2, -4, -4, -6, -5, -5, -3, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, 0, 0, 2, 0, 0, -2, -2, -3, -3, -1, -2, -2, -4, -4, -5, -3, -3, -1, 0, 0, 0, 0, 1, 0, 1, 0, -1, -1, 0, -1, -1, 0, 0, 1, 1, 0, 0, -2, -1, -3, -1, -1, -1, -1, -4, -3, -3, -4, -2, 0, 0, 0, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 2, 0, 0, -1, -1, 0, 0, 0, -1, -3, -2, -3, -2, 0, 0, 0, 3, 3, 4, 4, 3, 3, 2, 1, 1, 1, 2, 3, 3, 5, 4, 5, 4, 0, 0, -1, 0, 0, 1, -1, 0, -1, 0, -1, 0, 0, 1, 0, 3, 5, 6, 6, 5, 3, 3, 4, 3, 3, 4, 3, 3, 4, 4, 5, 3, 1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 1, 1, 2, 3, 3, 3, 2, 2, 3, 2, 2, 2, 1, 2, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 2, 1, 1, 1, 1, 1, 2, 1, 0, 0, -2, 0, 0, 0, 0, -1, -3, -2, -1, -2, -2, 0, 0, 0, 0, 1, 0, 0, 1, 2, 3, 2, 3, 2, 3, 1, 3, 3, 2, 1, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, 0, -1, -1, -2, -1, -2, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 2, 0, 0, -2, -1, -1, 0, -1, 0, 0, -1, -1, 0, -1, -1, -2, -2, -3, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, -2, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, -1, -2, -2, -2, -3, -1, -1, -1, 0, -2, -2, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, -2, 0, 0, -1, -1, 0, 0, 1, 2, 0, 0, 0, 0, -2, -2, -2, -1, -1, -1, 0, 0, -2, -2, 0, 0, 0, -1, -1, -1, 1, 0, 0, -2, 0, 0, 0, -1, 0, 0, 0, 2, 2, 1, 0, -1, -1, -2, -2, -1, -2, -1, 0, 0, -1, -2, -1, -1, 0, 0, -2, 0, 0, 0, 0, -3, -2, 0, 0, 0, 0, -1, 0, 2, 2, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, -2, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 2, 2, 1, 1, -1, -1, -1, -1, 0, -1, 0, -1, 0, -1, -2, -2, 0, 0, -1, -2, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 2, 1, 1, 1, 2, 1, 0, 0, 0, 0, 1, 0, 0, 1, -1, -1, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 1, 1, 2, 0, 0, 0, 0, 1, 1, 2, 2, 0, 1, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 1, -2, -1, 0, 0, 0, 1, 0, 2, 1, 3, 3, 2, 1, 0, 0, 1, 3, 3, 4, 1, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 2, 2, 2, 3, 1, 0, 0, 0, 0, 3, 3, 1, 0, -2, -3, -1, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, -1, -2, -1, 0, 0, 0, 1, 3, 2, 3, 3, 1, 0, 0, 1, 2, 3, 2, 0, -3, -2, -3, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 2, 4, 6, 6, 3, -1, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 2, 4, 5, 7, 5, 0, 0, -3, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, -1, -1, 0, 1, 1, 4, 5, 6, 4, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 2, 3, 3, 4, 1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, -2, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 3, 3, 2, 1, 0, -2, -1, 0, 0, 0, 0, 2, 0, 0, -3, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -2, -2, -1, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 1, 0, -2, -1, -2, -2, 0, -1, 0, 0, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -3, -1, -1, -2, -1, 0, 1, 2, 2, 2, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, -2, -2, -1, 0, 0, 0, 0, 3, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 2, 1, 2, 1, 2, 0, 0, 0, 0, 0, 1, 0, -1, -2, -1, 0, -1, 0, 0, 0, 2, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 1, 0, 0, 0, 0, 0, -2, 0, -1, 0, -1, 0, 0, 1, 2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 2, 1, 2, 2, 1, 1, 0, 0, 0, 0, -3, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 2, 2, 2, 2, 2, 0, 0, 0, 0, -3, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 3, 0, 1, 2, 3, 2, 2, 2, 2, 1, 0, 0, -2, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -1, 0, 2, 1, 1, 1, 0, 0, 1, 2, 2, 0, -1, 0, -2, -3, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 0, 0, -2, 0, -1, 0, 0, 0, 1, 1, 2, 2, 2, 1, 2, 1, 2, 0, 0, -2, -2, -1, -1, 0, 1, 1, 1, 0, -1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 2, 2, 3, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 3, 3, 3, 2, 1, 1, 1, 0, 1, 2, 1, 0, 2, 1, 2, 3, 3, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 1, 1, 2, 1, 2, 2, 1, 1, 0, 0, 1, 1, 0, 0, 0, 2, 1, 1, 2, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 0, 0, 2, 2, 2, 0, 2, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 1, 1, 0, 0, 1, 1, 2, 1, 1, 1, 1, 0, -1, -2, 0, -1, 0, -1, -1, -1, -2, 0, 0, 0, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 1, 0, 0, -2, -1, -1, -1, 0, -2, -2, -2, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, -3, -3, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 2, 0, 0, -3, -2, -2, -1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 2, 1, 2, 1, 0, 0, -1, -1, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 1, 3, 1, 1, 1, 0, 0, -1, -2, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 1, 0, 2, 2, 3, 2, 1, 0, 0, -1, -2, -3, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, -1, 1, 1, 2, 1, 2, 3, 2, 1, 1, -1, -2, -2, -3, -2, -2, -1, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, -2, -2, 0, 0, 1, 1, 2, 2, 1, 2, 1, 2, 0, -2, -1, -4, -4, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, -2, -1, -2, -2, 0, 1, 0, 2, 0, 0, 0, 1, 1, 0, -2, -1, -2, -2, -1, 1, 2, 1, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -2, -2, -2, -2, -1, 0, 2, 2, 2, 0, 1, 1, 0, 0, -1, -1, -4, -2, -1, 0, 2, 2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, -1, -1, -1, -1, 0, 2, 0, 1, 1, 0, 1, 1, 0, -1, -1, -2, -3, -3, 0, 1, 2, 0, 0, -1, 0, 0, -2, -1, 1, 0, 0, -1, -2, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, -1, -4, -4, -2, 0, 1, 1, 2, 0, 0, -1, 0, -1, 0, 0, 0, 0, -2, -1, 0, -1, 0, 0, 0, 2, 1, 0, 1, 1, 0, 0, -1, -3, -3, -3, -1, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 1, 1, 1, 1, 1, 0, 0, -1, -1, -3, -2, -2, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 0, 2, 1, 0, 0, 0, -2, -3, -3, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 2, 2, 0, 0, 0, 0, -1, -3, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, -2, 0, -1, 0, 0, 0, 0, 2, 0, 0, -1, -1, -1, -1, -2, -2, -1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, -2, 0, 0, -1, 0, 0, 1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 2, 1, 0, -1, -3, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -2, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 3, 1, 0, 0, -1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 1, 1, 0, 2, 2, 1, 1, 1, 0, 1, 2, 0, 0, 2, 3, 2, 2, 4, 4, 2, 1, -1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 1, 2, 2, 2, 3, 3, 1, 2, 2, 1, 3, 2, 3, 2, 4, 3, 2, 4, 3, 2, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 3, 1, 2, 2, 2, 2, 1, 1, 0, 1, 1, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 0, 1, 2, 1, 2, 2, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 1, 0, 2, 1, 2, 3, 2, 2, 3, 3, 1, 1, 1, 1, 2, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 2, 3, 3, 1, 1, 1, 3, 3, 3, 4, 4, 3, 3, 4, 5, 3, 3, 1, 0, 0, 0, 0, 1, 1, 1, -1, -1, -2, -3, -2, 0, 0, 3, 4, 2, 2, 3, 4, 4, 4, 5, 5, 5, 3, 4, 4, 3, 4, 4, 0, 1, 0, 1, 0, -2, -1, 0, 0, -1, -2, -2, -1, 0, 1, 2, 3, 3, 3, 4, 3, 6, 5, 7, 5, 6, 5, 3, 1, 2, 1, 0, 0, 0, 1, 1, 0, -3, -2, -3, -1, -1, -1, -1, 0, 1, 1, 3, 2, 3, 2, 2, 4, 4, 6, 5, 5, 6, 5, 4, 1, 1, 0, 0, -1, 0, -1, -1, 0, -3, -2, -2, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 3, 4, 4, 2, 3, 3, 3, 2, 2, 1, 2, 2, 1, 0, 0, 0, -1, 0, 0, -3, 0, 0, 2, 2, 1, 2, 1, 1, 3, 3, 3, 3, 5, 5, 4, 4, 3, 4, 4, 2, 2, 2, 3, 4, 2, 4, 2, 2, 0, 0, 0, 0, 0, 1, 3, 4, 3, 2, 3, 3, 4, 3, 2, 3, 3, 2, 3, 4, 4, 5, 4, 5, 5, 4, 4, 3, 1, 1, 1, 1, 0, 0, 0, 0, 1, 2, 2, 2, 1, 2, 4, 4, 6, 5, 6, 2, 1, 3, 3, 4, 5, 4, 3, 2, 1, 3, 2, 2, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 3, 3, 4, 4, 5, 6, 7, 7, 7, 6, 3, 2, 3, 2, 1, 0, 0, -1, -1, 0, 0, 1, 1, 1, 0, -1, -1, 0, 0, 0, 1, 1, 2, 4, 4, 6, 5, 7, 7, 5, 6, 6, 5, 3, 2, 1, 1, 0, -1, 0, 0, 0, 2, 2, 2, 2, 0, 0, -1, 0, 0, 1, 3, 3, 3, 4, 6, 6, 7, 5, 6, 4, 3, 4, 2, 0, 0, 1, 1, 2, 3, 1, 0, 0, 1, 2, 2, 3, 1, 0, 0, 0, 1, 1, 4, 4, 3, 4, 5, 7, 7, 7, 5, 1, 2, 0, 0, 1, 0, 0, 0, 1, 2, 2, 1, 1, 0, 0, 1, 2, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 5, 6, 8, 6, 4, 3, 2, 1, 0, 1, 1, 0, 0, 0, 0, 1, 2, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 3, 5, 7, 8, 7, 6, 5, 4, 3, 1, 1, 2, 1, -1, 0, 0, 2, 2, 2, 2, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 3, 3, 4, 4, 5, 6, 4, 4, 3, 3, 2, 2, 1, 0, 0, 0, 1, 1, 3, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 1, 2, 3, 4, 2, 4, 5, 4, 4, 3, 3, 3, 3, 4, 4, 2, 1, 1, 2, 1, 1, -1, 0, -1, 0, 0, -1, 0, 2, 0, 0, 0, 0, 0, 1, 1, 3, 5, 5, 5, 5, 3, 1, 2, 2, 3, 3, 3, 3, 1, 1, 2, 1, 1, 0, 0, -1, -1, -2, 0, 1, 2, 1, 0, 1, 1, 3, 3, 3, 4, 6, 6, 7, 5, 4, 4, 2, 4, 3, 4, 4, 4, 3, 2, 1, 1, 0, 0, 0, -1, -2, 0, 0, 1, 0, 1, 0, 3, 3, 3, 3, 3, 3, 5, 5, 6, 5, 5, 5, 5, 6, 6, 5, 4, 4, 3, 2, 2, 2, 1, 0, -1, -1, 0, 0, -1, 0, 1, 1, 2, 3, 3, 5, 2, 2, 3, 6, 5, 4, 4, 6, 6, 8, 6, 5, 4, 4, 3, 3, 2, 2, 1, 0, 0, 0, -1, -2, 0, -1, 0, 1, 0, 1, 3, 4, 3, 2, 4, 4, 3, 4, 3, 4, 3, 3, 3, 4, 2, 2, 1, 1, 1, 1, 1, 1, 1, -1, -1, -1, -1, 0, 0, 0, 0, 2, 3, 3, 4, 3, 2, 2, 3, 1, 2, 3, 1, 2, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 2, 2, 2, 3, 1, 1, 0, 2, 2, 1, 2, 3, 2, 2, 2, 2, 1, 0, 1, 1, 0, 0, -2, -2, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 2, 0, 1, 0, 0, 0, 0, 0, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -4, -3, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 3, 2, 3, 3, 3, 2, 3, 1, 2, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -2, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, -2, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -2, -1, 0, -1, -1, -1, -2, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, -1, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, -2, -2, 0, 0, -1, 0, 0, 1, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 2, 2, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 2, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 1, 2, 2, 2, 2, 1, 2, 0, 0, -1, -2, -2, -2, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 3, 2, 3, 2, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 3, 2, 3, 2, 2, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 4, 4, 3, 2, 2, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 2, 3, 3, 3, 4, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 3, 3, 3, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 3, 3, 2, 3, 2, 2, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 3, 3, 1, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 1, 2, 1, 1, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 2, 2, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 2, 2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 2, 2, 2, 1, 2, 1, 2, 1, 1, 1, 1, 3, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 2, 3, 1, 1, 1, 2, 2, 1, 2, 2, 2, 2, 4, 2, 3, 0, 0, -2, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 2, 2, 2, 1, 0, -1, -1, -2, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 1, 1, 2, 1, 1, 0, 0, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 1, 0, 1, 1, 1, 1, 1, 1, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 1, 1, 2, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -3, -1, -1, -2, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -2, 0, -1, -1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -2, -1, -2, 0, 0, 0, 0, 1, 1, 1, 2, 2, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 1, 2, 1, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 1, 1, 2, 2, 2, 1, 1, 1, -1, -1, -2, -2, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 2, 3, 2, 2, 1, 0, -1, -2, -1, -1, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 2, 1, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 2, 2, 1, 1, 0, 0, -1, -2, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, -1, -2, -2, -2, -1, 0, 0, 1, 1, 1, 1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, -2, -1, -1, -2, -1, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, -2, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, -2, -2, -1, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, -1, -1, -3, -1, -2, -1, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -2, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 1, 1, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 1, 2, 1, 2, 2, 2, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 1, 1, 1, 0, 1, 1, 1, 1, 1, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 2, 2, 1, 2, 2, 1, 1, 3, 2, 3, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 1, 1, 2, 0, 1, 1, 2, 1, 2, 3, 2, 2, 2, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 2, 3, 2, 0, 1, 1, 1, 1, 0, 0, 1, 0, 2, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, -2, -1, 0, 1, 2, 3, 4, 4, 3, 2, 1, 1, 1, 2, 2, 1, 1, 3, 2, 0, 0, 3, 1, 0, -1, -2, -1, -1, 0, -1, 0, -2, -2, -1, 0, 2, 1, 3, 3, 2, 2, 2, 1, 1, 2, 1, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, -1, 0, -2, -1, 0, 0, -1, -1, -1, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, -1, -1, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, -1, -2, 0, 1, 0, -1, -1, -1, 0, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 1, 0, -1, -2, -1, -1, -1, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 2, 1, -1, -1, 0, 1, 0, 0, -2, -2, -1, 0, 0, 0, -1, -2, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -2, -2, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -3, -2, -3, 0, 0, 0, 0, 2, 0, 0, 1, 2, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, -3, -3, -5, -4, -1, 0, 0, 0, 0, 2, 1, 1, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -4, -5, -5, -3, -3, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -5, -6, -5, -5, -2, -1, 0, 1, 1, 0, 0, 1, 1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, -2, -4, -4, -5, -6, -4, -2, 0, 1, 1, 2, 0, 0, 1, 1, 0, -1, 0, 1, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, -2, -1, 0, -2, -3, -6, -7, -5, -3, -2, 2, 4, 4, 3, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -3, -4, -6, -5, -3, 0, 2, 5, 6, 5, 3, 2, 0, 0, 0, -1, 0, 0, 0, -1, -2, -1, 0, 0, 1, 0, 1, 0, -1, 0, 0, -2, -2, -5, -6, -5, -3, -1, 2, 4, 5, 4, 2, 0, 0, 0, 0, -1, 0, 1, 0, -1, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -3, -5, -6, -5, -5, -1, 1, 4, 5, 5, 2, 1, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -2, -4, -5, -6, -4, -1, 1, 2, 3, 4, 2, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, -4, -4, -4, -4, -2, 0, 0, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, -1, -1, -4, -4, -6, -3, -4, -1, -1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, -1, -3, -2, -2, -5, -4, -3, -3, -1, 0, 1, 1, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, -4, -3, -2, -4, -3, -2, 0, -1, 0, 0, 1, 2, 0, 1, 0, -1, 0, 0, 1, 1, 0, 1, -1, -1, 0, 0, 0, 0, -1, -1, 0, -2, -3, -3, -2, -2, -3, -2, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -2, -2, -2, -3, -2, 0, -2, -2, -1, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, -2, -1, -2, -1, -2, 0, 0, -2, 0, -1, -1, 0, -2, -3, -1, 0, 0, 0, 0, -2, -1, 0, 1, 0, -1, -3, -1, -1, 0, 0, -1, -2, -2, -2, -2, -1, -1, -1, 0, 0, -1, 0, -1, 0, -2, -1, -2, -2, 0, 0, 0, -1, 0, 1, 0, 0, 0, -3, -1, -1, 0, 0, -2, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, -1, -1, -2, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -2, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 1, 2, 1, 1, 2, 1, 0, 1, 0, -1, 0, 0, 1, 1, 0, 1, 1, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 3, 3, 2, 3, 3, 2, 2, 2, 1, 1, 1, 1, 2, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 1, 1, 2, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 2, 1, 0, 0, 0, 0, -1, 0, -1, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 2, 1, 1, 2, 0, 0, 0, -2, -2, -1, -3, -2, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 1, 0, 0, -2, -2, -2, -4, -3, -3, -2, -1, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 2, 1, 1, 0, 0, -1, -2, -3, -3, -3, -3, -3, -2, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, 0, -2, -2, -3, -2, -2, -3, -2, -2, -1, 0, 1, 2, 1, 0, 1, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 1, 2, 1, 1, 1, 0, -1, -2, -2, -2, -2, -2, -3, -3, 0, 0, 0, 1, 2, 1, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 1, 0, 1, 0, -1, -2, -3, -4, -4, -3, -1, -1, 0, 1, 1, 3, 1, 2, 1, 0, 2, 2, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, -1, -2, -2, -1, -3, -3, -2, -3, 0, 0, 1, 1, 3, 2, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 2, 1, 0, 1, 0, -1, -2, -2, -3, -2, -3, -2, -1, -1, 0, 0, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -2, -2, -2, -3, -3, -3, -2, 0, 0, 1, 3, 3, 2, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, -2, -2, -2, -3, -2, -1, -2, 0, 0, 0, 1, 2, 1, 0, 1, 0, 0, 1, 0, 0, -1, -1, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, -2, -1, -1, -2, -2, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, -1, -2, -1, -1, -1, -3, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 2, 0, 0, 0, 0, 0, -1, 0, -2, -2, -2, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, -1, -2, -2, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -2, -2, -1, -1, -2, 0, 0, -1, 0, -1, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -2, -1, -1, -1, 0, -1, -2, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 2, 1, 1, 3, 3, 1, 1, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 2, 2, 0, 0, 0, 1, 1, 2, 1, 2, 2, 3, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 1, 0, 0, 0, 1, 2, 3, 0, 2, 1, 2, 2, 0, 0, 0, 0, -1, -1, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 2, 0, 0, 1, 0, 1, 0, 1, 1, 2, 2, 1, 1, 2, 1, 2, 1, 0, 0, -1, -3, 0, 0, -1, -1, 0, -2, -1, -1, -1, 0, 2, 2, 0, 0, 0, 0, 1, 0, 2, 1, 1, 1, 1, 2, 3, 1, 1, 1, 1, 0, -3, -3, -1, 0, -1, -1, 0, -3, -2, -1, -2, 0, 1, 3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 3, 1, 0, 1, 0, -1, -2, -4, -3, -2, -3, -1, -1, -1, -3, -2, -1, -1, 2, 2, 0, -1, 1, 0, 2, 0, 0, 0, 0, 1, 0, 1, 3, 0, 0, 0, 0, -3, -3, -4, -3, -3, -3, -2, -2, -2, -2, -1, -2, -2, 0, 2, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 3, 2, 1, 0, -1, -1, -1, -3, -2, -3, -3, -3, -1, -3, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, -2, 0, 0, 0, -2, -2, -2, -3, -2, 0, 0, -1, 0, 1, -2, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, -2, -1, -1, 0, -1, -1, -1, -2, -2, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 2, 1, 0, 1, 1, 0, 0, -1, 1, 0, -2, -2, -2, 0, 0, 0, 0, -1, -1, -2, -2, 1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 2, 1, 0, -1, 0, 1, 1, 0, 0, 0, 0, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 1, 0, -1, -2, -2, -2, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 2, 0, -2, -2, -2, -1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, -2, -2, -3, -2, -1, 0, 0, 1, 2, 0, 1, -1, 0, 0, -1, 0, 0, 0, -3, 0, 0, 0, 0, 1, 0, 0, 0, 2, 1, 2, 2, 0, -1, -4, -3, -3, -1, 0, 1, 1, 3, 2, 0, -1, 0, 1, 0, 0, 0, 1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 3, 0, 1, 0, -1, -3, -4, -3, -3, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 2, 3, 2, 1, 1, -1, -2, -2, -3, -2, -4, -2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, -2, -1, 0, 0, 0, 1, 0, 2, 3, 2, 1, 0, -1, -2, -1, -3, -1, -1, -3, -1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, -1, -3, 0, 0, -1, -1, -2, -1, 0, -1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, -1, -2, 2, 0, -1, -2, -1, 0, -1, -2, -1, 0, -2, -3, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 2, 2, 0, 1, 0, 1, 1, 1, 0, 0, 2, 0, -2, -2, -1, -1, -1, -3, -1, -1, -3, -2, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 4, 2, 0, 1, 0, 1, 2, 2, 1, 1, 2, 0, -3, -2, -1, -2, -2, -2, -2, -1, -1, -2, 0, -1, 0, 0, 0, -1, -1, 1, 0, 0, 3, 3, 0, 0, 1, 0, 1, 2, 3, 1, 2, 0, -2, -2, 0, -1, -2, -1, -2, 0, -3, -2, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 3, 2, 0, -1, 0, 1, 2, 3, 4, 3, 3, 2, -1, -1, 0, -2, -1, -1, -1, 0, -2, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 4, 2, 0, 0, 2, 2, 2, 2, 4, 4, 3, 3, 0, 0, -1, -1, -2, -1, 0, -1, 0, -1, 0, 0, -1, 0, 1, 0, -1, 1, 0, 0, 4, 0, 0, 0, 2, 3, 1, 2, 5, 4, 5, 3, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 1, 3, 3, 4, 3, 3, 3, 3, 2, 2, 0, 0, 0, 0, 0, -1, 0, 0, 2, 1, 0, 0, 1, 0, -1, 1, 1, 0, 1, 0, 0, 1, 1, 1, 3, 4, 4, 2, 1, 3, 3, 2, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 2, 1, 1, 0, 1, 2, 4, 3, 1, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 2, 2, 0, 0, -1, 0, 0, 0, 0, 2, 2, 2, 0, 0, 1, 0, 0, 0, -1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 2, 1, 1, 1, 0, 0, 1, 0, 1, 1, 1, 1, 1, 1, 2, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, -1, -1, 0, 0, 2, 1, 2, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, -2, -1, 0, 0, 0, 1, 2, 1, 2, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, -1, -1, -1, 0, -1, -2, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 2, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 1, 0, -1, 0, 0, 0, 2, 2, 1, 1, 2, 2, 2, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 1, 0, 1, 1, 0, 1, 2, 1, 2, 3, 2, 2, 2, 2, 1, 0, 1, 1, 1, 1, 2, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 1, 0, 1, 2, 2, 2, 4, 3, 3, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 2, 2, 2, 3, 5, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 2, 1, 3, 3, 3, 3, 2, 2, -1, 0, -1, 0, 0, -1, -1, -1, -2, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 1, 1, 1, 1, 0, 1, 3, 2, 2, 1, 1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -2, -1, 0, 1, 1, 1, 1, 0, 2, 2, 3, 1, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -1, -1, 0, 0, 1, 0, 0, 0, 2, 3, 3, 0, 0, 0, -1, -2, 0, 0, 0, 1, 0, 0, -1, 0, 0, -2, -1, 0, 1, 0, 0, -1, -2, -1, 0, 1, 1, 2, 1, 2, 2, 4, 2, 1, 0, -1, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, -1, -1, 0, 0, 0, 1, 2, 2, 2, 2, 2, 3, 4, 1, 0, 0, -2, -2, 0, 0, 0, 1, 0, -1, -1, -1, 0, -2, -1, -2, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 2, 3, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 1, 1, 0, 0, -1, 0, 0, 0, 1, 1, 2, 2, 1, 3, 3, 2, 0, 0, 0, 0, 0, 1, 1, 1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 2, 3, 1, 2, 1, 1, 2, 2, 1, 0, 0, 0, 0, 1, 1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 3, 1, 0, 1, 1, 1, 1, 0, 1, 1, 3, 2, 2, 2, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -2, -1, 0, 0, 1, 1, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 1, 0, -2, -1, 0, 0, 1, 0, 1, 1, 1, 0, 1, 1, 1, 2, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 1, 2, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 2, 2, 3, 2, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 2, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, 2, 1, 2, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, -1, -1, -2, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 2, 0, 1, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 2, 2, 1, 2, 2, 2, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 1, 1, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -2, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 2, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 1, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, -1, 0, 1, 0, -1, 0, 1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 2, 1, 2, 1, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 0, 2, 1, 2, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 1, 2, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, -1, -1, -2, -3, -2, -3, -2, -2, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, -3, -2, -4, -3, -2, -3, -2, -2, 0, 0, 0, 0, 2, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 0, 0, -1, -3, -3, -4, -3, -4, -3, -2, -2, 0, 0, 0, 2, 0, 2, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 2, 1, 2, 2, 2, 0, 0, 0, -1, -2, -2, -4, -3, -2, -1, -1, 0, 1, 2, 1, 2, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 3, 1, 2, 1, 1, -1, -2, -2, -2, -3, -3, -3, -2, 0, 0, 0, 0, 1, 1, 2, 2, 1, 1, 2, 1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 1, 0, 0, -2, -1, -2, -2, -2, -3, -2, -2, -1, 0, 1, 2, 3, 2, 3, 1, 2, 0, 1, 1, 0, 0, 0, -1, 1, 0, 1, 2, 1, 1, 1, 0, -1, -2, -2, -2, -3, -2, -1, -2, 0, -1, 1, 2, 3, 2, 3, 2, 2, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -3, -2, -3, -2, -2, -2, -1, 0, 1, 1, 2, 3, 3, 3, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -1, -2, -2, -1, -2, -1, -1, 0, 0, 1, 1, 3, 2, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -2, -2, -1, -2, -2, -1, -2, 0, 0, 0, 2, 2, 3, 3, 2, 2, 2, 0, 1, 1, 0, 0, 0, 1, 1, 2, 2, 0, 1, 0, 0, 0, -1, -2, -1, -3, -2, 0, -1, 0, 0, 0, 2, 1, 3, 3, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 2, 1, 0, 0, 0, -1, -1, -2, -1, -2, -2, 0, 0, 0, 1, 1, 1, 2, 2, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 0, 0, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 1, 1, 1, 0, 1, 1, 2, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 4, 4, 3, 3, 1, 2, 1, 2, 2, 0, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -2, -1, -1, 0, 2, 3, 5, 3, 3, 2, 2, 0, 1, 1, 0, 0, 1, 1, 1, 2, 1, 1, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, -2, -1, -1, 0, 0, 3, 4, 3, 4, 2, 2, 1, 0, 1, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, -2, -1, -1, -3, -1, 0, 0, 0, 1, 2, 1, 3, 3, 1, 1, 2, 1, 1, 1, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, -2, -3, -2, -3, -2, -1, 0, 1, 0, 1, 2, 0, 1, 2, 0, 1, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -3, -2, -2, -2, -1, -2, -3, -1, -1, 0, 1, 1, 2, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 2, 0, 0, 0, 0, -1, -3, -2, -3, -2, -1, -1, -1, -2, -1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, 0, 0, 0, 0, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -2, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 2, 1, 0, 0, 0, -1, -1, -2, -1, 0, 0, 1, 1, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 2, 2, 2, 3, 1, 2, 0, 0, -2, -2, -1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 3, 1, 1, 1, 2, 1, -2, -3, -3, -3, -2, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 2, 1, 1, 1, 2, 1, 0, -1, -3, -5, -4, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, -1, -2, -2, 0, 0, 0, 2, 0, 0, 0, 1, 1, 2, 0, -3, -3, -4, -2, 0, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -2, -1, -3, -1, 0, 0, 1, 2, 0, 0, 0, 1, 0, -1, -3, -4, -4, -1, 0, 2, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -3, -2, -2, -3, -1, 0, 1, 1, 1, 0, 2, 1, 1, -1, -3, -4, -4, -3, 0, 1, 2, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -1, -1, 0, 1, 0, 1, 1, 2, 2, 1, 0, -4, -4, -4, -2, 0, 0, 1, 3, 0, 0, -2, -2, -1, -1, -2, 0, 0, 0, -2, -1, 0, -2, 0, 0, 0, 0, 1, 1, 1, 2, 0, -1, -3, -5, -3, -2, 0, 0, 0, 2, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 1, 1, 0, 1, 1, 0, 0, -2, -2, -4, -4, -2, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, -2, -2, 0, 2, 2, 2, 2, 1, 1, 1, 0, -1, -2, -2, -3, -2, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, -2, -1, -2, -1, 0, 2, 1, 2, 3, 0, 0, 0, 0, -1, -2, -2, -3, -1, 0, 1, 0, 2, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -2, -1, 0, 2, 1, 1, 1, 0, -1, 0, 0, -1, -2, 0, 0, 0, 1, 1, 1, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -3, -1, -2, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, -3, -2, -2, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, -1, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -2, -2, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, -3, -2, -2, -1, -2, -2, -1, -1, -2, -1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 2, 0, 0, 0, 0, 0, -2, -3, -1, -1, -2, -1, -2, -2, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 1, 1, 1, 2, 1, 1, 0, 1, 0, 0, 0, 1, 3, 2, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 2, 2, 2, 3, 2, 2, 1, 3, 4, 3, 4, 4, 5, 4, 3, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 2, 3, 3, 3, 3, 2, 2, 2, 4, 2, 3, 3, 4, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -3, -2, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -3, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -2, -1, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, -1, -1, -3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, 0, -1, 0, 0, 0, 0, -1, -2, -1, -1, -1, -3, -1, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, -2, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -2, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, -1, -1, -2, -2, -2, -3, -2, -2, -2, 0, -1, -1, 0, 0, 0, -1, -1, -1, -2, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -2, -2, -1, -2, -3, -2, 0, 0, -2, 0, -1, -1, -1, 0, -1, 0, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -3, -3, -2, -1, -2, -2, -2, -1, -2, -1, -1, 0, -1, -1, -1, -1, -2, -1, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, -1, 0, 0, -2, -2, -2, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 2, 1, 1, 1, 0, 1, 0, 0, -1, -1, 0, 0, -2, -2, -1, -1, -2, 0, -1, -1, 0, -1, 0, -1, -2, -1, -2, -1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, 0, 0, 0, -1, -1, -1, -1, -2, 0, 0, 0, -1, -1, -1, -2, -3, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, -1, -1, 0, 0, -1, -1, -1, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, -1, -2, -1, -2, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, -2, -1, -1, -1, -1, -1, -1, 0, 0, 0, -2, -1, -1, 0, -1, -1, -1, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, -1, -1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, -2, -1, -1, -1, -1, -1, 0, 0, -1, 0, -1, -1, -1, -2, -2, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, -2, -1, -1, -1, -1, -1, -1, 0, -1, 0, 0, -1, 0, -1, -2, -1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -2, -2, -2, -1, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, -1, 0, 1, 1, 0, 0, 0, 0, -1, -2, -2, -2, -1, -1, 0, 0, -1, -2, -2, -2, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, -2, -1, -2, -1, -1, -1, -2, -1, -2, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, -2, -1, -1, -2, -1, -2, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, -1, -1, -2, -1, 0, 0, -1, -1, -1, -1, -2, 0, -2, -1, 0, -1, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -2, -1, -2, 0, -1, -2, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -2, -1, 0, 0, 2, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -3, -2, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 3, 3, 1, 2, 1, 0, 0, 1, 0, -1, 0, -1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, -2, 0, 1, 2, 2, 3, 3, 1, 1, 1, 0, -1, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -1, -1, 0, 3, 3, 2, 1, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, -2, 0, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, -2, 0, 2, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, -2, -2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 1, 2, 1, 0, 1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 2, 1, 2, 2, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 2, 1, 2, 2, 1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 2, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 2, 0, 1, 0, 0, 0, 1, 2, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 2, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 0, 0, -1, 0, 1, 1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -2, 0, 0, 1, 1, 0, 0, -1, 0, 0, 2, 0, 0, -1, 0, 1, 1, 1, 0, 0, -2, -2, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, -2, 2, 2, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 2, 2, 2, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -1, 0, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 2, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 2, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -3, 0, 3, 3, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -2, -2, -2, 1, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -3, -1, 2, 3, 3, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -2, -3, -1, 0, 4, 4, 1, 0, 1, 0, 0, 1, 1, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, -1, -1, -3, 0, 0, 3, 2, 2, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, -1, 0, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 2, 2, 2, 1, 0, 2, 1, 2, 1, 2, 1, 1, 0, 1, 2, 0, 0, -2, -1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 3, 3, 2, 4, 3, 4, 3, 2, 1, 2, 2, 1, 1, 1, 1, 1, 0, 1, 1, 1, 0, -2, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 2, 2, 3, 2, 3, 1, 3, 2, 0, 1, 2, 1, 1, 0, 1, 0, 1, 1, 0, -1, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 2, 3, 3, 2, 2, 1, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 3, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, -2, -2, -1, 0, 0, 0, 0, 0, 2, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, -2, 0, 0, -1, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, -2, -1, -1, -1, -2, -1, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -2, -1, -2, -3, -2, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -2, -2, -3, -2, -3, -4, -3, -2, -1, 0, 0, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, -3, -3, -5, -4, -5, -3, -3, -2, 0, 0, 2, 2, 1, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -2, -2, -2, -3, -4, -5, -4, -3, -3, -1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, -2, -2, -3, -4, -5, -5, -5, -3, -3, -1, 0, 1, 2, 3, 0, 2, 1, 0, 0, 1, 1, 0, 0, 0, 0, 2, 1, 2, 0, 1, -1, -2, -2, -3, -3, -3, -4, -5, -5, -4, -2, -1, 0, 2, 3, 2, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 2, 2, 0, 0, 0, -1, -1, -3, -3, -6, -6, -5, -3, -2, 1, 3, 5, 4, 4, 3, 1, 1, 0, 0, 1, 1, 0, -1, 0, 0, 1, 1, 2, 0, 0, 0, -2, -2, -3, -4, -3, -4, -6, -4, -3, -1, 1, 5, 6, 6, 4, 4, 1, 0, 0, 1, 3, 1, 0, 0, -1, -1, 0, 1, 1, 0, 0, 0, 0, -1, -3, -3, -4, -4, -6, -5, -2, 0, 2, 4, 6, 6, 5, 4, 1, 0, 0, 0, 2, 1, 0, -1, -1, 0, 0, 0, 2, 0, 0, 0, -2, -1, -1, -2, -5, -4, -5, -6, -4, -2, 1, 5, 5, 5, 4, 3, 2, 1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, -2, -3, -4, -6, -5, -6, -5, -2, 0, 3, 4, 4, 4, 2, 1, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, -2, -2, -3, -4, -5, -5, -6, -5, -2, 0, 2, 3, 4, 2, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -3, -4, -4, -4, -5, -5, -3, -2, -1, 1, 3, 3, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -3, -4, -4, -4, -4, -3, -3, -1, 0, 1, 2, 2, 2, 1, 1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -3, -4, -3, -2, -3, -2, -1, 0, 1, 2, 3, 3, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -2, -3, -2, -4, -2, -3, -2, -1, 0, 0, 0, 0, 2, 2, 2, 2, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, -1, -2, -2, -2, -3, -3, -3, -1, -2, -1, 0, 0, 1, 1, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, -2, -1, -2, -3, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 1, 0, -2, -1, 0, 0, 0, 0, -2, -3, -2, -2, -3, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -2, -1, 0, 0, 0, -2, -2, -1, -1, -2, -1, 0, 0, 1, 1, 0, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 1, 2, 0, -1, -2, -2, 0, 0, 0, -1, -2, -2, -2, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, 0, 0, 0, -1, -1, -3, 0, 0, 0, 0, 0, 1, 1, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 3, 3, 4, 3, 1, 1, 0, 1, 0, 1, 1, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 2, 1, 1, 1, 1, 2, 0, 2, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 2, 0, 1, 1, 1, 2, 0, 1, 0, 0, 0, 1, 1, 0, 0, 2, 1, 2, 2, 2, 2, 2, 3, 1, 0, 2, 1, 1, 2, 1, 0, 2, 1, 0, 0, 1, 1, 2, 0, 0, 0, 1, 0, 0, 0, 0, -1, 2, 2, 3, 2, 3, 0, 1, 4, 2, 0, 2, 0, 0, 2, 1, 0, 1, 2, 0, 0, 1, 0, 1, 0, -1, 0, 1, 0, 0, -1, 0, 0, 1, 2, 2, 3, 3, 1, 2, 1, 2, 1, 2, 1, 0, 1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, -1, 0, 0, 1, 2, 2, 3, 0, 2, 2, 2, 2, 1, 2, 2, 1, 0, -1, -1, 1, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, 1, 0, -1, -1, 0, 1, 1, 2, 2, 2, 1, 2, 2, 1, 1, 3, 2, 2, 0, -3, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 2, 2, 1, 0, 0, 1, 0, 2, 1, 2, 1, 2, 0, 0, -3, -2, -1, -3, -3, -1, -1, -1, 0, -1, -2, 0, 1, 1, 0, -1, 0, -1, 2, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, -1, -1, -1, -1, -1, -3, -1, -1, -1, -1, -1, -2, -2, -1, 0, 0, -2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 3, 2, 0, 0, 0, -1, -2, -2, 0, -2, -3, -2, -2, -2, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 2, 2, 1, 0, 0, -1, 0, -1, 0, -1, -1, -2, 0, -1, -1, 0, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 3, 0, 0, 2, 1, 0, 2, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, -2, 0, 1, 0, -1, 0, -1, -1, 0, 0, -1, 2, 3, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, -2, -1, 0, 0, 0, 1, 2, 1, -1, 0, 1, 2, 1, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, -2, 0, 0, -1, 0, 0, -1, 1, 2, 1, 0, 0, 1, 1, 2, 1, 0, -1, -2, -1, -1, 0, 1, 2, 1, 2, 1, 0, -1, 1, 1, 0, 0, -1, 0, -2, 0, 0, 0, 2, 4, 2, 0, 0, 0, 1, 1, 1, 0, -2, -3, -1, -1, 0, 2, 1, 1, 2, 0, 0, -1, 1, 0, 0, -1, 0, 0, -2, -1, 0, 0, 2, 2, 3, 0, 0, 1, 1, 1, 1, 0, -2, -4, -1, 0, 0, 2, 1, 2, 2, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 1, 3, 2, 0, 1, 2, 1, 1, 0, 0, -2, -3, -2, 0, 0, 2, 3, 3, 2, 1, 0, -1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 1, 1, 2, 2, 1, 2, 1, 1, 0, 0, -2, -3, -1, 0, 0, 2, 1, 3, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 1, 3, 2, 2, 0, -2, -2, -4, -2, -1, 0, 1, 2, 3, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 1, 0, 0, 2, 2, 3, 2, 0, -2, -1, -1, -3, -1, 0, 0, 1, 1, 2, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 2, 1, 2, 3, 2, 2, 2, 0, -2, -1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, -1, 0, 0, 0, 0, -2, 0, -1, 2, 3, 1, 2, 1, 1, 2, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -2, -1, 0, -2, -1, 0, 0, 0, 0, -2, 0, 0, 3, 2, 2, 1, 1, 2, 2, 1, -1, 0, 2, 0, -1, -2, 0, 0, 0, -1, -1, 0, -3, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 4, 3, 1, 0, 1, 1, 1, 1, 1, 0, 2, 0, -1, -1, -1, 0, 0, -1, -1, -2, -2, -1, 0, -1, 0, 0, -1, 0, -1, -1, -1, -1, 5, 3, 1, 0, 1, 2, 0, 2, 1, 0, 0, 0, 0, -2, -1, -1, -1, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 6, 2, 0, 1, 1, 2, 1, 1, 2, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, -3, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 5, 2, 0, 1, 1, 0, 1, 3, 3, 1, 2, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, -2, -2, 0, 0, 4, 0, 0, 1, 2, 2, 0, 2, 3, 3, 3, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 3, 1, 0, 1, 2, 2, 2, 4, 3, 2, 3, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, -2, -1, 0, 0, 4, 2, 1, 1, 2, 2, 3, 4, 2, 1, 2, 2, 2, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 3, 2, 2, 2, 0, 2, 3, 4, 4, 2, 1, 1, 0, 1, 1, 0, 1, 1, 2, 1, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 3, 1, 2, 1, 3, 2, 3, 1, 3, 2, 1, 2, 3, 3, 2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 2, 1, 1, 1, 0, 0, 1, 1, 1, 1, 0, 0, 1, 1, 1, 3, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 2, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 3, 2, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 2, 1, 3, 2, 1, 1, 3, 3, 2, 0, 0, 1, 1, 0, -1, -1, 1, 1, 0, -1, -1, -1, -1, 0, 0, 1, 1, 1, 0, 2, 2, 1, 2, 1, 1, 2, 1, 2, 2, 2, 1, 0, 1, 0, 2, 0, -2, -2, -1, 0, 0, -2, -2, -2, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 2, 3, 3, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 2, 1, 2, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, -2, -2, -1, 0, 1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -2, 0, 1, 2, 3, 2, 2, 2, 1, 1, 0, 0, 0, 1, 0, 2, 2, 3, 2, 2, 2, 1, 1, 2, 1, 3, 1, 2, 2, 0, 0, 0, 0, 0, 2, 2, 4, 3, 2, 2, 3, 2, 2, 1, 0, 0, 0, 1, 2, 4, 4, 2, 2, 2, 3, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 2, 1, 3, 3, 2, 4, 3, 5, 3, 2, 0, 0, 0, 1, 2, 2, 3, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 1, 2, 2, 3, 2, 3, 4, 4, 2, 0, 0, 0, 0, 0, 0, 1, 0, -2, 0, 0, 1, 1, 1, 0, 0, -1, -1, 0, -1, 0, 0, 2, 2, 3, 2, 2, 4, 2, 4, 3, 2, 1, 1, 0, 1, 1, 2, 3, 1, 0, -1, 0, 0, 2, 2, 1, 0, 1, 0, 0, -2, 1, 2, 2, 1, 3, 3, 4, 2, 3, 1, 2, 0, 0, 0, -1, 0, 2, 2, 4, 5, 2, 1, 0, 0, 1, 2, 2, 2, 1, 2, 0, -1, 0, 1, 2, 1, 3, 3, 5, 4, 2, 0, 0, -1, -2, -2, -2, 0, 0, 3, 4, 5, 4, 2, 1, 0, 0, 0, 1, 1, 1, 1, 0, -2, 0, 1, 1, 0, 1, 2, 3, 4, 1, 2, 1, 0, 0, -1, 0, -1, 1, 2, 3, 3, 2, 2, 0, 1, 0, 0, 0, 0, 2, 1, 0, -1, -1, 2, 1, 1, 2, 2, 2, 1, 2, 2, 1, 0, -1, -2, -1, -1, 0, 1, 1, 1, 3, 2, 1, 0, 0, 0, 0, 0, 2, 2, 0, -1, 0, 0, 0, 1, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 2, 1, 1, 1, 1, 1, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, 0, 0, 0, 0, 0, 0, 2, 0, 1, 2, 3, 2, 1, 3, 1, 2, 3, 2, 2, 4, 3, 3, 2, 1, 0, 0, 0, 1, 0, -2, -3, -2, -1, -1, 0, 0, 1, 1, 1, 0, 0, 0, 3, 4, 3, 3, 3, 2, 4, 4, 4, 4, 4, 3, 3, 1, 2, 2, 1, 2, 1, -1, -2, -1, -1, -1, -1, 1, 0, 0, 2, 1, 2, 1, 0, 1, 3, 3, 2, 4, 4, 3, 5, 5, 3, 2, 3, 2, 1, 0, 1, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 2, 0, 3, 2, 2, 2, 1, 1, 2, 2, 3, 1, 1, 2, 2, 3, 2, 2, 1, 1, 1, 2, 2, 0, -1, -2, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 3, 1, 2, 1, 2, 2, 1, 1, 1, 1, 1, 2, 1, 1, 1, 1, 0, 2, 0, -1, -2, 0, 0, 0, 0, -1, 0, 0, 1, 2, 2, 3, 1, 1, 2, 1, 0, 1, 1, 2, 2, 1, 1, 2, 2, 2, 1, 1, 0, 0, 0, -1, -3, -1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 0, 1, 0, 1, 0, 1, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, -2, 0, 0, 0, 0, 0, -1, 0, 1, 2, 1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 2, 1, 1, 1, 2, 1, 1, 3, 2, 3, 3, 2, 2, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 2, 2, 1, 1, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 2, 2, 2, 1, 2, 1, 0, 0, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 2, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 2, 1, 1, 2, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -1, 0, -1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, -1, -1, -1, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 2, 2, 1, 2, 2, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 1, 1, 1, 2, 0, 1, 0, 1, 0, 2, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 2, 2, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 1, 0, 1, 1, 1, 1, 0, 0, 1, 2, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 1, 0, 1, 1, 1, 1, 1, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 3, 2, 4, 3, 2, 2, 1, 2, 2, 1, 1, 2, 2, 1, 1, 2, 0, 0, -1, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 3, 4, 3, 4, 2, 1, 2, 1, 1, 0, 0, 0, 0, 0, 1, 3, 1, 0, -2, -1, -2, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 2, 2, 2, 2, 2, 1, 1, 1, 2, 1, 0, -1, 0, 0, 0, 2, 1, 0, -1, -1, -2, -1, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, 0, 1, 2, 2, 3, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, -1, -2, -2, -1, -2, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -2, -2, -1, -1, 0, 0, 0, 0, 1, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, -1, -1, -1, 0, 0, -2, -2, -2, -1, -1, 0, 0, 0, 1, 0, 1, 2, 2, 1, 1, 2, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -2, -3, -4, -2, -1, -2, 0, 0, 0, 0, 2, 2, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, -4, -3, -2, -2, -3, -2, -1, 0, 0, 1, 1, 3, 3, 1, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -4, -4, -4, -5, -5, -2, -3, 0, 0, 0, 0, 1, 3, 2, 2, 0, 0, 0, 1, 1, 0, 0, 0, 2, 2, 1, 0, 0, 0, -1, -2, -3, -4, -4, -5, -6, -5, -4, -5, -3, -2, 0, 0, 2, 2, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, -1, -1, -2, -3, -4, -5, -5, -5, -5, -5, -5, -4, -1, 0, 2, 2, 3, 3, 2, 0, 0, 0, 0, 0, 1, 0, 0, 3, 2, 1, 2, 1, 0, -1, -2, -4, -4, -5, -4, -6, -6, -7, -6, -3, -2, 0, 4, 4, 4, 3, 2, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 1, 1, 0, -2, -3, -4, -3, -4, -5, -4, -4, -5, -5, -2, -1, 1, 4, 6, 5, 5, 2, 0, 0, 2, 1, 1, 0, -1, 0, 0, 3, 3, 1, 2, 0, -2, -3, -3, -5, -4, -4, -3, -5, -6, -3, -2, 0, 3, 7, 8, 8, 6, 3, 2, 1, 2, 2, 1, 1, -1, 0, 0, 2, 2, 1, 1, 0, -1, -2, -3, -4, -4, -4, -4, -4, -5, -4, 0, 0, 3, 8, 8, 8, 6, 3, 2, 1, 1, 2, 1, 1, 0, 1, 0, 1, 3, 2, 2, 0, -2, -1, -3, -4, -3, -4, -4, -5, -5, -4, -3, 1, 3, 6, 7, 7, 6, 3, 0, 0, 1, 2, 1, 1, 0, 0, 1, 2, 2, 1, 1, -1, -1, -2, -3, -5, -4, -4, -5, -6, -7, -5, -3, 0, 3, 4, 7, 7, 5, 3, 0, 0, 0, 2, 2, 1, -1, 1, 1, 2, 1, 2, 0, 0, -1, -1, -2, -3, -5, -4, -4, -5, -6, -5, -3, 0, 2, 4, 5, 6, 5, 3, 0, 0, 1, 2, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, -2, -3, -3, -3, -3, -5, -6, -5, -6, -5, -3, -2, 2, 3, 5, 4, 5, 2, 1, 0, 1, 2, 2, 1, 0, 1, 2, 2, 1, 0, 0, 0, -1, -1, -3, -3, -4, -5, -4, -5, -6, -4, -3, -1, 1, 4, 4, 5, 4, 2, 0, 0, 1, 2, 2, 0, 0, 0, 3, 0, 0, 0, 0, -1, -1, -1, -3, -3, -5, -6, -5, -5, -4, -2, 0, 0, 1, 3, 3, 5, 5, 2, 0, 0, 0, 1, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, -2, -3, -4, -3, -5, -6, -4, -2, -3, -1, 0, 1, 3, 4, 4, 5, 4, 1, 1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, -1, -1, -2, -3, -4, -3, -3, -3, -2, -2, 0, 0, 0, 1, 2, 4, 4, 3, 2, 0, 1, 0, 0, 2, 1, 0, -1, 1, 0, 0, 0, 0, -1, -3, -4, -3, -4, -2, -2, -3, -1, 0, -1, 0, 1, 1, 2, 1, 1, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -3, -4, -3, -2, -2, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -3, -3, -2, -2, -1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, -1, -1, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -3, -2, -2, -1, -2, -1, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -2, -2, -2, -3, -1, -2, -1, 0, 0, 1, 1, 1, 2, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, -1, -1, -2, 0, -1, 0, 0, 0, 0, 1, 2, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, -1, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 3, 3, 3, 2, 2, 2, 1, 2, 1, 1, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 2, 0, 2, 1, 0, 1, 0, 0, 1, 2, 1, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 1, 1, 1, 0, 0, 0, -2, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -2, -2, -1, -3, -2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -3, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -2, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -2, -2, -1, -2, 0, 0, -2, -1, -1, 0, 0, 0, -1, -1, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -2, -3, -2, -4, -2, -3, 0, -1, -2, -2, -2, -2, -1, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, -2, -2, -3, -3, -5, -4, -4, -1, -2, -1, -2, -2, -2, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 1, 2, 1, 0, 0, 1, 0, 0, 0, -3, -4, -4, -3, -4, -4, -4, -2, -2, -3, -2, -2, -2, -2, -2, -1, -1, -1, 0, 0, 2, 0, 1, 0, 1, 1, 0, 1, 0, 1, 0, 0, -3, -4, -5, -2, -4, -3, -4, -2, -2, -2, -2, 0, -1, -2, -1, -2, -2, -1, 0, 0, 2, 0, 0, 1, 1, 4, 0, 0, 0, 0, -1, 0, -2, -3, -4, -2, -2, -4, -4, -3, -3, -3, -3, -2, -1, -1, -1, -3, -2, 0, 0, 0, 1, 1, 1, 0, 1, 3, 1, 0, 0, 0, -2, -1, -2, -3, -4, -3, -3, -2, -4, -3, -2, -3, -2, -1, -1, -1, -2, -3, -3, 0, 0, 0, 2, 1, 1, 0, 0, 2, 2, 1, 0, -1, -1, 0, -1, -2, -2, -2, -1, -3, -3, -3, -2, -1, -2, -1, 0, -2, -1, -2, -1, -1, 1, 0, 1, 3, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -2, -2, -2, -1, -2, -2, -3, -2, -2, -1, 0, -1, -1, -1, -1, 0, 0, -1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, -1, -2, -1, -2, 0, -2, 0, -1, -1, -1, -2, -3, -1, 0, -1, -2, -2, -2, -2, -2, 0, -1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, -2, -1, -1, -1, -1, -1, -1, 0, -1, 0, -3, -1, -2, 0, -1, -3, -3, -2, -2, 0, 0, -1, 0, 1, 1, 0, -1, 0, 0, 1, 1, 2, 0, -2, -2, -3, 0, -1, 0, 0, -1, -2, -1, -1, -1, -1, -1, -3, -3, -1, -1, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -3, 0, -1, 0, 0, 0, -2, -2, -1, 0, -1, -2, -1, -2, -2, -1, -1, 0, 0, 2, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, -2, -2, -1, -1, -2, -1, -1, -2, -1, -2, -1, 0, -1, 1, 1, 0, 0, 0, 0, -1, 0, -1, -2, -2, -1, -3, -2, -1, -1, -1, 0, 0, -2, -2, -2, -1, -2, -2, 0, -1, -2, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, -3, -2, -2, -3, -2, -1, 0, 0, -2, -2, -1, -2, 0, -1, -1, -1, -2, -1, -1, -1, 0, -1, -1, 0, 0, 1, 0, 0, -1, -1, -2, -3, -3, -2, -1, -3, -2, -1, 0, -1, -2, -2, -3, -3, -1, -2, -1, -1, -1, 0, 0, -2, 1, -1, 0, 0, 0, 2, 0, 0, 0, 0, -2, -3, -1, 0, -2, -2, -3, -1, -2, -2, -2, -1, -3, -2, -3, -1, -1, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -2, -2, -2, -1, -3, -3, -1, -3, -3, -3, -3, -2, -2, -1, -1, -1, -2, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 1, -1, -1, -2, -2, 0, -1, -2, -2, -2, -3, -3, -3, -3, -2, -2, -2, -1, 0, -1, -2, 0, 0, 0, -2, 0, 0, 0, 0, 0, -1, 0, 0, -2, -2, -2, -1, 0, 0, -1, -2, -2, -2, -3, -2, -3, -3, -3, -3, -1, 0, -1, -2, -1, 0, -1, -2, 1, 0, 1, 0, 0, 0, 0, 1, -1, -1, 0, 0, -1, 0, -2, -2, -2, -3, -3, -1, -1, -2, -1, -2, -1, 0, -1, -2, -2, 0, 0, -3, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, -3, -1, -1, -2, -2, -1, -1, 0, -1, -2, -1, 0, -1, -2, 0, 1, 2, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, -2, -1, -1, 0, -2, -1, -1, 0, 0, 0, -1, -1, 0, 0, -3, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -3, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, -1, 0, 0, 0, 0, -1, -2, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 1, 0, 2, 0, 0, 0, 1, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 3, 2, 1, 1, 1, 0, 0, 1, -1, -2, -1, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, -1, -1, -1, -1, -2, -2, -2, -3, -2, 0, 0, 4, 2, 2, 1, 1, 0, 0, 0, -2, -3, -1, -1, 0, 0, 1, 0, 1, 0, 1, 0, 0, -1, -1, -2, -2, -2, -2, -2, -3, -3, -1, 1, 2, 2, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -2, -1, -3, -4, -4, -1, 2, 3, 2, 1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -2, -2, -3, -2, -1, 0, 2, 2, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -2, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, -2, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 2, 1, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 2, 3, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 2, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 2, 0, 1, 1, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, -2, -1, 0, 1, 2, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 2, 1, 0, 0, -2, -2, -1, -1, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 1, 2, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 2, 0, 0, -2, -1, -1, 0, -1, 0, 1, 0, -1, 0, -1, 0, -2, 0, 0, 2, 1, -1, -2, 0, -1, -1, 0, 0, -2, -1, 0, 2, 1, 2, 1, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 2, 0, -1, -1, -2, -1, 0, 0, 0, 0, -1, 0, 2, 1, 1, 1, 1, -1, -1, -2, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, 0, 2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 2, 3, 1, 1, 1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 2, 2, 2, 2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 1, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 2, 2, 2, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 1, 2, 2, 1, 0, 0, -1, -1, 0, -1, 0, 1, 2, 0, 2, 1, 1, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 3, 3, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 2, 3, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -2, -1, 2, 2, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 2, 2, 2, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -2, -1, 1, 3, 0, 0, 0, 0, 0, -1, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, -4, -1, 2, 2, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -2, -3, -1, 1, 4, 2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, -2, -3, -4, -1, 1, 2, 2, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -2, -2, -2, -1, -2, -3, -4, -1, 1, 4, 2, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 1, 0, 0, 0, -2, -2, -1, -2, -2, -1, 2, 2, 3, 3, 1, 1, 0, 1, 1, 1, -1, 0, 0, 0, 0, 1, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, 0, 1, 2, 2, 3, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 1, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 1, 0, -1, 0, 1, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 2, 0, 2, 1, 0, 0, 1, 0, 1, 0, 1, 1, 0, 1, 0, 1, 1, 2, 2, 1, 0, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 3, 2, 1, 1, 1, 1, 3, 1, 1, 1, 2, 1, 2, 2, 1, 0, -1, -3, -2, -1, -1, -1, 0, 0, -1, 0, 1, 0, 1, 2, 3, 3, 4, 3, 2, 3, 3, 4, 3, 2, 3, 3, 4, 3, 5, 5, 2, 0, -2, -2, -3, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 3, 2, 2, 1, 1, 3, 3, 2, 2, 1, 3, 3, 3, 4, 5, 2, 1, -1, -3, -2, -2, 0, -1, 0, -1, -2, -1, -1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 1, 1, 1, 1, 2, 2, 0, 1, 3, 3, 1, -1, -4, -3, -1, -1, 0, -1, -1, -1, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 1, 1, -1, 0, 2, 2, 1, -2, -4, -2, -1, -1, -3, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 1, 0, -3, -3, -3, -1, -2, -3, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 2, 0, -3, -4, -3, -2, -1, -3, -3, 0, 0, 1, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -3, -3, -2, -2, -1, -2, -2, -1, 0, 1, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, -4, -4, -3, -2, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -2, -2, -2, -2, -2, -1, -2, -1, 0, -1, 0, 1, 1, 0, 0, 1, 0, 0, -2, -3, -2, -1, 0, -1, 0, 0, 1, 1, 1, 1, -1, -2, -2, -2, -1, -2, -3, -3, -1, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, 1, -1, -3, -2, -1, -1, 0, 1, 0, 1, 2, 2, 2, 1, -1, -3, -4, -2, -2, -3, -2, -2, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, 0, -1, -3, -2, -1, -1, 0, 0, 1, 2, 1, 2, 2, 0, -1, -4, -4, -2, -2, -2, -2, -2, -1, -1, 0, 1, 0, 0, 0, -2, 0, 0, 0, -1, -1, -2, -1, 0, 0, 1, 1, 1, 2, 3, 1, 1, 0, -4, -4, -4, -2, -2, -1, 0, -1, 0, -1, 0, 1, 0, -1, -1, 0, 1, 1, -2, -1, -2, 0, 1, 2, 1, 0, 0, 0, 1, 2, 0, -3, -4, -4, -3, -2, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -2, -3, -1, 0, 0, 0, 1, 2, 1, 0, 1, 0, -2, -3, -4, -5, -5, -2, 0, 1, 2, 3, 2, 1, 0, 1, 0, 1, 1, 0, 2, 0, -3, -2, -1, -1, 0, 1, 1, 0, 0, 1, 0, 0, -1, -3, -4, -5, -5, -2, -1, 2, 3, 4, 4, 3, 0, 0, 1, 1, 0, 2, 2, 0, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -4, -5, -4, -4, -2, 0, 1, 4, 3, 2, 1, 0, 0, 0, 0, 0, 2, 0, -2, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -2, -5, -5, -4, -5, -3, -1, 0, 2, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, -2, -2, 0, 0, 0, 0, -1, -1, 0, 1, 0, -1, -1, -3, -3, -5, -5, -4, -3, -2, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 2, 1, -1, -2, -2, -2, -1, 0, -1, -1, 0, 0, 0, 0, -1, -4, -5, -3, -6, -4, -3, -2, -1, 0, 0, -1, 0, -2, 0, 0, 0, 1, 1, 1, -1, -2, -3, -2, -2, -1, 0, -1, 0, 0, 0, 0, -2, -3, -3, -3, -4, -5, -3, -2, -2, 0, -1, -2, -2, -1, -1, 0, 0, 0, 1, 0, -2, -2, -1, -2, 0, 0, -1, 0, 1, 0, 0, -1, -2, -3, -3, -2, -2, -2, -1, -1, -1, 1, 0, -1, 0, 0, 0, -1, 0, 0, 2, 1, -2, -2, -3, -2, -1, 0, -1, 0, 0, 1, 0, -2, -2, -1, -2, -2, -1, -1, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 1, 2, 0, -3, -3, -2, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, -2, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 2, 2, 1, -3, -3, -3, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 2, 1, 0, -4, -4, -2, -1, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 3, 2, 1, -4, -3, -2, 0, 0, -1, -1, 0, -1, -1, -2, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 4, 2, 0, -3, -5, -3, 0, 0, 0, -1, -2, -1, -2, -1, -1, 0, 1, 0, 2, 2, 1, 1, 1, 1, 1, 0, 0, 2, 3, 1, 2, 3, 4, 2, 0, -3, -5, -4, -1, 0, 0, 0, 0, -2, -1, 0, 0, 1, 1, 2, 2, 2, 1, 2, 3, 2, 1, 1, 2, 2, 3, 3, 2, 2, 4, 2, 0, -2, -4, -2, 0, 1, 1, 0, 0, -1, 0, 0, 1, 2, 2, 1, 2, 2, 2, 3, 4, 3, 2, 2, 3, 2, 4, 4, 4, 3, 4, 1, 0, -1, -1, -1, 0, 1, 0, 1, 0, 0, -1, 0, 0, 2, 2, 1, 2, 1, 2, 1, 2, 1, 1, 2, 3, 2, 3, 3, 3, 3, 2, 1, 1, 0, 1, 0, 0, -1, -1, 0, -2, -1, -2, 0, 0, 0, -2, 0, -1, -1, -1, 0, 1, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -2, -2, -2, 0, -2, -3, -1, -1, -1, 0, 0, 1, 2, 0, 1, 1, 1, 0, 0, 1, 1, 1, 0, 0, -2, 0, 1, 0, -1, -3, -3, -1, -1, -2, -2, 0, -1, 0, 0, 0, 0, 0, 2, 2, 3, 2, 2, 2, 2, 1, 2, 1, 1, 1, 0, 0, -1, 0, 0, 0, -2, -1, -2, -2, -1, -2, -2, -2, -1, -2, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, -2, 0, -3, -3, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, -2, 0, 0, 0, 0, -1, 1, 0, 0, -1, -1, 0, 1, 2, 1, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, -2, -2, -1, 0, 0, -1, -3, -2, 0, 0, 0, 0, -1, 1, 1, 0, -1, -1, 1, 0, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -3, 0, 0, 0, -2, -2, -1, 0, 0, 0, -1, 1, 1, 0, -1, -1, 0, 2, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, -1, -2, -1, 0, 0, 0, -1, 1, 1, 0, 0, -1, 0, 1, 4, 3, 2, 0, 1, 1, 0, 1, 0, 0, 1, 1, 0, -1, -1, 0, -1, -2, -1, -2, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 1, 3, 4, 2, 0, 0, 0, 1, 1, 0, 1, 0, 2, 1, 0, 0, 0, 0, -2, -2, -1, -1, -1, 0, 0, -2, 0, 1, 1, 0, 1, 0, 2, 3, 3, 2, 1, 2, 0, 2, 4, 3, 2, 0, 0, 0, -1, -1, -2, -2, -2, -3, -1, -2, -1, 0, 0, -3, 0, 0, 1, 2, 3, 2, 1, 3, 2, 2, 2, 2, 1, 3, 6, 6, 4, 3, 3, 1, 0, 0, -2, -2, -2, -3, -1, -1, 1, 0, 0, -2, 0, 0, 0, 1, 2, 2, 1, 1, 3, 3, 3, 2, 1, 4, 5, 7, 6, 5, 3, 2, 1, 0, -2, -3, -3, -3, -2, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, 1, 1, 1, 2, 3, 4, 2, 4, 3, 4, 6, 6, 5, 4, 2, 0, 0, 0, -1, -2, -3, -1, -2, -2, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 1, 2, 2, 3, 5, 4, 4, 5, 5, 6, 6, 4, 0, -2, -3, -2, -1, 0, 0, 0, -1, -2, 0, -1, 0, 1, 0, -1, -2, 0, 0, 0, 1, 0, 2, 4, 4, 4, 4, 6, 6, 7, 7, 7, 2, 0, -3, -2, -1, 0, 1, 0, -1, -1, 0, 0, 0, 2, 1, -1, -1, -1, 0, 0, 0, 0, 0, 2, 2, 3, 4, 4, 6, 7, 9, 7, 4, 0, -2, -3, -3, 0, 0, 1, 0, -1, 0, 0, 0, 3, 2, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 3, 4, 4, 7, 6, 6, 5, 1, -2, -3, -1, 0, 0, 0, 0, 0, -1, -1, 0, 2, 1, -1, -2, -1, 0, 1, 0, 1, 0, 2, 1, 2, 3, 3, 4, 6, 5, 5, 5, 3, -1, -2, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -3, -2, 0, 1, 1, 0, 3, 4, 1, 1, 4, 4, 4, 5, 4, 4, 2, 2, 0, -1, -2, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -2, -3, -3, 0, 0, 0, 0, 4, 4, 2, 3, 4, 3, 3, 4, 3, 1, 1, 0, -1, -1, -2, 0, 0, -1, 0, 0, 0, 0, -2, -1, 0, -2, -2, -2, 0, 0, 1, 0, 2, 3, 2, 3, 4, 3, 3, 2, 2, 1, 2, 0, -1, -1, -3, 0, -1, -1, -1, 0, 0, 0, -2, -1, 0, -2, -2, -1, 0, 1, 1, 2, 1, 3, 2, 1, 1, 2, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, 0, 0, -1, 0, 0, 0, -4, 0, 0, -1, -1, -1, 0, 2, 3, 2, 1, 0, 0, 1, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -3, 0, 0, -2, -1, -1, 0, 1, 3, 1, 1, 0, -1, 0, 1, 1, 1, 0, 1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -3, 0, 0, -1, -1, 0, 0, 2, 3, 1, -1, -1, 0, -1, 1, 2, 1, 0, 0, 1, 2, 2, 3, 2, 2, 1, 0, 0, 0, 0, 0, -1, -3, 1, 0, -1, -2, -2, 0, 0, 2, 0, -1, 0, 0, -1, 0, 0, 1, 1, 1, 1, 0, 1, 2, 3, 2, 1, 2, 1, 0, 1, 0, 1, -2, 1, 0, -1, 0, -1, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 2, 3, 2, 0, 1, 2, 3, 2, 3, 2, 0, 0, 0, 0, -3, 0, 1, 0, 0, -1, -2, 0, 0, 0, 0, 0, -1, -1, -1, -1, 1, 0, 1, 2, 3, 2, 2, 3, 2, 2, 4, 2, 1, 0, 0, 0, -3, 0, 0, 0, -1, -1, -1, -1, -2, -2, 0, -1, 0, -2, -2, -2, -1, 0, 0, 1, 2, 2, 2, 1, 2, 1, 3, 2, 1, 1, 0, 0, -4, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, -1, -1, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, -2, 0, 0, 1, 1, 0, 0, -1, 0, 0, 1, 2, 0, 0, -1, -2, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 2, 1, 1, 1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 2, 2, 1, 0, 3, 3, 3, 0, 2, 1, 0, 1, 0, 1, 4, 2, 1, 1, 1, 1, 3, 2, 0, 0, 2, 1, -1, 0, 0, 0, 2, 0, 3, 3, 1, 1, 2, 2, 1, 0, 1, 2, 0, 0, -1, 0, 3, 2, 0, 0, 0, 0, 1, 2, 0, 0, 2, 1, 0, -2, 1, -1, 1, 0, 3, 3, 1, 0, 1, 1, 1, 0, 1, 1, 0, 0, -2, -2, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 2, 2, -1, -1, 0, 0, 0, 1, 3, 3, 1, 1, 1, 3, 1, 0, 1, 1, 1, 0, -4, -3, -1, -1, -1, 0, -1, -2, -2, -1, 0, 0, 2, 2, 0, -1, 0, 0, 0, 0, 3, 1, 2, 0, 1, 1, 2, 0, 1, 2, 1, -2, -4, -5, -4, -4, -2, -1, -2, -3, -1, -1, -2, 0, 1, 1, 0, 0, 0, 0, 1, 0, 2, 2, 1, 1, 2, 3, 3, 0, 0, 0, 0, -3, -6, -5, -4, -5, -4, -1, -3, -2, -2, -2, -1, 0, 2, 1, -1, 0, 0, 0, 2, 2, 1, 0, 2, 0, 0, 2, 4, 3, 0, -1, -1, -2, -4, -4, -4, -7, -6, -4, -3, -3, 0, -1, -2, 0, 0, 1, -2, 0, 0, 0, 1, 1, 2, 2, 3, 1, 1, 1, 4, 2, 1, 0, -2, -3, -3, -3, -2, -4, -6, -2, -4, -4, -1, 0, 0, -2, 0, 0, -2, 0, 0, -1, 0, 3, 2, 2, 2, 4, 3, 3, 4, 2, 0, 0, -3, -2, -2, -1, -2, -3, -4, -2, -3, -5, -1, 0, -1, -2, -1, 0, -3, 0, 0, 0, 1, 2, 1, 1, 3, 4, 4, 3, 1, 0, 0, 0, -3, -3, -1, 0, 0, -4, -2, -2, -2, -2, -1, 1, -2, -2, -1, -1, -3, -1, 0, 0, 0, 2, 1, 0, 1, 2, 5, 4, 2, -1, 0, 0, -3, -2, -1, 1, 0, 0, -2, -1, -2, -3, 0, 1, 0, -1, 0, -3, -3, -1, 0, -2, 3, 4, 2, 0, 1, 2, 5, 3, 2, 0, -1, -2, -4, -3, 0, 1, 1, 0, -1, -1, -2, -2, 0, 1, -2, -2, -1, -2, -2, -2, 0, -2, 1, 3, 2, 0, 0, 2, 3, 4, 3, 0, -2, -4, -4, -3, 1, 1, 3, 1, 1, 0, -1, -3, 0, 0, -2, 0, 0, 0, -3, -2, 0, -1, 1, 3, 2, 0, 0, 3, 4, 3, 4, 0, -3, -5, -3, -3, 0, 2, 3, 1, 1, 0, 0, -2, 0, 1, -2, -2, -1, -1, -2, -1, 0, -1, 2, 4, 3, 1, 1, 3, 3, 4, 4, 0, -4, -6, -3, -2, 0, 2, 4, 3, 1, 0, -1, -2, 0, 0, -1, -2, 0, 0, -3, -1, 0, -1, 2, 3, 4, 1, 2, 3, 3, 4, 1, 0, -4, -5, -3, -3, 0, 3, 4, 4, 3, 0, -2, -1, 1, 0, 0, -1, 0, 0, -2, -2, 0, -1, 1, 3, 2, 1, 3, 3, 2, 2, 0, 0, -4, -6, -4, -3, -1, 2, 4, 3, 3, 0, -1, -1, 0, 0, 0, 0, 0, 0, -2, -2, 0, -2, 0, 1, 1, 2, 2, 4, 3, 1, -1, -2, -4, -6, -4, -4, -1, 1, 2, 2, 1, 0, 0, -2, 1, -1, 0, 0, 0, 0, -2, -3, 0, -3, 0, 0, 2, 2, 1, 3, 2, 1, -1, -2, -2, -5, -4, -2, -2, -1, 1, 2, 0, 0, -2, -3, 0, 0, -1, 0, 0, 0, 0, -2, 0, -2, 0, 1, 2, 4, 1, 3, 3, 1, -2, -2, 0, -1, -3, -2, -3, 0, 0, 0, -1, 0, -3, -2, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, 2, 0, 1, 3, 2, 3, 3, 3, -1, 1, 2, 0, -3, -3, -1, 0, -2, -1, -1, -1, -4, -3, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 3, 2, 0, 2, 2, 2, 4, 1, 0, 2, 2, -1, -3, -3, -1, -2, -2, -3, -1, -3, -5, -3, 0, -2, 0, 0, 0, 0, -1, -1, 0, -1, 6, 3, 0, 1, 2, 2, 4, 2, 1, 1, 4, 0, -3, -3, -2, -1, -1, -2, -2, -1, -2, -3, -1, 0, -1, 0, 0, 0, -2, -2, 0, 0, 8, 2, 0, 2, 3, 3, 3, 4, 4, 2, 2, 1, -2, -2, 0, -1, -1, 0, -1, 0, -2, -1, -1, -1, 0, 0, 0, 0, -3, -2, 0, 0, 7, 2, 0, 2, 4, 4, 2, 3, 5, 4, 2, 1, 0, -1, 0, -1, -2, 0, 0, -1, -2, -2, 0, 0, 0, 0, 1, 0, -3, -2, 0, 0, 7, 2, 0, 2, 4, 4, 1, 3, 6, 4, 3, 3, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 1, 2, -1, 0, 1, 1, -2, -3, 0, 1, 6, 2, 1, 1, 5, 5, 3, 4, 3, 4, 3, 3, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 2, 2, 0, 0, 1, 0, -1, -2, 0, 0, 5, 2, 0, 3, 4, 4, 5, 6, 4, 3, 2, 3, 2, 2, 0, 0, 0, 1, 1, 0, 0, 1, 3, 2, 0, 0, 0, 1, -1, -1, 0, 0, 3, 2, 1, 0, 2, 3, 4, 6, 4, 1, 3, 2, 2, 1, 0, 0, 0, 1, 1, 0, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 2, 1, 3, 5, 5, 1, 1, 2, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 2, 0, 1, 1, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 1, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -2, 0, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, 1, 2, 2, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 1, 0, 2, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -2, -3, -2, -2, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, -2, -4, -2, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -2, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, -2, -3, -3, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, 0, 0, 0, -1, -2, -1, -1, 0, -1, -1, -2, -2, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, -2, 0, 0, -1, -1, 0, -1, -1, 0, 1, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, -1, -1, -1, -2, -2, -1, -2, -1, -1, -1, -1, -1, -1, -1, 0, -1, -1, 0, 0, -1, -1, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, -2, -1, -3, -3, -1, -2, -2, -2, -2, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -2, -3, -1, -1, 0, -2, -1, 0, -1, -1, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 2, 0, 0, 1, 1, 2, 1, 0, 0, 0, -2, -3, -2, -3, 0, -1, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, -1, -2, -1, 0, 1, 1, 2, 1, 2, 2, 1, 1, -1, -1, 0, -1, -1, -1, -2, -1, -1, -2, 0, -1, -1, 0, -1, -1, -1, -1, -1, 0, -1, -1, 0, 0, 1, 1, 1, 1, 2, 2, 1, 1, 0, 0, -1, -1, -1, -2, -2, -1, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, -1, -2, -1, -1, -2, 0, 1, 1, 1, 2, 1, 1, 1, 2, 0, 0, 0, -2, 0, -2, -1, -1, -1, 0, -1, -2, 0, -1, -1, 0, -1, -1, 0, -1, -1, -1, -1, 0, 1, 0, 0, 1, 1, 1, 0, 0, 1, 0, -1, -2, -2, -2, 0, -1, -1, -1, 0, 0, -2, -1, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 2, 0, 1, 0, 0, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, -1, -1, 0, 1, 0, 0, 0, 1, 2, 2, 1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -2, -1, 0, -2, -1, 0, 0, 0, 1, 0, 0, 2, 2, 2, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 1, 2, 0, 1, 0, 2, 1, 0, 1, 0, 0, -1, -2, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 1, 2, 2, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, -2, -2, -1, -1, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, -2, -1, -3, -3, -1, 0, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -2, -2, -3, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -2, -1, -2, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, 0, 0, -1, -1, 0, -1, -1, 0, -1, -2, 0, -2, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, -1, 0, 0, 0, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -3, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -2, -3, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 1, 0, 1, -1, 0, 1, 1, 2, 2, 0, 0, 0, 0, 1, 2, 0, 1, 2, 1, 0, 0, 1, 0, 0, 0, 0, -1, -2, -2, -2, -2, 0, -1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -4, -2, -1, 0, 0, 2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, -3, -1, -2, -1, 0, 2, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, -3, -1, -1, -1, 0, 1, 0, -1, 0, 0, 0, -1, -1, -1, -2, 0, 0, 1, 0, 1, 2, 2, 2, 0, 1, 1, 0, 0, -1, 0, -1, -2, -2, -3, 0, -1, 0, 2, 0, -1, 0, 0, -1, -1, -1, -3, -1, -2, 0, 0, 0, 0, 0, 2, 2, 1, 1, 1, 1, 1, 0, 0, 0, -1, -3, -1, -2, 0, 0, 2, 1, 1, 0, 1, 0, 0, -2, -2, -2, -2, -2, 0, -1, 0, 0, 1, 2, 3, 2, 3, 3, 1, 1, 0, 0, -1, 0, -2, -2, 0, 0, 2, 2, 1, 1, 1, 0, 0, 0, -2, -2, -1, -2, -1, -1, 0, 0, 2, 3, 3, 3, 4, 4, 3, 1, 1, 0, 0, 0, -2, -2, 0, 1, 2, 4, 1, 1, 2, 1, 0, -1, -2, -3, -2, -2, -1, -1, -1, 0, 0, 0, 3, 2, 3, 4, 2, 1, 0, 0, -1, 0, -1, -2, 0, 0, 2, 3, 1, 2, 2, 0, 0, -2, -2, -1, -1, -2, -2, -2, -1, -2, -2, -1, 1, 1, 2, 1, 2, 2, 1, 0, -1, 0, -1, 0, 0, 1, 3, 3, 3, 2, 2, 0, 0, -1, -2, -2, -4, -4, -2, -3, -3, -4, -4, -3, -2, 0, 1, 2, 2, 2, 1, 0, 0, 0, -2, 0, 0, 0, 3, 3, 1, 2, 1, 1, 0, -1, -3, -3, -4, -3, -3, -2, -3, -4, -4, -4, -2, 0, 1, 3, 2, 3, 1, 1, 0, 0, 0, 0, 0, 0, 2, 2, 2, 3, 1, 1, 0, -1, -3, -4, -5, -5, -2, -3, -4, -4, -4, -3, -1, 2, 4, 5, 5, 4, 3, 1, 1, 1, 0, 0, -1, 0, 0, 1, 2, 1, 1, 0, 0, -1, -3, -5, -5, -4, -3, -2, -3, -2, -2, -1, 0, 2, 4, 6, 7, 4, 4, 2, 0, 2, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, -1, -3, -4, -4, -4, -3, -2, -2, -2, -2, -2, 0, 2, 5, 6, 6, 4, 3, 1, 1, 1, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, 0, 0, -2, -3, -3, -3, -1, -1, -2, -3, -3, -1, 0, 1, 4, 5, 7, 4, 3, 2, 1, 0, 0, -1, 0, 0, 2, 2, 1, 1, 1, 0, -1, -1, -2, -3, -2, -3, -2, -1, -1, -2, -2, -2, 0, 1, 3, 6, 5, 5, 2, 1, 1, 0, 0, 0, 0, 1, 2, 3, 1, 1, 1, 0, 0, -3, -3, -2, -3, -2, -3, -2, -1, -2, -3, -1, -1, 2, 3, 3, 4, 5, 2, 1, 0, 0, 0, 0, 0, 0, 2, 3, 2, 1, 0, -1, -1, -1, -3, -3, -2, -3, -3, -2, -1, -2, -2, -1, 0, 1, 2, 3, 4, 4, 2, 1, 2, 0, 0, 0, 0, 0, 3, 3, 2, 2, 0, 0, 0, -2, -3, -3, -3, -4, -3, -3, -1, -1, -1, 0, 1, 4, 4, 4, 5, 5, 3, 3, 1, 1, 1, 0, 0, 0, 2, 2, 2, 1, 0, 0, -1, -3, -3, -4, -5, -4, -4, -2, -1, -2, 0, 1, 2, 4, 7, 7, 7, 5, 4, 1, 1, 0, 0, 0, 0, 0, 2, 3, 0, 0, 0, -1, -2, -3, -4, -5, -5, -4, -4, -2, 0, 0, 2, 3, 2, 5, 5, 4, 4, 3, 3, 2, 1, 0, 0, 0, 0, 0, 1, 3, 1, 0, 0, -2, -3, -5, -3, -3, -4, -2, -2, 0, 0, 0, 2, 1, 2, 3, 4, 3, 3, 3, 2, 1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, -1, -1, -2, -4, -3, -4, -2, -2, -1, 0, 0, 0, 0, 1, 1, 2, 1, 1, 0, 2, 2, 0, 0, 0, -1, -1, 0, 0, 1, 2, 0, -1, -1, -1, -3, -4, -4, -3, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, -1, -1, 0, -2, -1, -3, -1, -3, -2, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, 1, 1, 0, 0, 0, -1, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -2, -1, -1, 0, 0, -1, -1, -1, 1, 2, 3, 0, 0, 0, 0, -2, -1, -1, -1, -1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, 0, -1, -1, 0, 2, 4, 1, 1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 2, 1, 2, 2, 2, 1, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 3, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 1, 1, 2, 2, 2, 2, 2, 1, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, -1, 0, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 1, 0, 0, -2, 0, -2, -2, -3, -2, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 1, 1, 0, 0, -1, -1, -3, -3, -3, -3, -1, -1, -1, 0, -1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 1, 2, 0, 0, -1, -1, -3, -2, -2, -2, -2, -1, -1, -1, 0, 0, 1, 2, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 0, -1, -1, -2, -3, -3, -2, -2, 0, 0, 0, 0, 0, 1, 1, 2, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 2, 2, 2, 0, 0, 0, -1, -1, -2, -2, -3, -1, -1, -1, 0, 0, 1, 1, 0, 1, 1, 2, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, -3, -3, -2, -2, -1, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 2, 0, 0, -1, 0, -2, -2, -2, -2, -1, -2, 0, 0, 0, 0, 1, 1, 2, 2, 1, 1, 0, 2, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -2, -2, -2, -2, -1, 0, 0, 2, 2, 1, 2, 2, 1, 1, 1, 2, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, -1, -1, -3, -2, -2, -1, -1, -1, 0, 0, 0, 2, 2, 2, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, -2, -1, -3, -3, -1, 0, -1, 0, 0, 2, 1, 2, 1, 3, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -2, -1, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, -2, -2, -2, -2, -1, 0, -1, 0, 0, 1, 0, 2, 2, 1, 2, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, -2, -1, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, 1, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 2, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, -1, -1, -3, -1, 0, -2, -1, -1, 0, -1, 0, 0, 0, 1, 0, -1, 0, 1, 0, 0, -1, 0, 1, 1, 0, -1, 0, 0, 2, 1, 0, -1, -1, -2, -2, -2, -1, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 1, 2, 1, 0, 0, 0, 1, 1, 0, 1, -1, -1, -2, -1, -2, -1, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -2, 0, 0, 1, 2, 0, 0, 0, 1, 1, 1, 0, -1, 0, -2, -1, -2, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 1, 0, -2, 1, 1, 2, 2, 2, 1, 0, 1, 1, 1, 0, -1, 0, -2, -1, -1, 0, -1, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 2, 1, 3, 2, 2, 0, 1, 2, 0, 1, -1, -2, -2, -2, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 2, 1, 1, 1, 2, 1, 2, 1, 1, 1, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 2, 1, 1, 1, 3, 1, 2, 2, 1, 1, 0, -2, -2, -2, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 1, 0, 2, 3, 2, 2, 2, 1, 2, 2, 0, 0, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, -1, 0, 0, 2, 2, 1, 3, 1, 2, 1, 2, 2, 1, -1, -2, -1, 0, 0, 1, 0, 0, 0, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 3, 3, 1, 1, 1, 0, 1, 0, -1, -2, -1, 0, 0, 2, 2, 1, 0, -1, -1, 0, 1, 0, 0, -1, -1, 0, 0, -1, 1, 1, 1, 1, 2, 3, 1, 0, 0, 0, 0, -1, -2, -2, -1, 0, 0, 1, 1, 1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 1, -2, 2, 2, 1, 1, 2, 2, 3, 1, 0, 0, 0, 0, -3, -2, -1, 0, 0, 0, 2, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 2, 1, 2, 2, 0, 0, 1, 0, -1, -2, -1, -1, 0, 0, 2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 2, 0, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 2, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, -1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, -2, -1, -1, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, -1, -1, 1, 0, -2, 0, 2, 0, 1, 1, 2, 1, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 3, 1, 2, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, 2, 2, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, 1, 1, 2, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -2, 0, 1, 2, 1, 2, 3, 3, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, 0, 0, 1, -1, 0, 2, 1, 0, 2, 2, 4, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 2, 2, 0, 1, 2, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, 2, 1, 1, 1, 2, 2, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 1, -1, 1, 0, 0, -1, 0, 0, 1, 2, 2, 3, 2, 1, 0, 0, 1, 2, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 1, 2, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 1, 1, 0, 1, 1, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 2, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 1, 1, 1, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, -2, -1, -1, -1, 0, 0, 0, 1, 1, 2, 3, 3, 3, 2, 2, 1, 1, 2, 1, 2, 3, 3, 2, 1, -1, 0, -1, -1, -1, -2, 0, -1, -2, -3, -1, -1, 0, 0, 0, 1, 2, 1, 2, 3, 3, 3, 2, 2, 3, 3, 3, 2, 2, 4, 1, 0, -1, -2, -1, 0, -2, -1, -2, -1, -2, -1, -3, 0, 0, -2, -1, 0, 0, 1, 1, 0, 0, 1, 2, 1, 1, 2, 1, 1, 2, 4, 2, 0, -2, -1, -2, 0, -1, -1, 0, -1, -1, -3, -1, -1, -3, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 2, 2, 1, 3, 1, 0, 0, 0, 0, -2, -2, -1, 0, -1, 0, -1, 0, -3, -2, -4, -3, -1, -1, 0, -1, 0, 0, 0, 1, 1, 2, 1, 0, 0, 2, 2, 1, 0, 0, -1, -2, -2, -2, 0, -1, 0, 0, 0, -1, -1, -2, -2, -1, -2, -1, -1, -1, 0, -1, 0, 0, 1, 0, 0, 1, 0, 1, 3, 1, 0, -3, -2, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, -2, -1, -1, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 2, 0, 0, -4, -2, -1, 0, 0, 0, 1, 2, 2, 2, 1, 0, 0, -1, -2, -2, -2, -1, -3, -3, -2, -2, -1, -1, -1, -1, 0, 0, -1, 0, 1, -1, -4, -3, -2, 0, 0, 1, 2, 2, 3, 3, 1, 1, 0, 0, -1, -2, -1, -3, -3, -4, -3, -2, 0, -1, 0, -1, 0, 0, 0, 1, 1, -1, -4, -3, -1, -1, 0, 0, 1, 4, 3, 3, 3, 3, 2, 0, 0, 0, -1, -3, -3, -3, -3, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -4, -2, -1, 0, 0, 1, 1, 2, 4, 4, 3, 3, 1, 1, 0, 0, -1, 0, -3, -3, -2, -2, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, -3, -3, -3, -3, 0, 0, 1, 3, 4, 4, 5, 4, 1, 0, 0, 0, -1, -1, -2, -1, -3, -2, -2, 0, -2, 0, 0, -1, -1, 0, 0, 0, -2, -3, -2, -2, -1, 0, 1, 2, 5, 5, 6, 5, 2, 2, 0, 0, -1, -2, -3, -2, -2, -2, -2, -1, -1, -1, 0, -1, -1, -2, 0, -1, -1, -2, -3, -3, 0, 1, 2, 3, 5, 5, 4, 4, 2, 1, 1, -1, -1, -1, -2, -2, -3, -2, -2, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, -2, -3, -2, 0, 2, 2, 4, 4, 4, 2, 4, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -3, -1, -1, 0, 0, -1, -2, -1, 0, 0, -1, -2, -1, 0, 0, 1, 2, 3, 2, 3, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, -1, -1, 0, 0, 0, -3, -3, -2, -2, 0, 0, 1, 2, 2, 3, 1, 1, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, -4, -3, -1, -1, -1, 1, 2, 1, 2, 2, 1, 1, 1, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -4, -3, -3, -2, 0, 0, 1, 2, 2, 2, 1, 1, 0, -1, 0, -1, -2, -2, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -3, -3, -2, -2, -1, -1, 0, 1, 1, 3, 2, 2, 0, -1, 0, 0, -1, -2, -1, -2, -2, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -4, -2, -3, -3, -3, -1, 0, 0, 1, 4, 3, 2, 0, 0, -1, -1, -2, -3, -2, -1, -2, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, -3, -4, -1, -2, 0, 0, 0, 1, 3, 2, 2, 3, 1, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -2, -3, -2, -1, 0, 1, 1, 3, 2, 2, 2, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, -1, -3, -1, 0, 1, 0, 2, 1, 3, 2, 1, 0, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 1, -2, -2, -1, 0, 1, 1, 2, 1, 1, 1, 0, 0, -1, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 2, 0, 0, 0, -2, -2, 0, 0, 0, 2, 1, 1, 1, 1, 0, 0, 0, -2, -1, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 2, 0, 0, -1, -1, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 2, 1, 2, 1, 1, 1, 2, 1, 0, -1, -2, -1, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 1, 2, 2, 2, 2, 3, 1, 2, 2, 4, 2, 0, -3, -3, -1, -1, 0, 0, 1, 0, 0, -1, 0, -1, -1, -1, -1, -1, -1, 0, 1, 2, 1, 1, 2, 1, 2, 2, 2, 2, 2, 4, 2, -1, -3, -1, -1, 0, 0, 2, 2, 1, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 2, 2, 2, 3, 3, 3, 2, 3, 3, 2, 2, 4, 1, -1, -1, -2, -2, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 2, 2, 3, 4, 4, 3, 3, 3, 3, 4, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, -1, -1, 0, 0, -1, -1, -1, -1, -1, -2, -2, -2, 0, 0, 1, 1, 2, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, 0, -1, 0, -1, -2, -2, -2, -1, 0, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -1, 0, 0, -1, -1, -2, -2, 0, 1, 1, 2, 2, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -2, 0, 0, 0, -1, 0, 0, -1, -1, 1, 3, 2, 2, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, 0, -1, 0, -2, -1, -2, 0, 1, 2, 3, 3, 2, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -2, 0, 0, 2, 2, 3, 2, 2, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, -2, -2, 0, 0, 0, 2, 1, 3, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, -2, -1, -1, -1, 0, 2, 1, 2, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -2, -1, 0, 0, 1, 3, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 2, 3, 1, 2, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, -2, -1, -1, 0, 0, 1, 2, 1, 2, 1, 2, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, -2, 0, -2, -2, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 2, 2, 2, 1, 2, 0, 1, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 2, 2, 1, 1, 1, 2, 0, 1, 0, 1, 1, 0, 1, 1, 1, 0, -3, -1, 0, 1, 0, 0, -1, -2, -2, -2, 0, 2, 2, 2, 3, 2, 2, 1, 3, 4, 3, 3, 1, 1, 3, 4, 4, 4, 4, 5, 2, 0, -6, -1, 0, 0, 0, 0, -1, -4, -3, 0, 0, 2, 5, 4, 3, 4, 3, 4, 3, 4, 4, 3, 1, 3, 4, 3, 4, 5, 8, 6, 1, 0, -7, -3, -2, 0, 1, 0, -1, -2, 0, 0, 1, 1, 3, 3, 2, 4, 3, 2, 4, 4, 4, 2, 1, 3, 2, 2, 3, 4, 7, 7, 2, 0, -6, -3, -2, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 2, 0, 0, 1, 1, 0, 0, -1, 1, 1, 0, -1, 0, 2, 6, 2, 0, -7, -2, 0, 0, 0, 0, 0, 1, 2, 1, 2, 0, -1, -3, -2, 1, 1, 1, 1, 0, 0, -2, -4, -1, 0, -1, -2, -4, 0, 3, 1, -1, -5, -3, -1, -1, -2, -3, 0, 3, 3, 3, 3, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, -2, -4, -1, 0, 0, -1, -4, -2, 2, 1, 0, -6, -3, 0, 0, -1, -3, -1, 1, 4, 4, 3, 1, 0, -1, 0, -1, 0, 2, 1, 2, 0, -1, -4, -3, 0, 0, -1, -4, -2, 1, 2, 0, -6, -3, -1, 0, 0, -3, -2, 1, 3, 3, 3, 0, 0, -1, -1, 0, 1, 1, 1, 0, 0, -2, -4, -2, 1, 0, -1, -2, -1, 3, 1, 0, -5, -3, 0, 0, 0, -1, -2, 0, 3, 4, 1, -1, -3, -3, -2, 0, 0, 0, 0, 0, 0, -2, -3, -3, 1, 1, 0, -1, 0, 2, 0, 0, -4, -3, 0, 1, 0, 0, -1, 1, 3, 2, 1, 0, -3, -3, -2, -2, 1, 0, -1, -1, 0, 0, -1, -2, 0, 0, 1, -1, 0, 2, 2, 0, -3, -2, 0, 1, 0, 0, 0, 1, 1, 1, 0, -1, -4, -4, -4, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 0, -4, -2, 0, 1, 0, 0, 2, 0, 2, 0, 1, -1, -3, -4, -4, -1, 0, 3, 0, 1, 3, 1, 1, 0, 1, 1, 1, -1, 0, 4, 2, 1, -3, -1, -1, 1, 0, 2, 2, 1, 1, 2, 0, -1, -3, -4, -5, -1, 1, 2, 3, 3, 2, 2, 0, 1, 3, 0, 0, -1, 0, 2, 2, 0, -3, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, -3, -4, -4, -6, -3, 1, 4, 3, 5, 4, 0, -1, 0, 3, 3, 1, 1, 2, 3, 1, 1, -1, 0, 0, 0, 2, 2, 1, 0, -1, -1, -1, -4, -5, -5, -4, -2, 2, 5, 7, 10, 7, 3, 0, 0, 3, 4, 3, 2, 4, 4, 1, 0, -3, -1, 0, 2, 0, 1, 1, 0, 0, -2, -2, -5, -7, -6, -4, -2, 2, 6, 10, 13, 13, 7, 2, 0, 3, 5, 5, 4, 4, 6, 2, 0, -3, 0, 2, 3, 2, 0, 0, 0, 0, -2, -4, -5, -8, -8, -5, -2, 1, 4, 9, 14, 13, 9, 4, 2, 2, 2, 2, 3, 4, 6, 2, 0, -3, 0, 2, 1, 1, 0, 0, 0, 0, -3, -3, -6, -6, -7, -5, -3, 0, 3, 7, 10, 11, 9, 6, 3, 0, 2, 2, 0, 3, 5, 3, 0, -4, -1, 2, 2, 0, -2, -1, 0, 0, -1, -3, -4, -5, -8, -4, -4, -1, 1, 5, 7, 8, 7, 4, 2, 0, 1, 1, 1, 2, 4, 2, 0, -4, -2, 0, 1, 0, -2, 0, 0, -1, 0, -2, -2, -3, -5, -3, -2, -1, 0, 1, 3, 3, 2, 1, 0, 0, 0, 0, 0, 1, 4, 2, 0, -2, -2, 0, -1, 0, -3, -1, 0, 0, -1, -2, -1, -2, -4, -3, -2, -2, 0, 0, 0, 0, 1, -1, -3, -2, 0, 0, -1, 0, 3, 2, 0, -4, -2, -1, 0, 0, -2, -1, 0, 0, 0, -2, 0, -1, -3, -4, -2, -1, -2, 0, 0, 0, 0, 0, -2, -2, 0, 0, -1, 0, 3, 1, 1, -3, -2, -2, -1, 0, -1, 0, 0, 0, 0, -1, -2, -1, -3, -3, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 2, 2, 0, -4, -2, -1, -1, -1, 0, 0, 0, 2, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 3, 1, 0, -5, -2, -1, -2, -2, -1, 0, 0, 2, 1, 0, -1, -1, -1, 0, 1, 2, 0, 1, 0, 0, 0, 0, 1, 3, 1, 0, 0, 2, 3, 0, 0, -5, -3, -2, -1, -1, -2, -1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 1, 2, 2, 0, 0, 4, 4, 0, 0, -6, -2, 0, 0, 0, -1, -2, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, -1, -2, 1, 3, 1, 2, 1, 3, 4, 1, 0, -8, -3, -1, 1, 0, 0, -2, -1, 0, 0, -1, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, -1, -1, 0, 2, 2, 2, 3, 4, 4, 2, 0, -8, -3, 0, 1, 1, 0, -1, -2, -2, -1, 0, 0, 2, 2, 2, 1, 2, 2, 2, 2, 2, 0, -1, 0, 1, 0, 2, 2, 4, 4, 1, 0, -9, -6, -1, 2, 3, 1, 0, 0, -2, -2, -1, 0, 2, 3, 1, 2, 1, 3, 1, 1, 2, 0, 0, 0, 1, 0, 2, 3, 4, 2, 0, -1, -5, -5, 0, 2, 3, 3, 1, 1, -2, 0, 0, 2, 5, 5, 5, 2, 3, 3, 2, 2, 2, 2, 1, 3, 3, 1, 1, 2, 4, 4, 1, 0, -2, -4, 0, 1, 2, 2, 2, 0, 0, 0, 0, 2, 4, 4, 3, 2, 2, 1, 2, 2, 1, 0, 1, 2, 2, 1, 1, 3, 3, 2, 2, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 2, 3, 3, 3, 2, 0, 0, 1, -1, -1, -2, 0, -1, 0, 1, 1, 0, 2, 1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 4, 3, 0, 0, 0, 0, 0, -1, -3, -4, -3, -1, 0, 0, 2, 2, 3, 1, 1, 0, 0, 0, -1, -2, -1, 0, -1, 0, 0, -1, 0, 2, 4, 2, 0, 0, 0, -2, 0, -1, -2, -1, -1, 0, 1, 1, 1, 1, 2, 1, 0, -1, 0, -1, -1, -1, 0, 0, 0, -2, -2, 0, -1, 3, 3, 1, 0, 0, 0, -2, -2, -2, -2, -2, 0, 1, 0, 1, 0, 0, 1, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, 1, 3, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -2, -1, -1, 1, 3, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, 0, -2, -1, 0, 0, -1, -2, -1, 0, 2, 2, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, -1, -1, -1, -1, 2, 2, 0, 0, 0, 1, 1, 1, 2, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 3, 1, 0, 1, 0, 2, 2, 3, 1, 2, 1, 1, 2, 2, 0, 0, -1, 0, 0, -2, 0, 0, 0, 1, 1, 0, 0, 1, 0, -1, -1, -1, 2, 2, 2, 1, 2, 1, 1, 2, 2, 2, 3, 2, 4, 4, 2, 2, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 2, 2, 2, 1, 1, 1, 3, 3, 3, 4, 3, 4, 5, 4, 2, 0, 0, 0, 0, -1, -1, 0, -1, 0, -2, -2, 0, 0, -1, -1, -1, 1, 2, 1, 0, 0, 2, 2, 3, 3, 3, 3, 4, 5, 5, 6, 4, 1, 0, -2, -3, -2, -1, -1, 0, -1, -2, -2, 0, 0, 0, -1, -1, 2, 1, 0, -1, -1, 0, 1, 2, 3, 3, 3, 3, 3, 4, 4, 3, 0, -2, -4, -2, -2, 0, 0, -1, -2, -1, -1, 0, 0, -1, -1, 0, 0, 0, -1, -3, -3, 0, 2, 1, 3, 2, 1, 2, 3, 4, 5, 2, 0, -2, -4, -4, -3, -1, 0, 0, 0, -1, 0, 0, -1, -2, -1, 0, 0, 0, -2, -2, -3, -3, 0, 1, 3, 1, 2, 0, 2, 5, 4, 2, 0, -1, -4, -4, -3, -1, 1, 0, 0, 0, 0, 0, 0, -2, 0, -2, 1, 0, -1, -2, -3, -2, 0, 1, 1, 3, 1, 1, 2, 5, 4, 2, 0, -2, -4, -4, -2, -2, 1, 1, 0, 0, 0, -1, -1, -1, -1, -2, 0, 1, -1, -1, -2, -2, 1, 2, 3, 3, 3, 3, 3, 6, 5, 2, 0, 0, -2, -3, -3, -1, 0, 0, 0, -1, -1, -1, -1, -2, -3, -1, 1, 0, -1, 0, -1, 0, 1, 2, 2, 2, 4, 3, 5, 4, 5, 2, 1, 0, -1, -2, -2, -1, 0, 1, 0, -1, 0, -1, -3, -3, -2, -1, 1, 2, 1, -1, 0, 0, 1, 3, 3, 3, 4, 3, 4, 4, 3, 3, 1, 0, -2, -2, -1, 0, 0, 0, 0, -1, -1, -1, -2, -1, -2, -2, 1, 2, 1, 0, -1, 0, 3, 3, 3, 4, 4, 5, 3, 4, 3, 1, 1, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, -1, -2, -1, -1, -1, 2, 2, 0, 0, 0, 1, 3, 4, 3, 4, 4, 5, 3, 2, 1, 2, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, -1, 0, 1, 1, 0, 1, 0, 2, 3, 2, 4, 4, 4, 4, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 2, 2, 0, 0, 0, 0, 1, 3, 2, 2, 3, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, 0, -2, 0, 2, 3, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -2, -1, -3, -1, 0, 3, 2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, -1, -2, -1, 0, -1, -2, -3, -1, -1, 1, 1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 1, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, 2, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 0, 0, 0, 0, -1, -2, -1, 0, 0, -1, -1, -2, 2, 4, 1, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 2, 5, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 2, 1, 1, 0, 2, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 3, 5, 4, 1, 1, 1, 1, 1, 0, 0, -1, -1, -1, 0, 1, 1, 2, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 2, 3, 2, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 3, 1, 1, 1, 0, 0, 0, -1, -1, -2, 0, -1, 0, 2, 1, 1, 0, 0, 0, -1, 0, -1, -2, 0, -2, 0, 0, -1, -1, 0, 0, 2, 3, 1, 1, 1, -1, -1, 0, -2, -3, -2, -2, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, -1, -2, -1, -1, -1, -1, -1, -2, -1, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -2, -1, 2, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 1, 2, 1, 0, 0, 0, 0, 0, 0, -1, 1, 2, 2, 1, 1, 1, 0, 2, 1, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, -2, -1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, -1, -1, -1, 1, 1, 1, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 1, 2, 2, 2, 2, 1, 1, 0, 2, 2, 2, 1, 2, 2, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 1, 2, 1, 2, 1, 2, 1, 2, 3, 4, 4, 4, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 2, 0, 1, 1, 1, 1, 2, 2, 3, 2, 4, 3, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 0, 0, 0, 0, 2, 1, 2, 1, 2, 1, 2, 3, 4, 4, 2, 1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 2, 2, 1, 1, 3, 3, 3, 2, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 1, 2, 1, 0, 0, 2, 4, 4, 2, 0, 0, -1, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 1, 0, -1, -1, 0, 0, 0, 2, 1, 0, 0, 3, 3, 3, 2, 1, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, -1, -2, -2, -1, 0, 2, 2, 3, 1, 1, 2, 5, 4, 3, 0, 0, -1, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, -1, 0, 1, 2, 3, 3, 3, 2, 3, 3, 4, 2, 2, 1, 0, -1, -1, 0, 1, 2, 0, 0, -1, 0, 0, -2, -2, -1, 1, 1, 0, 0, 0, 1, 2, 3, 2, 2, 3, 3, 3, 4, 4, 2, 2, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 1, 1, 1, 0, 0, 0, 2, 2, 3, 2, 3, 3, 3, 3, 4, 2, 2, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 2, 1, 2, 0, 0, 0, 2, 1, 3, 2, 4, 3, 2, 2, 3, 2, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 3, 1, 1, 0, 1, 0, 1, 3, 3, 3, 4, 3, 1, 0, 1, 1, 1, 0, 1, 1, 0, 1, 0, 1, 2, 0, 0, 1, 0, 0, -2, 0, 3, 1, 0, 1, 1, 0, 2, 2, 3, 3, 4, 2, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 1, 1, 1, 0, 0, -1, 0, 0, 2, 2, 0, 0, 0, 1, 1, 1, 1, 1, 2, 0, 1, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 1, 2, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 2, 2, 0, 1, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 2, 2, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 2, 1, 1, 1, 1, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, -2, 0, 0, 0, -2, -2, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 2, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 2, 3, 3, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 4, 4, 3, 3, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -2, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, -2, -1, -1, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, -1, 0, 1, 0, 0, -1, -2, 0, 0, 0, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 2, 0, 1, 2, 1, 0, 1, 1, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 2, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, 0, -1, 0, -1, 0, 0, -2, -2, -3, -2, -1, 0, -1, -1, -1, 0, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -3, -2, -1, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, -1, -3, -2, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 3, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -2, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 2, 1, 0, 2, 4, 3, 3, 1, 1, 0, 2, 0, 1, 0, 1, 0, -1, -3, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 1, 2, 2, 2, 1, 1, 1, 2, 1, 2, 2, 1, 0, -1, -3, -1, -3, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 1, 1, 1, 1, 0, 2, 0, 1, 2, 2, 1, 1, 0, -1, -2, -2, -2, -3, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 3, 2, 2, 2, 2, 0, 2, 1, 1, 0, 0, -1, -1, -2, -2, -2, -2, 0, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 2, 2, 3, 3, 2, 3, 2, 1, 3, 2, 1, 0, -1, -1, -2, -2, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 2, 3, 4, 2, 2, 3, 2, 4, 3, 3, 0, -1, -2, -3, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 2, 3, 1, 2, 2, 2, 3, 4, 3, 1, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 2, 3, 2, 1, 0, -2, -2, -2, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 2, 1, 1, 1, 1, 0, 1, 1, 2, 2, 2, 0, -2, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, -1, 0, 1, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 1, 3, 0, 2, 0, 0, 0, -1, -1, 0, -1, -1, 0, 1, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 2, 2, 2, 0, 1, 1, 1, 2, 0, 0, 0, 0, -1, -1, -2, -2, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 2, 2, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, -1, -1, -1, -3, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 2, 2, 1, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 2, 2, 1, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 1, 2, 2, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, -1, -1, -1, 0, -1, 0, -1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 1, 1, 1, 0, 1, 1, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 2, 2, 0, 1, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 1, 0, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, -2, -2, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, -1, -2, -2, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -2, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 0, 0, -1, -1, 1, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, -1, 1, 2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, -1, 0, 1, 1, 0, -1, -1, 0, 0, 0, -2, 0, 2, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, -1, 0, -2, 0, -2, -1, -2, 0, -1, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, -2, -1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, -2, -2, -1, -2, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 1, 0, 2, 1, 0, 0, 1, 1, 2, 0, 0, -1, -2, -1, -1, -1, -2, -1, 0, -1, -1, -1, -1, 0, 0, -1, -2, 0, -1, 0, -3, -1, 0, 0, 1, 3, 1, 1, 2, 3, 1, 0, 0, 0, -2, -2, -1, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, -2, 0, 0, 1, 2, 2, 1, 1, 3, 3, 1, 0, 0, -2, -1, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, -1, 0, 1, 2, 1, 2, 1, 2, 1, 1, 1, 0, -1, -2, -2, -1, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -2, 0, 0, 1, 0, 1, 1, 2, 2, 3, 2, 2, 0, -1, -1, -3, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 2, 2, 2, 2, 1, 1, 0, -2, -3, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -2, 0, -1, 0, -2, 0, 0, 0, 0, 2, 2, 2, 0, 2, 1, 1, 1, -1, -2, -3, -1, 0, 0, 3, 1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 2, 2, 2, 1, 0, 0, 1, 0, -1, -1, -3, -1, 0, 1, 1, 4, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -2, -3, -2, -1, 0, 0, 1, 2, 3, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, 0, 0, 1, 1, 1, 1, 0, -1, -1, 0, -2, -3, -2, -2, -1, 0, 2, 1, 3, 1, 0, 0, 0, 1, -1, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 1, 2, 0, -1, 0, 0, -2, -2, -1, -3, -1, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -3, -3, -1, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, 0, 0, -2, -2, 0, -1, 0, 0, 0, 0, 0, -1, -3, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 1, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 2, 1, 1, 2, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 1, 1, 2, 2, 1, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 1, 1, 2, 2, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, -2, 1, 0, 0, 0, 1, 1, 2, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -2, -2, 1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, -1, 1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -2, 0, 1, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 2, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -2, -2, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -3, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -3, -4, -2, 0, -1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -2, -2, -4, -3, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, -2, -3, -3, -5, -3, -2, -1, -1, -1, 0, 0, -1, 0, -1, 1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, -2, -3, -3, -4, -4, -4, -3, -4, -1, -2, -3, -1, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 2, 2, 1, 1, 0, 0, -2, -3, -4, -2, -2, -2, -4, -4, -2, -3, -2, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 3, 2, 2, 0, 0, 0, -2, -2, -3, -2, -2, -2, -2, -4, -2, -2, -2, -1, 0, -1, -2, -1, -2, 0, -1, 0, 0, 1, 1, 1, 1, 2, 2, 2, 2, 1, 1, 0, 0, -3, -2, -3, -1, 0, -2, -4, -1, -3, -1, -1, 0, -1, 0, -2, -2, 0, 0, 0, 0, 1, 2, 0, 0, 2, 3, 3, 1, 2, 0, 0, -2, -2, -2, -1, -1, 0, -1, -2, -2, -2, -2, -1, 0, -1, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 2, 2, 3, 1, 0, -1, -2, -3, -1, -2, 0, 0, -1, -1, -3, -2, -3, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 2, 2, 2, 1, 1, -1, -2, -2, -2, 0, 0, 0, 0, 0, -2, -2, -2, -1, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 2, 0, 1, 0, 1, 2, 4, 3, 1, 0, -2, -3, -2, -2, 1, 1, 1, 0, -1, -2, -3, -1, 0, -1, -1, -2, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 2, 2, 3, 2, 2, 0, -1, -2, -1, 0, 0, 2, 2, 1, 0, -1, -2, -1, 0, -1, -2, -2, -1, -1, 0, 0, 0, 0, 1, 2, 2, 2, 3, 3, 2, 2, 2, 0, -3, -1, -2, -1, 0, 1, 1, 1, -1, -1, -2, 0, -1, -1, -2, -1, -1, 0, -1, 1, 0, 1, 0, 1, 1, 1, 3, 2, 1, 1, 0, -1, -3, -2, -3, -2, 0, 2, 0, 1, 0, -2, -2, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, -1, -3, -3, -3, -1, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -2, 0, 0, -2, 0, -1, -1, 0, 0, 0, 1, 0, 1, 1, 0, -2, 0, -1, -3, -4, -1, -1, 0, 0, -1, -1, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, -3, -3, -2, -2, 0, 0, 0, -1, -1, -2, -2, 0, -1, -1, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -2, -2, -2, -1, 0, -2, -1, -2, -2, -2, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, -2, -3, -1, -2, 0, 0, -2, -1, -1, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, -1, -2, -1, -2, 0, -1, 0, -2, -2, -3, 0, -1, 0, -1, 0, 0, 0, -2, 0, -1, 1, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, -1, -1, -2, -1, 0, -1, -1, -1, -2, -1, -1, 0, -1, -1, -1, 0, 0, -2, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, -1, -2, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 1, -1, 0, 0, 2, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -2, 0, 0, 0, -2, 0, 0, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, -2, 0, 0, 3, 0, 0, 0, 1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 1, 2, 2, 1, 1, 1, 0, 2, 1, 2, 3, 3, 2, 0, -1, -3, -2, -2, 0, -1, 0, -1, 0, 0, 0, 1, 1, 1, 2, 2, 2, 2, 2, 1, 2, 2, 3, 2, 2, 1, 3, 3, 4, 4, 4, 2, -1, -3, -2, -2, -2, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 2, 1, 1, 2, 1, 2, 1, 1, 1, 0, 2, 2, 1, 2, 2, 2, 0, -1, -3, -2, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 2, 1, 2, 2, 2, 2, 3, 2, 0, -3, -2, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 1, 1, 1, 0, 2, 2, 3, 1, -1, -4, -2, -1, -2, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 3, 2, -1, -4, -3, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, -4, -3, -1, -2, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -4, -2, -1, -1, -1, -1, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, -2, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, -1, -2, -1, -1, -2, -3, -2, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, -1, -1, -1, -1, -1, -2, -1, 0, 0, -1, 0, 0, 0, -2, -2, -1, -2, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -1, -1, -1, -2, 0, 0, 0, -1, 0, -1, -1, -1, -2, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -3, -1, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, -1, -1, 0, 0, -1, -1, 0, 0, 1, 0, 1, 1, 1, 1, 0, 1, 2, 1, 1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, 0, 0, 1, 0, 2, 2, 2, 2, 2, 0, 0, 0, 1, 1, 2, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -2, -1, -1, 0, 0, 0, 1, 1, 2, 2, 1, 1, 1, 0, 0, 1, 1, 2, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, -2, 0, 0, -1, 0, 0, 0, 0, 2, 2, 3, 1, 0, 1, 0, 0, 1, 3, 1, 0, -3, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -3, -1, -2, -1, 0, 0, 1, 1, 2, 3, 3, 1, 0, 1, 1, 1, 1, 2, 0, 0, -1, -2, 0, -1, -1, -1, 0, -1, 0, 0, -2, -1, -1, -2, -2, -1, -2, 0, 0, 1, 2, 1, 2, 1, 1, 0, 1, 0, 1, 2, 0, -1, -2, 0, -1, -1, -1, -2, -1, -1, 0, -1, 0, -2, -3, -2, -1, -2, -2, -2, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 2, 3, 0, 0, -1, -2, -1, -2, -2, 0, -1, -1, 0, -1, -2, -2, -2, -3, -1, -2, -1, -1, -1, 0, 0, 1, 1, 0, 0, 1, 1, 1, 2, 3, 1, 0, -1, -1, 0, -1, -2, -1, 0, 0, 0, 0, -2, -3, -3, -1, -2, -1, 0, -1, 0, 0, 0, 1, 2, 1, 0, 1, 0, 1, 2, 2, 1, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 1, 0, -1, -2, -2, 0, -1, -2, 0, 0, 0, -1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 1, 3, 1, -1, -2, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, -2, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, -1, -2, -2, -2, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 3, 4, 2, 0, -2, -3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 3, 2, 4, 1, 0, -2, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 2, 1, 0, 2, 3, 3, 4, 1, -1, -2, -3, -1, 0, 0, 1, 0, 0, 0, -1, 0, 1, 2, 2, 2, 1, 1, 2, 2, 1, 0, 2, 2, 1, 3, 3, 2, 2, 4, 5, 2, 0, -2, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 2, 2, 3, 3, 2, 2, 2, 3, 2, 2, 2, 1, 2, 2, 2, 2, 3, 3, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -2, -1, -1, 0, 1, 3, 4, 4, 4, 3, 2, 1, 1, 2, 1, 2, 1, 2, 1, 1, 2, 2, 2, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 2, 2, 3, 4, 3, 2, 1, 0, 1, 2, 1, 0, 0, 1, 1, 1, 1, 2, 2, 0, -1, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 2, 3, 2, 3, 3, 2, 1, 2, 1, 1, 0, 0, -1, 0, 1, 1, 0, 0, 1, 2, 0, 0, -2, -1, 0, -1, 0, -1, 0, 0, -2, 0, 1, 2, 1, 1, 2, 2, 2, 2, 1, 1, 1, 1, 0, 0, 0, 1, 0, -1, 0, 1, 0, -1, -1, -2, 0, 0, 0, 0, -1, -2, -1, 0, 1, 0, 0, 2, 1, 3, 1, 1, 2, 2, 2, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -2, -1, -2, -1, 0, -1, -1, -2, -1, 0, 0, 1, 1, 2, 0, 2, 1, 1, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, -2, 0, 1, 0, -1, -3, -2, -2, -1, -1, -1, -1, 0, 0, 1, 0, 1, 0, -1, 1, 1, 1, 0, 1, 1, 2, 1, 0, 0, 1, 0, 0, -2, 1, 2, 0, -1, -3, -3, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 1, 2, 1, 0, 1, 0, 0, 0, -1, 1, 1, 0, 0, -2, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, 1, 2, 4, 2, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, -2, 0, 0, 0, -1, -1, -1, 0, -2, -3, -2, -1, -1, 0, 1, 3, 2, 3, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -2, 0, -1, -2, -3, -4, -2, -2, 0, 0, 2, 3, 2, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -3, -2, -5, -6, -6, -5, -5, -2, 0, 2, 1, 2, 1, 2, 2, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -3, -5, -8, -7, -7, -5, -2, 0, 3, 3, 2, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, -1, -2, -2, -1, -1, -4, -5, -7, -7, -6, -4, 0, 2, 4, 6, 4, 2, 1, 1, 0, 0, 1, 1, 0, 0, -2, -1, 0, 1, 2, 2, 1, -1, -1, 0, -1, -2, -4, -4, -6, -6, -4, -1, 0, 4, 7, 6, 6, 3, 2, 1, 0, 0, 1, 1, 0, -2, -1, 0, 0, 2, 1, 2, 0, 0, -1, -1, 0, -2, -3, -5, -6, -5, -4, -3, 2, 4, 6, 6, 4, 3, 2, 0, 0, -1, 1, 1, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -4, -5, -6, -7, -6, -4, 0, 4, 4, 5, 4, 1, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 2, 1, 2, 0, 0, 0, -1, -2, -3, -6, -8, -8, -6, -4, 0, 2, 5, 4, 4, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, -2, -4, -5, -7, -6, -4, -3, 0, 3, 3, 4, 2, 1, 1, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, -2, -1, -3, -5, -5, -6, -4, -3, -1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 2, 1, 0, 1, 1, -1, -2, -3, -3, -6, -5, -5, -5, -1, 0, 0, 2, 2, 2, 1, 0, 1, 0, 0, 1, 2, 1, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, -1, -3, -4, -4, -4, -5, -4, -2, 0, 2, 2, 3, 2, 3, 1, 2, 1, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -3, -3, -4, -2, -4, -2, -1, 0, 1, 1, 2, 2, 2, 1, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -3, -2, -2, -2, -3, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -3, -4, -3, -2, -3, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, -1, 0, 1, 1, 0, -1, -2, -2, 0, 0, 0, -2, -2, -3, -3, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -1, 0, 0, 0, 0, 1, 2, 0, -1, -3, -3, 0, -1, -1, -1, -2, -4, -4, -3, -1, -1, -1, 0, 0, 0, 0, 0, -1, -2, -2, -2, -2, 0, 0, 0, 0, 0, 0, 2, 0, -2, -2, -3, -1, 0, 0, -1, -2, -2, -2, -2, -2, -1, 0, 0, 0, -1, 0, 1, -1, 0, -1, -1, -2, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, -2, -2, 0, -1, 0, -2, -2, -3, -2, -1, 0, 0, 0, 2, 1, 1, 1, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -2, 0, 0, 0, -1, -2, -2, -2, -1, -1, 1, 1, 3, 2, 3, 2, 2, 0, 0, -1, 0, 0, 1, 3, 1, 1, 2, 3, 2, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 2, 1, 3, 2, 3, 2, 2, 2, 2, 1, 2, 1, 2, 2, 1, 2, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, -2, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 3, 1, 1, 0, 2, 2, 1, 0, 1, 2, 0, 1, 2, 2, 2, 2, 3, 2, 2, 0, -3, -2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 3, 3, 2, 2, 1, 2, 0, 0, 1, 2, 1, 0, 0, 1, 1, 2, 3, 3, 2, 0, -2, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 2, 2, 2, 2, 1, 0, 0, -1, 0, 0, 0, 1, 1, 2, 2, 1, 0, -3, 0, 0, 0, 1, 1, 0, 1, 0, 2, 0, 1, 1, 1, 1, 1, 2, 1, 2, 1, 0, 0, -1, 0, 0, 0, -1, -2, 0, 2, 1, 0, -3, -1, 0, 0, 1, 1, 1, 3, 2, 2, 1, 0, 0, 0, 0, 2, 1, 2, 2, 1, 0, -1, -2, 0, 0, -1, -2, -2, -2, 1, 1, -1, -1, 0, 0, 0, 0, 0, 2, 2, 4, 3, 1, 0, 0, 0, 0, 1, 2, 3, 2, 1, 0, -2, -3, -2, 0, -2, -3, -3, -2, 0, 0, -1, -1, 0, 0, 1, 0, -1, 1, 2, 3, 3, 1, 0, 1, 1, 0, 2, 3, 3, 2, 3, 1, 0, -3, -1, 0, 0, -2, -3, -2, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 1, 3, 2, 3, 1, 1, 0, -2, -2, 0, 0, -1, -2, 0, 0, 0, 0, -1, 1, 1, 1, 0, 0, 0, 1, 1, 1, 0, -1, -1, -1, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 2, 0, 0, 0, 1, 2, 1, 0, -1, -1, -1, 0, 0, -2, -2, -3, -4, -2, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 2, 0, 0, 0, 0, -2, -2, -3, -3, -3, -4, -3, -1, 0, 0, 0, 0, 2, 1, 0, 0, 1, 1, 1, 0, 1, 3, 2, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, -2, -4, -3, -5, -5, -4, -3, 0, 0, 0, 1, 1, 1, 1, 2, 1, 0, 0, 0, 0, 2, 2, 0, 0, 0, 1, 1, 1, 1, 2, 0, -2, -1, -3, -4, -4, -4, -5, -2, 0, 0, 0, 2, 3, 1, 1, 1, 2, 2, 1, 1, 1, 3, 3, 0, 0, 0, 0, 1, 2, 2, 2, 0, -2, -2, -4, -6, -5, -6, -4, 0, 0, 1, 3, 3, 3, 2, 2, 2, 2, 2, 1, 3, 3, 3, 2, 0, 0, 0, 1, 1, 1, 1, 1, -1, -2, -3, -5, -7, -8, -5, -3, 0, 3, 5, 4, 4, 5, 4, 2, 2, 4, 4, 4, 3, 3, 3, 3, 0, 0, 0, 1, 1, 1, 0, 0, -2, -1, -4, -4, -6, -7, -5, -3, -1, 2, 4, 4, 7, 5, 4, 4, 2, 3, 3, 4, 4, 3, 4, 4, 0, 0, 1, 1, 3, 2, 1, 0, 0, 0, -2, -4, -5, -7, -5, -2, 0, 0, 3, 4, 7, 5, 6, 4, 4, 4, 3, 2, 3, 2, 4, 3, 0, -1, 0, 2, 3, 2, 0, 0, 0, 0, -2, -3, -4, -5, -4, -3, 0, 0, 0, 3, 4, 4, 6, 4, 3, 2, 1, 2, 2, 2, 3, 2, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -2, -4, -4, -5, -2, 0, 0, 0, 2, 2, 4, 3, 3, 2, 1, 2, 2, 2, 0, 2, 3, 0, 0, 0, 1, 2, 1, 0, -1, 0, -1, 0, -2, -3, -3, -3, -3, -1, 0, 0, 2, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 1, 2, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -3, -3, -2, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 1, 2, 3, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, -1, -3, -2, -3, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 3, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 1, 0, 0, -1, -1, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 2, 1, -1, -2, 0, 0, 0, 1, -1, -1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 1, 1, 2, 0, -3, -1, -1, 1, 1, -1, -1, -2, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -2, -3, -1, 0, 0, 0, 0, 1, 1, 2, 0, -3, -1, 0, 0, 1, 0, 0, -2, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -3, -2, -2, -1, 0, -1, 0, 0, 2, 0, 0, -2, 0, 0, 2, 1, 1, 0, -1, -2, -1, -1, 1, 1, 0, 2, 1, 0, 1, 1, 0, 0, -1, -2, 0, -1, 0, 0, 0, 1, 0, 0, 0, -2, 0, 1, 1, 1, 2, 0, -1, -2, 0, -1, 0, 1, 1, 1, 2, 0, 2, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0,
    -- filter=0 channel=8
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, -2, -1, -1, -1, -1, -2, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, 0, -1, -1, -2, -2, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, -1, -1, -2, -2, -1, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, -1, -1, 0, -2, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, -2, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -2, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -2, -1, 0, -1, -2, -2, -2, -2, -1, -2, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, -1, -1, -2, -3, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -2, -2, -2, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -2, 0, 0, -1, -1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 1, 1, 2, 0, 0, 2, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 2, 2, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 2, 1, 1, 0, 1, 2, 0, 1, 1, 1, 2, 2, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 2, 2, 0, 1, 0, 1, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 2, 2, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, -1, 0, 1, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -1, -1, 0, 0, -1, 0, 0, 1, 0, 2, 1, 1, 2, 1, 0, 0, 0, 0, -1, 0, 4, 3, 1, 0, 0, 0, -1, -1, -2, -4, -3, -4, -3, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, -1, 0, 4, 4, 0, 1, 0, 0, 0, -1, 0, -1, -3, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 3, 1, 0, 1, 0, -1, 0, 0, 3, 4, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 2, 1, 2, 1, 1, 1, 0, -1, -2, 0, 2, 3, 2, 3, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, -1, 1, 0, 1, 0, 1, 0, -1, 0, -2, 0, 4, 4, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, -2, -1, 0, 1, 0, 0, 0, 0, 0, -2, -3, 0, 2, 2, 2, 2, 2, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 1, 0, 0, 0, -1, -3, -2, 0, 3, 2, 3, 1, 2, 1, 0, 0, 1, 1, 0, 0, 0, 2, 2, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -2, -2, -3, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 2, 2, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, -1, 0, -2, -1, -3, -2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 1, 2, 1, 2, 1, 0, 0, -1, -1, -2, -1, -3, -3, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 2, 3, 2, 1, 0, 2, 1, 0, 0, 1, 1, 2, 2, 1, 0, 0, -1, -2, -2, -2, -3, -4, 0, 1, 0, 0, 0, 0, -1, 0, 0, 2, 2, 3, 1, 1, 0, 0, 0, 0, 0, 0, 2, 1, 2, 1, 0, 0, -1, -1, -2, -2, -3, -3, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 2, 3, 2, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 1, 0, 0, 0, -1, -1, -2, -2, -4, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 2, 2, 0, 0, 0, -2, -2, -1, -1, -3, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, -1, -1, 0, 0, 0, 2, 1, 3, 1, 1, 0, 0, -1, 0, -1, -1, -2, -4, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 1, 1, 3, 2, 2, 3, 2, 1, 0, -1, -2, -2, -2, -2, -4, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 2, 3, 2, 3, 2, 2, 0, 0, -1, -3, -2, -1, -4, -3, -1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, -1, 0, 1, 2, 2, 2, 1, 2, 1, 0, 0, -1, -1, -2, -3, -3, -3, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 2, 1, 1, 2, 1, 1, 0, 0, -1, -1, -1, -3, -3, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 2, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, -3, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, -1, -3, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 2, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 2, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, -1, -2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -2, -3, 0, 1, 0, 0, 0, 1, 0, -1, 1, 1, 1, 1, 1, 0, 0, 0, 2, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -3, -3, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, 0, 1, 2, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, -2, -1, -1, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 2, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -2, -1, 0, -2, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, -1, -1, 0, 1, 2, 0, 0, 0, -1, 0, 0, -1, -2, -2, -1, -3, -2, -1, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, -1, 0, -1, 0, -2, -2, -2, -3, -2, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -1, -1, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 3, 1, 0, -1, 0, -3, -2, -4, -4, -5, -4, -2, -1, 0, 1, 0, 0, 1, 2, 2, 2, 2, 2, 2, 1, 1, 1, 1, 0, 0, 1, 3, 4, 3, 2, 1, 0, -1, -1, 0, -2, -1, -1, 0, 1, 1, 3, 1, 0, 1, 2, 4, 4, 3, 5, 2, 3, 3, 4, 4, 2, 0, 0, 4, 5, 3, 4, 2, 2, 1, 0, 0, 1, 0, 0, 2, 3, 3, 2, 0, 0, -1, 0, 0, 0, 2, 3, 3, 3, 3, 4, 2, 1, 0, 0, 3, 5, 3, 4, 2, 2, 1, 0, 1, 2, 2, 1, 2, 2, 2, 1, -1, -1, -2, -3, -1, -2, 0, 1, 2, 3, 2, 2, 2, 0, -2, 0, 2, 6, 5, 3, 4, 2, 1, 0, 1, 0, 0, 2, 2, 2, 2, 0, -1, -2, -2, -5, -4, -4, -2, 0, 1, 2, 1, 1, 1, -1, -3, 0, 2, 4, 5, 5, 2, 1, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, -1, -1, -3, -4, -5, -3, -1, 0, 1, 0, 0, 0, 0, -2, -2, 0, 2, 5, 4, 4, 2, 1, 0, 1, 0, 0, 1, 1, 1, 2, 1, 0, -1, -1, -3, -4, -3, -2, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 2, 4, 3, 3, 2, 0, 0, 0, 1, 2, 1, 2, 1, 2, 1, 0, -1, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, -1, -2, 0, 0, 3, 3, 1, 2, 0, 0, 0, 2, 3, 1, 2, 2, 2, 1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, -1, -1, 0, -2, -2, 0, 0, 2, 3, 2, 1, 0, 0, 1, 1, 2, 3, 2, 2, 0, 0, 0, -1, -1, 0, 0, 0, 2, 2, 1, 1, 0, 0, 0, 0, -2, -2, 0, 0, 1, 3, 2, 1, 1, 0, 2, 2, 3, 2, 1, 0, 0, -2, -1, -1, -1, -1, 0, 0, 2, 3, 2, 2, 0, 0, 0, -2, -2, -3, 0, 0, 2, 2, 1, 1, 0, 0, 1, 2, 3, 3, 2, 0, -1, -2, -2, -2, -1, -1, 0, 1, 2, 3, 4, 1, 0, 0, 0, -2, -2, -3, -1, 0, 1, 2, 1, 1, 1, 2, 1, 2, 1, 2, 0, 0, -2, -2, -1, -1, 0, 0, 0, 2, 3, 3, 3, 2, 1, 1, 0, -1, -2, -3, 0, 0, 2, 2, 3, 2, 1, 2, 1, 0, 0, 1, 0, -2, -3, -4, -2, -1, -1, 0, 1, 2, 4, 3, 4, 3, 0, 0, -1, 0, -2, -3, 0, 2, 2, 3, 2, 3, 2, 1, 2, 2, 0, 0, 0, -1, -3, -2, -2, -1, 0, 1, 1, 4, 5, 4, 3, 2, 0, 0, 0, -2, -3, -4, 0, 2, 4, 4, 4, 2, 0, 0, 1, 1, 0, 1, 0, -2, -3, -3, -2, 0, 1, 3, 3, 3, 3, 5, 2, 2, 0, -1, -2, -2, -3, -4, 0, 2, 2, 2, 2, 2, 1, 0, 2, 1, 1, 0, 1, 0, -1, -3, -2, 0, 1, 2, 3, 4, 4, 3, 1, 0, -1, -2, -2, -2, -3, -4, -1, 1, 1, 2, 2, 0, 0, 0, 1, 0, 0, 1, 0, 0, -2, -3, -2, 0, 1, 3, 4, 4, 4, 2, 0, 0, -2, 0, -2, -2, -3, -4, -1, 0, 1, 1, 0, 0, 1, 0, 1, 1, -1, 0, 0, 0, -1, -3, -2, 0, 1, 3, 2, 2, 2, 0, 0, 0, 0, -1, 0, -1, -1, -3, -1, 0, 0, 1, 1, 2, 1, 1, 3, 0, 0, 1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -2, -2, 0, 0, -1, -1, -2, 0, 1, 1, 1, 1, 1, 2, 3, 2, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, -1, -1, -1, 0, -2, -2, 0, -1, 0, 0, 1, 1, 1, 1, 1, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -2, -2, -2, 0, -1, -2, -2, -1, -1, 0, 1, 1, 0, 1, 0, 1, 1, 3, 1, 2, 1, 1, 0, 0, 0, 1, 0, -1, -2, -1, -2, -3, -2, -2, -2, -1, 0, -2, -2, -1, -1, 0, 0, 0, 1, 1, 0, 1, 2, 3, 2, 1, 1, 0, 0, 0, -1, -1, 0, -2, -3, -2, -3, -2, -2, -2, -2, 0, -1, -3, -4, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 2, 3, 0, 0, 0, -1, -2, -3, -4, -3, -3, -3, -3, -2, -3, -1, -1, -1, 0, 0, -2, -3, -1, 1, 1, 3, 1, 3, 1, 1, 0, 1, 2, 2, 0, -1, 0, -1, -2, -4, -5, -3, -4, -3, -1, -2, -2, -1, -1, 0, 0, -1, -2, -2, 0, 0, 2, 2, 2, 3, 1, 1, 2, 1, 1, 0, -1, 0, 0, -2, -3, -4, -4, -4, -3, -1, -1, -2, 0, 0, 0, 1, 0, 0, -2, -1, 0, 2, 3, 3, 3, 2, 1, 0, 1, 1, 1, 0, 0, -1, 0, -1, -2, -1, -2, -1, -2, 0, 0, 0, 1, 1, 1, 0, 2, 0, 0, -2, 0, 2, 4, 2, 1, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 2, 2, 2, 1, 2, -1, -2, 0, 1, 3, 0, 0, -1, -2, -1, -1, -1, -2, -1, -1, 0, 0, 2, 1, 3, 3, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, -1, 0, 1, 0, 0, -2, -2, -2, -3, -2, -4, -3, -3, -1, -1, -1, 1, 0, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 1, 1, 0, 1, 2, 1, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 2, 4, 4, 5, 3, 3, 3, 3, 4, 3, -1, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 1, 1, 4, 4, 4, 4, 5, 4, 3, 3, 5, 4, 2, -1, 1, 1, 0, 0, 1, -1, -1, 0, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 2, 4, 3, 4, 3, 3, 3, 2, 0, 0, 1, 0, 0, 1, -1, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 2, 3, 3, 2, 3, 2, 2, -1, 0, 1, 0, 1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 2, 3, 2, 2, 2, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -2, 0, 1, 0, 1, 1, 2, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 2, 1, 1, 0, 1, 0, 1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 2, 0, 1, 0, 0, -1, 0, 0, 1, 2, 1, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 1, 3, 0, 1, 0, 0, -1, 0, 1, 0, 1, 1, 1, 1, 2, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 1, 0, 2, 0, 0, 0, 1, 3, 3, 2, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 2, 1, 0, 1, 2, 1, 1, 0, 2, 3, 1, 2, 3, 0, 0, -1, -1, 0, 0, 1, 0, 1, 1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 3, 1, 0, 1, 1, 2, 1, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 2, 1, 1, 1, 2, 1, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -2, 0, 1, 0, 0, 0, 1, 2, 1, 2, 3, 2, 2, 2, 3, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, 0, 1, 0, 1, 0, 2, 3, 2, 2, 2, 1, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, 0, 0, 1, 0, 0, 0, 0, 2, 2, 1, 2, 0, 1, 1, 2, 2, 1, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 1, 0, 0, 2, 2, 2, 2, 1, 0, 0, 1, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 0, 1, 2, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 2, 2, 1, 0, 0, 1, 0, 0, 1, 2, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 1, 1, 2, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 2, 0, 0, -1, -1, 1, 0, 0, 0, 1, -1, 0, 0, 1, 2, 2, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 2, 2, 0, 1, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, -2, -2, -1, -1, 0, 0, 0, 1, 2, 0, 2, 2, 0, 0, -1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 2, 0, 2, 1, 2, 0, -2, -1, -1, 0, 0, 0, 0, 1, 1, 1, 2, 3, 1, 1, -1, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 2, 1, 0, 1, 2, 1, 0, 0, -1, -1, 0, 1, 0, 1, 1, 1, 1, 3, 2, 4, 2, 0, 0, 1, 1, 2, 1, 0, 0, 0, 1, 2, 0, 1, 1, 1, 4, 2, 2, 1, 1, 0, 1, 1, 0, 1, 3, 1, 3, 2, 3, 4, 2, -2, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 2, 3, 3, 3, 2, 2, 1, 2, 1, 1, 3, 3, 2, 2, 4, 3, 4, 3, -2, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 1, 1, 1, 2, 2, 2, 2, 2, 2, 3, 3, -1, -2, 0, 0, -1, -2, -2, -2, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 2, 2, 2, 2, 1, 2, 1, 1, 2, 1, -2, -1, 0, 0, -1, -1, -3, -3, -2, -1, -3, -3, -2, -1, 0, 1, 1, 0, 0, 0, 2, 4, 4, 5, 6, 7, 4, 4, 6, 6, 5, 3, -2, 0, 2, 0, 0, 0, -2, -2, -2, -1, -1, 0, 0, 0, 2, 2, 2, 1, -1, 1, 2, 4, 4, 5, 6, 7, 7, 7, 7, 8, 7, 3, -1, 0, 2, 2, 1, 1, 0, -1, 0, 1, 1, 3, 3, 4, 3, 3, 1, 0, -1, -2, 0, 0, 0, 0, 2, 5, 5, 5, 6, 5, 4, 2, -2, 0, 2, 1, 2, 1, 0, 0, 0, 2, 2, 3, 4, 4, 3, 1, 0, 0, 0, -2, -2, -3, -3, -3, -1, 2, 3, 4, 4, 3, 3, 1, -2, 0, 2, 2, 3, 1, 1, 0, 1, 2, 1, 2, 2, 3, 1, 0, 0, 0, 0, -2, -4, -5, -5, -6, -3, 0, 1, 1, 1, 1, 0, 0, -3, 0, 1, 3, 3, 1, 0, 0, 0, 1, 1, 0, 1, 2, 1, 0, 0, 0, 0, -1, -4, -4, -4, -4, -2, 0, 0, 0, 0, 0, -1, -2, -2, 0, 2, 2, 2, 1, 1, 0, 2, 2, 1, 0, 1, 1, 0, 1, -1, -1, 0, -2, -3, -3, -4, -4, -1, -1, -1, -1, -1, -2, -3, -3, -2, 0, 2, 3, 3, 1, 1, 1, 3, 3, 3, 0, 0, 0, 0, 1, 0, -1, -1, -2, -2, -2, -1, -3, 0, 0, 1, -1, -2, -3, -3, -2, -1, 0, 1, 2, 3, 3, 2, 1, 2, 3, 3, 2, 0, 0, 0, 0, -1, -2, -2, -1, -2, 0, 0, -1, 0, 0, 0, 0, -2, -3, -4, -3, -1, 0, 1, 3, 3, 2, 2, 1, 3, 4, 4, 2, 2, 0, 0, 0, -2, -1, -1, -1, -1, 0, 1, 1, 1, 0, 1, 0, -1, -2, -3, -3, -1, 0, 2, 2, 4, 2, 2, 2, 5, 5, 4, 2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, -2, -3, -3, -2, 0, 1, 4, 4, 3, 2, 2, 6, 5, 3, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 3, 1, 1, 2, 0, 0, 0, 0, -1, -2, -2, 0, 0, 1, 3, 2, 2, 4, 3, 4, 0, 0, 0, -1, -1, -1, 0, 1, 2, 0, 2, 3, 2, 2, 1, 1, 2, 0, 0, -1, -1, -3, -2, 0, 0, 3, 3, 2, 3, 3, 4, 1, 0, 0, 0, -2, -2, -2, -1, 2, 1, 1, 2, 3, 4, 3, 2, 0, 1, 1, 0, -1, -2, -1, -3, -1, 1, 1, 2, 2, 1, 3, 3, 2, 0, 0, 0, 0, -2, -3, -1, 1, 1, 2, 3, 4, 4, 3, 2, 0, 0, 0, 0, -2, -2, -2, -2, -2, 0, 2, 2, 3, 1, 1, 3, 2, 0, 0, 0, 0, -2, -1, 0, 0, 3, 4, 3, 5, 5, 3, 2, 0, 0, 0, -1, -2, -3, -3, -2, -2, 0, 1, 0, 1, 0, 2, 2, 2, 1, 0, 1, 1, 0, -2, 0, 0, 2, 4, 4, 4, 3, 2, 1, 0, 0, -1, -3, -4, -2, -2, -3, -2, 0, 1, 0, 0, 0, 1, 2, 2, 0, 0, 1, 2, 0, -1, -1, 0, 1, 3, 3, 3, 3, 0, 0, 0, 0, -1, -1, -1, -2, -2, -3, -2, 0, 1, 0, 0, 0, 0, 4, 3, 0, 0, 3, 3, 0, -1, -1, 0, 0, 2, 1, 2, 0, 0, -3, -1, -1, -1, -1, -2, -2, -2, -3, -2, 0, 0, 0, 0, 0, 0, 2, 2, 1, 2, 3, 4, 2, 0, 0, 0, 1, 0, 0, 0, 0, -1, -3, -2, 0, 0, -1, 0, 0, -1, -2, -3, -1, 0, 1, 0, 0, 0, 3, 2, 3, 2, 4, 4, 1, 1, 0, -1, 0, 0, 0, -1, 0, -1, -1, -2, 0, -2, -1, 0, -2, -1, -2, -2, -1, 0, 0, 0, 0, 0, 1, 3, 4, 4, 4, 3, 3, 0, -1, -1, 0, 0, -2, -2, -1, -1, -1, -2, -2, -2, 0, 0, -1, -2, -3, -2, -1, 0, 0, 0, 0, -1, 1, 2, 3, 4, 3, 2, 3, 0, 0, -1, 0, -2, -3, -2, -2, -1, -2, -3, -2, -2, -1, -1, -1, -3, -3, -2, 0, 1, 1, 2, 1, 0, 1, 2, 3, 2, 3, 2, 2, 0, -1, -3, -2, -3, -4, -3, -3, -2, -1, -1, -2, -1, 0, 0, 0, -1, -3, -2, 0, 0, 3, 2, 2, 1, 0, 1, 2, 4, 4, 2, 1, 0, -1, -3, -4, -4, -4, -6, -4, -2, -2, -1, -1, -1, 0, 0, -1, -1, -2, 0, 1, 1, 3, 3, 3, 2, 1, 2, 2, 3, 2, 1, 1, 0, -1, -3, -4, -6, -6, -4, -3, -1, -1, 0, 1, 0, 2, 1, -1, 0, -2, 0, 3, 2, 2, 2, 2, 2, 1, 2, 3, 2, 3, 2, 1, 2, 0, -2, -3, -5, -4, -4, -1, 0, 1, 3, 3, 2, 2, 1, 1, 0, -1, 0, 3, 3, 2, 2, 1, 0, 0, 0, 2, 1, 2, 3, 3, 5, 5, 2, 1, 0, -1, 0, 0, 0, 3, 4, 4, 4, 3, 3, 2, 2, -1, 0, 2, 2, 0, 0, 0, -1, -1, 0, 0, 1, 1, 2, 3, 5, 5, 5, 4, 4, 2, 2, 2, 3, 5, 5, 4, 4, 5, 4, 4, 2, -2, 0, 2, 1, 0, -2, -3, -4, -3, -3, -1, 0, 0, 1, 2, 5, 6, 5, 7, 5, 4, 3, 2, 2, 3, 6, 6, 4, 5, 4, 5, 2, -2, 0, 0, 0, -2, -2, -4, -4, -4, -4, -3, -2, -2, -2, 0, 1, 2, 2, 3, 4, 2, 1, 3, 2, 1, 3, 3, 2, 3, 2, 3, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -4, -4, -3, -4, -2, -2, -2, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, 0, 0, 1, 0, 0, 0, 0, -2, -1, -2, -3, -3, -4, -4, -3, -2, -2, -2, -3, -2, -1, -1, -1, 0, -1, -1, -1, -2, -4, -4, -4, -3, 0, 1, 3, 0, 1, 1, 1, 0, 0, 0, -2, -2, -3, -4, -2, -1, -3, -2, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, -3, -4, -5, -3, 1, 1, 3, 3, 2, 2, 2, 2, 2, 1, 1, 0, -2, -2, -3, -1, -1, -1, -2, -1, -1, 0, -1, 0, 1, 1, 2, 0, -2, -3, -4, -3, 0, 1, 3, 1, 3, 4, 3, 2, 2, 2, 0, 0, 0, -2, -2, -2, -1, -2, -3, -1, -2, -1, 0, 0, 0, 2, 2, 0, 0, -2, -4, -2, 1, 0, 3, 3, 3, 3, 4, 4, 2, 2, 0, 0, 0, 0, 0, -1, 0, -2, -1, -2, -2, -4, -3, -1, 0, 1, 0, 0, 0, -2, -5, -2, 0, 0, 5, 3, 3, 3, 4, 3, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -4, -2, 0, 0, 0, 0, -2, -4, -4, -1, 0, 1, 3, 2, 3, 3, 2, 1, 1, 1, 1, 2, 2, 1, 2, 2, 1, 0, 0, 0, 0, -3, -3, 0, 0, -1, 0, 0, -2, -3, -4, -1, 0, 0, 3, 2, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 1, 1, 0, 1, 1, 1, 0, 0, -1, -1, 0, 0, -2, -2, -4, -5, -3, 1, 0, 3, 2, 1, 0, 0, 0, 0, 0, 1, 3, 1, 1, 0, 1, 0, 1, 0, 2, 2, 0, 1, 0, -1, -2, -2, -2, -2, -4, -4, -3, 0, 0, 2, 1, 0, -1, -1, 0, 0, 0, 1, 4, 3, 1, 1, 1, 2, 1, 0, 2, 2, 3, 1, 0, 0, 0, -1, -2, -4, -4, -6, -3, 0, 1, 1, 0, 0, 0, -2, -1, 0, 1, 2, 3, 3, 2, 1, 0, 1, 0, 1, 3, 2, 1, 2, 2, 0, 0, -1, -2, -3, -5, -4, -3, 0, 0, 1, 0, 0, -1, -2, -2, 0, 0, 1, 2, 2, 0, 0, 0, 0, 1, 0, 2, 1, 1, 1, 1, 1, 0, 0, -2, -2, -4, -6, -2, 0, 0, 1, 0, 0, -1, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 3, 2, 1, 1, 1, 1, -1, -2, -4, -5, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 0, 2, 1, 0, 0, -2, 0, 0, 0, 1, 2, 2, 4, 2, 1, 0, 0, 0, -2, -4, -4, -2, 0, 0, 2, 0, 1, 0, 0, 0, 2, 1, 1, 0, 1, 0, -1, -2, 0, 1, 1, 1, 3, 3, 3, 3, 2, 1, 0, 0, -2, -4, -4, -2, 0, 0, 2, 2, 1, 0, 0, 1, 2, 2, 1, 0, 1, 0, 0, -1, -1, 2, 3, 4, 3, 5, 4, 2, 1, 1, 0, -1, -2, -4, -4, -2, 0, 0, 3, 2, 0, 0, 0, 0, 1, 2, 1, 2, 0, 0, -3, -1, -2, 1, 2, 3, 5, 3, 3, 4, 2, 0, 1, -1, -1, -2, -3, -2, 0, 0, 2, 1, 1, 2, 1, 0, 2, 1, 1, 1, 1, -2, -2, -3, -1, 0, 1, 3, 4, 4, 3, 2, 1, 1, 0, 0, -2, -3, -3, -2, 0, 0, 2, 2, 1, 1, 1, 2, 0, 1, 1, 1, 0, -1, -1, -1, -1, 1, 2, 4, 4, 1, 1, 2, 2, 0, 1, 0, -1, -2, -4, -3, 0, 0, 1, 1, 0, 1, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 3, 3, 0, 0, 1, 0, 0, 0, 0, -1, -3, -5, -2, -1, 0, 0, 1, 0, 0, 2, 2, 2, 1, 0, 0, 0, 1, 1, 1, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, -4, -4, -2, -1, -1, 0, 0, 0, 0, 2, 1, 2, 0, 0, 0, 0, 1, 2, 3, 3, 2, 1, 1, 2, 0, 0, 0, 0, -1, 0, 0, -1, -4, -4, -3, 0, -1, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 1, 0, 0, 0, 0, -1, -1, -2, 0, -2, -3, -5, -4, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 1, 2, 2, 1, 0, 1, 0, -1, 0, -2, -1, -2, -3, -6, -4, 0, 0, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 0, 1, 1, 0, 0, 0, -1, 0, -1, -3, -5, -3, 0, 0, 3, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, -2, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -4, -5, -2, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -3, -3, -3, -2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -3, -4, -2, 0, 0, 4, 2, 0, 0, 0, -1, 0, 0, -1, -1, -2, -3, -3, -4, -4, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -5, -2, 0, 0, 4, 2, 0, 0, -1, 0, 0, 0, 0, -1, -2, 0, -2, -3, -2, -3, -1, -2, -1, 0, 0, 0, 0, -2, 0, -1, -3, -3, -4, -3, 0, 0, 2, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, -2, 0, -3, -2, -1, -1, -1, -1, 0, 0, 0, -2, -2, -3, -3, -3, -3, -5, -2, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, -1, -1, -1, -1, -1, 0, -1, -1, -2, -1, -1, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, -2, -1, -2, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, -2, -1, -3, -3, -3, -3, -3, -1, 0, 0, 0, -1, -2, -1, -1, 0, 0, -2, -1, -2, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -2, -2, -3, -2, -4, -4, -3, -5, -3, -3, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -3, -4, -4, -3, -1, -1, 0, 0, -1, 0, -1, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, -1, -3, -3, -4, -1, -1, 0, 0, -1, -1, -1, -1, -1, -2, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 3, 1, 0, -1, -3, -2, -1, 0, 1, -1, -2, 0, -1, -1, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 2, 3, 3, 1, 2, 0, -2, -2, 0, 0, 1, 0, -2, -2, -2, -1, -2, 0, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 2, 3, 2, 3, 3, 3, 0, 0, -1, 0, 0, 1, 0, -2, -2, 0, -2, 0, 0, 0, -1, -2, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 3, 3, 1, 2, 2, 3, 2, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, -1, -1, 0, -1, -1, 0, -1, -1, -2, -2, -2, -1, 0, 0, 0, 0, 1, 3, 3, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -1, 0, -2, -2, -1, -1, -1, -2, -3, -1, -1, 0, 0, 1, 1, 0, 1, 2, 1, 1, 2, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, -2, 0, -1, 0, -1, -1, -1, -2, 0, -2, -2, 0, -1, 0, 0, 0, 2, 1, 2, 1, 1, 1, -1, 0, 0, 0, -1, -1, 0, -1, -2, -1, -1, -1, 0, -1, -2, -2, -1, 0, -1, -1, -2, -1, 0, -1, 1, 0, 1, 2, 1, 1, 0, 0, -1, -1, -1, 0, 0, -1, -1, -2, -1, -2, -1, -1, 0, 0, -2, -2, -1, -1, -1, -2, -1, -2, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, -2, -1, -1, 0, 0, -1, -2, -1, -2, -1, -2, -2, -1, 0, -1, -1, -1, 0, -1, -3, -2, -2, -3, -2, -2, 0, 0, 2, 1, 2, 0, 1, -2, -1, 0, 0, 0, -1, -1, 0, -2, -1, -1, -2, -1, -1, 0, 0, 0, -1, -2, -3, -1, -2, -2, -2, -2, 0, 0, 1, 1, 2, 2, 0, 0, -1, 0, 0, 0, 0, -1, -1, -3, -2, -2, -2, -1, 0, 0, 1, 0, -1, -1, -1, -1, -2, 0, -1, 0, -1, 0, 1, 1, 1, 2, 0, 0, -2, 0, 0, 0, -1, -1, -2, -2, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 2, 2, 0, -1, -1, -1, 0, 0, -2, -1, -2, -3, -3, -2, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 2, 0, 0, -2, -1, -1, 0, 1, 0, -2, -2, -1, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, -1, -1, 0, -1, 0, -2, -2, -2, -2, -2, -2, -1, 0, 0, 0, -1, 0, 0, -1, -2, -1, 0, 1, 0, 0, 0, 0, 1, 2, 2, 2, 0, -2, -2, 0, -1, -1, -1, -2, -2, -3, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, 0, 0, 2, 2, 3, 1, 2, 0, -3, -1, -1, 0, 0, -2, -2, -1, -1, -3, -3, -1, -2, -1, 0, 0, 0, 0, -1, -2, -2, -1, -2, 0, 0, 0, 0, 1, 3, 2, 2, 0, -2, -3, -1, 0, 0, -2, -1, -3, -2, -1, -3, -3, -2, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 1, 0, -2, -2, -1, 0, 0, -2, -2, -1, -2, -1, -1, -2, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 1, 1, 2, 2, 1, 2, -1, -1, -3, -1, 0, 0, -1, -2, -1, -2, -2, -1, -1, -2, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, -2, -2, -2, 0, 0, -1, -1, -1, -1, -1, -2, 0, 0, 0, -3, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, -1, -3, -3, -2, -1, 0, -3, -1, -2, -1, -2, -1, 0, 0, -1, -2, -2, -1, -1, 0, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, -4, -3, -2, 0, -1, -2, -2, -1, -1, -1, -1, -1, -2, -2, -2, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -3, -5, -2, 0, -1, -2, -2, -1, -1, -2, -2, -1, 0, -1, -2, -3, 0, 0, -1, -1, 0, -1, 0, 0, -1, -2, -2, -2, -2, -2, -2, -3, -5, -3, -2, -1, 1, -1, -3, -2, -1, -2, -1, -1, 0, -1, -2, -1, -2, -1, -1, -1, 0, -2, -1, -2, -1, -2, -2, -3, -3, -4, -3, -5, -5, -5, -3, -1, 2, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, -1, -1, -2, -2, -2, -3, -2, -2, -2, -3, -3, -4, -4, -4, -6, -3, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -3, -1, -2, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, -2, 0, -1, -1, -2, 0, 2, 1, 2, 0, 0, 1, 0, 0, 0, -1, -3, -3, -3, -1, -1, -1, -1, -2, 0, 0, 0, 0, -1, 0, -1, 0, 0, -2, -1, -2, -2, -2, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -2, -1, -1, -2, -3, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -3, -4, -2, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -3, -2, 0, 2, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, -3, -3, -1, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, -1, -2, -3, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 1, 1, 1, 1, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -2, -3, -1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -3, -3, -2, 0, 0, 2, 1, 1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 2, 0, 0, 0, 1, 1, 0, -1, -1, 0, -1, -3, -1, 0, 1, 0, 0, 0, -2, -2, -1, -1, 0, 0, 0, 1, 2, 2, 1, 2, 1, 1, 2, 1, 2, 2, 2, 1, 0, -1, 0, 0, -3, -4, -2, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, 1, 0, 2, 2, 2, 2, 2, 2, 1, 1, 2, 2, 2, 2, 2, 0, 0, 0, -1, -2, -4, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 1, 1, 3, 1, 1, 2, 2, 2, 2, 1, 1, 3, 2, 2, 1, 0, -1, -2, -1, -4, -4, -2, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 2, 1, 3, 2, 3, 3, 2, 1, 0, 0, -2, -4, -5, -2, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 3, 2, 3, 1, 0, 1, -1, -2, -4, -4, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 1, 2, 1, 0, 2, 1, 3, 1, 3, 1, 1, 0, 0, -2, -3, -4, -1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 2, 2, 2, 3, 3, 2, 1, 1, 0, 0, 0, -3, -4, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 2, 0, 0, 1, 0, 0, 2, 4, 3, 2, 3, 3, 1, 1, 0, 0, 0, -2, -5, -2, 1, 1, 0, 0, 0, 0, -1, 0, -1, 1, 1, 0, 2, 1, 0, 0, 0, 2, 3, 3, 3, 3, 2, 1, 1, 1, 0, 0, -1, -2, -5, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 1, 2, 3, 2, 1, 1, 0, 0, 1, 1, -1, 0, -1, -3, -1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 3, 2, 2, 1, 2, 1, 0, 1, 0, 1, 0, 0, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 3, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, -2, -3, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 2, 0, 2, 0, 0, 1, 1, 0, 0, 0, 0, -2, -3, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 1, 0, 1, 1, 0, 1, 0, 0, 0, -1, -4, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 3, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, -4, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 1, 1, 2, 0, 0, 0, 1, 0, 0, 0, 0, -3, -4, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 1, 0, 1, 1, 1, 1, 0, 0, 0, -1, -2, -4, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 1, 2, 1, 1, 1, 2, 2, 1, 0, 0, -2, -2, -5, -1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, -1, -1, -1, -2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -2, -4, -5, -2, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -2, -2, -1, -1, -2, -2, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, -1, -2, -6, -1, 2, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, -2, -2, -1, -2, -2, -1, -2, -1, -1, 0, 0, 0, -1, -1, -2, -1, -2, -2, -4, -6, -2, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -2, -1, -2, -1, -1, -1, -2, -1, -1, -1, -1, -2, -3, -3, -3, -3, -4, -5, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, -1, -1, 0, -2, -1, -1, -1, -2, -3, -3, -2, -4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -1, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, -1, -2, -1, 0, 0, -2, -3, -4, -3, -5, -7, -9, -9, -9, -9, -7, -7, -3, -3, -3, 0, 1, 1, 3, 1, 1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, -3, -3, -4, -5, -5, -5, -7, -6, -6, -6, -6, -4, -3, -2, -2, 0, 1, 2, 2, 2, 2, 2, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, -3, -4, -4, -5, -4, -4, -4, -5, -4, -5, -4, -3, 0, 0, 0, 1, 3, 3, 1, 2, 3, 2, 0, 0, 1, 0, 0, -1, 0, 0, 0, -3, -2, -3, -4, -3, -4, -4, -5, -4, -5, -4, -4, -3, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 1, 2, 0, 0, 0, -2, -1, 0, 0, -2, -3, -3, -2, -2, -4, -4, -5, -6, -6, -4, -5, -3, -2, -2, -1, -1, 0, -2, -2, 0, 0, 1, 1, 2, 2, 0, -1, -2, -1, 0, 1, -2, -1, -3, -2, -1, -3, -4, -5, -5, -5, -3, -2, -4, -1, -1, -2, -2, -3, -3, -4, -3, -3, 0, 0, 0, 0, -1, 0, -2, -2, 0, 0, -1, 0, 0, -2, -1, -1, -2, -3, -4, -4, -1, -2, -1, -1, 0, -1, -3, -4, -4, -4, -5, -2, -1, -1, 0, -2, 0, -1, -1, -1, -1, 0, -1, -2, -2, -2, -3, -3, -2, -2, -4, -3, -2, -2, -1, -1, -1, 0, -1, -2, -4, -4, -4, -3, -2, -2, -2, -2, -1, 0, -1, 0, 0, 0, -1, -2, -2, -2, -4, -3, -3, -3, -4, -4, -5, -2, -1, -1, -1, 0, 0, 0, -3, -5, -4, -4, -4, -3, -1, -1, 0, 0, -1, -1, -1, -1, -2, -3, -2, -3, -4, -3, -3, -3, -3, -2, -3, -2, 0, -1, -1, -3, -1, -2, -3, -4, -4, -4, -4, -4, -4, -3, -2, -1, -2, -1, 0, -2, -2, -2, -4, -3, -4, -2, -3, -1, -2, -2, -1, -2, 0, 0, -3, -2, -4, -5, -6, -5, -2, -3, -4, -5, -5, -4, -3, -2, -2, -2, 0, 0, -2, -3, -5, -4, -6, -6, -5, -3, -4, -2, -1, -2, -2, -2, -1, -2, -3, -5, -7, -8, -6, -5, -5, -4, -4, -4, -4, -2, -4, -2, 0, -1, -2, -3, -4, -3, -4, -3, -4, -3, -3, -3, -2, -3, -4, -3, -3, -3, -5, -8, -10, -10, -8, -7, -6, -5, -3, -4, -3, -2, -3, -1, 0, -1, -3, -3, -3, -3, -3, -3, -2, -2, 0, -1, -3, -4, -5, -4, -2, -4, -4, -6, -8, -9, -6, -6, -5, -4, -4, -2, -1, -2, -2, -3, 0, 0, -3, -1, -3, -3, -2, -2, -1, -2, 0, -2, -2, -2, -2, -3, -2, -3, -6, -5, -6, -7, -5, -6, -5, -3, -4, -2, -3, -1, -4, -3, -1, 0, -1, -2, -1, -2, -2, -3, -2, -2, -2, -2, -1, -2, -2, 0, 0, -2, -3, -5, -5, -5, -6, -5, -4, -3, -3, -3, -3, -3, -4, -3, 0, 0, -1, -2, -3, -3, -3, -4, -3, -2, -2, -2, -1, 0, 0, -1, -1, -3, -3, -4, -4, -4, -4, -3, -4, -4, -4, -4, -3, -4, -4, -2, 0, 0, -2, -2, -4, -4, -5, -5, -3, -2, -2, -1, 0, -1, -2, -2, -1, -3, -3, -3, -3, -2, -4, -4, -3, -2, -3, -2, -3, -4, -4, -3, 0, 0, -2, -2, -5, -4, -3, -5, -4, -4, -2, -2, -2, -3, -4, -5, -3, -1, -2, -3, -4, -2, -3, -3, -2, -1, -1, 0, -2, -2, -4, -1, 0, -1, -3, -3, -3, -4, -4, -3, -4, -4, -2, -2, -2, -1, -3, -3, -2, -2, -2, 0, -1, -1, -2, -2, -1, -1, -1, -1, -1, -1, -2, 0, 0, 0, -1, -3, -4, -4, -5, -5, -4, -4, -5, -3, -3, -1, -2, -2, 0, 0, -1, 0, -1, -2, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, 0, -1, -3, -3, -2, -4, -4, -5, -4, -4, -4, -3, -4, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -3, -3, -3, -4, -4, -5, -5, -5, -4, -5, -3, -3, -3, -2, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, -4, -4, -3, -4, -6, -6, -5, -5, -4, -5, -3, -2, -1, 0, 0, 1, 2, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, -1, -1, 0, -2, -3, -4, -3, -4, -5, -5, -4, -5, -2, -3, -3, -1, 0, 0, 0, 0, 1, 0, 2, 1, 1, 2, 1, 2, 1, 0, 0, -1, -3, -2, 0, -2, -3, -4, -3, -2, -5, -4, -5, -3, -4, -3, -4, -2, 0, 0, 0, 0, 0, 1, 3, 2, 2, 3, 2, 2, 1, 0, -1, -1, -3, -2, 0, -1, -3, -3, -2, -3, -3, -3, -3, -3, -4, -4, -5, -4, -4, -4, -2, -3, -1, 1, 2, 2, 2, 1, 2, 0, 1, 0, -1, -1, -3, -1, 0, 0, -2, -2, -2, -2, -2, -2, -2, -3, -3, -4, -5, -5, -4, -3, -4, -2, -1, 0, 1, 3, 3, 2, 2, 1, 0, 0, 0, -1, -2, -1, 0, 2, 2, 1, 2, 1, 1, 1, 0, 1, 1, 0, 0, -2, -1, -2, -3, -1, 0, 0, 1, 1, 1, 1, 0, 0, -1, -2, -2, -1, -1, -2, 3, 6, 3, 1, 1, 0, 0, -1, 0, 0, 0, -3, -3, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, -1, 0, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -2, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, -2, -2, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, -2, -1, -1, -2, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, -2, -1, 0, -1, -2, -2, -1, -1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -2, -2, -2, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -1, 0, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -2, -1, -2, -1, -2, -1, -1, 0, 1, 0, 0, -1, -1, 0, 2, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, -1, 0, -2, -2, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -2, -2, -1, -1, 0, 0, 0, -1, -1, 0, 1, 0, 0, -1, -1, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, -1, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -2, -1, -1, -1, -1, -2, -2, -2, -3, -2, -3, -1, -3, -4, -1, -2, -1, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, -2, -2, -2, 0, -2, -1, -2, -3, -1, -2, 0, -1, -1, -1, -3, -2, -2, -3, -4, -4, -2, 0, 2, 0, 0, 0, -1, 0, -1, 0, 0, -1, -2, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -3, -4, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 0, -1, -1, -3, -2, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, -2, -2, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, -2, -1, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 0, -1, 0, -2, -2, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 2, 2, 1, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, -1, -2, -1, -1, -1, -1, 0, 0, 1, 0, 1, 2, 1, 1, 2, 2, 1, 2, 1, 2, 0, 0, 0, 0, -2, -2, -1, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 2, 1, 2, 3, 2, 2, 1, 0, 1, 0, 0, -1, -1, -2, -3, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 2, 0, 0, 2, 2, 1, 0, 1, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 2, 1, 2, 1, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 2, 0, 1, 1, 0, 0, 0, 0, -1, -2, -2, 0, 0, -1, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, -2, -1, -2, -1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, -1, -1, -1, -2, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, -2, -2, -2, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 2, 0, 0, 0, 2, 1, -1, -1, -1, -2, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 1, 0, -1, -1, -1, -1, 0, 0, 0, -1, -1, -1, 0, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 1, 1, 1, 0, 0, -1, -2, -2, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 1, 2, 2, 2, 2, 2, 1, 1, 0, 1, 0, 0, -2, -2, -3, 0, 0, -1, 0, -1, -1, -1, 0, 0, -2, 0, -2, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 0, -1, -1, -1, -3, -3, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, -3, -2, -3, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -2, -2, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, -2, -3, -3, -3, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, -1, -1, -2, -2, -2, -2, -1, -1, -1, -2, 0, 0, 0, -2, 0, -2, -2, -2, -3, -3, -1, 0, 0, 0, 0, -1, -1, -2, -2, 0, -1, 0, 0, -1, -3, -2, -1, -2, -3, -3, -1, -3, -2, -2, -1, -2, -2, -4, -4, -3, -4, -4, -4, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, -2, -2, -2, -2, -1, -1, -3, -2, -3, -3, -2, -3, -1, 1, 0, 0, 0, 0, 0, -1, -1, -1, -2, -3, -3, -2, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -2, 0, 2, 1, 0, 0, 0, 0, -1, -1, 0, -2, -2, -1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -2, -2, -1, -2, -2, -1, -3, -4, 0, 1, 0, -1, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, -2, -3, -3, 0, 2, 0, 0, 0, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -4, 0, 2, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -2, 0, 1, 1, 0, 1, 1, 2, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, -1, 0, 1, 0, -2, 0, 1, 0, 1, 0, 0, 0, -1, -2, -3, 0, 2, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, -1, -1, -1, -2, 0, 2, 2, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, 0, 2, 1, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 2, 2, 0, 1, 1, 2, 2, 1, 2, 2, 0, 0, 0, 0, 0, 0, -1, -3, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 2, 0, 0, 1, 1, 3, 1, 3, 2, 1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 2, 0, 1, 1, 0, 0, 0, 2, 2, 3, 3, 2, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, 1, 0, 0, -1, -1, 0, -1, 0, 1, 1, 2, 1, 0, 1, 0, 1, 1, 0, 1, 1, 3, 3, 2, 1, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 1, 1, 2, 1, 0, 0, 1, 0, 0, 2, 3, 3, 2, 3, 2, 1, 0, 0, 0, 0, -1, -3, 0, 1, 0, -1, 0, -1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 1, 1, 1, 0, 1, 1, 3, 2, 2, 1, 0, 0, 0, 1, 0, -2, -3, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 2, 3, 3, 3, 2, 1, 0, 1, 1, 0, 0, -1, -3, 0, 2, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 2, 1, 1, 3, 3, 4, 4, 3, 0, 1, 1, 0, 0, 0, -2, -3, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 3, 4, 3, 2, 2, 2, 2, 0, 0, 0, 1, 0, -2, -4, 0, 1, 2, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, 0, 1, 2, 3, 2, 2, 2, 2, 3, 1, 0, 1, 0, 0, 0, -2, -4, 0, 2, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, -2, -1, 1, 3, 3, 3, 3, 1, 0, 0, 1, 0, 0, 0, 1, -2, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, -2, 0, 1, 2, 3, 1, 1, 2, 0, 1, 2, 0, 1, 0, 0, -1, -4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 1, 3, 2, 3, 3, 1, 0, 0, 1, 2, 0, 0, -1, -3, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 3, 1, 0, 1, 2, 2, 1, 1, 0, -1, -3, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 2, 1, 1, 1, 0, 3, 2, 1, 0, 1, 1, 1, 0, 0, -3, -2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 2, 1, 1, 1, 2, 0, 2, 1, 2, 0, 0, 0, 0, 0, -1, -2, -4, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 3, 3, 1, 1, 2, 0, 2, 2, 0, 0, 0, 1, 1, 0, -1, -4, -4, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 2, 0, 1, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, -2, -3, -4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 1, 1, 0, 1, 1, 0, 0, 0, -1, -3, -3, 0, 2, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 1, 0, -1, 0, 0, 2, 1, 1, 2, 1, 1, 1, 0, 0, -1, -2, -4, -4, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 0, 0, 0, -1, 0, -1, 0, -3, -5, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, -2, -1, -3, -4, 0, 3, 2, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, -3, -3, -3, -3, -3, -2, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, 0, 2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 2, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 1, 1, 0, 2, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 1, 1, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 0, 1, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 1, 2, 0, 0, 1, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 3, 3, 1, 2, 0, 1, 0, 1, 1, 2, 0, 1, 0, 0, 1, 1, -1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 4, 3, 2, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 3, 2, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, -1, -1, -1, 0, 0, 3, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 2, 2, 2, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 1, 2, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 2, 2, 0, 1, 3, 1, 1, 1, 2, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 1, 0, 4, 2, 3, 3, 2, 1, 0, 1, 2, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 2, 2, 1, 3, 2, 3, 3, 3, 2, 3, 3, 2, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 2, 3, 2, 1, 2, 2, 3, 4, 3, 2, 2, 2, 3, 0, -1, 1, 2, 1, 0, 0, 1, 0, -2, 0, 0, 0, 0, 0, -2, -1, 0, 0, 1, 4, 2, 1, 2, 2, 2, 3, 3, 4, 3, 3, 3, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 2, 3, 2, 2, 1, 1, 3, 2, 3, 4, 4, 2, 3, 1, 0, 1, 2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -2, 0, 0, 1, 2, 1, 2, 3, 1, 2, 1, 1, 2, 3, 2, 3, 3, 2, 0, 2, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 1, 3, 2, 1, 2, 3, 2, 1, 2, 4, 3, 2, 3, 4, 2, 1, 1, 1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 2, 3, 1, 1, 4, 3, 2, 2, 3, 5, 3, 1, 3, 4, 1, 2, 1, 1, 0, -1, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 3, 2, 3, 3, 0, 3, 3, 2, 3, 4, 6, 3, 1, 3, 4, 1, 2, 2, 1, 0, -2, 0, 0, 0, -1, 0, 0, -1, -2, 0, -1, 0, 2, 2, 4, 4, 2, 5, 4, 1, 2, 3, 4, 4, 2, 3, 4, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -2, 0, 1, 1, 4, 4, 3, 3, 2, 2, 3, 2, 5, 3, 2, 3, 4, 3, 2, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 4, 4, 4, 2, 1, 2, 2, 2, 5, 4, 1, 3, 3, 3, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, 0, 0, 0, 2, 2, 4, 3, 2, 2, 4, 1, 2, 4, 1, 1, 1, 4, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 1, 1, 3, 3, 3, 3, 3, 3, 2, 3, 2, 1, 2, 2, 0, -1, 0, 1, 0, 0, 1, 0, -2, 0, -2, -1, -2, 0, 0, 0, -1, 1, 0, 0, 0, 2, 3, 2, 4, 3, 2, 2, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -2, -2, -2, -2, 0, 0, 0, -1, 0, 0, 1, 0, 1, 4, 4, 4, 2, 2, 2, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, -1, 1, 0, 0, 0, 0, 1, 0, 3, 4, 4, 4, 2, 2, 3, 1, 1, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 1, 1, 3, 5, 4, 3, 2, 3, 1, 0, 2, 2, 2, 0, 0, 1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 4, 4, 4, 3, 1, 2, 3, 0, 2, 3, 1, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 3, 2, 3, 2, 3, 1, 1, 1, 2, 2, 1, 0, 0, -2, -2, 0, 1, 0, -1, 1, 1, 0, -1, 0, -1, 0, 2, 0, 0, 1, 2, 1, 0, 2, 3, 3, 2, 1, 0, 1, 1, 0, 0, 0, 0, -2, -3, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, -2, 0, 3, 0, 0, 0, 1, 3, 2, 2, 0, 1, 1, 0, -1, 0, 0, 0, -2, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, -1, 0, 1, 0, -2, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, -2, 0, 2, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -1, 0, -2, 0, 1, 0, 1, 0, 1, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -1, -2, 0, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -2, -1, -2, -1, 0, 0, 0, 2, 2, 1, 1, 0, 0, -1, -1, -1, -3, -3, -2, -1, -1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 2, 2, 1, 1, 0, 0, 0, 0, 0, -2, -2, -2, -2, -1, 0, 0, 0, 0, 1, 1, 2, 1, 2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 2, 0, 1, 1, 1, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 2, 2, 1, 1, 0, 0, 0, -1, -1, -1, 2, 2, 2, 1, 1, 1, 2, 0, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 2, 0, 0, -1, -2, 0, 2, 3, 2, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, 1, 0, 1, 1, 1, 0, 0, -2, -1, 0, 1, 2, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, 3, 3, 3, 1, 1, 1, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, -2, 0, 2, 3, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, -2, -1, 0, 1, 1, 2, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 2, 3, 2, 1, 1, 0, 0, -1, -1, 0, -2, -3, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, -2, -2, -2, -2, -2, -1, 0, 1, 1, 0, 0, -1, 0, -1, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 2, 3, 1, 1, 1, 0, -1, -2, -1, -1, -3, -1, 0, 0, 0, 1, -1, -1, -1, -1, -1, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 1, 1, 2, 2, 2, 0, 0, 0, -1, 0, -2, -1, -1, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 2, 2, 2, 1, 1, 0, 0, 0, -2, -2, -1, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -2, -1, 0, -1, 0, 0, 1, 2, 2, 2, 2, 0, 0, 0, -2, -1, -2, -1, 0, 0, 2, 1, 2, 1, 0, 0, 0, 0, 0, 1, 1, 0, -1, -2, -1, -1, 0, 0, 1, 3, 1, 3, 1, 0, -1, -1, -2, 0, -1, -3, 0, 2, 2, 2, 1, 1, 0, -1, -1, 0, 1, 0, 1, 0, -1, -2, -1, 0, 1, 2, 2, 2, 2, 1, 0, 0, -1, 0, -1, 0, -1, -2, -1, 1, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, -2, 0, 0, 0, 1, 2, 1, 2, 1, 1, 1, 0, -1, 0, -1, 0, -2, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, 1, 2, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 1, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, -2, 0, 0, 1, 1, 0, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 3, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -3, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, -1, -1, -1, 0, 0, -2, 0, -2, -1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -3, -2, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, -3, -2, -2, -3, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -2, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -2, -1, -2, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 1, 3, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 1, 2, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, -2, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -2, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -2, -1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, -1, -1, -1, 0, -1, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, -1, 0, -1, -1, -1, -3, -3, -1, -1, -1, -1, 0, 0, 1, 0, 2, 1, 3, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -3, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, -1, 0, -1, -2, -1, -2, -1, 0, 0, 0, 0, 1, 0, 1, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -1, -1, -1, 0, 0, 3, 3, 1, 1, 0, -1, -1, -2, -2, -5, -5, -5, -2, -2, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, -2, -2, -2, 0, 2, 3, 1, 1, 0, -1, -1, -1, -3, -4, -4, -5, -3, -2, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -4, -2, 0, 1, 4, 2, 0, 0, 0, 0, 0, 0, -1, -3, -2, -2, -1, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -2, 0, 1, 3, 3, 2, 2, 2, 0, 0, 0, 0, -2, -2, -2, -1, -1, 0, 0, -2, -2, -1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -3, -2, 0, 2, 3, 2, 3, 2, 1, 0, 1, 0, 0, -2, -2, -1, 0, 0, 0, 0, -2, -2, -2, -1, -1, 0, 2, 1, 0, 1, -1, -1, -4, -4, -1, 1, 3, 3, 3, 3, 1, 2, 0, 0, -1, -2, 0, 0, -1, 0, 0, 0, -2, -1, -3, -4, -2, 0, 1, 0, 1, 0, -2, -3, -4, -2, 0, 1, 5, 3, 3, 3, 1, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, 0, -1, -2, -3, -3, -1, 0, 0, 0, 0, -2, -3, -4, -2, -1, 2, 4, 2, 3, 3, 1, 0, 0, 0, 1, 0, 0, 1, 2, 1, 0, 1, 1, 2, 1, 0, -1, 0, 0, 0, -1, -2, -2, -2, -5, -4, 0, 1, 3, 2, 1, 0, 0, -1, -2, 0, 0, 0, 1, 1, 1, 1, 2, 1, 1, 4, 2, 1, 1, 1, 0, 0, -1, -1, -2, -3, -5, -4, 0, 1, 2, 0, 1, 0, -2, -1, -1, 0, 1, 1, 2, 1, 0, 1, 2, 1, 2, 3, 3, 2, 3, 1, 0, 0, -2, -3, -4, -3, -4, -3, -1, 0, 1, 0, 0, -1, -1, -1, 0, 0, 1, 4, 2, 2, 0, 2, 1, 1, 1, 3, 2, 2, 3, 2, 1, 0, -2, -3, -5, -3, -4, -4, 0, 1, 1, 0, 0, -1, -1, -1, 0, 0, 2, 3, 2, 2, 1, 0, 0, 1, 2, 2, 2, 3, 2, 3, 2, 0, 0, -2, -4, -3, -4, -4, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 2, 2, 3, 2, 4, 2, 1, 1, 1, -2, -3, -4, -5, -4, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 2, 1, -1, 0, 1, 1, 1, 1, 2, 4, 4, 2, 2, 1, 0, 0, -3, -4, -4, -4, -1, 0, 2, 1, 0, 0, 0, -1, 0, 0, 0, 2, 1, 0, -1, -1, 0, 1, 1, 2, 4, 4, 4, 3, 2, 1, 0, -1, -4, -4, -5, -5, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 1, 2, 3, 5, 6, 4, 3, 3, 0, 0, -2, -3, -3, -4, -4, -1, 1, 3, 2, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, -2, 0, 3, 3, 4, 6, 5, 5, 2, 2, 1, -1, -1, -2, -2, -5, -3, -1, 0, 2, 1, 0, 1, -1, -1, 0, 1, 1, 1, 0, 1, 0, -2, 0, 2, 3, 3, 3, 3, 4, 2, 2, 1, 0, -2, -4, -3, -4, -4, -1, 1, 2, 2, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 2, 3, 4, 3, 3, 3, 2, 0, 1, 0, 0, -2, -2, -2, -4, -1, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 2, 2, 5, 3, 2, 3, 1, 1, 1, 1, -1, -1, -2, -3, -2, 0, 0, 1, 1, 1, 1, 0, 2, 2, 1, 0, 0, 2, 2, 1, 1, 2, 3, 3, 2, 1, 0, 1, 1, 1, 0, 0, 0, -2, -2, -3, -3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 2, 1, 2, 3, 2, 3, 0, 2, 1, 0, 1, 0, 0, -2, -1, -2, -2, -3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 2, 2, 3, 2, 3, 4, 2, 2, 1, 1, 0, -1, -2, 0, -1, -1, -3, -3, -4, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 1, 2, 1, 3, 3, 3, 3, 2, 1, 1, 0, 0, -1, 0, 0, -1, -1, -3, -3, -4, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 1, 2, 3, 3, 2, 1, 1, 0, 0, -1, -2, -2, -3, -2, -3, -3, 0, 0, 2, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 0, 0, 0, -1, -1, -2, -3, -4, -4, 0, 1, 3, 1, 1, 1, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, -2, 0, -2, -3, -3, -4, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, -1, -1, -2, -4, -3, -3, -3, -3, 0, 0, 0, 1, 2, 2, 0, 0, 0, -1, -2, -3, -3, -3, 0, 2, 2, 1, 1, 0, 0, 0, -1, -1, 0, -2, -1, -4, -2, -3, -2, -2, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -2, -2, -4, -3, 0, 2, 4, 1, 0, 0, 0, 0, -1, -1, 0, -2, -3, -3, -2, -2, -2, -1, -1, 0, 0, 0, 1, 0, 0, -2, -3, -3, -4, -2, -4, -3, 0, 1, 2, 1, 0, 0, -1, 0, -2, -2, -3, -2, -2, -3, -2, -1, -1, -1, 0, 0, -1, -1, 0, 0, -1, -3, -1, -3, -3, -3, -2, -2, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, -1, -1, -1, -2, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, -2, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 3, 3, 4, 3, 3, 3, 2, 2, 2, 1, 1, -1, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 2, 2, 2, 2, 3, 4, 3, 3, 2, 3, 3, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 1, 3, 4, 3, 3, 3, 5, 4, 3, 0, 0, 1, 1, 1, 1, -1, 0, 0, 1, 1, 2, 2, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 3, 3, 2, 3, 3, 3, 2, -1, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 1, 0, 0, 0, -2, -1, 0, 1, 2, 2, 2, 2, 2, 0, -2, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -2, -1, 0, 1, 0, 1, 2, 2, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 1, -1, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 0, 0, 0, 0, -1, -1, 0, 1, 1, 1, 2, 1, 0, 0, 0, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 2, 1, 2, 1, 0, 0, 0, -1, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, -1, -2, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 1, 1, 1, 2, 2, 1, 0, 1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, -2, -1, -2, 0, 0, 0, 0, 1, 2, 1, 0, 1, 2, 0, 0, 2, 1, 1, 1, 2, 1, 0, -1, 0, 0, 1, 2, 1, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 2, 3, 2, 1, 2, 2, 0, 0, 2, 1, 1, 1, 0, 1, -1, -2, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 3, 1, 2, 1, 3, 2, 0, 0, 0, 0, 0, 0, 0, 2, 0, -1, 0, 0, 0, 2, 2, 0, -1, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 2, 1, 1, 1, 0, 1, 0, 0, 0, 0, -2, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 0, 1, 0, 1, 2, 1, 1, 2, 1, 2, 1, 0, 0, 0, 0, 1, 0, -2, -1, 0, 0, 0, 1, 0, 0, 0, -1, -2, 0, 0, 2, 2, 0, 0, 0, 1, 2, 1, 2, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 1, 1, 2, 1, -1, 0, 0, 1, 0, 1, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 1, 0, -1, -1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, -1, 0, 0, 0, 0, 1, 2, 0, -1, -1, 0, 0, 0, -2, -1, 0, 0, 0, 0, -1, 1, 3, 1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 1, 2, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 1, 1, 0, -1, 0, 0, 0, 1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -2, 0, 0, 1, 2, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 0, -1, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 2, 0, 1, 1, 1, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 1, 1, 2, 0, 0, 3, 0, -1, -2, -2, -1, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 2, 0, 2, 2, 0, 2, 3, 2, 0, -1, -2, -1, 0, 0, 0, 1, 1, 1, 1, 2, 3, 2, 0, -1, 0, 1, 2, 2, 0, 0, 0, 0, 0, 2, 1, 1, 0, 1, 4, 2, 1, 0, -1, 0, 0, 0, 0, 1, 2, 2, 1, 3, 3, 4, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 3, 3, 2, 1, 1, 0, 1, 1, 0, 1, 3, 2, 1, 1, 3, 3, 0, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 1, 2, 0, 2, 2, 2, 2, 1, 0, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 2, 1, 3, 2, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 2, 2, 1, -1, 0, 0, -1, 0, -1, -2, -3, -1, 0, 1, 2, 0, -1, 0, 1, 1, 1, 2, 2, 1, 1, 0, 1, 2, 1, 0, 0, 4, 3, 3, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 3, 1, 0, -1, 0, 1, 1, 0, 2, 3, 2, 2, 1, 1, 2, 3, 1, 0, 3, 3, 3, 2, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 2, 2, 0, -2, -1, 0, -1, -1, 1, 1, 2, 1, 2, 1, 1, 1, 0, 0, 2, 3, 3, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 2, 3, 1, 0, 0, 0, -2, -1, -2, 0, 0, 1, 1, 2, 1, 1, 1, 0, 0, 3, 3, 4, 3, 1, 0, 0, 0, 0, 1, 0, 2, 1, 1, 2, 0, 0, 0, -2, -3, -2, -3, -2, 0, 1, 0, 1, 0, 1, 0, -1, 0, 3, 3, 4, 3, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, -1, -2, -3, -3, -3, -1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 3, 2, 2, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 1, 0, 0, -2, -1, -3, -1, 0, 2, 2, 2, 2, 1, 1, 1, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 1, 0, -2, -1, 0, -2, -3, 0, 0, 2, 2, 2, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 2, 0, 0, 0, 0, -3, -3, 0, 2, 2, 2, 2, 0, 0, 0, 1, 2, 1, 1, 2, 1, 1, 0, 0, 0, 0, -1, 0, 0, 2, 0, 0, 0, 0, 0, -2, -2, -2, -2, -1, 1, 1, 2, 2, 1, 1, 1, 2, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, -2, -2, 0, 1, 1, 1, 2, 1, 1, 1, 1, 1, 2, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, -1, -1, -2, -1, 0, 1, 0, 2, 1, 2, 0, 1, 2, 2, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 2, 1, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 2, 1, 1, 1, 1, 2, 0, 1, 0, 0, -2, -1, 0, 0, 0, 0, 2, 3, 2, 1, 2, 1, 0, 0, 0, -1, -2, -1, 0, 1, 1, 2, 1, 1, 0, 1, 2, 2, 2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 2, 1, 2, 1, 2, 1, 0, -1, -2, -1, -2, -1, 0, 1, 0, 1, 1, 2, 1, 0, 2, 2, 1, 0, 0, 0, 0, -2, -1, 0, 1, 2, 2, 2, 2, 2, 2, 0, 0, -2, -1, -2, -3, -2, -1, 0, 1, 1, 1, 0, 0, 0, 2, 0, 1, 0, 2, 0, 0, 0, -2, 0, 1, 2, 1, 3, 1, 2, 1, 0, 0, -1, -2, -3, -2, -3, 0, 1, 0, 0, 1, 0, 0, 0, 2, 2, 1, 0, 1, 1, 0, -2, 0, 1, 1, 1, 3, 2, 1, 0, 1, 0, 0, -1, -1, -1, -3, -1, -1, 1, 0, 1, 0, 1, 0, 2, 3, 2, 0, 1, 1, 1, 0, -2, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 2, 1, 1, 0, 0, -2, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -2, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 3, 2, 2, 1, 1, 2, 1, 0, 0, 1, 1, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, 1, 2, 3, 3, 3, 1, 1, 1, 0, 0, 1, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, -1, -2, -1, -1, 0, 0, 1, 0, 0, 1, 2, 1, 3, 3, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, -1, 0, -2, -1, -1, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 3, 2, 3, 2, 0, 0, -1, 0, 0, 0, 0, -1, -1, -2, -1, -2, -1, -1, -1, -1, 0, -2, -2, 0, 0, 1, 1, 1, 1, 0, 0, 0, 2, 2, 1, 0, 1, 0, 0, -1, -1, -1, -2, -1, -2, -3, -1, -1, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 2, 2, 2, 0, 0, 0, 1, 2, 1, 2, 0, 1, 0, -2, -1, -1, -3, -3, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 1, 2, 0, 1, 2, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 1, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 0, 2, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, 1, 1, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, -1, -1, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, -1, -1, -1, -3, -3, -2, -1, -1, -1, 0, 1, 1, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, -2, -2, -1, -3, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, -1, -3, -2, -3, -2, -3, -4, -3, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, -2, 0, -2, -2, -1, -1, -3, -4, -5, -4, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -3, -3, -4, -3, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, -3, -2, -2, 0, 0, 1, 0, 0, 1, 0, 1, 2, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -3, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 2, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -2, -3, -2, 0, 0, 0, 1, 0, 0, 1, 2, 2, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -3, -2, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 2, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -3, -2, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, -2, 0, 0, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, -1, 0, -1, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 1, 0, 0, 0, -2, -3, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, -1, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 1, 1, 1, 1, 0, -2, -2, -3, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 1, 2, 0, 1, 0, 0, 0, 0, -2, -3, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 2, 0, 0, 0, 0, -1, 0, 0, 1, 1, 2, 1, 1, 0, 0, 1, 1, 0, 0, -1, -2, -2, 0, 0, 0, 1, 1, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 2, 2, 2, 1, 2, 0, 0, 0, 0, 0, 0, -1, -1, -3, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 2, 0, 0, 0, 0, -1, -1, 0, 1, 1, 2, 2, 1, 0, 1, 1, 1, 0, 0, 0, -1, -3, 0, 0, 0, 0, 1, 0, 1, 1, 1, 2, 1, 1, 0, 0, -1, -1, -1, 0, 1, 0, 1, 2, 0, 0, 1, 1, 1, 0, 0, -1, -3, -2, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 1, 1, 0, -1, -2, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, -3, -2, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 2, 2, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -3, -3, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 1, 1, 0, 1, 2, 0, 0, 0, 0, -1, -1, 0, -2, -3, -3, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 2, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -2, -2, -4, -3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 2, 1, 1, 2, 2, 0, 0, 1, 0, 0, -1, -1, 0, -1, -2, -3, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -2, -2, -1, -2, -2, -3, -3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -2, -1, -1, -2, -2, -2, -2, -4, -3, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, -3, -2, -3, -3, -3, -3, -3, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, -1, 0, 0, -1, -1, -1, -2, -2, -2, -2, -1, -1, -2, -3, -3, -4, -3, -2, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, -2, -1, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 2, 2, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 1, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 3, 2, 2, 1, 0, -2, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 1, 1, 1, 0, 0, 2, 1, 0, 0, -1, 0, 3, 0, 1, 4, 2, 1, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 2, 0, -1, 0, 3, 1, 0, 0, -1, 1, 2, 0, 1, 2, 1, 1, 0, 0, -1, -2, -1, 0, -1, 0, 1, 1, 0, 0, 1, 2, 0, 2, 1, 0, -1, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -2, -2, -1, 0, -1, -1, 0, 2, 0, 0, 0, 2, 0, 2, 1, 0, -1, -1, 2, 1, 2, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, -1, 0, -2, -1, 0, 2, 2, 0, 1, 2, 2, 2, 1, 0, -1, 0, 2, 2, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 1, 1, 1, 0, 0, 2, 1, 2, 1, 0, 0, 2, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 0, 1, 0, 2, 2, 0, 1, 1, 3, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 1, 2, 3, 1, 0, 0, 1, 2, 1, 1, 2, 3, 3, 3, 1, 1, 1, 1, 0, 0, 0, 1, -1, 0, 0, -1, 0, -1, -1, -2, -1, 1, 1, 1, 2, 0, 0, 1, 2, 0, 1, 1, 2, 2, 3, 3, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, -2, 0, 0, -1, -1, 1, 0, 2, 1, 0, 0, 2, 1, 0, 1, 2, 1, 1, 3, 3, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 1, 0, 1, 1, 2, 0, 1, 1, 1, 0, 3, 3, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 2, 0, -1, 1, 1, 1, 1, 1, 1, 0, 0, 2, 2, 2, 1, 1, 2, 0, 0, 0, -1, -2, 0, 0, 0, -1, 0, 0, -1, 1, 0, 1, 1, -1, 0, 1, 1, 0, 1, 2, 4, 1, 1, 4, 4, 2, 1, 0, 1, 0, 0, 0, -1, -2, 0, 1, 0, -1, -2, -2, 0, 2, 1, 0, 2, 0, 1, 2, 0, 0, 2, 2, 3, 1, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 2, 1, 2, 0, 1, 1, 0, 2, 3, 1, 3, 3, 4, 3, 2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 1, 1, 2, 3, 1, 0, 2, 1, 1, 4, 3, 4, 5, 4, 3, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, 0, 0, 0, 1, 1, 2, 0, 1, 1, 2, 0, 2, 2, 2, 4, 3, 3, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -2, -1, 0, -1, -2, 0, 0, 1, 0, 1, 1, 2, 3, 3, 2, 2, 4, 2, 2, 2, 2, -1, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -2, 0, 0, 0, -2, 0, 0, 1, 0, 0, 0, 3, 2, 2, 1, 2, 2, 2, 1, 2, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, 0, 1, 1, -1, -1, 1, 0, 0, 0, 0, 2, 2, 1, 1, 3, 1, 2, 1, 3, 1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 2, 3, 2, 2, 2, 1, 2, 1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 2, 1, 0, 3, 1, 1, 2, 1, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, -1, 0, 2, 1, 0, 0, 0, 2, 3, 2, 3, 1, 3, 1, 0, 2, 2, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, -1, 0, 2, 0, 0, 1, 0, 2, 3, 0, 1, 1, 2, 0, 0, 1, 2, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 1, 1, 1, 1, 0, 0, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 1, 1, 0, -1, 2, 2, -1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 0, 0, 1, 1, 1, 1, 0, -2, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, 1, 0, 0, 0, 2, 1, 1, 2, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, -3, -1, 0, 1, 2, 0, 1, 4, 1, 1, 2, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -2, 0, 2, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -1, -1, 1, 1, 0, -1, 0, -1, -1, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, -1, 0, -2, -1, -2, -3, -2, -2, -2, -2, 0, 0, 0, -1, -2, -1, -2, 0, -1, -2, -2, -2, -2, 0, -2, 0, -2, -1, -1, 0, 0, -1, -1, -2, -2, -3, -3, -4, -4, -4, -5, -4, 0, 2, 0, 0, -1, -3, -2, -2, -4, -5, -5, -6, -4, -4, -4, -2, -2, -2, 0, 0, 1, 1, 0, 0, 0, -2, -3, -4, -5, -4, -3, -3, 0, 2, 0, -1, -2, -3, -2, -3, -2, -3, -5, -5, -3, -3, -3, -3, -2, -1, 0, 1, 2, 2, 1, 3, 2, 0, 0, -2, -3, -3, -4, -2, 0, 2, 0, 0, -2, -2, -2, -2, -1, -1, -3, -3, -2, -2, -3, -2, 0, 0, 0, 2, 1, 1, 2, 3, 3, 3, 1, 0, -2, -2, -2, -3, 0, 2, 0, -1, -1, -1, -2, -2, -1, -1, -3, -2, -2, -1, -3, -2, 0, 0, 2, 1, 2, 1, 2, 3, 3, 2, 2, 0, 0, -2, -2, -2, 0, 2, 0, -1, -2, -2, -2, -1, -2, -3, -3, -2, -1, -2, -2, -2, -2, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 1, 0, -1, -3, -3, 0, 2, 1, 0, -2, 0, -2, 0, -1, -1, -3, -2, -1, -1, -2, -2, -2, -1, -1, -1, -3, -1, 0, 0, 0, -1, 0, 0, -1, -2, -4, -2, 0, 1, 0, 0, 0, -1, -1, -2, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -2, -2, -1, 0, 0, -1, 0, -1, 0, -1, -3, -3, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, -2, -1, -2, -1, 0, 0, -1, 0, 0, 1, -1, -2, -2, -1, -1, -1, -1, 0, -1, -2, -3, -1, 0, 0, -1, 0, -2, -2, -1, -2, -3, -2, -1, -2, -2, -2, -2, 0, 0, -2, 1, 1, 0, 0, 0, -3, -3, -2, -1, -2, -2, -3, -2, -2, 0, 0, 0, 0, -1, -2, -3, -3, -2, -1, 0, -2, -2, -2, 0, -1, -1, -1, -1, -1, -1, -1, 0, -1, -2, -1, -2, -4, -3, -3, -4, -3, 0, 1, -1, -1, -2, -2, -3, -2, -2, -1, 0, 0, -2, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -2, -1, -2, -3, -3, -4, -5, -4, -4, 0, 1, -2, -1, -2, -3, -4, -2, -2, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -2, -4, -4, -4, -2, -2, -2, -2, -2, -4, -4, -2, 0, 0, -1, -2, -2, -3, -2, -1, -1, -1, 0, 0, 0, 0, 0, -2, -1, -2, -2, -2, -3, -4, -6, -6, -5, -4, -3, -2, -3, -3, -5, -4, 0, 1, 0, -1, -2, -3, -2, -1, 0, 0, 0, 0, 0, 1, -1, -2, -1, -2, -2, -1, -4, -4, -5, -5, -5, -2, -2, -2, -2, -4, -3, -4, -1, 1, 0, -1, -2, -1, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, -2, -2, -3, -3, -2, -2, -3, -4, -5, -2, -2, -2, -2, -2, -3, -3, 0, 2, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -3, -3, -3, -4, -3, -2, -2, -3, -3, -4, -2, 0, 1, 0, -1, -1, -3, -2, -3, 0, 0, 0, 0, -1, 0, 1, 1, 1, 1, 0, 0, -1, 0, -1, -3, -3, -1, -1, -2, -3, -4, -4, -3, 0, 1, 0, 0, -2, -2, -3, -2, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, -3, -3, -2, -1, -2, -2, -3, -5, -4, 0, 0, 0, -2, -3, -2, -4, -3, -1, -1, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -2, -1, -1, -2, -4, -4, -3, 0, 0, 0, -2, -2, -3, -4, -3, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, -2, -3, -4, -3, -2, 0, 1, 0, -2, -1, -2, -3, -4, -2, -2, -2, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, -2, -3, -3, -3, 0, 0, -1, -2, -2, -2, -2, -4, -2, -3, -2, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, -1, -2, -4, -3, -2, -1, 0, -1, -3, -3, -2, -2, -4, -2, -2, -3, -3, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -3, -3, 0, 1, -2, -2, -2, -1, -3, -3, -3, -2, -2, -2, -2, -1, 0, 1, 0, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, -1, -3, -4, -3, 0, 1, -1, -1, -2, -3, -3, -4, -2, -2, -1, -3, -2, 0, 0, 1, 1, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, -1, -1, -5, -5, -3, 0, 0, -2, -1, -2, -1, -2, -2, -3, -3, -2, -3, -2, -1, 0, -1, -1, 0, 0, 0, 2, 1, 1, 0, -1, 0, 0, -1, -3, -4, -5, -2, 0, 0, -3, -3, -2, -1, -2, -3, -3, -2, -3, -2, -4, -2, -2, -2, -2, -2, -1, -1, 0, 1, 0, 0, -1, -1, -1, -1, -1, -2, -4, -3, 0, 1, -1, -3, -2, -1, -2, -2, -2, -2, -3, -4, -4, -4, -4, -4, -3, -2, -2, -2, 0, 0, 0, 0, -1, 0, -2, -1, -2, -3, -3, -3, 0, 3, 1, 0, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, -1, -1, -1, -2, -1, -1, 0, 0, -1, 0, -1, -2, -2, -3, -2, -2, -3, -3, -1, 2, 4, 2, 0, 0, 0, 0, 1, 0, -1, 0, -2, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -2, -3, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 2, 0, 0, 0, 0, -1, -1, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, -1, -1, 0, 0, 1, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 1, 0, -1, -1, 0, -1, 1, 0, 1, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -2, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 0, 0, 1, 0, 0, -1, -2, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 2, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, -2, -2, 0, -1, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 2, 1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, -1, -1, 0, 0, -1, 0, -2, -1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -2, 0, -1, -1, -1, 0, 0, -1, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -2, -1, -1, 0, -2, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, 0, -1, -1, -2, 0, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, -1, 0, 0, -2, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -2, -1, -1, 0, -1, -1, -1, 0, -1, -1, 0, -2, -1, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -2, -2, -2, -1, 0, 0, -1, -2, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 1, -1, 0, -1, -1, -1, -2, -1, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, 1, 0, 0, 0, -1, -1, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, 0, -1, 0, -2, -2, -1, -2, -2, -1, -2, -1, -2, -1, -1, -3, -2, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -1, -2, 0, -1, -1, -1, -2, -2, -2, -1, -1, -1, -2, -2, -3, -5, -3, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, -1, -2, -1, 0, -2, -2, -1, -1, -2, -2, -1, 0, 0, -2, -2, -5, -2, -1, 0, 0, 0, 0, 2, 1, 3, 2, 1, 2, 1, 1, 0, -1, 0, -1, 0, -1, -2, 0, 0, -2, -1, -1, 0, 1, 0, -1, -2, -3, -2, -1, 0, 0, 0, 2, 1, 1, 2, 1, 2, 3, 1, 0, 1, 0, -1, -1, 0, -1, -2, -1, -1, -1, 0, -2, 0, 0, 0, 0, -2, -3, -3, -1, 0, 0, 1, 2, 2, 2, 2, 1, 1, 1, 1, 2, 1, 0, 0, 0, -1, 0, -2, -1, -2, -1, -2, -1, -1, 0, 0, 0, 0, -3, -2, -1, 0, 0, 1, 1, 2, 2, 3, 1, 2, 2, 2, 1, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, -2, -3, -2, -2, 0, 1, 2, 1, 1, 1, 1, 0, 0, 1, 1, 1, 1, 2, 1, 0, 0, -1, -2, 0, -1, -1, -2, -2, -1, -1, 0, -1, 0, -2, -3, 0, 0, 0, 1, 1, 2, 2, 0, 0, 1, 1, 2, 3, 2, 1, 0, 0, 0, -1, 0, 0, 0, -1, -2, -2, -1, 0, 0, -1, -2, -2, -2, -2, 0, 0, 2, 1, 2, 1, 0, 0, 1, 1, 2, 2, 2, 1, -1, 1, 0, -1, -1, 0, 0, 0, -1, -2, -2, 0, 0, -1, -1, -3, -2, -1, 0, 0, 1, 2, 0, 2, 1, 0, 1, 1, 2, 2, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -3, -2, -2, -1, 0, 2, 0, 2, 0, 0, 0, 1, 1, 1, 3, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -3, -2, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 2, 2, 1, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -3, -2, -2, -1, 0, 0, 1, 0, 2, 1, 1, 1, 2, 1, 2, 0, 1, 0, -2, -1, -2, -2, 0, 0, 0, 1, 0, 0, 0, 2, 0, -1, -1, -2, -1, 0, 0, 0, 1, 0, 2, 1, 1, 2, 1, 1, 1, 0, 0, 0, -2, -1, 0, -1, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, -1, -2, -1, 0, 0, 1, 1, 1, 1, 1, 3, 2, 1, 1, 0, 0, 0, 0, -3, -3, 0, 0, 0, 1, 0, 2, 0, 2, 1, 1, 1, 0, -2, -1, 0, 0, 0, 1, 1, 2, 1, 2, 1, 2, 2, 2, 2, 0, -1, -1, -2, -1, -1, 0, 0, 1, 0, 1, 2, 1, 2, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 2, 3, 3, 1, 2, 0, 1, 0, -2, -1, -2, -1, 0, 0, 0, 0, 1, 0, 1, 1, 2, 0, 0, 0, -2, -2, -2, -1, 0, 0, 0, 0, 1, 3, 2, 1, 2, 1, 1, 0, -2, -3, -3, -1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 1, 1, 1, -2, -1, -1, -1, 0, 0, 1, 1, 1, 2, 2, 3, 3, 1, 1, 0, -1, -2, -1, -2, -1, 0, 1, 0, 0, 1, 0, 1, 0, 1, 1, 0, -1, -1, -1, 0, 0, 1, 0, 1, 1, 3, 2, 2, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -2, -1, 0, 0, 1, 0, 1, 1, 2, 1, 2, 2, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -2, -2, 0, -1, 1, 1, 1, 2, 2, 2, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -3, -1, -1, 0, 1, 0, 0, 1, 2, 2, 2, 1, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -2, 0, 0, 1, 0, 0, 0, 2, 2, 2, 2, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -3, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, -1, -2, -2, -2, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -3, -1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 2, 1, 1, 1, 1, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, -2, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, -1, -2, -1, 0, -1, 0, 0, 0, -2, -3, -2, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 1, 0, -1, 0, -1, -1, 0, -1, -1, 0, -1, -1, -2, -2, -1, -3, -3, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, -2, -2, -2, -2, -2, -3, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 4, 2, 3, 3, 5, 4, 2, 2, 2, 3, 2, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 2, 3, 1, 2, 4, 4, 3, 2, 4, 4, 3, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 3, 0, 1, 1, 0, 0, 1, 0, 0, -1, 0, 1, 2, 0, 1, 3, 2, 3, 2, 3, 4, 4, 0, 0, 1, 1, 0, 1, 1, -1, -1, 1, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 3, 3, 3, 2, 2, 3, 3, 0, -1, 1, 0, 0, 1, 1, 0, -1, 1, 2, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, -2, -2, 1, 2, 1, 2, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, -1, 0, 1, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 1, 2, 2, 1, 0, -1, 0, 0, 2, 1, 2, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 2, 1, 0, -2, -1, 0, 0, -1, 0, 2, 1, 1, 2, 2, -1, 0, 2, 3, 2, 0, 0, 3, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -2, -1, -2, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 2, 2, 0, 1, 2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -2, -3, 0, 0, 0, 0, 0, 1, 2, 2, 0, 2, 0, 3, 3, 1, 1, 0, 2, 0, 0, 0, 1, 0, 0, 2, 1, 0, 0, 0, -2, -2, -3, -4, -2, 0, 0, 0, 0, 1, 1, 0, 1, 2, 2, 3, 3, 3, 1, 1, 3, -1, 0, 0, 2, 0, 1, 1, 1, 0, 1, 0, -1, -2, -3, -3, 0, 0, 1, 0, 3, 2, 2, 1, 1, 1, 1, 2, 4, 2, 2, 1, 3, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, 1, 1, 3, 4, 2, 3, 3, 1, 0, 1, 4, 1, 2, 3, 3, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, -2, -2, -1, -2, 0, 0, 0, 2, 2, 3, 3, 3, 4, 2, 1, 2, 2, 2, 2, 3, 2, 0, 0, 0, 0, -1, 0, 2, 0, -1, 0, -1, -2, -1, -1, 0, 2, 0, 0, 3, 3, 3, 2, 4, 6, 4, 1, 3, 2, 1, 2, 3, 3, -1, -1, -1, 1, 0, 0, 1, 0, -2, -1, -1, -1, -2, -1, 0, 1, 0, 1, 2, 2, 3, 2, 4, 4, 4, 1, 2, 1, 2, 1, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -2, -1, -1, -1, 0, 2, 1, 0, 1, 1, 2, 2, 2, 5, 4, 1, 2, 3, 3, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, -1, 0, 0, 0, 1, 2, 1, 0, 1, 2, 1, 4, 4, 2, 3, 2, 3, 3, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, 0, 0, 0, 0, 2, 1, 1, 1, 1, 1, 4, 3, 1, 2, 2, 4, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -1, 1, 2, 2, 1, 0, 2, 1, 1, 0, 3, 3, 1, 2, 1, 3, 2, 0, 1, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 2, 1, 1, 0, 1, 1, 1, 0, 3, 3, 1, 1, 1, 2, 1, 1, 2, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 1, 3, 2, 1, 0, 2, 3, 1, 0, 2, 0, 0, 1, 3, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 2, 3, 2, 1, 2, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 1, 1, 0, 1, 2, 3, 1, 0, 0, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 1, 0, 0, 0, 1, 2, 1, 0, 2, 1, 1, 2, 2, 3, 0, 0, -1, 0, 1, 1, 1, 2, 0, -1, 0, 0, 0, 1, 0, 0, 1, 2, 0, 0, 0, 0, 1, 1, 1, 0, 2, 3, 2, 3, 3, 3, 1, -1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 2, 0, 0, 3, 4, 0, 0, 0, -1, 1, 0, 1, 1, 2, 3, 3, 2, 3, 4, 2, 0, 0, 0, 0, 2, 2, 1, 0, 0, 0, 0, 2, 2, 1, 0, 2, 4, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 2, 1, 5, 4, 2, 0, -1, 0, 1, 2, 2, 2, 0, 0, 2, 1, 2, 2, 1, 1, 3, 3, 2, 0, 0, 0, 2, 1, 2, 1, 3, 2, 1, 2, 4, 5, 3, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 2, 3, 1, 0, 0, 1, 1, 1, 2, 1, 3, 2, 2, 2, 4, 5, 2, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 1, 2, 0, 0, 0, 0, 2, 2, 2, 2, 1, 2, 0, 1, 1, 2, 3, 0, -1, 1, 0, 1, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 2, 1, 2, 1, 2, 0, 1, 2, 3, 2, -1, -1, -1, 0, -2, -2, -1, -2, -2, -1, -2, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, -2, -2, -1, -1, -3, -4, -3, 0, 1, 0, 0, 1, 1, 4, 5, 5, 5, 4, 5, 4, 3, 5, 5, 3, 0, 0, 1, 3, 2, 0, 0, 0, -2, -1, -1, -2, -2, -1, -1, 0, 1, 0, 0, -1, 1, 2, 3, 4, 4, 6, 6, 4, 6, 6, 6, 3, 1, 0, 0, 3, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 3, 3, 4, 3, 3, 5, 5, 2, 1, 0, 0, 1, 3, 2, 0, 0, 0, 1, 0, 2, 1, 0, 1, 1, 1, 0, 0, -1, -2, -2, -2, -3, -1, 2, 3, 3, 4, 3, 2, 1, 0, -1, 1, 2, 3, 3, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, -3, -4, -4, -1, 0, 2, 3, 3, 2, 2, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -2, -4, -4, -1, 0, 1, 0, 1, 2, 0, 0, -1, -1, 0, 1, 3, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -2, -2, -2, -2, -1, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, 2, 2, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, -2, 0, 0, 2, 2, 2, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, -2, -1, 0, 0, 1, 0, 0, 2, 2, 2, 0, 0, 0, -1, -1, -1, 0, 2, 2, 2, 1, 0, 1, 1, 1, 1, 0, 1, 0, 0, -1, 0, -1, 0, -1, 0, 1, 1, 1, 2, 2, 1, 1, 0, 0, -1, -2, -1, -1, 1, 2, 2, 1, 0, 1, 1, 2, 1, 1, 0, 1, 1, -1, 0, -1, 0, 0, 0, 1, 2, 3, 2, 3, 1, 1, 0, 1, 0, -1, -1, -1, 0, 2, 2, 1, 1, 2, 3, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 3, 3, 1, 1, 1, 1, -1, -2, 0, 0, 1, 2, 3, 0, 1, 0, 1, 1, 1, 0, 1, -1, 0, 0, 0, 1, 0, 0, 1, 2, 3, 2, 3, 2, 3, 2, 1, 0, -1, -1, 0, 0, 2, 1, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 2, 3, 4, 3, 3, 3, 1, 2, 1, 0, -2, -1, -1, 1, 2, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 2, 2, 2, 4, 3, 3, 2, 2, 0, 0, 0, -1, -2, 0, -1, 1, 1, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 1, 3, 3, 3, 4, 2, 2, 0, 0, 0, 0, -2, -1, -1, -1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, -1, -2, 0, 1, 3, 4, 3, 3, 2, 3, 1, 0, 0, 0, 0, -3, -2, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 1, 4, 3, 3, 2, 2, 2, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, -1, -1, 0, 0, 2, 2, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -2, -2, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 4, 3, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 2, 3, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 1, 0, -1, -1, -1, -2, 0, 0, 0, -1, 0, 0, 1, 2, 1, 1, 2, 2, 1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 2, -1, -2, -1, -2, 0, 1, 0, 0, -1, 0, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 1, 1, 0, 0, 0, 0, 2, 1, 3, 0, 0, -1, -1, -2, -3, -3, -3, -1, -1, -1, -1, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 1, 2, 1, 0, 0, 0, 3, 2, 1, 0, 0, 0, -2, -4, -4, -4, -3, -2, 0, -1, 0, 0, 2, 1, 2, 0, -1, -2, -1, 0, 2, 2, 1, 1, 1, 0, 0, 1, 1, 2, 0, 0, 1, 0, -1, -3, -4, -4, -2, -1, 0, 0, 1, 1, 2, 3, 3, 1, 1, -1, 0, 1, 2, 2, 1, 1, 0, -1, 0, 0, 1, 1, 2, 2, 2, 1, 0, -1, 0, 0, 0, 0, 1, 1, 2, 4, 4, 4, 4, 4, 1, 0, 0, 0, 3, 2, 1, -1, 0, -1, -1, 0, 0, 1, 0, 1, 1, 2, 2, 2, 2, 2, 1, 3, 3, 1, 4, 4, 3, 5, 4, 5, 3, 0, -1, 0, 0, 0, -1, -1, -3, -2, -1, -2, 0, 0, -1, 0, 0, 1, 1, 2, 3, 3, 3, 1, 2, 2, 3, 2, 2, 2, 4, 3, 2, 0, 0, 0, 0, 0, -2, -1, -3, -3, -2, -2, -3, -1, -1, 0, 0, 1, 1, 2, 1, 2, 0, 0, 1, 0, 1, 1, 2, 2, 1, 1, 1, 0, 0, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 1, 0, -2, -2, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, -1, -1, -2, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, -1, 0, 1, 1, 1, 1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 1, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -2, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -2, 0, -1, -2, -1, -1, 0, 0, -1, -2, -1, 0, -1, -1, -1, -1, -3, -3, -3, -2, -3, -5, -3, -2, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -2, -1, 0, 0, 0, -1, -3, -2, -1, -1, -2, -3, -4, -3, -4, -3, -4, -6, -6, -7, -3, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, -1, -2, -3, -1, -1, 0, -2, -2, -3, -4, -2, -4, -5, -5, -7, -9, -4, -2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -4, -7, -8, -3, -2, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, 1, 0, 1, 0, 1, 0, 0, -1, -3, -4, -6, -4, -2, 1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 2, 3, 2, 0, 0, 0, -3, -5, -4, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 1, 2, 2, 2, 0, 0, 0, -3, -5, -2, 0, 1, 1, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, -3, -3, -2, 0, 1, 1, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, 0, 2, 1, 0, 0, 0, 0, -2, -4, -1, -1, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, -2, -1, 0, 0, 1, 0, 0, 0, 2, 0, 0, 2, 3, 1, 0, 0, 0, 0, -2, -3, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 2, 2, 1, 3, 2, 1, 1, 0, 0, 0, 0, -2, -4, -2, 0, 0, 0, -1, 0, -2, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 1, 1, 2, 2, 2, 0, 0, -1, -1, -3, -4, -2, 0, 0, 1, 0, 0, -2, -2, -2, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 2, 1, 1, 2, 0, 1, 0, -1, -1, -3, -5, -2, 0, 0, 0, -1, -1, -2, -2, -2, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, -1, -4, -5, -2, 0, 0, 0, -1, -2, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -5, -2, 0, 0, 0, -1, -2, -1, -3, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -2, -3, -2, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -2, -3, -3, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 2, 1, 1, 1, 2, 1, 1, 1, 1, 1, 2, 0, 0, 0, 1, 0, 2, 0, 0, 0, -4, -3, -1, 0, 1, 0, -1, 0, -2, -1, 0, 0, 1, 2, 1, 1, 1, 0, 1, 2, 2, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, -1, -4, -3, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 2, 1, 1, 0, 1, 0, 1, 0, -1, -4, -3, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 1, 1, 1, 1, 0, 0, -1, -3, -3, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 3, 3, 1, 1, 2, 1, 0, 0, -1, -4, -2, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, -1, -2, 0, 0, 0, 1, 0, 0, 1, 2, 3, 2, 2, 1, 1, 2, 1, 0, -2, -4, -3, -1, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 2, 1, 2, 3, 3, 1, 1, 2, 1, 1, 0, -3, -6, -3, 0, 0, 0, 0, -1, -1, 0, -1, -2, 0, 0, -1, -1, 0, 0, 2, 1, 1, 1, 1, 2, 3, 3, 2, 2, 2, 1, 0, -2, -3, -6, -4, -1, 0, -1, 0, 0, 0, 0, -2, -1, 0, -1, -1, 0, 0, 1, 1, 1, 1, 1, 3, 3, 3, 2, 2, 0, 1, 1, -1, -2, -4, -6, -4, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 3, 2, 2, 1, 1, 0, 1, 0, -1, -3, -5, -6, -3, -1, 0, -1, 0, 0, -1, -1, -2, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 1, 2, 1, 2, 1, 0, -1, -1, -2, -3, -4, -5, -6, -5, -2, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -2, -2, -4, -4, -5, -5, -7, -7, -4, -1, 0, 0, -2, -1, -1, -2, -1, -1, 0, 0, -1, -1, -1, -2, -1, -2, -1, 0, -1, -2, -2, -3, -2, -4, -5, -6, -6, -7, -7, -7, -4, -1, 1, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, -2, -2, -1, -1, -2, -1, -2, -3, -2, -3, -3, -3, -4, -6, -6, -6, -6, -7, -8, -5, -3, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, -2, -1, -2, -2, -3, -3, -4, -4, -4, -5, -5, -4, -3, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, -2, -2, -2, -1, -2, -2, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, -1, -1, -1, -2, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 0, -1, 0, 0, -1, 0, 0, 0, -1, -2, -1, -1, -1, -3, -3, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -2, -2, -3, -2, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, 0, -3, -2, -2, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 1, 0, 0, 2, 1, 1, 0, 1, 1, 0, 2, 2, 2, 1, 0, 0, 0, -1, -3, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, -1, 0, 0, 1, 0, 0, 0, 1, 1, 2, 3, 3, 2, 2, 2, 0, 0, -2, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 3, 3, 2, 2, 1, 2, 2, 2, 1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 3, 4, 2, 0, 1, 1, 3, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, -1, -1, -1, -1, -2, -2, 0, 0, 1, 1, 2, 3, 0, 0, 1, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, -1, -2, -2, -2, -1, -2, -4, -1, 0, 2, 0, 0, 2, 2, 2, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, -1, -1, -1, -2, -3, -2, 0, 0, 1, 2, 2, 0, 2, 2, 0, 0, 1, 0, 0, 1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -3, -1, -2, -1, -1, 0, -1, 0, 0, 2, 2, 2, 2, 1, 0, 0, 0, 0, -1, 1, 1, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, -3, -2, -3, -2, 0, 0, -1, 0, 0, 0, 2, 2, 2, 2, 0, -1, 0, -2, 0, 1, 1, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, -3, -2, -1, -1, -2, -3, -1, -1, 0, 0, 1, 2, 1, 0, 0, -1, -1, 0, 1, -1, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, -1, -2, -2, -3, -2, 0, -1, -1, -2, -2, 0, 0, 3, 3, 2, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -3, -2, -1, 0, 0, 0, -1, -1, 0, 2, 2, 2, 0, 0, -1, -1, 1, 1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, -2, -1, 0, 0, 0, 0, -2, 0, 1, 2, 0, 2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, -2, -1, 0, 1, 1, 0, 0, -1, 0, 2, 1, 2, 0, 0, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -2, -1, 0, 1, 0, 0, 0, 0, 0, 2, 1, 2, 0, 0, -2, -1, 0, 0, -1, -2, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, -1, -1, -1, 0, 0, 0, -1, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 2, 3, 2, 2, 0, -2, -1, 0, 0, -2, -2, -1, -2, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, -1, -1, 1, 0, -1, 0, 0, 0, 0, 0, 1, 2, 0, -1, -2, -2, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, -1, -1, 0, 1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, -1, -1, 0, 1, -1, -2, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 1, 1, 0, 0, 2, 1, 1, 0, 1, 0, 0, 0, -3, -1, 0, 1, -1, -1, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, 0, 1, -3, -1, -2, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, -2, -2, 0, 0, -2, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -2, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, -1, -2, -2, 0, 0, -2, -2, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, 0, -1, -2, -2, -1, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, -1, -2, -1, -3, -1, 0, 0, -1, -2, -1, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, -2, 0, 0, -1, 0, -1, -2, -3, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 1, 0, 1, 1, 0, 0, 1, 2, 1, 1, 0, 0, 0, 1, 0, -1, -1, 0, 1, 1, 0, 0, 1, 0, 0, -1, -1, 0, 2, 0, 0, 6, 2, 2, 2, 0, 0, 1, 3, 4, 1, 0, 0, 0, 1, 1, 1, -1, -2, 0, 1, 1, 1, 2, 2, 2, 0, -2, -1, 0, 4, 0, 1, 5, 3, 1, 0, 0, -2, 0, 1, 1, 1, 0, 1, 0, 1, 2, 1, -1, 0, 0, 2, 2, 0, 1, 3, 2, 0, -1, 0, 0, 4, 0, 1, 4, 1, 1, 0, 0, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 1, 1, -2, 0, 3, 2, 0, 0, 0, 1, 3, 0, 0, 3, 2, 1, 0, -2, -2, -2, 0, 0, -2, 0, 1, 1, 0, 0, 3, 3, 2, 2, 3, 2, -2, 0, 2, 2, 1, 1, 0, 0, 0, 0, 0, 3, 0, 0, 0, -1, -4, -3, -1, 0, -3, -1, 0, 1, 0, 0, 3, 3, 2, 5, 4, 0, -1, 0, 4, 2, 1, 2, 0, 1, 0, 0, 0, 2, 0, -1, 0, 0, -3, -2, -1, 0, -2, -3, 0, 2, 1, 0, 2, 4, 3, 5, 4, 1, 0, 2, 5, 3, 1, 1, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, -1, -1, 0, -1, -2, -3, 0, 2, 3, 0, 0, 3, 2, 5, 5, 1, 2, 4, 5, 3, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -2, -1, 0, 3, 3, 0, 0, 0, 1, 5, 3, 2, 3, 5, 6, 4, 1, 1, 2, 1, -1, 0, 0, 1, -2, -1, 0, -2, -1, -1, -1, -1, -3, 0, 0, 2, 4, 0, 0, 1, 2, 4, 2, 1, 5, 5, 5, 6, 1, 0, 1, 0, 0, 0, 0, 0, -2, 0, 0, -2, -2, -1, 0, -2, 0, 0, 0, 1, 4, 1, 0, 3, 4, 4, 1, 2, 4, 3, 6, 6, 2, 1, 1, 1, -2, 0, 0, 0, -2, 0, 0, -2, -3, -2, -1, -4, -2, 0, 0, 1, 2, 2, 2, 4, 4, 2, 3, 2, 3, 1, 5, 7, 4, 2, 1, 1, -2, 0, 0, 0, -3, 0, 1, -2, -3, -1, 0, -2, 0, 0, 1, 2, 2, 1, 3, 5, 3, 2, 4, 5, 2, 1, 3, 5, 4, 2, 1, 1, -2, 0, 0, -1, -3, 0, 1, 0, -1, 0, 0, -2, 0, 1, 3, 3, -1, 0, 3, 4, 2, 3, 6, 6, 2, 1, 4, 4, 2, 2, 1, 1, -1, 0, 0, -1, -3, -1, 0, 0, -1, -2, -1, -1, 2, 1, 2, 5, 0, 1, 4, 3, 1, 3, 6, 6, 2, 2, 5, 5, 4, 3, 1, 0, -1, 0, 0, 0, -2, -1, 0, 0, -1, -1, -3, -2, 0, 0, 2, 5, 2, 3, 2, 2, 2, 3, 4, 7, 3, 4, 6, 5, 3, 2, 1, 0, -1, 0, 0, 0, -2, 0, 0, 0, -1, -1, -2, -2, 1, 0, 1, 5, 4, 5, 2, 1, 1, 3, 4, 6, 4, 4, 7, 5, 5, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -2, -2, -2, 0, -1, 0, 1, 3, 4, 6, 3, 0, 3, 2, 3, 5, 4, 5, 5, 5, 5, 2, -1, 0, -1, 0, -1, 0, -1, -1, -1, -1, -3, -1, 0, 0, -1, 0, 0, 2, 4, 6, 2, 1, 4, 1, 2, 4, 4, 3, 4, 4, 4, 0, 0, 0, 0, 0, -1, 0, -2, -3, -1, -2, -2, 0, 0, 0, -3, 0, 1, 1, 0, 3, 2, 3, 2, 2, 2, 3, 5, 2, 3, 4, 3, 0, 0, 0, 0, 0, 0, 0, -1, -4, -3, -3, -2, 0, 0, 1, -2, -2, 0, 1, 1, 0, 3, 4, 3, 3, 3, 4, 4, 3, 2, 3, 2, -1, 0, 0, 0, 0, 0, 0, -2, -2, -3, -2, -2, -1, 0, 1, -2, -3, -1, 0, 0, 1, 3, 4, 4, 4, 2, 3, 4, 3, 4, 5, 1, -2, -1, 1, 0, 0, -1, 0, -2, -1, -1, -2, -2, -2, 0, 0, 0, 0, -1, 0, 0, 1, 2, 5, 2, 3, 3, 4, 3, 3, 4, 3, 1, -2, 0, 1, 0, 0, 0, 0, -1, -1, -1, -2, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 4, 2, 2, 4, 4, 1, 4, 3, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -3, -2, -1, 1, 3, 1, 0, 1, 0, 3, 3, 4, 2, 3, 3, 3, 2, 3, 3, 2, -1, 0, 0, -2, 0, 0, 1, -1, -1, 0, 1, -1, -1, -2, -2, 0, 3, 0, 0, 2, 3, 1, 3, 2, 2, 4, 3, 3, 2, 4, 3, 1, 0, 0, 0, -1, 0, 0, 2, 0, 0, 2, 2, -1, -2, -1, -3, 0, 0, -1, -2, 1, 2, 0, 0, 1, 0, 2, 2, 2, 2, 1, 1, 0, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, -1, -1, 0, 0, 0, 1, -1, -3, 2, 3, -2, -1, 0, 0, 1, 1, 1, 1, 0, 0, -1, -1, 0, 1, 0, 0, 0, 3, 0, 2, 1, 2, 0, 0, 0, 0, 0, 0, -3, -3, 0, 1, -3, 0, 0, 0, 0, 0, 1, 0, 0, 0, -4, -4, -1, 2, 2, 0, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, -1, -4, -3, 0, 0, -2, -1, -1, -1, 0, -1, 1, 0, 0, -2, -4, -4, -2, 2, 2, 0, 0, 2, 1, 1, 1, 1, 0, 0, 2, 0, 0, 0, -3, -4, -1, -1, -3, -1, 0, 0, 0, 1, 1, 0, 0, -2, -5, -3, -2, 1, 2, -1, 0, 2, 1, 2, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, -2, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -2, 0, 0, 1, 1, 0, 0, 1, 2, 3, 2, 4, 3, 3, 1, 1, 2, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 2, 1, 3, 3, 2, 2, 2, 2, 2, 0, 0, 2, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -2, -1, -2, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, -1, -2, -3, -2, -2, -1, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 1, 0, 2, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, -1, -2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -2, -3, 0, 0, 0, 0, 2, 1, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -2, -2, -1, 0, 0, 0, 2, 1, 0, 0, 1, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, 0, -1, -2, -2, 0, 0, 0, 1, 1, 0, 1, 0, 2, 1, 2, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 2, 0, 1, 0, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, -1, -2, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 1, 2, 1, 1, 0, 0, -1, -1, 0, -2, -1, -2, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 1, 0, 0, 0, -1, -2, -2, -2, -1, -2, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, 0, -1, -2, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 0, 0, 1, 1, 0, 0, 1, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, -1, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, -2, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, 0, -1, 0, 0, 1, 1, 0, 1, 1, 0, -1, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 2, 1, 2, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 2, 2, 3, 3, 3, 4, 4, 3, 4, 3, 3, 4, 2, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 4, 4, 5, 4, 4, 4, 4, 5, 4, 2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 1, 0, 0, -1, 0, 0, 3, 2, 3, 4, 4, 4, 3, 4, 4, 2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 3, 3, 3, 2, 1, -2, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 1, 1, 2, -2, 0, 1, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, -1, -1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -2, -1, 0, 0, 0, 0, 1, 1, 0, 2, 1, 0, 1, 1, 0, 0, 0, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 2, 1, 0, 0, 1, 1, 0, 1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, -2, -1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 1, 2, 0, 1, 1, 1, 0, -1, -2, -2, -2, 0, 0, 2, 0, 2, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, -2, -1, 0, 0, 1, 1, 1, 1, 0, 0, -1, -2, -1, -1, -1, -1, 0, 0, 1, 1, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 1, 1, 1, 2, 2, 1, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 1, 0, 0, 0, 0, -1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, -2, 0, -1, 0, -1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -2, 0, 0, 0, -1, -1, 0, 1, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, -1, -1, 0, -1, 0, 1, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 1, -1, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, -1, 0, 1, 1, 1, 0, -1, -1, 0, 0, 1, 1, 0, 0, 1, 0, -2, -2, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 1, 1, 2, 2, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, -1, -3, -2, 0, 0, 0, 0, 1, 1, 1, 0, 2, 2, 2, -1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, -2, -2, -1, 0, 0, 1, 1, 2, 2, 0, 1, 3, 1, 0, -1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 0, 0, 0, 0, 0, 1, 2, 2, 1, 2, 3, 3, 4, 3, -1, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 3, 2, 3, 2, 2, 1, 2, 0, 0, 0, 3, 2, 3, 1, 3, 5, 2, -2, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, -1, 0, 1, 2, 1, 1, 2, 1, 2, 1, 2, 0, 2, 1, 2, 2, 3, 3, 3, -1, -1, 0, -1, 0, -1, -2, -1, -1, 0, -1, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, -1, 0, 0, 0, 0, -1, -2, 0, 0, 0, -2, -1, -2, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 1, 1, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, -1, 0, -1, -1, -2, -3, -2, -1, -3, -1, -2, -2, 0, 0, 2, 1, 1, 1, 3, 3, 2, 3, 1, 0, 0, 0, -3, -1, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, -3, -2, -1, -2, -1, -1, -2, -1, 1, 0, 1, 2, 2, 3, 2, 2, 2, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, -2, -1, -1, 0, 0, -1, -1, 0, 0, 0, 1, 3, 3, 3, 2, 0, 0, -2, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -3, -1, -2, 0, 0, 2, 2, 3, 2, 2, 1, -2, 0, -2, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -3, -3, -2, 0, 1, 1, 1, 2, 0, 0, -1, -1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -2, -1, 0, 0, 0, 1, 1, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 2, 0, 1, 1, 0, -2, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, -3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -3, -1, -1, 1, 0, 0, 0, 0, 0, 2, 2, 2, 3, 2, 0, 0, 0, 0, -1, -2, -3, -1, -1, 0, 0, 1, 0, 1, 1, 0, 0, -1, -3, 0, -1, 0, 0, 1, 2, 0, 0, 1, 3, 2, 2, 1, 1, 1, 1, 0, -1, -2, -1, -2, -1, 0, 0, 1, 1, 2, 2, 1, 1, 0, -2, -1, -1, 0, 1, 0, 0, 0, 1, 1, 1, 2, 1, 1, 1, 0, 0, 1, -1, -1, -1, -1, 0, 0, 1, 1, 2, 1, 1, 2, 0, 0, -2, -1, -1, 0, 0, 0, 2, 2, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, -3, -1, 0, 0, 0, 0, 2, 0, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, 2, 1, 1, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 0, 2, 1, 1, 1, 0, -2, -1, -2, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 0, -2, -2, -1, 1, 0, 0, 1, 0, 1, 1, 1, 2, 1, 0, 0, 0, -3, 0, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, -1, -2, 0, 0, 1, 0, 0, 0, 1, 1, 2, 1, 1, 2, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 4, 4, 3, 1, -2, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 1, 3, 3, 3, 3, 2, -2, 0, -1, 0, 0, 0, 1, 0, 0, 0, 2, 1, 0, 1, 0, 0, -1, -1, -2, -2, 0, 0, 0, -1, 0, 0, 0, 2, 3, 2, 3, 2, -2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, -1, -2, 0, -1, -1, 0, 0, 0, 0, 1, 1, 3, 3, 1, -3, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 1, 1, 1, 2, 2, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 2, 2, 1, 0, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 3, 1, 0, -3, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -2, -2, -1, -1, 0, 0, 0, 1, 0, 0, 2, 3, 3, 2, 1, -3, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -3, -3, -2, -1, 0, 0, 0, 0, 1, 1, 3, 3, 4, 3, 0, -3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -3, -1, -1, -1, 0, 0, 2, 1, 3, 3, 4, 4, 2, 1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 2, 3, 4, 4, 4, 3, 4, 2, -1, 0, 0, 1, 0, -1, -1, -1, -2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 3, 4, 5, 4, 3, 2, 0, -1, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 3, 2, 1, 3, 1, 3, -2, 0, -1, 0, 0, -1, -2, -1, -2, 0, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -2, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 2, 0, 0, 1, 0, 1, 1, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 2, 2, 0, 0, 0, 0, -1, -1, 0, -2, -2, -1, -1, 0, 0, 2, 0, 0, 0, 2, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 2, -1, 0, 0, 0, -1, 0, 0, 0, -1, -2, -1, 0, 0, 0, 1, -1, 0, 1, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, -1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 3, 2, 1, 2, 0, 0, 0, -2, 0, 1, 3, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 1, 2, 1, 1, 0, 0, -1, 0, 2, 3, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 0, 0, 1, -2, 0, 1, 2, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 2, 0, 1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, -2, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 2, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 2, 1, 0, 0, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 1, 1, 2, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 1, 0, -1, 0, -1, -2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, -1, -1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 1, 0, -1, 0, -1, -2, -1, 1, 0, 0, -1, -1, -1, -2, -1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -3, 0, 2, 1, -2, -1, 0, -1, 0, -1, 0, 0, 2, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, -2, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 2, 1, 2, 1, 2, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, -2, -1, -1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 2, 1, 2, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, -1, -1, 0, -1, 0, -1, 0, -1, 1, 0, 1, 0, 0, 1, 2, 2, 2, 2, 1, 0, 0, -1, 0, 0, -1, 0, -1, 0, -2, -1, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, -1, 0, 0, 1, 1, 3, 2, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, -2, -1, 0, 1, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 1, -1, -2, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 2, -1, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 1, 1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, -1, -1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 1, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -2, 0, -1, -1, -2, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 2, -1, 0, 0, 0, 0, -1, 0, -1, -1, -2, -1, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 2, 1, -2, -1, 0, 0, 0, -1, 0, 0, 0, -2, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, -1, -2, -1, 2, 3, -1, 0, 0, 1, 0, 0, 0, 1, 1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -2, 0, 1, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, -1, -2, -2, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 0, -1, -1, -1, -1, -1, 0, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, -2, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, -1, -1, -1, -1, -1, -1, -1, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -1, -2, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, -2, -2, 0, 0, -1, -1, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -2, 0, 0, 0, 0, -2, -1, 0, -1, -1, -1, 0, -1, -2, -1, -2, -1, -3, -4, -2, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, -3, -1, -1, 0, 0, 0, -1, -3, -2, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -4, -5, -2, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -4, -4, -2, 2, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 3, 2, 1, 0, 0, -3, -4, -2, 1, 2, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 4, 3, 3, 2, 0, -2, -4, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 2, 3, 4, 4, 4, 2, 0, -2, -4, -2, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 4, 4, 2, 3, 3, 1, 0, -3, -2, 0, 1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, 1, 2, 3, 4, 3, 1, 0, 1, -2, -4, -1, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 2, 1, 2, 1, 1, 0, 1, 0, 2, 4, 5, 4, 2, 2, 2, 1, 0, -3, -1, 0, 0, 0, 0, 0, -2, -2, -2, -2, -2, 0, 0, 1, 2, 1, 2, 1, 1, 2, 1, 2, 2, 4, 5, 4, 3, 2, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 2, 1, 2, 2, 1, 2, 2, 2, 4, 4, 5, 4, 2, 2, 2, 0, -1, -4, -1, 0, 0, -1, 0, 0, 0, -2, -2, -1, -1, 0, 0, 1, 2, 2, 2, 2, 1, 0, 1, 1, 4, 5, 5, 4, 4, 1, 0, -1, -3, -5, -1, 0, 0, 0, -1, -1, -2, -2, -1, -2, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, 0, 2, 3, 3, 4, 4, 3, 3, 2, -1, -2, -5, -2, 0, 0, -1, 0, 0, -1, -1, -3, -2, -1, 0, 1, 1, 0, 0, 0, 2, 0, 0, 0, 2, 3, 2, 3, 3, 4, 3, 1, -1, -3, -5, -2, 0, 0, 0, -1, 0, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 2, 2, 3, 3, 3, 2, 0, -2, -4, -2, -1, 0, 0, -1, 0, -1, -2, -1, -1, 0, 0, 1, 1, 0, 0, 1, 1, 2, 0, 0, 1, 2, 2, 3, 4, 2, 2, 1, 0, -1, -4, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 2, 1, 1, 2, 2, 2, 2, 3, 3, 1, 2, 0, -1, -3, -2, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 2, 3, 2, 2, 1, 1, 2, 3, 2, 2, 0, 0, -2, -3, -2, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 3, 3, 2, 2, 1, 2, 1, 2, 2, 1, 2, 0, -1, -3, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, 0, 0, 1, 0, 0, -1, 0, 2, 2, 1, 2, 2, 3, 3, 2, 4, 4, 3, 1, 0, -1, -3, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 2, 0, 1, 0, 2, 2, 4, 5, 5, 3, 1, 0, -1, -2, -1, 0, -1, -1, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, -1, 1, 0, 1, 0, 2, 3, 3, 4, 4, 4, 2, 1, 0, -2, -3, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, -2, -2, 0, 0, 0, 1, 0, 0, 1, 1, 3, 3, 4, 3, 2, 2, 0, -1, -4, -1, 0, -1, -1, -1, 0, -1, -2, -2, 0, -1, 0, -1, -1, -2, 0, 0, 0, 0, 1, 2, 1, 1, 2, 3, 4, 4, 3, 1, 0, -2, -5, -2, 0, 0, -1, 0, 0, -1, -1, -3, -3, -2, -2, -1, -2, -1, -2, -1, 0, 0, 1, 1, 0, 2, 3, 4, 4, 4, 3, 2, 0, -3, -5, -2, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -3, -1, -2, -1, -1, 0, 1, 1, 1, 1, 2, 3, 4, 3, 3, 1, 0, -2, -4, -3, 0, 0, 0, 0, 0, 0, -2, -1, -1, -2, -1, -3, -3, -3, -1, -2, -1, 0, 0, 1, 2, 1, 3, 3, 2, 3, 1, 0, -1, -3, -5, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -3, -3, -4, -2, -1, -2, -2, -1, -1, 0, 0, 1, 0, 1, 1, 0, 0, -1, -1, -3, -5, -3, 0, 0, -1, -1, 0, 0, 0, 0, -2, -1, -2, -3, -4, -4, -3, -3, -4, -2, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -2, -5, -6, -3, 1, 1, -1, 0, 0, 0, -1, 0, -1, -1, -2, -2, -4, -4, -3, -3, -4, -2, -3, -2, -2, 0, -1, 0, -2, -1, -3, -2, -3, -5, -5, -2, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, -1, -2, -1, -3, -2, -1, -2, -2, -2, -1, -2, -1, -1, -2, -1, -3, -4, -2, -3, -4, -5, -3, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -2, -1, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, -2, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 1, 1, 2, 1, 2, 2, 0, 0, 0, 2, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, -2, -1, 0, -2, -2, -2, -1, 0, 0, 0, -1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, -2, -1, -1, 0, 0, 0, -1, -1, 0, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -2, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -2, -2, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -2, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -2, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -2, -2, -1, 0, -1, -1, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, 0, -2, -1, -3, -1, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -2, -1, 0, -1, -1, -1, -1, -2, -2, -1, -1, 0, 0, -2, -3, -3, -3, -2, -3, -2, -1, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -3, -4, -7, -8, -7, -6, -7, -9, -8, -8, -6, -4, 0, -1, -1, -3, -4, -4, -4, -3, -1, -2, -1, -1, 0, 0, 0, 0, -2, -1, -1, -3, -4, -7, -9, -9, -9, -9, -10, -12, -12, -14, -12, -5, -2, -1, -1, -3, -3, -4, -4, -2, -1, -1, -1, 0, 1, 1, 1, 0, -1, 0, -2, -3, -4, -8, -8, -8, -9, -8, -10, -12, -13, -14, -13, -7, -3, 0, -2, -3, -5, -4, -2, -3, -2, -2, 0, 0, 1, 1, 1, 1, 1, 0, -1, 0, -4, -5, -5, -4, -6, -5, -6, -7, -10, -13, -13, -7, -2, -1, -2, -1, -4, -3, -2, -2, -2, -1, 0, 0, 1, 2, 2, 1, 1, 3, 1, 0, -1, -2, -1, 0, -1, 0, -2, -4, -6, -10, -10, -6, -1, 0, 0, -2, -4, -3, -1, -1, 0, 0, -1, 0, 1, 2, 2, 1, 1, 2, 2, 1, 0, -1, 0, 1, 2, 1, 0, -2, -2, -6, -7, -4, -2, 0, -2, -4, -3, -3, -2, -1, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 1, 2, 3, 4, 3, 2, 1, -1, -3, -5, -2, 0, 0, -1, -3, -3, -3, -3, -1, 0, -1, -2, -2, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 5, 4, 4, 2, 2, 2, 0, -1, -3, -2, -1, 0, -1, -3, -3, -4, -3, -1, 0, -1, -1, -3, -1, 0, 0, -1, -3, -2, 0, 0, 0, 1, 5, 5, 4, 3, 2, 2, 0, 0, -1, 0, 0, 0, 0, -1, -3, -4, -4, -2, 0, 0, -2, -2, -3, -1, -1, -2, -3, -3, -2, 0, 0, 0, 4, 4, 2, 1, 1, 2, 0, -1, -1, -1, 0, 0, 0, -2, -4, -4, -4, -3, -2, -1, -2, -4, -3, -3, -3, -3, -5, -4, -1, 0, 1, 0, 3, 4, 4, 1, 2, 0, 0, 0, -2, 0, 0, 0, -1, -4, -4, -4, -3, -3, -2, 0, -3, -5, -4, -4, -3, -3, -4, -4, -2, 0, 0, 0, 2, 2, 3, 3, 1, 0, 0, -3, -3, 0, 0, 0, -1, -4, -4, -5, -4, -3, -2, -1, -3, -4, -4, -4, -2, -2, -4, -5, -4, -1, -1, 0, 1, 2, 2, 2, 1, 0, 0, -5, -4, 0, 0, -2, -3, -4, -4, -3, -5, -3, -2, 0, -2, -4, -3, -4, -3, -4, -4, -4, -4, -3, -2, -1, 0, 1, 3, 2, 1, 2, 0, -4, -5, -1, 0, -1, -2, -3, -3, -3, -3, -3, -2, -1, -2, -3, -1, -1, -2, -4, -6, -5, -3, -3, -4, -2, -2, 0, 2, 3, 2, 2, 0, -2, -5, -2, 0, -1, -2, -3, -3, -4, -4, -3, -2, -1, -1, -1, 0, 0, -1, -3, -6, -6, -4, -3, -2, -4, -2, -1, 1, 3, 3, 2, 0, -1, -3, -2, 0, -1, -2, -4, -4, -4, -3, -3, -2, -1, 0, -1, 0, 1, 1, -2, -5, -4, -3, -1, -1, -4, -3, -1, 0, 4, 4, 3, 2, -1, -4, -2, 0, 0, -1, -2, -3, -5, -4, -3, 0, 0, 0, 0, 0, 0, 0, -1, -5, -5, -3, 0, 0, -2, -3, -1, 0, 4, 4, 3, 3, -1, -4, -3, -1, 0, -2, -4, -3, -4, -5, -2, 0, 0, 0, -1, -2, 0, -1, -3, -4, -3, 0, 0, 0, -1, -3, 0, 1, 4, 4, 2, 2, -3, -5, -1, -1, 0, -2, -3, -4, -5, -4, -2, 0, 0, 0, -1, -2, 0, -1, -3, -4, -3, 0, 1, 2, 0, 0, 0, 1, 3, 4, 3, 0, -3, -5, -3, -1, 0, -4, -4, -4, -4, -4, -3, -2, 0, 0, 0, -1, 0, -1, -3, -5, -3, 0, 2, 1, 2, 1, 2, 1, 2, 4, 2, 0, -3, -5, -3, -1, 0, -4, -3, -4, -4, -5, -5, -1, -1, -1, -1, -2, 0, 0, -1, -2, -3, -1, 1, 2, 4, 2, 2, 3, 2, 3, 2, 0, -4, -5, -3, -1, 0, -4, -3, -4, -5, -5, -4, -3, -1, -1, -1, -3, 0, 0, 0, 0, -1, -1, 0, 4, 4, 4, 3, 2, 4, 3, 1, -1, -5, -6, -3, 0, 0, -4, -4, -4, -3, -5, -5, -3, -1, -3, -2, -2, 1, 1, 0, 0, 0, 0, 1, 3, 4, 4, 3, 2, 3, 1, 1, -2, -7, -7, -4, -1, 0, -1, -4, -3, -3, -4, -4, -4, -1, -3, -2, -2, 1, 2, 0, 0, 0, 2, 3, 4, 3, 4, 4, 0, 1, 0, -2, -5, -8, -8, -6, -1, -1, -1, -2, -4, -3, -4, -4, -3, -2, -1, -2, -2, 1, 1, 2, 0, 0, 3, 2, 2, 3, 2, 2, 0, -1, -1, -5, -7, -11, -9, -5, -1, -1, -3, -3, -4, -3, -2, -3, -3, 0, -1, -2, -2, 1, 2, 1, 0, 2, 2, 3, 2, 1, 1, 1, -1, -3, -3, -7, -9, -11, -12, -6, -2, -1, -4, -4, -4, -4, -3, -2, -2, -1, 0, -2, -1, 1, 2, 1, 1, 0, 0, 1, 2, 1, 0, -1, -3, -6, -5, -8, -11, -12, -14, -7, -2, -2, -4, -4, -3, -4, -4, -4, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, -1, -2, -3, -6, -7, -8, -8, -10, -13, -14, -14, -8, -3, -1, -4, -3, -5, -4, -3, -4, -2, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -4, -5, -8, -10, -10, -11, -13, -14, -14, -16, -14, -9, -3, -2, -4, -4, -4, -3, -2, -1, -2, 1, 1, 0, 0, 0, -1, 0, 0, -1, -3, -5, -6, -9, -9, -12, -13, -13, -15, -16, -15, -16, -15, -11, -3, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, -1, -3, -4, -5, -6, -6, -7, -9, -9, -9, -10, -9, -11, -9, -5, -2, -2, 0, 0, 0, 0, 0, -1, -2, -2, -3, -3, -3, -5, -4, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -1, 0, 2, 2, 2, 0, 0, 0, -2, -2, -4, -4, -5, -5, -3, 0, 0, 0, 0, 0, 1, 2, 2, 1, 3, 2, 0, 0, 1, 0, -1, -1, -2, 0, 5, 5, 3, 2, 1, 0, 0, -1, -1, -1, -3, -4, -1, 0, 0, 1, 0, 0, 0, 2, 2, 2, 3, 4, 2, 2, 1, 2, 0, -1, 0, 1, 3, 4, 4, 3, 1, 1, 0, 1, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 3, 2, 2, 0, -2, -1, 0, 3, 5, 5, 3, 3, 2, 1, 1, 1, 0, 0, 0, 0, 2, 1, 0, -1, -2, -2, -2, -2, -1, 0, 0, 3, 3, 2, 1, 0, -1, -3, 1, 4, 6, 5, 5, 3, 2, 0, 1, 0, 1, 0, 2, 1, 2, 0, 0, -1, -2, -3, -4, -4, -3, -2, 1, 2, 2, 2, 1, 0, -4, -4, 1, 3, 6, 6, 5, 3, 1, 1, 0, 0, 0, 0, 1, 2, 3, 1, 0, 0, -1, -3, -3, -6, -4, -1, 0, 1, 0, 0, 0, -2, -4, -3, 0, 2, 5, 6, 4, 3, 2, 0, 0, 1, 1, 1, 1, 3, 4, 2, 2, 1, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, -1, -2, -4, -4, 0, 3, 4, 4, 4, 1, 1, 0, 0, 0, 1, 1, 2, 3, 2, 2, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, -3, -5, -4, 0, 2, 2, 3, 1, 1, 0, 0, 0, 1, 1, 2, 3, 2, 3, 1, 1, 0, 1, 3, 3, 3, 3, 1, 1, 1, 0, -1, -1, -3, -5, -5, 0, 1, 1, 2, 1, 0, -1, 0, 0, 0, 3, 3, 3, 2, 1, 1, 0, 0, 0, 0, 2, 3, 4, 4, 2, 1, 0, -2, -1, -3, -4, -4, 0, 1, 2, 2, 0, 0, -1, -1, 0, 2, 3, 3, 4, 2, 0, 0, 0, 0, 0, 0, 2, 2, 5, 5, 2, 1, 0, -2, -2, -2, -4, -5, 0, 1, 1, 2, 1, 0, -1, 0, 0, 0, 2, 4, 2, 0, 0, 0, -1, 0, 1, 1, 2, 4, 5, 5, 3, 2, 1, 0, -2, -3, -4, -5, -1, 0, 0, 2, 1, 0, -1, 0, 1, 1, 2, 2, 2, 0, 0, -1, -1, 0, 0, 0, 3, 3, 5, 4, 3, 2, 0, 0, -1, -3, -4, -4, 0, 1, 1, 1, 1, 2, 1, 0, 1, 2, 2, 1, 0, 0, -2, -2, 0, 0, 1, 2, 3, 4, 6, 5, 3, 3, 0, 0, -2, -3, -4, -4, 0, 1, 2, 3, 3, 1, 0, 0, 0, 0, 1, 1, 0, -1, -3, -3, 0, 0, 1, 3, 4, 5, 7, 5, 3, 2, 0, -2, -2, -3, -4, -4, 0, 2, 3, 3, 3, 2, 1, 0, 0, 1, 2, 1, 0, 0, -2, -3, 0, 0, 3, 4, 5, 5, 6, 6, 3, 0, 0, -2, -3, -3, -5, -4, 0, 2, 2, 3, 3, 2, 0, 0, 0, 1, 1, 0, 1, 0, -2, -2, -1, 0, 3, 5, 4, 7, 5, 4, 3, 0, 0, -2, -2, -3, -5, -4, 0, 1, 2, 2, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -1, 0, 3, 4, 4, 4, 4, 3, 2, 1, 0, -1, -1, -2, -5, -4, 0, 0, 2, 2, 2, 2, 1, 1, 2, 0, 0, 0, 0, 0, -1, -2, 0, 2, 3, 4, 4, 4, 2, 2, 0, 0, 0, 0, -1, -2, -3, -4, 0, 0, 1, 2, 1, 1, 1, 2, 3, 1, 0, 0, 2, 0, 0, -1, 0, 1, 2, 3, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, -2, -4, 0, 0, 0, 1, 1, 1, 2, 2, 2, 3, 0, 1, 1, 1, 0, 0, 1, 2, 2, 1, 0, 0, 1, 0, 0, -1, 0, 0, -1, -2, -4, -4, 0, 0, 0, 1, 0, 1, 1, 1, 3, 2, 1, 0, 2, 0, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, -2, -3, -2, -2, -1, -4, -3, -1, 0, 0, 0, 1, 0, 0, 1, 1, 2, 3, 0, 0, 2, 1, 2, 2, 2, 3, 1, 0, -1, 0, 0, 0, -1, -2, -3, -1, -1, -5, -5, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 2, 1, 1, 2, 0, 1, 2, 2, 2, 1, 0, -1, -1, -2, -2, -2, -2, -2, -2, -2, -5, -5, 0, 0, 1, 2, 2, 2, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, -1, -2, -1, -2, -2, -2, -4, -3, 0, 0, 1, 3, 1, 3, 2, 1, 0, 2, 2, 1, 0, -2, -2, -1, -3, -3, -2, 0, 0, -1, 0, -2, -1, -1, 0, 0, -1, -2, -4, -3, 0, 2, 3, 3, 3, 2, 1, 0, 0, 1, 1, 0, -1, -3, -3, -2, -3, -3, -3, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -3, -3, 0, 3, 2, 3, 1, 1, 2, 0, 0, 0, -1, -1, -2, -3, -2, -2, -2, -3, 0, 0, -1, 0, 1, 0, 2, 1, 0, 1, 1, 0, -2, -3, 1, 4, 3, 4, 2, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, -1, 0, 0, 1, 2, 1, 2, 3, 2, 2, 1, 1, 0, 1, -1, -2, -3, 0, 2, 4, 2, 0, 0, 0, -1, -1, -3, -1, -1, -3, -2, -1, -1, 0, 2, 2, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, -1, -3, -3, 0, 0, 1, 0, 0, -2, -1, -1, -1, -1, -2, -2, -2, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 0, 0, 0, 0, -2, -2, -3, -4, -3, -2, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 3, 2, 2, 0, 0, -1, 0, 0, -1, -2, -3, -2, -1, 0, 0, 1, 0, 0, 0, 0, 1, 2, 2, 1, 1, 0, 0, 1, 1, 1, -1, 1, 4, 4, 3, 2, 1, 1, 0, 0, 0, 0, -1, -1, 0, 2, 2, 1, 0, -1, 0, 1, 1, 2, 2, 2, 1, 0, 1, 0, 1, 0, 0, 1, 3, 3, 3, 3, 2, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, -1, -2, -2, -2, 0, -1, 0, 1, 1, 1, 2, 1, 0, 0, -1, 1, 3, 4, 3, 3, 1, 0, 1, 0, 0, 0, 0, 2, 1, 2, 2, 1, 0, -3, -2, -2, -3, -1, -1, 1, 0, 0, 0, 0, 0, -1, -2, 1, 4, 5, 4, 3, 1, 2, 1, 0, 0, 0, 0, 2, 2, 1, 0, 0, -1, -2, -2, -3, -5, -3, -2, 0, 1, 0, 1, -1, 0, -3, -2, 1, 3, 4, 3, 4, 2, 1, 0, 1, 0, 0, 1, 2, 2, 2, 0, 0, -1, -1, -1, -4, -3, -4, 0, 0, 0, 0, -1, -1, -1, -3, -1, 0, 3, 4, 4, 3, 2, 0, 1, 0, 0, 1, 1, 1, 2, 2, 2, 1, 0, 0, 0, -2, -2, 0, 0, 0, 0, -1, 0, -1, -2, -2, -2, 0, 1, 1, 2, 2, 1, 0, -1, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -2, -1, -1, -3, -1, 0, 2, 2, 2, 2, 0, 0, -1, 0, 0, 1, 1, 1, 0, 1, 0, -1, 0, 0, 0, 1, 1, 2, 1, 0, 0, -2, -1, -2, -1, -2, -1, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 2, 3, 1, 1, 0, 0, -2, -1, 0, 0, 0, 0, 2, 2, 1, 0, -2, -2, -1, -2, -3, -1, 0, 0, 2, 2, 0, 0, 0, 0, 0, 1, 1, 3, 2, 1, -1, 0, -1, -1, -1, 0, 0, 0, 2, 2, 0, 0, 0, -2, -2, -1, -2, -2, -1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, -2, -2, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, -1, -2, -3, -2, -1, 0, 1, 2, 1, 1, 0, 0, 1, 1, 1, 1, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, 2, 3, 1, 1, 0, 0, 0, -2, -3, -3, -1, 0, 1, 2, 2, 2, 1, 0, 1, 1, 0, 2, 0, 0, -1, -3, -2, 0, -1, 0, 0, 1, 3, 4, 1, 1, 0, 0, -1, -2, -3, -4, -2, 0, 1, 3, 2, 3, 0, 0, 1, 1, 1, 1, 1, 0, 0, -3, -3, 0, 0, 0, 0, 2, 3, 2, 4, 1, 0, -1, -3, -3, -2, -3, -2, 0, 2, 2, 3, 2, 2, 0, 1, 0, 0, 0, 0, 0, -1, -2, -2, -1, 0, 2, 2, 3, 2, 3, 2, 1, 0, -2, -2, -4, -4, -4, -3, 0, 2, 2, 2, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, -2, -1, 1, 1, 3, 3, 4, 3, 2, 0, 0, -2, -1, -3, -3, -3, -2, 0, 1, 1, 2, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, -2, 0, 1, 2, 1, 3, 2, 2, 0, 0, -1, -1, -1, -1, -1, -3, -1, -1, 0, 2, 1, 1, 2, 1, 1, 2, 1, 0, 0, 1, 0, -1, -1, 0, 1, 2, 1, 2, 1, 0, 0, -1, -1, -2, -1, -1, -1, -3, -2, -1, 0, 1, 1, 1, 1, 2, 2, 2, 0, 0, 2, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, -1, -2, -1, -2, -2, -2, -1, -1, 0, 0, 1, 0, 0, 2, 1, 2, 2, 1, 1, 2, 0, 0, 0, 2, 1, 1, 1, 0, 0, 0, -1, -2, -1, -1, -1, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -2, -2, -2, -4, -3, -2, -2, -3, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, 2, 1, 0, 0, 1, 2, 2, 2, 0, 0, 0, 0, -1, -1, -2, -4, -2, 0, -1, -3, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 2, 2, 1, 1, 0, 0, 1, 0, 1, 1, 0, 0, -1, -2, -2, -2, -2, -3, -2, -1, -2, -4, -2, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, -1, -1, -1, -1, -1, -2, -2, -2, -1, -1, -1, -2, -2, -2, -1, 0, 0, 1, 1, 1, 2, 0, 1, 1, 1, 1, 0, -1, -2, -1, -1, -2, -3, -3, -2, -2, 0, -1, -1, -1, -2, -1, -1, 0, -2, -3, -1, 0, 1, 2, 3, 2, 1, 0, 0, 1, 1, 0, -1, -1, -1, -1, -3, -2, -3, -1, -2, -1, -1, 0, -1, 0, -1, 0, 0, 0, -2, -2, 0, 0, 2, 3, 3, 1, 1, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 4, 3, 3, 2, 0, 0, 0, -1, -2, -1, -1, -1, -1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 1, 2, 2, 0, 0, 0, -1, -2, -1, -2, -2, -2, 0, 0, 0, 2, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, -1, -1, 0, 0, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 2, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 2, 1, 1, 1, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, -1, 0, -1, -1, 1, 1, 2, 1, 1, 0, 0, 1, 1, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -2, -1, 0, -2, -2, -1, 0, 0, 1, 1, 1, 0, 1, 0, 1, 1, 0, 2, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -2, -2, -1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -2, -2, -1, -2, 0, -1, 0, 0, 2, 2, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -2, 0, 0, 0, 0, 1, 1, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -3, -1, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 2, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -2, -1, 0, 1, 0, 0, -1, 0, 0, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 2, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, -1, 0, 1, 2, 1, 1, 0, 0, -2, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, -1, -1, 0, 0, 2, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 2, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -2, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 1, 0, 1, 0, -1, 0, -1, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, -2, -2, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 2, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, -1, 0, 0, -1, -2, -2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, -1, -1, 0, -2, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, -1, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, -1, -1, 1, 1, 1, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 2, 1, 2, 1, 1, 0, 0, 0, 0, -1, 0, -1, -2, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 1, 2, 1, 2, 1, 0, 0, 0, 0, 0, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 1, 0, 0, -1, 0, 0, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -2, 0, -2, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, -1, 0, 0, 0, -1, -1, -1, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 3, 0, 0, 1, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 4, 2, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 2, 1, 0, 1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 3, 1, 1, 1, 0, 0, 0, 0, 0, 0, 4, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 3, 1, 1, 1, 0, 0, 0, -2, -2, 0, 4, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 2, 1, 0, 2, 0, 0, 0, -1, -1, 0, 2, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 1, 0, 0, 0, -2, 0, 2, 1, 0, 0, 0, 0, -1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 2, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, -1, 0, 1, 0, 0, 0, 1, 2, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 2, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, -1, 1, 2, 3, 1, 2, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, -1, 0, -1, -1, -1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 2, 3, 2, 2, 1, 0, 1, 0, 0, -2, -1, -2, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 1, 3, 2, 2, 2, 0, 0, -1, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 2, 3, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 2, 2, 0, 1, 0, -1, 0, -1, -1, 0, 0, 2, 0, 0, 0, -1, -1, 0, -1, 0, 1, 2, 1, 0, 0, 1, 1, 0, 1, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 1, 0, -1, 0, -1, -2, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 2, 2, 3, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 0, -1, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 3, 2, 3, 1, 2, 0, 0, 0, 0, -1, 0, -1, -1, -2, 0, 3, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 3, 2, 3, 2, 2, 2, 1, 1, 0, 0, 0, -1, 0, -1, -2, 0, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 3, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 2, 2, 1, 2, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 2, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 2, 2, 1, 0, 2, 1, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 2, 2, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 3, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 2, 3, 2, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 0, 0, 0, -1, -1, -2, -1, 0, 0, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -2, -1, -1, 0, 0, 1, 0, -1, -1, 1, 0, 0, 0, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, -1, -2, -1, -1, 0, -1, -2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 1, 1, 1, 1, 1, 1, 2, 2, 4, 0, -1, 3, 1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 2, 2, 2, 3, 2, 1, 1, 0, 1, 3, 0, 0, 2, 2, 1, 1, 0, 0, 0, 0, 1, 2, 1, 2, 1, 0, 1, 2, 1, 0, 0, 1, 2, 0, 1, 3, 2, 2, 1, 1, 1, 3, 0, 0, 1, 0, 0, 2, 1, -1, -1, 0, 2, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 2, 1, 0, 0, 2, 2, 1, 2, 0, 1, 3, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 2, 1, 0, 2, 1, 0, -1, -1, 0, 2, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 3, 2, 2, 2, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 1, 1, 1, 1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 1, 1, 1, 1, 1, 2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 2, 3, 2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 1, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, -2, 0, -2, -2, 0, 0, 0, 2, 2, 1, 2, 0, 0, 1, 1, 1, 1, 2, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 2, 3, 2, 2, 2, 1, 0, -1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 2, 3, 2, 2, 3, 3, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, -1, -2, -1, -1, 0, 0, 0, 0, 1, 2, 1, 2, 3, 2, 0, 1, 2, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, -1, -1, 0, -1, 0, -1, 0, 1, 1, 0, 0, 0, 1, 1, 1, 4, 1, 1, 2, 2, 1, 1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, 0, 1, 1, 2, 1, 0, 1, 2, 1, 2, 2, 1, 1, 2, 2, 0, -2, -2, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 2, 2, 1, 2, 0, 0, 1, 2, 2, 3, 1, 1, 0, 0, 0, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, 0, 2, 1, 1, 2, 1, 1, 1, 1, 2, 2, 0, 0, 0, 0, 1, -2, -1, 0, -1, -1, -2, 0, 0, -2, 0, -1, 1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 1, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -2, -2, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 1, 1, 0, 0, 2, 0, 2, 1, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 1, 1, 0, 0, 2, 1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, -1, -1, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, -1, 0, 0, 0, 1, 0, -1, 0, 3, 0, -1, -1, -2, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 2, -1, 0, 1, 1, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 2, 0, -1, 0, 1, 1, 2, 1, 0, 0, 0, -1, -1, -1, -2, -3, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 4, 0, -1, 1, 0, 1, 2, 1, 0, -1, 0, 0, 0, 0, -2, -1, 0, 1, 0, -1, 0, 0, 1, 0, 0, 1, 1, 1, 0, -1, 0, 2, 4, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 1, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -2, 0, -1, -1, -1, 0, -1, 0, 0, -1, -2, -1, -2, -1, -2, -2, -4, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, -2, -2, -3, -4, -3, -4, -3, -4, -5, -5, -5, -6, -5, -5, -3, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, -1, -3, -3, -3, -3, -4, -4, -4, -4, -6, -4, -5, -2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, -1, -1, -2, -3, -3, -2, -3, -2, -4, -3, -4, -4, -5, -2, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -1, -1, -2, -1, -3, -3, -4, -4, -1, 0, 0, 0, -2, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -2, 0, -1, -3, -3, -3, -2, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -3, -1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, -1, -2, -2, -2, -1, 0, -1, -1, -2, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 0, 0, 0, -2, -2, -2, -2, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 1, 0, 0, 0, -1, 0, -3, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 2, 0, 0, 0, -2, -2, -2, 0, 0, 0, -1, -1, -1, -2, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, -1, -1, -2, -1, 0, 0, 0, -1, -1, -2, -1, -2, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, -1, -1, -2, -2, -1, 0, -1, -1, -1, 0, -1, -2, -1, -1, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, -2, -2, -1, -1, -1, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, -1, 0, -1, 0, -1, -2, -1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, -1, -3, -3, -1, 0, 0, 0, 0, -1, -1, -2, -1, 0, -1, 0, -1, 0, 0, 0, -1, -1, -2, 0, 0, 0, 1, 0, 1, 1, 2, 1, 0, 0, -1, -2, -2, 0, 0, -1, -2, 0, -2, -1, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, -2, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, -1, -1, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, -1, -1, -2, 0, 0, -1, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -2, -1, 0, 0, 0, -1, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, -1, -2, 0, -1, 0, -1, 0, -2, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, -2, -2, -2, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, -2, -1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 2, 0, -1, -2, -3, -2, -2, -1, -1, 0, -2, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 0, 0, 0, -1, -1, -3, -1, 0, -1, -1, -2, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, 1, 2, 1, 0, -2, -2, -4, -1, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 2, 1, 1, 2, 0, 0, 0, -2, -3, -3, -1, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, -2, -3, -3, -5, -2, 0, -1, -1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -3, -3, -5, -3, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -4, -4, -4, -2, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, -1, -1, -2, -2, -3, -3, -5, -4, -5, -5, -5, -3, -1, -1, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -2, -4, -4, -6, -5, -7, -6, -5, -6, -3, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, -3, -2, -3, -4, -5, -5, -6, -7, -6, -7, -6, -6, -3, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -1, -2, -2, -2, -2, -3, -3, -2, -2, 0, 3, 3, 0, 0, 0, 0, -1, -1, -1, -1, -3, -4, -2, -1, 0, 0, -2, -2, -1, 0, -1, -1, 0, -1, -2, -2, -1, -3, -3, -3, -3, 0, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -4, -5, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, -1, -2, -2, -2, -2, 0, 0, 0, -1, -2, -2, -2, -2, -2, -2, -3, -5, -4, 0, 1, 1, 0, 1, 2, 1, 1, 1, 1, 1, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, -1, -3, -4, 0, 1, 1, 0, 0, 2, 2, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, -2, 0, 0, 0, 0, 0, -1, -1, -3, -3, 0, 1, 1, 1, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -2, 0, 0, 0, -1, -1, -2, -1, -3, -3, 0, 2, 2, 0, 1, 0, 1, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -2, -2, -2, -4, -3, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, -2, -1, 0, -3, -2, 0, 1, 0, 1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 1, 2, 1, 1, 0, 1, 0, -1, 0, -1, 0, 0, -2, -3, 0, 1, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 2, 2, 2, 0, 1, -1, -1, 0, 0, -1, -2, -2, 0, 0, 0, 0, 0, 0, -2, -1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, -3, -3, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 1, 2, 2, 2, 1, 0, 0, 0, 0, 0, -1, -1, -4, -4, 0, 0, 1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, -2, -3, 0, 0, 1, 0, 0, 0, -2, 0, 0, 0, 0, 0, -1, -1, -2, 0, 1, 0, 0, 0, 1, 3, 3, 1, 1, 0, 0, 0, 0, 0, -2, -3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 1, 1, 3, 3, 0, 0, 0, 0, 0, 0, -2, -4, 0, 0, 1, 1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 3, 3, 1, 0, -1, 0, -1, 0, -2, -4, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, -1, 0, 0, 1, 3, 3, 3, 2, 2, 0, 1, 0, 0, 0, 0, -1, -3, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 2, 2, 2, 2, 1, 0, 1, 0, 0, 0, 0, 0, -1, -3, 0, 1, 1, 0, 0, 0, 0, 0, 2, 2, 1, 1, 0, -1, -2, -2, -2, 0, 2, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 1, -2, -3, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, -2, -1, 0, 1, 0, 2, 0, 1, 0, 0, 0, 1, 0, 1, 1, -1, -4, -1, 0, 1, 1, 0, 1, 0, 1, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -5, 0, 0, 2, 0, 0, 0, 1, 1, 2, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, -2, -4, -1, 0, 1, 0, 0, 1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 1, 2, 1, 0, 0, 1, 0, 1, 0, 0, -3, -5, 0, 0, 2, 0, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 2, 3, 0, 0, 1, 1, 2, 2, 1, 1, 0, 1, 0, 0, -2, -4, -3, 0, 1, 0, 2, 1, 1, 0, 0, 1, 0, 1, 0, -1, -1, 0, 1, 0, 0, 0, 1, 1, 2, 2, 0, 0, 0, 1, 0, -1, -3, -3, -5, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 2, 2, 0, 0, -1, -1, -3, -5, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 2, 1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, -1, -2, -4, -5, 0, 3, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -5, -5, 0, 3, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -2, -2, -2, -2, -4, -4, -4, -4, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, -2, 0, -1, -1, -1, -3, -2, -2, -3, -4, -4, -3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -2, -1, 0, 0, -1, -2, -1, -2, -3, -2, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, -2, -2, -4, -5, -7, -6, -5, -6, -7, -7, -6, -6, -4, -3, -2, -1, -2, -3, -3, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -3, -5, -5, -8, -8, -8, -7, -8, -8, -9, -10, -10, -7, -3, -1, -2, -3, -3, -1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, -2, -3, -6, -7, -7, -7, -7, -8, -9, -8, -9, -10, -6, -3, 0, -2, -2, -2, -2, -1, 0, 0, 0, 0, 1, 2, 2, 1, 0, 1, 0, 0, 0, -3, -4, -6, -5, -5, -5, -6, -6, -6, -7, -8, -5, -2, 0, -3, -1, -1, -1, -1, 0, 0, 0, 0, 2, 1, 2, 1, 1, 1, 2, 0, -1, -3, -4, -3, -3, -2, -3, -4, -5, -5, -6, -6, -3, -2, 0, -2, -2, -2, 0, -1, 0, 0, 0, 1, 1, 2, 2, 0, 0, 1, 1, 0, 0, -3, -3, -2, -1, 0, -1, -1, -1, -2, -4, -3, -4, 0, 0, -1, -1, -1, -1, 0, 0, 1, 0, 1, 0, 2, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -3, -2, 0, 0, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, -1, -1, -1, 0, 1, 2, 2, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -2, -2, -2, -1, 1, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, -1, -1, -2, -2, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -3, -4, -3, -1, -2, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -2, -2, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -5, -4, -2, -1, -1, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, -1, -2, -1, 0, -1, 0, 0, -2, -3, -1, -2, -3, -4, -4, -2, -3, -2, -1, 0, 0, 0, 1, 2, 0, 0, 0, -1, 0, 2, 0, 0, -2, -2, -1, 0, 0, 0, -1, -1, -3, -2, -3, -2, -3, -4, -5, -4, -2, -3, -2, 0, 1, 1, 1, 2, 0, 0, 0, -1, 0, 1, 0, 0, -2, 0, -2, 0, 0, -1, 0, -2, -3, -2, -2, -3, -4, -5, -5, -5, -2, -3, -2, 0, 0, 1, 2, 1, 1, 1, 0, -1, -1, 0, 0, -2, -1, -2, -1, -1, 0, 0, -1, -1, -1, -3, -2, -2, -4, -4, -5, -5, -4, -3, -2, -2, -1, 0, 2, 2, 2, 2, 0, -1, -1, 1, 0, -2, -2, -1, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, -4, -6, -5, -4, -4, -3, -3, -3, -1, 0, 2, 2, 1, 1, 0, -1, 0, 1, 0, -1, 0, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -5, -5, -5, -4, -4, -2, -3, -3, 0, 0, 3, 2, 3, 2, 2, 0, 0, 0, 0, -2, 0, -1, 0, -1, 0, 0, 1, 0, 0, -1, 0, -2, -4, -6, -5, -3, -2, -1, -2, -2, -1, 0, 1, 3, 1, 3, 1, -1, 0, 1, 0, -1, 0, -1, -1, -1, 0, 0, 1, 0, 0, -2, -2, -3, -4, -7, -5, -4, -2, -1, -1, -2, 0, 1, 2, 2, 2, 1, 0, -1, 0, 1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, -1, -2, -2, -4, -6, -5, -3, 0, 0, 0, 0, 0, 1, 1, 3, 1, 2, 0, 0, 0, 1, 0, 0, -1, -2, -1, -2, -1, 0, 0, 0, 0, -2, -2, -3, -4, -5, -4, -1, -1, 0, 0, 0, 0, 0, 2, 2, 2, 0, 0, -2, 0, 0, 0, -2, -2, -2, -2, -1, 0, 0, 0, 1, 0, 0, -1, -1, -2, -3, -2, -1, -1, 0, 1, 1, 0, 0, 2, 2, 2, 0, -1, -2, -1, 0, 0, -1, -1, -2, -2, -2, -1, 0, 0, 0, 0, -1, 0, 0, -2, -2, -1, -1, 0, 0, 1, 0, 1, 0, 2, 2, 0, 0, -2, -4, -3, 0, -1, -1, -1, -1, -2, -2, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 1, 2, 1, 1, 0, 1, 1, 0, 0, -2, -4, -3, -1, 0, -1, -1, -1, -2, -2, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, -2, -3, -3, -3, 0, 0, -2, -2, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -2, -5, -5, -5, -5, -2, 0, -2, -2, -2, -1, -2, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -2, -1, -2, -4, -4, -5, -7, -5, -2, 0, -2, -2, -2, -1, -1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 1, 0, -1, 0, -2, -2, -3, -4, -5, -5, -5, -8, -7, -5, -1, -1, -2, -2, -3, -1, -2, 0, 0, 1, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, -2, -3, -2, -5, -5, -7, -6, -6, -8, -9, -9, -7, -2, 0, -3, -2, -2, -1, -3, -1, -1, 0, 1, 0, 0, 1, 1, 2, 0, 0, -1, -1, -3, -4, -6, -7, -8, -9, -9, -8, -9, -9, -9, -7, -4, 0, -1, -2, -2, -2, -2, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -2, -3, -5, -7, -7, -9, -9, -9, -9, -9, -10, -9, -7, -3, 0, 0, -1, -1, -1, 0, -1, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, -1, -1, -2, -2, -4, -4, -4, -5, -5, -6, -4, -4, -4, -5, -3,
    -- filter=0 channel=9
    1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 2, 2, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 1, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -2, -2, -2, -2, 0, -1, -1, -1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -1, -3, -1, -2, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, -2, -3, -2, -1, -2, -3, -2, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -3, -2, -2, -2, -2, -2, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, -2, -2, -2, -1, -1, -2, -1, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -2, -2, -2, -1, -1, -2, -2, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, -2, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 2, 2, 0, 1, 0, -1, -1, -1, -2, -2, -2, -1, -2, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, -1, -1, -1, 0, -2, -2, -1, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 2, 1, 2, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 2, 2, 1, 1, 1, 0, 0, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 2, 1, 1, 0, 0, 0, -1, -1, -2, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 2, 1, 1, 1, 0, 1, 0, -1, -1, -1, 0, -2, -1, -1, 0, -1, -1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -2, -2, -2, -1, -2, -1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -2, -2, -2, -1, -2, 0, 0, 1, 0, 0, 1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, -1, 0, -1, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -3, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -2, -3, -3, -1, -2, -2, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -2, -1, -2, -2, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -2, -1, -1, -2, -3, -2, -1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -2, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 3, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 3, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, -1, 0, -1, -1, 0, 0, -1, 1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 2, 2, 1, 0, 1, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 2, 0, 0, 0, -1, -1, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 2, 1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, -2, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, -1, -1, -2, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 2, 2, 0, -1, 0, 0, 0, -1, -1, 0, -2, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -2, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -2, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -2, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 3, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 2, 1, 1, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 1, 2, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 2, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 2, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -2, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, -2, 0, -1, -2, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, -1, -2, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, -1, -1, 0, 0, 0, -1, 0, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, -2, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 1, 1, 1, 0, 2, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 2, 1, 0, 1, 0, 2, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 1, 2, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 3, 1, 1, 1, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, -2, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 4, 3, 3, 1, 1, 1, 0, 0, 0, 0, -1, -2, -2, -2, -3, -3, -4, -2, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 2, 1, 2, 0, 4, 3, 2, 1, 0, 1, 0, 0, 0, 0, 0, -1, -2, -2, -1, -2, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 2, 3, 0, 3, 1, 2, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 1, 0, 1, 1, 0, 0, 1, 1, 2, 1, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 2, 1, 0, 1, 1, 1, 1, 1, 2, 1, 0, -1, 0, 0, 0, -1, -2, -1, -1, -1, -1, 1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -2, -1, 0, 0, -2, -1, -1, -1, 0, 0, 0, 1, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, 0, -1, -1, 0, 0, -1, 1, 0, 0, 0, -2, -2, 0, -1, -2, -2, -1, -1, -1, 1, 0, 0, -1, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, -2, 0, -1, -2, -2, -2, 0, -1, 0, 1, 0, 0, -2, -3, -3, -2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, -2, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 1, 2, 0, -2, 0, 0, 0, 0, 0, 0, -1, 0, 2, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, -2, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -3, -2, 0, 0, 0, 0, 0, 1, 2, 3, 1, 2, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, 2, 3, 1, 2, 1, 0, 0, 0, 0, 0, 2, 2, 2, 1, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, -2, -1, 0, 0, 0, 0, 1, 1, 2, 2, 0, 2, 1, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 1, 0, 2, 2, 1, 1, 0, -1, -2, 0, 0, 0, 1, 0, 0, 0, 2, 0, 2, 1, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 3, 1, 1, 0, -1, -1, 0, -1, 0, 0, 0, 1, 1, 3, 0, 3, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 2, 0, -1, -1, -2, -1, -1, 0, 0, 1, 1, 1, 1, 1, 0, 3, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -2, -2, -2, 0, 0, 0, 0, 0, 1, 1, 2, 0, 1, 0, -1, -1, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 2, -1, -2, -1, -2, -1, 0, 1, 1, 1, 0, 0, -1, 0, 0, 2, 2, 1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, -1, -1, -1, 0, 1, 0, 1, 0, 0, -1, 0, 0, 2, 3, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, 1, 1, 1, 1, 0, 0, 0, -1, 1, 3, 2, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, -1, -1, 0, 0, 1, 2, 1, 1, -1, -1, -1, -2, -2, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -2, -2, -3, -1, -2, -2, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, -1, -4, -3, -3, -1, -2, -3, -1, -2, 0, 0, 2, 0, 3, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -3, -5, -3, -3, -1, -1, -2, 0, -1, 0, 2, 0, 3, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, -3, -3, -3, -2, 0, 0, 0, 0, 0, 1, 1, 0, 2, 2, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, -3, -3, -3, -1, -1, -1, 0, 0, 0, 1, 3, 0, 2, 2, 1, 2, 3, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -3, -3, -3, -2, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 3, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -3, -4, -2, -2, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 1, 1, 1, 0, 2, 2, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 2, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 2, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, -1, -1, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 3, 3, 2, 2, 1, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 8, 7, 4, 3, 1, 0, 1, 0, 0, 0, -1, -2, -4, -4, -5, -5, -4, -3, -3, -3, -4, -5, -4, -3, -2, -1, -1, 0, 0, 1, 4, 8, 8, 6, 4, 2, 1, 1, 2, 1, 0, 0, 0, -2, -3, -3, -4, -4, -3, -4, -5, -6, -7, -6, -6, -6, -4, -3, -3, -2, 0, 2, 5, 7, 8, 5, 2, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, 0, -2, -1, -1, -2, -2, -4, -6, -5, -3, -4, -4, -3, -4, -4, -2, 0, 4, 7, 5, 3, 1, 1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, -1, -3, -4, -4, -3, -3, -3, -4, -3, -5, -2, 0, 3, 4, 3, 2, 1, 2, 1, 1, 1, 3, 2, 2, 2, 1, 1, 1, 1, 0, 2, 0, 0, -1, -3, -3, -3, -2, -4, -4, -4, -4, -2, -1, 3, 5, 3, 2, 1, 1, 2, 0, 1, 3, 2, 2, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, -2, -2, -1, -3, -3, -4, -3, -5, -2, -1, 3, 5, 2, 2, 1, 1, 2, 1, 2, 1, 1, 1, 0, 0, 0, 1, 2, 1, 0, 0, 1, 0, 0, -1, -2, -3, -4, -4, -4, -5, -2, -1, 3, 4, 0, -1, 0, 1, 1, 1, 1, 2, 1, 0, 0, -2, 0, 0, 0, 0, 0, 2, 1, 1, -1, -1, -2, -3, -2, -4, -3, -4, -3, 0, 3, 2, 0, -2, -2, 0, 1, 1, 1, 1, 1, 0, -1, -2, 0, 0, 0, 0, 0, 2, 1, 0, 0, -2, -4, -2, -1, -2, -2, -3, -1, 0, 2, 0, -1, -5, -4, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 2, 2, 0, 0, -2, -2, -3, -3, -1, -1, -2, -1, -1, 0, 1, 0, -2, -3, -4, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -2, -3, -3, -2, -1, -1, -1, -2, 0, 1, 1, 2, 0, -3, -2, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, -4, -4, -2, -3, -2, -1, -1, -1, 0, 2, 2, 3, 2, 0, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, -4, -5, -4, -3, -2, 0, 0, 0, 2, 2, 2, 4, 3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 3, 3, 2, 0, -2, -5, -4, -2, -2, 0, 0, 0, 2, 3, 4, 5, 4, 1, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 1, 4, 3, 4, 2, -1, -3, -4, -3, -1, 0, 0, 0, 1, 3, 4, 5, 4, 2, 0, 0, 2, 1, 1, 0, 1, 1, 1, -1, 0, 1, 0, 2, 3, 3, 3, 1, 0, -2, -4, -3, 0, 0, 0, 0, 0, 1, 3, 6, 3, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, 0, -3, -4, -3, -2, 0, 0, 0, 0, 0, 2, 3, 5, 2, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -2, -4, -4, -2, -1, 0, 0, 0, 1, 2, 3, 2, 0, -2, -2, -2, -1, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 1, 0, 0, 0, -2, -2, -2, -1, -1, 0, 0, 0, 0, 2, 2, 2, 0, -2, -3, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, -1, -2, -1, 0, 0, -1, 0, 0, 1, 1, 2, 2, 0, -1, -2, -1, 0, 1, 1, 2, 2, 1, 0, 0, 0, 1, 3, 3, 3, 2, 0, 0, -1, -1, -1, -2, -1, -2, -2, -2, 0, 1, 2, 2, 0, -1, 0, -1, 0, 1, 1, 3, 2, 0, 0, 0, 0, 0, 1, 4, 3, 1, 0, -1, -2, -3, -1, -1, -3, -2, -1, -1, 0, 1, 2, 3, 2, 0, 1, 0, 0, 1, 1, 2, 0, 0, -1, 0, 0, 1, 3, 1, 2, 1, -1, -1, -4, -4, -4, -2, -3, -3, -4, -2, -1, 0, 3, 4, 2, 1, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 1, 1, 2, 2, 0, 0, 0, -2, -3, -4, -4, -3, -3, -4, -4, -3, -1, 0, 2, 3, 3, 3, 3, 3, 2, 2, 1, 0, 0, 0, 0, 2, 1, 1, 0, 0, 2, 0, 0, -2, -4, -5, -4, -4, -5, -5, -4, -4, -2, 0, 2, 4, 4, 3, 2, 1, 2, 3, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, -1, -4, -5, -4, -3, -3, -4, -3, -3, -2, 0, 3, 4, 6, 4, 1, 3, 1, 1, 2, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, -4, -4, -3, -2, 0, -1, -2, -2, 0, 2, 4, 7, 5, 4, 3, 3, 2, 1, 2, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, -2, -4, -6, -6, -4, -2, -1, 0, 0, -1, 0, 1, 4, 7, 8, 6, 5, 4, 3, 2, 1, 1, 0, -2, -2, -1, -1, -2, -1, -2, -2, -4, -4, -4, -5, -6, -4, -1, -1, -1, 0, 0, 0, 3, 4, 7, 8, 7, 5, 5, 3, 3, 0, 1, 0, -2, -1, -1, -2, -3, -2, -3, -4, -4, -6, -4, -5, -4, -3, -2, -1, 0, 0, 0, 2, 3, 5, 5, 5, 5, 4, 4, 4, 1, 0, 1, 0, 0, -2, -1, -2, -2, -3, -3, -4, -5, -5, -4, -3, -3, -2, -2, -1, 0, 0, 0, 2, 2, 1, 1, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -2, -2, -1, -2, -2, 0, -1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, -2, -1, 0, 0, 0, -1, 0, 1, 1, 1, 2, 1, 0, -2, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -2, -2, -3, -2, -2, -1, -1, 0, 0, 0, -1, 0, 0, 1, 3, 1, 1, 0, -2, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, -1, 0, 1, 1, 0, 0, 0, -1, 0, -1, 1, 2, 2, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 2, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, 1, 3, 3, 2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 2, 1, 0, 0, 1, 1, 1, 0, 0, 1, 0, 1, 0, 0, 1, 2, 3, 1, 2, 1, 0, -1, 0, 0, 0, 1, 0, 1, 0, -1, -1, 0, 1, 2, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 2, 3, 1, 0, 1, 0, -1, 0, 1, 0, 2, 1, 1, 0, 0, -2, 0, 1, 2, 1, -1, 0, 0, 1, 0, 0, 2, 2, 1, 1, 1, 2, 3, 3, 0, 0, 2, 1, 0, 0, 0, 2, 1, 1, 2, 2, 0, -1, 0, 1, 2, 0, -1, -2, 0, 0, 0, 1, 2, 2, 2, 0, 0, 1, 2, 2, 0, 0, 2, 1, 0, 1, 0, 1, 0, 1, 1, 0, 1, -1, 0, 2, 1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 2, 2, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 1, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 3, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 2, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 2, 2, 2, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 1, 0, 0, 1, 2, 2, 1, 2, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 2, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 2, 0, 2, 2, 2, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 3, 1, 0, 0, 0, -1, 0, 0, 1, -1, 0, 2, 0, 0, 0, 0, 0, 0, 0, -3, -1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 2, 2, 2, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 2, 0, 0, 0, 0, 1, 0, -1, -2, 0, 0, 0, 0, 1, 0, 0, 3, 3, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 2, 3, 4, 3, 2, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, -1, 0, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 2, 2, 1, 0, 2, 3, 2, 1, 0, 1, 1, 0, 2, 1, 1, 0, 0, 0, -1, -1, 1, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 1, 1, 3, 4, 1, 0, 1, 2, 2, 1, 2, 0, 1, 0, -1, -1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 0, 0, 0, 1, 2, 2, 0, 0, 1, 1, 2, 1, 1, 1, 2, 0, 0, -1, 0, 1, 2, 0, 0, 0, -1, -1, 0, 0, 0, 2, 1, 1, 0, 0, 0, 1, 2, 2, 1, 0, 1, 1, 1, 0, 0, 1, 1, 0, -1, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, -2, -1, 2, 2, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 2, 0, 0, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 0, 0, -1, 0, 2, 1, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 1, 0, 1, 0, 0, -1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, -2, -2, -2, 0, 0, -1, -1, 0, 0, -2, -1, 0, 2, 3, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, -2, -1, -2, -2, -2, -2, -1, 0, -1, -2, -1, -1, -1, -2, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, 0, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 3, 4, 4, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, -1, -1, -1, -3, -2, -3, -2, -2, -1, -1, -1, -1, 0, -1, 0, 4, 8, 10, 7, 4, 1, 0, 0, 0, 0, 0, -3, -4, -4, -4, -4, -4, -4, -5, -6, -7, -6, -7, -7, -7, -6, -3, -4, -2, -1, -1, 1, 5, 9, 10, 7, 2, 0, 0, 0, -1, 0, -2, -2, -4, -4, -5, -5, -3, -3, -4, -5, -8, -8, -9, -8, -8, -6, -3, -4, -3, -3, 0, 1, 7, 8, 8, 6, 2, 0, 0, 0, 0, -1, -2, -2, -2, -3, -2, -1, 0, 0, -1, -3, -6, -7, -7, -7, -6, -3, -2, -3, -3, -3, -2, 1, 6, 7, 7, 4, 3, 0, 0, 1, 1, 1, 1, 0, -1, 0, 0, 2, 2, 2, 0, 0, -4, -4, -4, -4, -3, -2, -2, -2, -4, -5, -3, 0, 6, 7, 6, 4, 3, 1, 2, 2, 2, 1, 1, 1, 2, 0, 2, 5, 4, 3, 2, 0, -3, -3, -3, -4, -3, -2, -3, -3, -3, -5, -3, -1, 6, 6, 5, 5, 3, 3, 3, 1, 1, 3, 2, 2, 1, 0, 3, 5, 4, 3, 2, 0, 0, -3, -2, -4, -3, -1, -2, -3, -3, -4, -4, -1, 6, 6, 6, 4, 3, 2, 2, 2, 2, 3, 4, 2, 2, -1, 1, 4, 3, 2, 0, 0, 0, -3, -3, -2, -3, -1, -2, -3, -3, -3, -3, 0, 4, 4, 2, 1, 0, 0, 1, 0, 2, 2, 3, 3, 0, 0, 2, 4, 2, 1, 1, 1, 0, 0, -2, -3, -2, -2, -3, -3, -2, -4, -4, -1, 5, 3, 1, -2, -4, -1, 0, 1, 2, 3, 3, 1, 1, 1, 3, 3, 3, 2, 1, 1, 0, -1, -4, -3, -4, -3, -2, -3, -2, -4, -2, -1, 3, 3, 0, -3, -5, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 3, 5, 4, 3, 3, 0, -2, -4, -6, -4, -4, -4, -3, -2, -3, -3, 0, 4, 2, 0, -3, -5, -2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 4, 3, 3, 2, 0, -1, -4, -5, -6, -2, -4, -2, -2, -2, -2, 0, 3, 2, 0, -2, -4, -2, -1, -2, -2, -1, -1, 0, 0, 1, 2, 2, 3, 2, 3, 3, 2, -1, -5, -5, -5, -3, -3, -3, -2, -3, -1, 0, 4, 3, 1, -2, -1, -3, -1, -2, -3, -2, -1, 0, 1, 2, 3, 3, 2, 3, 6, 5, 4, 0, -3, -5, -4, -2, -4, -3, -2, -3, 0, 1, 5, 4, 2, -1, -1, -1, -2, -1, -2, -1, 0, 2, 4, 4, 3, 3, 3, 5, 6, 8, 6, 2, 0, -4, -4, -4, -4, -3, -1, -1, 0, 2, 4, 5, 3, 0, -2, -1, 0, -1, -2, -1, 1, 3, 3, 3, 2, 2, 2, 6, 6, 8, 6, 4, 0, -4, -5, -4, -3, 0, 0, 0, 0, 1, 5, 5, 2, 0, -1, 0, 0, 0, -2, -1, 0, 1, 3, 2, 3, 4, 4, 6, 8, 8, 6, 2, -1, -4, -4, -4, -2, -1, -1, -1, -1, 1, 5, 4, 2, 0, 0, -1, 0, 0, -1, -1, 0, 2, 2, 2, 2, 5, 6, 7, 7, 6, 3, 1, -1, -3, -3, -3, -2, -1, -1, 0, -1, 0, 3, 4, 2, -1, -1, 0, 0, 0, -2, 0, 2, 2, 4, 4, 4, 3, 4, 6, 7, 5, 0, 0, -2, -4, -2, -1, -1, -1, 0, 0, 0, 0, 3, 3, 1, -1, -3, 0, -1, 0, 0, 1, 3, 3, 5, 4, 3, 3, 3, 5, 5, 2, 0, -1, -1, -2, -1, 0, 0, 0, -1, -1, -1, 0, 3, 3, 1, -1, -2, -2, 0, 1, 1, 2, 3, 4, 4, 4, 3, 3, 4, 7, 5, 2, 0, -1, -1, -1, -1, 0, 0, -2, -2, -3, -1, 0, 4, 3, 0, -1, -2, -2, -1, 0, 1, 3, 5, 3, 3, 2, 2, 2, 4, 6, 6, 3, 0, 0, -1, 0, 0, 0, -1, -1, -4, -4, -2, 1, 4, 4, 3, 1, -2, -2, 0, 0, 2, 3, 3, 3, 1, 1, 1, 2, 4, 5, 4, 1, 0, -1, -2, -3, 0, 0, -2, -2, -4, -4, -3, 0, 4, 4, 2, 0, 0, 0, 0, 0, 0, 1, 3, 2, 1, 1, 1, 0, 1, 3, 3, 0, -2, -3, -4, -4, -3, -2, 0, -3, -5, -4, -2, 0, 5, 3, 3, 2, 1, 0, 0, 0, 1, 0, 0, 1, 2, 1, 1, 0, 1, 3, 3, 0, -1, -3, -4, -4, -3, -2, -1, -3, -6, -6, -3, 0, 5, 4, 2, 2, 0, 0, 0, 1, 1, 0, 0, 1, 1, 2, 1, 0, 0, 0, 1, 0, -1, -3, -5, -6, -5, -3, -1, -2, -6, -6, -3, 0, 4, 5, 3, 3, 1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -2, -2, -5, -6, -3, -2, -2, -2, -4, -5, -3, 0, 6, 6, 4, 2, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, -3, -2, -1, 0, -2, -3, -5, -6, -6, -4, -3, -1, -2, -3, -4, -2, 1, 5, 7, 6, 3, 1, 2, 0, 0, 0, 0, 0, -1, -1, -2, -1, -4, -3, -3, -3, -5, -5, -6, -6, -6, -4, -5, -4, -2, -3, -3, -2, 1, 5, 6, 6, 5, 4, 3, 2, 0, 0, 0, -1, -1, -1, -3, -2, -4, -5, -5, -5, -7, -7, -7, -7, -7, -7, -4, -3, -4, -3, -4, -1, 1, 5, 8, 8, 5, 4, 4, 2, 2, 0, -1, -1, -3, -3, -1, -3, -4, -5, -7, -7, -10, -9, -8, -7, -7, -5, -5, -6, -4, -2, -2, 0, 1, 4, 6, 6, 4, 3, 3, 3, 0, 1, 0, 0, 0, -2, -1, -2, -3, -3, -5, -5, -5, -7, -6, -4, -3, -3, -4, -2, -2, -2, 0, 0, 0, 3, 5, 4, 3, 4, 2, 0, 0, 1, -1, 0, 0, -3, -4, -3, -4, -4, -3, -3, -1, -2, -2, 0, 0, 0, 2, 1, 2, 4, 5, 3, 1, 2, 6, 5, 4, 3, 2, 0, 0, 0, -1, -2, -3, -4, -4, -4, -5, -4, -4, -5, -2, -3, -3, -1, 0, 2, 1, 2, 4, 6, 6, 6, 2, 3, 5, 4, 5, 2, 1, 0, 0, -1, 0, -1, -2, -1, -1, -2, -2, -1, -3, -4, -4, -4, -4, -1, 0, 1, 0, 0, 2, 4, 5, 4, 1, 3, 4, 4, 2, 1, 0, -1, -1, -1, 0, -2, 0, 0, 0, 0, 0, 0, -2, -2, -2, -4, -4, -3, -3, 0, -1, 0, 1, 2, 4, 5, 2, 2, 3, 5, 2, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 2, 2, 1, -1, 0, -2, -4, -6, -5, -4, -4, -2, -3, -1, 0, 2, 3, 2, 2, 4, 3, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, -2, -1, -4, -5, -6, -6, -5, -4, -6, -4, -1, 1, 4, 2, 2, 2, 4, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, -2, -4, -7, -7, -6, -7, -7, -6, -4, -2, 0, 2, 1, 2, 1, 3, 1, 1, 0, 0, 1, 2, 2, 0, 0, -1, 0, 0, 0, 1, 0, -1, -3, -5, -5, -7, -7, -8, -8, -8, -7, -3, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 1, 3, 2, 0, 0, 0, 0, 1, 2, 0, -1, -2, -5, -6, -6, -7, -8, -7, -8, -6, -3, 0, 3, 2, 2, 0, 1, 0, -1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 2, 2, 1, 0, -2, -5, -6, -8, -6, -6, -6, -8, -7, -4, 1, 3, 2, 2, 0, 0, -2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, -3, -5, -6, -7, -6, -5, -7, -6, -5, -3, 1, 2, 2, 1, 1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 2, 3, 2, 2, 0, -2, -4, -7, -6, -6, -6, -6, -5, -4, -3, 1, 4, 3, 1, 0, 0, 0, 0, 0, -1, 0, 2, 3, 1, 2, 0, 0, 2, 4, 4, 4, 1, -1, -3, -7, -6, -7, -6, -4, -4, -4, -1, 2, 4, 3, 2, 2, 0, 0, 0, 0, -1, 1, 1, 4, 3, 3, 1, 2, 2, 5, 4, 5, 2, 1, -3, -5, -6, -5, -4, -4, -4, -4, -1, 1, 3, 3, 1, 1, 1, 0, 0, 0, 0, 0, 3, 4, 3, 4, 2, 1, 3, 5, 5, 5, 4, 1, -2, -4, -6, -6, -4, -3, -4, -2, 0, 3, 3, 3, 3, 3, 1, 0, 0, 1, 1, 1, 3, 3, 3, 3, 2, 3, 5, 6, 6, 7, 5, 2, 0, -3, -5, -4, -3, -2, -4, -2, 0, 2, 3, 3, 2, 1, 2, -1, -1, 0, 0, 1, 1, 2, 3, 2, 2, 3, 5, 7, 7, 7, 5, 2, -1, -4, -6, -5, -3, -2, -3, -1, 1, 2, 4, 2, 1, 1, 1, 0, -1, -1, -1, 0, 0, 1, 1, 2, 4, 4, 5, 6, 6, 5, 3, 0, -4, -6, -7, -5, -4, -1, -1, -1, 0, 2, 4, 4, 3, 1, 1, 0, -2, -2, -1, 0, 0, 0, 1, 1, 3, 5, 5, 4, 5, 4, 0, -1, -4, -6, -7, -6, -5, -3, -1, 0, 0, 1, 3, 3, 3, 2, 0, -1, -3, -4, -2, -1, -2, 0, 0, 0, 3, 2, 4, 4, 3, 2, 0, -1, -3, -3, -5, -6, -5, -3, -3, -1, -1, 1, 3, 3, 3, 2, 1, -2, -3, -2, -3, -1, -1, -1, 0, 0, 0, 1, 2, 3, 2, 3, 2, -1, -3, -3, -6, -5, -6, -5, -5, -3, -1, 1, 3, 2, 2, 2, 1, -1, -2, -2, 0, -1, 0, 0, 0, 1, 0, 0, 0, 3, 2, 1, 0, 0, -3, -6, -6, -7, -6, -6, -6, -4, -3, 1, 3, 3, 2, 2, 0, -1, -1, 0, 0, 1, 1, 1, 2, 0, 0, 0, 1, 0, 2, 1, 0, -2, -4, -6, -7, -8, -7, -7, -7, -7, -2, 0, 3, 2, 3, 2, 1, -1, 0, 0, 0, 0, 2, 1, 2, 0, 0, 0, 0, 0, 1, 0, -1, -3, -6, -7, -8, -9, -8, -9, -7, -7, -3, 0, 3, 2, 2, 3, 2, 0, 0, 0, 0, 1, 0, 1, 2, 0, 0, 0, 1, 1, 1, 0, -2, -4, -6, -8, -10, -9, -9, -7, -8, -8, -4, 0, 3, 3, 2, 4, 2, 0, 1, 2, 1, 1, 1, 2, 1, 2, 0, 0, 1, 0, 1, 0, -1, -5, -7, -10, -9, -11, -8, -8, -7, -7, -3, 1, 4, 2, 3, 5, 5, 2, 3, 3, 2, 0, 0, 2, 2, 1, 0, 1, 0, 0, -1, 0, -2, -6, -7, -8, -8, -10, -9, -6, -6, -5, -1, 1, 4, 1, 3, 5, 6, 3, 3, 4, 1, 0, 1, 1, 3, 2, 0, 0, 0, 0, 0, -1, -2, -5, -6, -8, -8, -7, -5, -4, -3, -1, 0, 3, 4, 2, 2, 5, 7, 4, 4, 2, 1, 2, 0, 1, 2, 2, 0, 0, -1, -1, 0, -2, -3, -4, -5, -6, -4, -4, -2, -1, 0, 1, 3, 4, 6, 3, 4, 5, 7, 5, 3, 2, 2, 2, 0, 0, 0, 0, -1, -1, -2, -1, -2, -3, -3, -6, -6, -5, -4, -2, 0, 1, 2, 6, 7, 6, 5, 4, 3, 4, 6, 6, 4, 3, 2, 2, 0, 0, 0, 0, -1, -4, -3, -5, -4, -4, -5, -5, -6, -4, -1, 0, 0, 2, 3, 4, 7, 7, 5, 4, 1, 2, 4, 3, 3, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -2, -2, -1, -1, 0, 0, 0, 2, 1, 3, 4, 3, 2, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 1, 2, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 4, 3, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -2, -3, -1, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, -1, 1, 1, 2, 3, 3, 3, 3, 1, 1, 3, 1, 0, -1, 0, 0, 0, -1, -2, -2, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -3, -3, -1, 0, 0, 0, 1, 1, 0, 0, -1, -1, -1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 2, 1, 1, 0, 0, -1, -1, -2, -1, 0, -1, 0, 1, 1, -1, -1, -2, -1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 0, -1, -2, -3, -1, -1, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 2, 2, 3, 1, 1, 0, -2, -3, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 3, 3, 3, 1, 0, 0, -1, -2, 0, 1, 0, 0, -1, 0, -2, 0, 1, 0, 1, 0, 2, 2, 0, 0, 0, 1, 1, 2, 1, 1, 1, 1, 2, 3, 0, 0, 1, 0, -2, -2, 0, 0, 1, -1, -1, 0, -1, -1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 1, 3, 3, 1, 2, 1, 0, -1, 0, -1, -3, -1, -1, 1, 1, -1, 0, 0, -1, 0, 2, 1, 0, 1, 1, 1, 0, 1, 1, 1, 1, 2, 2, 3, 3, 2, 1, 0, -1, -2, 0, -1, -2, -2, -2, 0, 0, 0, 0, -1, -1, 0, 1, 1, 0, 1, 2, 1, 0, 0, 0, 0, 2, 0, 2, 2, 3, 2, 1, 1, -1, -1, -1, -1, -3, -3, -2, -2, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 2, 2, 0, 0, 0, 0, 1, 1, 1, 2, 3, 2, 2, 0, 0, 0, 0, -2, -3, -3, -3, -3, -1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 2, 1, 0, 1, 0, 1, 2, 1, 0, 2, 2, 3, 3, 1, 0, 0, 0, -1, -4, -3, -2, -3, -1, 0, -2, -1, -1, 0, 1, 2, 1, 2, 2, 2, 1, 2, 1, 2, 3, 1, 1, 3, 3, 2, 3, 4, 1, 0, 0, -2, -1, -2, -3, -4, -2, -1, -2, -1, 0, 0, 0, 2, 2, 1, 2, 1, 0, 1, 1, 2, 2, 2, 2, 3, 4, 3, 2, 3, 1, 0, -1, -1, -1, -1, -1, -2, -1, -1, -1, -1, -1, 0, 0, 2, 2, 2, 2, 1, 0, 1, 2, 2, 3, 4, 3, 3, 3, 2, 3, 1, 0, -1, -2, 0, -2, -1, -1, 0, -1, 0, -1, 0, -1, 0, 1, 2, 2, 2, 2, 3, 1, 1, 1, 0, 1, 2, 3, 4, 3, 2, 2, 0, 0, -1, -1, -1, -1, -1, -2, -1, -1, -1, 0, 0, -1, 0, 1, 2, 2, 3, 2, 2, 0, 0, 0, 0, 1, 2, 2, 4, 1, 2, 1, 1, 0, -1, -2, 0, -2, -2, 0, -2, 0, -1, 0, 0, 0, 1, 1, 0, 2, 2, 2, 2, 0, 1, 0, 0, 0, 1, 3, 2, 1, 1, 0, 0, 0, 0, 0, -1, -2, -1, -2, 0, -1, -1, 0, 0, 0, 0, 1, 1, 2, 2, 3, 2, 0, 0, 0, 0, 0, 0, 2, 3, 2, 1, 1, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 2, 4, 3, 0, 0, 1, 0, 1, 1, 3, 2, 1, 0, 0, 0, 0, 2, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 2, 3, 2, 1, 1, 0, 1, 0, 2, 3, 1, 0, -1, 0, 0, 1, 1, 1, -1, -1, -1, 0, 0, 0, -1, 0, -1, -1, 1, 1, 1, 1, 2, 3, 1, 1, 0, 1, 1, 1, 3, 3, 3, 0, 0, -1, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, -1, -2, 0, 0, 1, 0, 2, 3, 1, 0, 1, 0, 0, 0, 1, 3, 2, 1, 0, 0, -1, 0, 0, -1, -2, -3, -3, -1, -1, -1, -1, 0, -1, -2, 0, 1, 0, 2, 1, 3, 4, 3, 2, 1, 1, 0, 1, 3, 3, 1, 0, 0, -1, 0, 0, 0, -2, -4, -3, -3, -2, 0, -1, 0, -2, -2, 0, 1, 2, 2, 1, 3, 3, 1, 2, 2, 2, 1, 3, 3, 3, 2, 2, 0, 0, 0, 2, 1, 0, -2, -2, -3, -1, -1, 0, -1, -2, -3, -2, 0, 0, 2, 0, 1, 1, 2, 2, 2, 1, 1, 2, 3, 3, 3, 4, 4, 3, 3, 3, 3, 2, 0, -1, -1, 0, -1, -1, -1, 0, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 3, 4, 4, 5, 3, 2, 3, 3, 2, 2, 1, 0, 1, -1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 2, 3, 0, 2, 1, 2, 1, 1, 1, 0, 0, -1, 0, -1, -3, -4, -3, -3, -2, -3, -3, -1, 0, -2, -1, 0, 0, 1, 1, 1, 2, 2, 4, 4, 3, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, -2, -2, -1, -3, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 3, 5, 2, 2, 1, 1, 0, 0, 0, -1, 0, -2, -2, 0, -1, -2, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 4, 1, 1, 1, 0, 0, 0, -1, -1, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, -1, -1, 0, 0, 2, 1, 1, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -3, -3, -2, -1, -1, -2, -1, 3, 1, 1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -2, -2, -3, -4, -3, -2, -3, -3, 0, 2, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, -2, 0, 0, -1, -1, -1, 0, -1, -1, -2, -3, -1, -3, -3, -2, -3, -1, -1, 1, 0, 2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, -2, -2, -1, -2, -3, -3, -2, -2, 0, 1, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, -2, -2, -2, -1, -3, -3, -1, -1, 0, 3, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, -2, -1, -1, 0, -2, -3, -2, -2, -2, -3, -3, -2, -1, 1, 2, 1, 1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, -2, 0, -1, -1, -2, -2, -1, 0, 3, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 2, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -3, -2, -1, -2, -1, -2, -1, 0, 1, 4, 1, 1, 0, 0, 0, 0, -1, -1, 0, 1, 2, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, -1, -3, -4, -2, -2, -2, -1, 0, -1, 1, 3, 1, 2, 1, 1, 1, 0, 1, 0, 1, 1, 2, 1, 1, 0, 0, -1, -1, 0, 1, 2, 1, 0, -2, -2, 0, -1, -2, -2, -1, 0, 1, 3, 0, 2, 0, 0, 1, 0, 0, 0, 1, 1, 1, 2, 1, 1, 0, -1, 1, 2, 2, 1, 1, 0, -2, -2, -2, -2, -2, 0, -1, -1, 1, 3, 1, 2, 1, 0, 0, 0, 1, 1, 1, 2, 2, 2, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 1, 2, 2, 2, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, -2, -3, -3, -1, -2, 0, 0, 0, 0, 0, 3, 0, 2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -3, -1, -1, -1, -1, 0, -1, -1, 1, 3, 0, 2, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -2, -2, -2, -2, -1, -1, 1, 3, 1, 2, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, -1, -1, 0, 0, 0, -2, -3, -2, -1, -3, 0, 0, 1, 0, 2, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 1, 1, 0, 0, 0, -1, -1, -2, -2, -1, -3, -2, -1, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, -1, -1, 1, 0, -1, 0, -1, -1, -2, -3, -3, -3, -2, -2, -1, 0, 2, 0, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, -2, -1, -3, -3, -2, -3, -4, -4, -2, -1, -1, 2, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 1, 1, -1, -1, -3, -3, -3, -2, -4, -4, -3, -2, -2, -1, 2, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, -1, -1, -3, -3, -2, -4, -3, -4, -2, -2, 0, 3, 0, 2, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -2, -3, -3, -3, -2, -1, -2, -2, -1, 0, 3, 0, 2, 2, 1, 2, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, -1, -2, -2, -3, -4, -2, -1, -1, 0, -1, -1, 1, 3, 0, 3, 1, 0, 2, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 2, 0, 0, 0, -1, -2, -3, 0, 0, 0, 1, 0, 0, 2, 4, 2, 3, 2, 1, 2, 1, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 1, 1, 2, 2, 3, 2, 5, 2, 1, 1, 2, 1, 0, 1, 1, 0, 0, 0, -2, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, -1, -1, 0, 2, 1, 2, 3, 3, 3, 4, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 2, 2, 3, 3, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, -3, -3, -1, 0, 1, 2, 0, 0, 0, 1, 2, 4, 4, 3, 4, 3, 3, 1, 2, 0, 0, 0, 0, 1, 1, 2, 4, 4, 4, 4, 1, 1, 0, 0, 0, -1, 0, 2, 2, 0, 0, 1, 2, 3, 2, 3, 3, 3, 2, 2, 0, -1, -2, -1, 0, 1, 1, 0, 0, 1, 3, 1, 0, 1, 1, 1, 0, 1, 0, 2, 2, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 2, 0, 1, 2, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 2, 1, 0, 1, 0, 1, 2, 1, 2, 2, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, 2, 1, 0, 1, 2, 1, 0, 1, 1, 0, 2, 1, 2, 0, 3, 2, 1, 0, 1, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 1, 3, 2, 2, 1, 1, 0, 0, 0, -1, 0, 0, -1, -3, 0, 0, 0, 0, 0, 3, 4, 2, 1, 0, 1, 1, 1, 1, 0, 0, 0, 1, 1, 1, 2, 1, 1, 0, -1, 0, 0, 0, -1, -2, -2, -4, -3, 0, 0, 1, 1, 0, 2, 2, 3, 3, 3, 3, 3, 2, 2, 2, 2, 0, 0, 1, 2, 2, 2, 1, 0, -1, 0, -1, -2, -2, -5, -4, -4, -2, 0, 0, 0, -1, -1, -1, 0, 1, 1, 2, 2, 2, 2, 1, 0, 0, 0, 1, 2, 2, 4, 2, 3, 2, 0, -1, -2, -3, -3, -3, -4, -1, 1, -2, -1, -1, -2, 0, 2, 0, 2, 1, 2, 2, 2, 2, 2, 2, 3, 3, 3, 2, 2, 1, 0, 0, 0, -1, -2, 0, -1, -2, -1, 0, 0, -3, -2, -2, 0, 0, 2, 2, 2, 2, 4, 4, 4, 3, 3, 4, 5, 4, 4, 3, 1, 1, -2, -2, 0, -1, -2, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 1, 0, 2, 3, 3, 3, 5, 4, 4, 5, 6, 5, 3, 3, 3, 0, -1, -1, -1, 0, -2, -2, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 2, 3, 1, 4, 4, 3, 3, 3, 3, 1, 1, 0, 1, 1, 0, 0, -1, -1, -2, -3, -1, 0, 0, 1, -1, 0, 0, -1, -1, 0, 0, 0, 2, 4, 3, 4, 5, 4, 2, 1, 1, 3, 3, 3, 3, 0, -1, 0, -1, -2, -2, -3, -2, -1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 4, 5, 5, 7, 7, 5, 4, 3, 4, 5, 6, 5, 4, 1, 0, 0, -1, 0, -3, -3, -2, 0, 0, 1, 0, 0, 1, 0, 1, 1, 3, 3, 4, 4, 5, 5, 5, 4, 4, 4, 5, 7, 6, 6, 4, 2, 0, 1, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 4, 5, 4, 4, 5, 4, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 2, 1, 2, 2, 3, 2, 3, 4, 4, 4, 3, 1, 0, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 1, 0, 0, 1, 2, 2, 2, 2, 2, 3, 3, 3, 3, 3, 2, 1, 0, 0, 0, -2, -1, -1, 0, 0, -2, -1, -2, 0, 1, 0, 0, 1, 0, 0, 0, 1, 3, 3, 2, 1, 1, 1, 2, 3, 2, 2, 2, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, -2, -2, -2, 0, 0, 1, 0, 1, 1, 1, 1, 2, 3, 1, 2, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 2, 0, 0, 0, 0, 0, -2, -3, 0, -1, 0, 0, 1, 2, 2, 2, 3, 2, 3, 2, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 1, 1, -1, -1, -2, -1, -2, -1, 0, 1, 0, 1, 2, 3, 2, 2, 2, 2, 3, 2, 2, 2, 0, 2, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, -2, -1, 0, 0, 0, -3, 0, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, -1, 0, 0, 0, -1, -3, -2, -3, -3, -2, -1, -1, 0, -1, -3, -1, 0, 0, 0, 0, 2, 4, 2, 0, 1, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, -1, -3, -5, -3, -3, -3, -2, 0, -1, 0, -1, 0, 0, 1, 1, 2, 3, 4, 5, 2, 1, 1, 1, 0, 0, 1, 2, 0, -1, -1, -1, -1, -3, -3, -6, -5, -4, -3, -2, 0, 0, 0, -1, 0, 2, 0, 1, 2, 3, 5, 4, 3, 2, 2, 2, 1, 1, 0, 1, 1, 1, -1, -2, 0, -2, -3, -3, -3, -3, -2, -2, 0, 0, 0, -1, 0, 1, 0, 1, 2, 4, 5, 4, 3, 3, 4, 3, 2, 3, 2, 3, 3, 2, 1, 0, -2, -2, -2, -2, -2, -1, -1, -2, 0, 0, -2, -3, -4, -2, -2, -2, -1, -2, 0, 0, 0, 0, 0, 1, 1, 2, 4, 2, 1, 0, 0, -2, -4, -4, -1, 0, 0, 0, 0, -3, -1, 1, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, -2, -2, -2, -2, -3, -2, -2, -1, -2, -2, -1, -2, -3, -3, 0, 0, 0, 0, 0, 1, 1, 3, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 2, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 2, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -2, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, 0, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, -2, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 2, 1, 1, 3, 2, 3, 3, 1, 1, 0, 0, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -2, -2, -2, -2, -1, -1, 0, 0, 1, 1, 0, 0, 1, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -2, -2, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, 0, 0, 1, 0, 0, 0, 1, 2, 2, 1, 2, 1, 0, 0, 1, 1, 2, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 2, 2, 0, 0, 0, 1, 1, 0, 1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -2, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -2, -2, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -2, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 2, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 3, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 2, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, -1, -2, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, 0, -1, -2, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 1, 2, 1, 1, 1, 2, 1, 1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, -2, -2, -1, -2, -1, 0, 0, 0, 0, 1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, -1, 0, -1, 0, -2, -2, -1, -2, -2, -2, -1, -2, -2, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, 0, 0, 0, -1, -1, -3, -3, -3, -3, -3, -3, -3, -2, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -2, -2, -2, -1, -2, -2, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -2, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -1, -1, -1, -2, -2, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -2, -3, -1, -2, -1, -1, -1, 0, 0, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 0, 1, 1, 0, 0, 0, 0, 0, -2, -2, -3, -3, -2, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, -1, 1, 0, 1, 0, 1, 1, 2, 2, 1, 1, 0, 1, 0, 0, 0, 0, -1, -3, -3, -1, -1, -1, -1, -1, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 2, 2, 2, 1, 2, 1, 1, 0, 0, 1, 1, 0, -1, -2, -2, -3, 0, 0, -1, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 2, 1, 1, 0, 0, 0, 1, 2, 3, 1, 0, -1, -1, -2, -1, 0, -2, -2, -1, -1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 1, 0, 1, 1, 2, 1, 3, 1, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 2, 0, -1, 0, 0, 1, 0, 0, 2, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, -1, 0, 2, 1, 1, 0, 0, 0, 1, 1, 0, 2, 1, 0, 1, 0, 0, -1, -3, -2, -2, -2, -1, -1, 0, -2, 0, 0, 2, 1, 2, 1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, -1, -2, -2, -1, -1, -1, -1, -2, -1, 0, 0, 1, 0, 1, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, -1, -1, -1, -2, -1, -1, -2, -2, -1, -1, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, -1, 0, -2, -2, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, -2, -2, -2, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, -1, 0, -1, -1, -2, 0, -2, -1, 0, 1, 2, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -2, -2, -1, -2, -1, -2, -2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -1, -1, -1, -2, -1, -2, -1, -2, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, -1, -2, 0, -1, -2, -2, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, -2, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 2, 2, 2, 1, 2, 0, 0, 1, 1, 2, 2, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 2, 2, 1, 0, 0, 1, 1, 1, 2, 2, 2, 1, 1, 3, 3, 3, 2, 1, 0, 1, 0, 0, 0, 0, 0, -1, -2, -2, -1, -3, -1, -1, -1, 0, 0, 0, 0, 0, 2, 2, 2, 2, 2, 1, 0, 4, 2, 1, 1, 1, 0, 0, -1, 0, 0, 0, -2, -3, -3, -2, -3, -2, 0, 0, -1, 0, 0, 0, 1, 3, 4, 5, 4, 3, 5, 3, 0, 2, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 2, 3, 3, 4, 2, 3, 3, 2, 0, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 1, 0, 1, 3, 1, 1, 2, 2, 4, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -2, -2, -1, 0, 0, 0, 1, 0, 1, 1, 2, 2, 0, 3, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, -1, -1, -1, 0, 0, 1, 2, 4, 0, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, -3, -2, -2, -3, -2, -2, 0, 1, 2, 2, 0, 1, 0, -1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, -3, -3, -3, -3, -3, -2, -1, 0, 2, 3, 0, 0, -1, -2, 0, 0, 1, 2, 1, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, -1, -1, -3, -2, -2, -4, -3, -3, 0, 0, 2, 3, 0, 1, -2, -1, 0, 1, 0, 2, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, -2, -1, -2, -3, -3, -2, 0, 2, 3, 2, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, -1, -4, -3, -1, -3, -3, -1, 0, 1, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, -3, -4, -2, 0, -3, -1, -3, 0, 1, 4, 4, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 1, 0, 0, 0, 2, 1, 0, 0, -1, -3, -2, -1, -1, -3, -1, 0, 2, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 1, 1, 0, 0, 0, 3, 3, 1, 1, 0, -2, -4, -1, -1, -1, -1, -1, 0, 2, 3, 2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 2, 3, 2, 2, 0, -2, -4, -1, -1, -1, -2, 0, 0, 0, 3, 2, 0, 2, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 1, 0, 1, 3, 5, 3, 1, 0, -3, -3, -3, 0, -1, -1, 0, 0, 0, 1, 2, 0, 2, 0, -1, -1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 2, 2, 2, 4, 2, 0, 0, -2, -4, -1, -1, -1, 0, 0, 0, 0, 2, 3, 0, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 3, 1, 0, 0, -3, -2, -3, 0, 0, 0, 1, 0, 1, 1, 2, 0, 2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, -3, -3, -2, -1, 0, 0, 0, 0, 0, 2, 2, 0, 2, -1, -1, -2, -2, 0, 0, 0, -1, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, -2, -3, -2, -1, 0, 0, 0, 0, 1, 3, 3, 0, 3, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, -3, -3, -2, -1, -1, -1, 0, 1, 2, 1, 0, 2, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 1, 0, 1, 2, 0, -1, 0, -3, -3, -3, -2, -1, -2, -1, 0, 1, 2, 2, 0, 1, 0, 0, -1, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, -2, -3, -3, -3, -2, -1, 0, 0, 0, 2, 3, -1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, -1, 0, -1, 0, 1, 0, 0, -1, -2, -4, -4, -4, -2, -2, -1, -1, 0, 0, 1, 2, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -2, -4, -4, -3, -3, -2, -2, -2, -1, 0, 3, 3, 0, 3, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, -2, -4, -5, -3, -2, -2, -2, -1, 0, 2, 4, 4, 0, 3, 2, 0, 1, 0, 0, 0, 0, 2, 0, 0, 0, 0, -1, -1, 0, 1, 0, -1, -3, -3, -5, -3, -3, 0, -2, 0, 0, 1, 4, 3, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 1, 0, 0, -1, -3, -3, -4, -3, -2, 0, 0, 0, 1, 1, 3, 4, 0, 3, 1, 0, 0, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -3, -1, 1, 2, 3, 2, 1, 2, 4, 3, 0, 4, 2, 0, 0, 0, 0, 1, 1, 0, -2, -1, -1, 0, 0, -1, 0, 0, 0, -2, 0, -1, -1, -1, 2, 3, 4, 4, 3, 2, 4, 4, -1, 3, 2, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, -1, -2, -1, -1, 0, 0, -2, -1, -1, 0, 1, 2, 4, 3, 4, 3, 3, 5, 4, 0, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 3, 2, 3, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 0, 0, 2, 1, 1, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 1, -1, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, -1, 1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, -2, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -2, -2, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, -1, -1, -1, -1, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 3, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 2, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 2, 2, 1, 1, 1, 3, 0, 0, 0, 0, 1, 1, 1, 0, 0, 2, 3, 0, 0, 1, 0, 2, 4, 2, 1, 0, 0, 2, 2, 2, 2, 2, 3, 3, 0, 0, 0, 2, 0, 2, 1, 0, 1, 0, 2, 0, 1, 0, 2, 0, 1, 0, 0, 2, 3, 3, 1, 0, 0, 3, 2, 3, 2, 1, 5, 3, 0, 1, 1, 1, 0, 1, 1, 1, 0, 1, 1, 2, 0, 1, 2, 1, 0, 0, 0, 2, 2, 2, 1, 1, 0, 2, 2, 2, 1, 2, 5, 4, 2, 0, 0, 1, 0, 1, 0, 0, 0, 1, 2, 1, 0, 0, 1, 0, 0, 0, 0, 3, 1, 0, 2, 1, 0, 3, 4, 2, 2, 3, 4, 3, 0, 0, -3, 1, 0, 0, 0, 0, 0, 2, 3, 1, 0, 0, 1, 0, 0, 0, 0, 2, 2, 0, 2, 4, 0, 3, 3, 1, 2, 3, 3, 2, 2, 1, -2, 0, 0, 1, 0, 0, 1, 2, 3, 1, 0, 0, 1, 1, 1, 0, 0, 2, 1, 0, 3, 2, 2, 3, 4, 1, 2, 3, 2, 3, 2, 1, -3, 0, 0, 1, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 1, 2, 2, 3, 3, 4, 2, 3, 1, 0, -2, 0, 0, 1, 0, 0, 1, 1, 2, 1, 0, 0, 0, 1, 0, -1, 0, 0, -1, -1, 1, 0, 0, 4, 3, 2, 3, 3, 2, 4, 3, 1, -3, 0, 0, 3, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, 0, 0, 0, 1, 2, 1, 4, 4, 4, 5, 3, 2, -2, 0, 0, 2, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, -1, -2, 0, 0, -1, -1, -1, 0, 0, 2, 2, 1, 6, 3, 3, 4, 3, 0, 0, 0, 0, 2, 0, 2, 2, 1, -1, 0, 0, 0, -1, -1, -1, -2, -2, -1, -1, -1, 0, 0, 1, 2, 1, 1, 4, 4, 2, 4, 3, 1, 0, 1, 0, 1, 0, 2, 3, 0, 0, 0, 0, -1, 0, -2, -2, -3, -3, -3, -1, 0, 0, 0, 0, 1, 0, 1, 3, 3, 1, 2, 1, 0, 1, 1, 0, 1, 0, 2, 4, 0, 0, 0, -1, -1, 0, -2, -3, -4, -2, -4, -3, 0, -1, 0, 1, 0, 0, 2, 3, 3, 1, 1, 2, 0, 0, 1, 0, 1, 1, 2, 4, 1, 0, 0, -1, -1, -2, -3, -2, -3, -4, -3, -4, -1, 0, 0, 0, 0, 0, 0, 2, 2, 1, 2, 2, 0, 0, 1, 0, 1, 2, 3, 2, 1, 1, 1, 0, -1, -3, -1, -2, -5, -4, -2, -3, -2, -2, 0, 0, 0, -1, 0, 1, 2, 2, 0, 1, 0, -2, 1, 0, 3, 1, 2, 2, 1, 1, 0, 0, -1, -3, -3, -3, -5, -5, -3, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, -1, -1, 2, 0, 2, 0, 2, 2, 1, 2, 0, 0, 0, -2, -3, -3, -5, -7, -3, -1, -1, 0, -2, 0, 0, 0, 1, 2, 2, 1, 0, 1, 0, -1, 1, 0, 3, 1, 1, 2, 1, 0, 1, -1, -1, -2, -3, -5, -4, -4, -2, 0, -1, 0, -2, 0, 2, 0, 2, 3, 2, 0, 0, 1, 0, -1, 0, 0, 4, 0, 2, 5, 3, 1, 2, 1, 1, 0, -2, -4, -5, -3, 0, -1, -1, 0, -3, -1, 2, 2, 4, 3, 2, 0, 0, 0, 0, -2, 1, 0, 2, 0, 1, 4, 3, 1, 1, 1, 0, 0, 0, -2, -3, -4, -1, -1, 0, 0, -2, 0, 4, 3, 4, 4, 1, 2, 1, 1, 0, -2, 0, 0, 2, 0, 1, 4, 3, 0, 1, 1, 0, 1, 0, 0, -3, -2, -2, -2, 0, 0, 0, 1, 4, 4, 5, 3, 2, 2, 2, 0, 0, -4, 0, 0, 3, 0, 3, 4, 2, 0, 0, 0, 1, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 2, 3, 4, 5, 4, 3, 4, 3, 0, 0, -3, 0, 0, 2, 0, 1, 3, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 3, 4, 4, 2, 1, 3, 2, 1, 0, -3, 0, 0, 1, 0, 1, 3, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 1, 2, 3, 1, 0, 2, 3, 3, 4, 2, 2, 2, 2, 2, 0, -3, 0, 0, 0, -1, 1, 1, 0, 0, 1, 1, 2, 0, 0, 0, -1, 0, 1, 2, 1, 1, 1, 0, 2, 3, 5, 2, 2, 2, 2, 2, 0, -1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 2, 1, 1, 0, 0, 0, 1, 1, 2, 3, 3, 1, 1, 2, 3, 3, 3, 3, 3, 2, 1, 1, -2, 0, 0, 1, 1, 1, 3, 0, 0, 2, 1, 2, 0, 0, 0, 0, 1, 0, 3, 4, 1, 1, 2, 0, 2, 1, 1, 2, 2, 1, 0, 0, -2, 0, 0, 1, 2, 0, 2, 1, 0, 2, 1, 1, 0, 0, 0, 0, 1, 0, 1, 2, 2, 2, 1, 2, 1, 0, 1, 0, 2, 3, 1, -1, -1, 2, 0, 1, 1, 0, 1, 1, 0, 2, 0, 0, 1, 0, 0, 0, 1, 0, 1, 3, 1, 1, 1, 1, 3, 1, 1, 1, 2, 2, 0, -1, 0, 3, 0, 1, 2, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 3, 2, 2, 1, 0, 1, 1, 1, 1, 0, -1, 3, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 2, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 2, 3, 3, 1, 2, 1, 1, 0, 0, -1, 0, -2, -2, -3, -4, -3, -4, -3, -3, -2, 0, -1, 0, -1, 1, 0, 1, 1, 2, 2, 3, 3, 1, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -2, -2, -1, -1, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 3, 3, 1, 2, 1, 2, 1, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 1, 2, 3, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, 1, 2, 2, 3, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, 1, 0, -1, -2, 0, 0, -1, -1, 0, -1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, -2, -1, -1, 0, -1, 0, 0, 2, 1, 2, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -1, -1, -1, -1, 0, 1, 1, 0, 0, -1, -1, 0, 1, 0, 0, 0, 1, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, -2, -2, -2, -1, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 2, 0, 0, 0, 0, -2, -1, -1, -1, -1, 0, 1, 2, 1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 2, 0, -2, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, -1, -3, -2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, -1, -2, -2, -1, 0, 0, -1, 0, 0, 1, 3, 1, 0, 0, -1, -1, 0, 0, -1, 0, 1, 1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, -2, -3, -2, 0, 0, 0, 0, 2, 3, 3, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 2, 1, 0, -1, 0, 0, 0, 1, 1, 1, 0, -1, -1, -1, -1, -1, 0, 1, 1, 2, 4, 0, 3, 1, 0, 0, 0, 1, 1, 1, 3, 3, 2, 0, 0, -1, -1, -1, 0, 1, 1, 1, 0, -1, -1, -1, 0, 0, 0, 1, 1, 1, 2, 2, 3, 0, 0, 0, 1, 2, 2, 2, 2, 2, 2, 1, 0, 1, 0, 0, 1, 2, 1, 1, 1, 0, -1, -1, 0, 0, 0, 0, 2, 3, 3, 1, 1, 0, -1, 0, 0, 1, 1, 1, 0, 2, 2, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, -1, -2, -1, 0, 1, 1, 2, 2, 1, 2, 0, 3, 0, 0, -2, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, 0, 0, 1, 2, 1, 3, 2, 0, 2, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, -1, -2, -2, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 2, 2, 3, 2, 1, 2, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, -1, -2, 0, 0, 2, 2, 3, 2, 2, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 3, 1, 2, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -2, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 1, 2, 2, 1, 2, 0, 1, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, -3, -2, -1, -1, -1, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -3, -3, -3, -2, -2, 0, 0, 1, 0, 1, 0, 0, 1, 0, 2, 1, 0, 0, 0, -1, -1, 0, 0, -1, 1, 0, 0, 0, -1, -1, -2, -3, -3, -2, -2, -3, 0, 0, 1, 2, 1, 1, 2, 1, 0, 2, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, -3, -3, -2, -1, -1, 0, -1, 0, 0, 2, 2, 1, 3, 2, 2, 1, 0, 2, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -2, -1, 0, 0, 1, 0, 0, 2, 2, 1, 3, 3, 3, 1, 1, 2, 1, 2, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, -1, -1, -3, -2, -1, 0, 1, 1, 1, 1, 2, 2, 2, 3, 2, 1, 2, 2, 1, 2, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 1, 2, 3, 3, 3, 3, 2, 0, 3, 2, 2, 2, 2, 0, 0, 1, 0, -1, -1, -1, -1, -2, -2, -2, -1, -2, -1, -2, -1, 0, -1, -1, 0, 0, 0, 2, 3, 2, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, -2, -1, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -2, -1, 0, -1, 0, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, -1, 0, 0, 0, -2, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 2, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, -2, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, -1, -1, -1, -1, -2, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 1, 1, 0, -1, -1, 0, 0, 0, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 2, 2, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 2, 1, 2, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 1, 0, 1, 0, 2, 2, 1, 1, 1, 2, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 3, 1, 1, 2, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 2, 2, 3, 3, 1, 2, 3, 1, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 2, 2, 1, 2, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 2, 1, 2, 1, 2, 2, 2, 2, 2, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 3, 1, 1, 2, 3, 4, 3, 3, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 2, 3, 2, 1, 2, 2, 3, 2, 2, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 3, 3, 2, 2, 4, 2, 2, 1, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 1, 1, 1, 2, 0, 2, 1, 1, 2, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 2, 2, 3, 3, 3, 1, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 1, 1, 1, 2, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -2, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, -1, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, -1, -1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 2, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 2, 1, 0, 1, 2, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 1, 0, 2, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 2, 1, 2, 1, 2, 2, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 1, 2, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 2, 1, 3, 1, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 1, 0, 1, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 2, 1, 1, 3, 1, 1, 1, 1, 0, 0, 0, 0, -1, -2, -1, -1, -1, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 1, 1, 1, 2, 2, 3, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 1, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, 3, 3, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 3, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 1, 1, 1, 1, 1, 0, 0, -1, -1, 0, -1, -1, -1, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 3, 6, 5, 3, 2, 2, 0, 0, 0, -1, -1, -2, -3, -4, -5, -6, -5, -4, -4, -2, -1, 0, 0, 0, 1, 1, 3, 3, 5, 3, 4, 1, 4, 5, 4, 2, 1, 2, 0, 0, 0, 0, 0, -1, -2, -4, -4, -2, -1, -3, -3, -1, -2, -2, -1, 0, 0, 1, 1, 2, 2, 2, 3, 2, 3, 4, 4, 3, 2, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, -2, -2, -1, -2, -2, -1, 0, 0, 0, 0, 2, 2, 3, 2, 4, 3, 5, 3, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, -2, -1, -2, -1, 0, 0, 0, 0, 0, 2, 3, 2, 3, 3, 1, 0, 0, 0, 0, -1, -1, 0, 1, 1, 0, 1, 2, 1, 0, 0, 0, 0, -1, -3, -2, -3, -2, -3, -3, -1, 0, 0, 1, 3, 2, 4, 2, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, 1, -1, -1, -1, -3, -3, -3, -4, -3, -4, -4, -3, -1, 0, 1, 2, 1, 4, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, -3, -3, -3, -5, -5, -4, -5, -3, -2, -1, 1, 1, 2, 3, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, -2, -2, -2, -1, -3, -2, -4, -4, -5, -5, -7, -3, -1, 0, 1, 2, 1, 2, 0, -2, -2, -1, 0, 1, 1, 1, 0, 1, -1, -1, -1, 0, 0, -1, 0, 0, -2, -2, -3, -4, -3, -5, -6, -5, -1, 0, 2, 3, 1, 2, -1, -3, -2, -2, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -3, -2, -5, -6, -3, -4, -4, -4, -1, 0, 2, 4, 1, 0, -2, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -2, -2, -2, -5, -5, -2, -4, -5, -3, -1, 0, 3, 4, 0, 1, 0, -2, -2, -2, -1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, -5, -4, -3, -4, -3, -3, 0, 1, 4, 4, 1, 1, 0, -2, -2, -1, -1, 0, 0, 2, 2, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, -3, -4, -6, -4, -1, -3, -1, 0, 1, 3, 3, 2, 2, 0, -1, 0, 0, 0, 0, 2, 3, 2, 1, 0, 0, 0, 0, 0, 1, 1, 0, -1, -1, -4, -4, -4, -2, -3, 0, 1, 3, 3, 4, 1, 5, 2, 0, 1, 1, 1, 0, 3, 3, 3, 1, 1, 0, 1, 1, 0, 3, 2, 2, 0, -2, -3, -4, -3, -3, -1, 0, 2, 2, 3, 5, 3, 4, 2, 0, 1, 2, 2, 1, 3, 4, 3, 2, 0, 1, 3, 3, 3, 2, 3, 1, 0, 0, -3, -2, -1, -2, 0, 1, 2, 3, 4, 5, 1, 5, 2, 1, 0, 0, 1, 0, 2, 1, 1, 1, 0, 1, 1, 3, 2, 1, 1, 0, -1, -1, -3, -4, -2, -1, -1, 0, 1, 3, 3, 4, 1, 5, 2, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 1, -1, -1, -3, -4, -3, -4, -3, -2, -1, 0, 2, 3, 3, 3, 2, 4, 1, -1, -1, 0, -1, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, -1, -3, -2, -3, -3, -2, -2, -2, 0, 0, 2, 4, 4, 2, 4, 0, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, -1, -1, -1, -2, -2, -2, -1, -2, -2, 0, 3, 2, 4, 2, 4, 0, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, -1, -2, -2, -3, -4, -4, -4, -3, 0, 1, 4, 2, 2, 3, 0, -1, -1, -1, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 2, 0, -1, -1, -1, -3, -4, -4, -4, -5, -3, -1, 1, 3, 3, 3, 5, 0, 0, 0, 0, -1, 0, 0, 1, 1, -1, -1, 0, 0, 0, 0, 1, 0, -1, -2, -2, -4, -6, -4, -5, -4, -5, -2, 1, 1, 3, 2, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, -1, -2, -4, -5, -6, -7, -5, -5, -5, -5, -3, 0, 1, 2, 1, 3, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -3, -4, -5, -5, -7, -6, -6, -7, -5, -2, 0, 2, 2, 3, 3, 0, 2, 2, 1, 1, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -2, -4, -5, -6, -8, -7, -7, -7, -4, -2, 1, 1, 3, 2, 4, 2, 1, 1, 1, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -2, -5, -5, -7, -8, -5, -4, -3, -3, 0, 2, 1, 2, 2, 6, 4, 3, 2, 1, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -3, -3, -5, -5, -6, -4, -2, -1, 0, 0, 1, 2, 4, 3, 5, 4, 3, 4, 3, 2, 1, 2, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, -2, -3, -3, -3, -4, -3, -1, 0, 2, 3, 2, 4, 5, 3, 7, 5, 4, 3, 2, 3, 0, 0, 1, 0, 0, -2, 0, -1, -1, -1, -2, -3, -3, -4, -2, -2, -1, 0, 2, 1, 3, 6, 4, 4, 5, 3, 6, 4, 3, 5, 4, 2, 1, 0, 0, 0, 0, -1, -1, -1, -3, -3, -2, -3, -2, -3, -2, -2, -1, 0, 0, 1, 2, 4, 5, 4, 4, 1, 1, 2, 2, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 2, 1, 2, 1, 1, 2, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, -1, -1, 0, 0, 0, -1, -1, -2, -1, -1, -2, -2, -3, -3, -2, -2, -3, -1, -2, 0, -1, -1, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, -1, -1, -2, 0, 0, 0, -2, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, -1, -1, -2, -2, -2, -1, -2, 0, -2, 0, 1, 0, -1, -1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 1, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 2, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 0, 1, 1, -1, 0, 1, 0, -1, 0, 1, 1, -1, -2, -2, 0, 2, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 1, 2, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, -2, -1, 2, 1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 1, 0, 2, 1, 3, 1, 1, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, -2, -2, 0, 2, 1, 0, -1, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 2, 2, 2, 0, 0, 2, 1, 0, 0, 0, 1, 0, 1, 1, 1, 0, -1, -1, 2, 1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 2, 3, 0, 0, 2, 1, 1, 0, 0, 0, 0, 1, 2, 1, -1, 0, -1, 2, 2, 0, -1, -3, -2, -1, 0, 0, 1, 0, 0, 0, 0, 1, 2, 3, 0, 0, 2, 0, 1, -1, 0, 0, 1, 1, 0, 1, 0, -1, 0, 1, 0, 1, 0, -1, -1, -1, -1, 0, 0, 1, 0, 0, 1, 1, 2, 1, 1, 2, 0, 0, 1, -1, -1, 0, 0, 0, 1, 2, 0, -1, 0, 2, 1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 2, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 2, 1, 0, -1, 1, 0, -1, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 2, 2, 2, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 2, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 1, 1, 0, 2, 1, 3, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, -1, 0, -1, -2, 0, -1, 0, -1, 0, 0, 0, 1, 1, 0, 1, 2, 1, 1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, -1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, -1, 1, 2, 2, 1, 1, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 2, 3, 2, 2, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -2, 0, 2, 1, 0, -1, 0, 0, 1, 0, 0, 0, 1, 2, 1, 0, 0, 0, 1, 2, 2, 1, 1, 1, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 1, 0, -1, 0, 1, 2, 3, 2, 0, 0, 0, 1, 1, 3, 2, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 2, 2, 1, 0, -1, 0, 0, 2, 2, 1, 0, 0, 1, 2, 2, 2, 2, 1, 0, -1, -2, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 0, 0, 0, 0, 1, 3, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, -2, -1, 0, 2, 2, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 2, 1, 1, 0, -2, -2, 0, 1, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, 0, 0, 0, 1, 1, 2, 1, -1, -2, 0, 2, 2, -1, -1, 0, -1, -2, 0, 1, -1, 0, 0, 0, -1, 0, -1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, -2, 0, 2, 2, 0, -1, -1, -1, -2, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 2, 2, 0, 0, -1, 0, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -2, -1, -1, -1, -1, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, -2, 0, 1, 3, 1, 0, 0, 0, 0, 0, -1, -2, 0, -2, -1, -1, 0, -1, -1, -2, -2, -2, -2, -1, -1, 0, -1, 0, -1, -1, 0, -1, -1, 1, 1, 2, 0, 0, 0, 1, 0, -1, -1, 0, 0, -1, 0, -1, 0, -1, -2, -2, -1, -1, -1, -2, -1, -1, -1, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, 0, 1, 2, 2, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 5, 5, 4, 3, 3, 2, 0, 1, 1, 0, 0, 0, -2, -2, -3, -1, -3, -2, -3, -4, -4, -2, -2, -2, -3, -2, -1, 0, 0, 2, 2, 3, 6, 5, 4, 3, 2, 1, 1, 1, 0, 0, -1, -2, -2, -2, -2, -1, -2, -1, -2, -4, -3, -3, -5, -3, -3, -3, -2, -2, -1, 0, 1, 2, 5, 5, 3, 1, 1, 2, 1, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, -3, -2, -3, -3, -3, -2, -1, -1, -1, -2, -1, 1, 3, 4, 4, 2, 2, 2, 1, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 2, 0, 0, 0, -2, -1, -3, -2, -1, 0, -1, -2, -3, 0, 0, 1, 2, 3, 1, 2, 2, 1, 1, 1, 2, 1, 2, 0, 0, 1, 2, 2, 2, 1, 0, 0, -1, -1, -1, -1, -1, -1, -2, -2, -2, -2, 0, 1, 3, 3, 1, 1, 3, 1, 2, 1, 3, 3, 1, 0, 0, 0, 2, 1, 2, 2, 0, 0, -1, -2, -1, 0, -2, -1, -1, -2, -4, -1, 0, 2, 3, 1, 0, 1, 2, 2, 1, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, -2, -1, -3, -3, -3, 0, 2, 1, 0, 0, 0, 1, 1, 0, 0, 2, 1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 1, 0, -3, -2, -2, -1, -2, -1, -2, -4, -2, 0, 1, 1, 0, -1, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, -2, -2, -2, -2, -1, 0, -1, -3, -1, 1, 0, 2, -1, -4, -4, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -2, -3, -2, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 2, 0, 0, -4, -3, -1, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, -2, -3, -1, -1, 0, -1, -1, -1, 0, 1, 0, 1, 0, -1, 0, 0, 0, -1, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 3, 1, 0, -2, -4, -1, -1, -2, 0, 0, -1, 0, 2, 1, 3, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 3, 1, 0, -2, -2, -2, -1, -1, 0, 0, 0, 0, 2, 2, 4, 3, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 1, 1, 2, 1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 2, 2, 3, 3, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 2, 2, 2, 0, -1, -1, -2, -2, 0, 0, 0, 0, 0, 2, 2, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 1, 0, -2, -2, -3, -1, -1, 1, -1, -1, 0, 2, 2, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 1, 1, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 2, 2, 3, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, -1, -2, 0, -1, 0, 0, 0, -1, -1, 0, 1, 1, 1, 0, -1, -1, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, -2, 0, 2, 2, 2, 1, 0, 0, -2, 0, 0, 1, 2, 1, 1, 0, -1, 0, 0, 2, 1, 2, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, -1, -1, 0, 1, 2, 1, 0, 0, 0, -1, 0, -1, 0, -1, -1, -2, -1, -1, 0, 2, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, -1, -1, -1, 0, -1, -1, -3, -3, -1, 0, 1, 1, 1, 1, 0, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -3, -3, -1, -2, -2, -1, -2, -4, -1, 1, 1, 0, 1, 2, 0, 1, 0, 0, 1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -3, -3, -1, -1, -2, -4, -3, -2, 0, 0, 1, 2, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, -2, -2, -3, -2, -2, 0, -2, -2, -2, -1, 0, 2, 3, 3, 1, 2, 0, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -3, -3, -3, -2, -1, -1, -2, -1, -1, 0, 1, 2, 4, 4, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -2, -2, -3, -4, -3, -3, -2, 0, -1, -1, -1, 0, 2, 1, 5, 5, 3, 2, 3, 0, 0, 1, 0, 0, -2, 0, 0, -2, 0, -1, -1, -1, -3, -4, -2, -4, -3, -3, -1, -1, 0, -1, 0, 0, 0, 1, 4, 4, 3, 3, 3, 3, 2, 0, 0, -1, 0, -1, 0, -1, -2, -2, -2, -2, -3, -3, -2, -2, -2, -3, -1, -1, -1, -1, 0, 0, 2, 0, 4, 4, 3, 3, 2, 1, 1, 1, 0, 0, -1, 0, 0, 0, -2, -1, -2, -2, -4, -4, -3, -2, -1, -1, -1, -1, 0, 0, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 2, 2, 1, 1, 2, 1, 2, 3, 1, 0, 0, 4, 2, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, -2, 0, 0, 0, 0, 0, 1, 2, 3, 4, 3, 4, 3, 4, 3, 1, 0, 2, 2, 1, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, -2, 0, 0, 0, 0, -2, -2, 0, 1, 2, 2, 2, 3, 2, 3, 3, 5, 2, 0, 2, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -3, -1, 0, 0, 1, 3, 2, 2, 3, 4, 4, 2, 0, 3, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, -1, 0, 0, 0, 1, 3, 3, 2, 0, 3, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -2, -1, -1, -2, -1, 0, 0, 0, 2, 2, 3, 0, 3, 1, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -2, -2, -3, -2, -1, 0, 0, 2, 2, 3, 0, 2, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -4, -4, -4, -4, -1, 0, -1, 1, 2, 3, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, -5, -4, -4, -3, -4, -1, 0, 0, 3, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 2, 1, 0, -1, -1, -3, -4, -3, -2, -2, -4, -3, -1, 0, 2, 2, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 2, 0, 0, -2, -4, -4, -3, -3, -2, -2, -1, -1, 0, 2, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 2, 3, 0, 0, -1, -3, -3, -3, -2, -3, -2, -2, -2, 0, 2, 2, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 3, 3, 1, 0, -1, -3, -4, -2, -1, -2, -1, -2, -2, 0, 3, 2, 0, 3, 0, 0, 0, -1, 0, -1, 0, 1, 2, 1, 0, 0, 0, 2, 4, 4, 1, 0, -2, -4, -3, -3, -2, -2, -2, -1, -1, 0, 1, 1, 0, 2, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 1, 0, 1, 1, 4, 4, 2, 0, -1, -3, -3, -3, -2, -2, -1, -2, -2, 1, 2, 2, 0, 2, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 2, 4, 4, 2, 1, -1, -3, -3, -3, -1, -1, -1, -2, -1, 0, 1, 2, 0, 2, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 2, 2, 3, 4, 4, 1, -1, -2, -2, -3, 0, -1, 0, -1, 0, 0, 2, 1, 0, 3, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 1, 1, 0, 2, 4, 3, 2, 0, 0, -2, -2, -3, -2, 0, 0, -1, 0, 0, 2, 2, 0, 2, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 2, 2, 3, 1, 1, 0, -1, -4, -3, -3, -1, 0, 0, 0, 0, 0, 1, 2, 0, 2, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 3, 2, 1, 0, 0, -1, -3, -2, -2, -1, -1, -1, 0, 0, 0, 1, 2, 0, 2, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, -2, -2, -2, -1, -2, -2, -1, 0, -1, 0, 0, 2, 0, 3, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 0, -1, -2, -3, -3, -2, -2, -2, -1, -1, -1, 0, 0, 1, 0, 2, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, -1, -2, -3, -4, -3, -3, -2, -1, -1, -1, 1, 1, 0, 3, 0, 0, -2, -1, -1, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -2, -3, -3, -4, -3, -3, -1, -3, -2, 0, 2, 3, 0, 4, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, -1, -2, -3, -4, -3, -2, -3, -2, -2, -1, 0, 2, 2, 0, 4, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, -3, -3, -4, -4, -3, -3, -3, -1, 0, 1, 1, 2, 0, 4, 0, 1, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, -1, -1, 1, 0, 0, -2, -3, -4, -4, -4, -3, -1, -2, -2, -1, 0, 1, 3, 0, 4, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 1, -1, -2, -4, -4, -4, -4, -2, -1, -1, 0, 0, 0, 2, 2, 0, 3, 2, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, -3, -3, -2, -1, 0, 0, 0, 0, 1, 3, 3, 1, 0, 3, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -2, -1, -1, 0, -1, -1, -2, 0, -1, 0, 1, 2, 1, 1, 2, 4, 4, 3, 0, 2, 1, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, -1, -2, -2, 0, 0, -1, 0, 0, -1, 0, 0, 2, 1, 2, 2, 3, 4, 4, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 2, 2, 3, 3, 2, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 1, 1, 1, 1, -1, 1, 2, 1, 3, 2, 3, 2, 0, 0, 1, 2, 1, 2, 2, 0, 1, 1, 1, 0, 0, 2, 1, 1, 1, 0, 0, 2, 2, 0, 1, 2, 0, 0, 4, 2, 3, 1, 1, 2, 0, 0, 1, 2, 0, 0, 0, 0, 1, 3, 1, 0, 1, 1, 2, 3, 1, 0, 1, 3, 2, 0, 0, 2, 0, 0, 3, 3, 3, 3, 2, 3, 2, 1, 1, 1, 0, 0, -2, 0, 2, 2, 2, 1, 1, 1, 2, 2, 1, 0, 1, 2, 2, 0, 0, 0, 0, 0, 2, 2, 2, 3, 1, 2, 3, 0, 1, 1, 0, 0, -2, 0, 2, 0, 1, 2, 2, 0, 2, 2, 0, 2, 0, 2, 3, 1, 0, -1, 0, 0, 3, 0, 2, 2, 1, 2, 3, 0, 0, 0, 0, 0, -1, 0, 2, 1, 0, 3, 1, 0, 2, 2, 0, 2, 0, 3, 3, 1, 0, 0, 0, 0, 1, 0, 1, 3, 3, 3, 1, 0, 0, 0, 0, 0, -1, 1, 3, 0, 0, 4, 1, 1, 2, 3, 1, 3, 0, 2, 2, 1, 0, -1, 0, 0, 2, 0, 2, 3, 3, 3, 0, 1, 1, 0, 2, -1, 0, -1, 0, 0, 0, 1, 0, 1, 2, 2, 1, 2, 1, 1, 3, 2, 0, 0, 0, 0, 1, 0, 1, 0, 2, 2, 1, 1, 0, 1, 0, 0, -2, 0, 0, -1, 0, 1, 0, 0, 2, 0, 2, 3, 1, 3, 4, 0, 1, 0, 0, 0, 2, 0, 0, 0, 0, 2, 1, 0, 0, 0, -1, -1, -2, -1, 0, -2, -1, 1, 1, 0, 2, 0, 2, 3, 2, 1, 3, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 2, 0, -1, -1, 0, -2, -3, -3, 0, -2, -3, 0, 0, 0, 0, 0, 1, 3, 1, 1, 2, 2, 1, 1, 0, -1, 1, 0, 1, 0, 0, 0, 1, 0, 0, -1, -2, -3, -3, -3, -2, -2, -1, 0, 0, 0, 1, 1, 2, 2, 1, 1, 1, 2, 0, 1, 0, 0, 0, 1, 2, 1, 0, 0, 0, -2, -1, -2, -3, -2, -3, -4, -1, -1, -1, -1, 0, 0, 0, 1, 1, 2, 1, 0, 1, 1, 0, 3, 0, 0, 2, 2, 3, 2, -1, 0, 0, -1, -1, -3, -3, -3, -4, -4, -4, -2, -2, -2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 2, 0, 2, 0, 0, 1, 1, 3, 3, 0, -1, 0, -1, -1, -2, -3, -3, -4, -4, -3, -4, -2, -2, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 3, 1, 2, 2, 0, 0, 0, 0, -1, -2, -3, -3, -4, -4, -3, -4, -4, -2, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 2, 1, 1, 0, 1, 0, -1, 0, -4, -2, -3, -4, -4, -3, -2, -4, -1, -2, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, 1, 1, 1, 1, -1, -2, -2, -3, -4, -4, -6, -4, -2, -1, -2, -3, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 3, 1, 0, 1, 1, 2, -1, -1, -2, -4, -4, -4, -6, -3, -3, -1, -1, -2, -2, 0, 1, 0, 1, 2, 0, -1, 1, 2, 0, 1, 0, 0, 2, 1, 1, 2, 0, 1, 0, 0, -1, -2, -3, -1, -4, -2, -2, -1, -1, 0, -2, 0, 1, 1, 2, 2, 0, -1, 0, 0, 1, 0, 0, 0, 2, 1, 2, 2, 0, 0, 0, 0, 0, -1, 0, -1, -4, -3, -2, -2, 0, -1, -2, 0, 2, 2, 2, 2, 0, 0, 1, 0, 0, -1, -1, 0, 2, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -3, -3, -2, -2, 0, 0, 0, 1, 2, 2, 3, 2, 2, 3, 2, 0, 0, -1, 0, 0, 3, 1, 1, 2, 1, 0, 0, -1, 0, 0, 0, -1, -3, -2, -2, -1, 0, 0, 0, 2, 3, 3, 3, 2, 1, 3, 3, 1, 0, -1, 0, 0, 2, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, -2, -2, -1, 0, 0, 1, 0, 0, 1, 3, 2, 2, 2, 1, 3, 4, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -2, -2, -1, 0, 1, 1, 0, 1, 0, 2, 2, 3, 1, 0, 0, 2, 3, 2, 0, -1, 0, 0, 0, 0, 1, 2, 0, 0, 1, 0, 1, -1, -1, -2, 0, 0, 1, 0, 0, 0, 0, 3, 3, 2, 1, 1, 1, 2, 3, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 3, 1, 0, 0, -1, -1, 0, 1, 1, 1, 1, 0, 0, 1, 2, 1, 1, 1, 1, 3, 3, 0, 0, -1, 0, 0, 1, 1, 3, 1, 0, 0, 2, 1, 1, 0, 0, 0, 0, 1, 0, 2, 1, 0, 2, 2, 1, 0, 0, 1, 0, 2, 2, 0, 0, 0, 0, 0, 2, 1, 2, 2, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 2, 3, 0, 1, 2, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 2, 0, 0, 1, 1, 0, 0, 0, 1, 1, 2, 2, 2, 2, 2, 1, 2, 0, 0, 0, 1, 2, 1, -1, 1, 0, 0, 2, 1, 1, 1, 1, 1, 0, 0, 1, 2, 0, 0, 0, 1, 2, 0, 0, 0, 1, 0, 1, 2, 0, 0, 0, 0, 1, 1, -1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 1, 0, 1, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 2, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 3, 1, 3, 2, 0, 2, 2, 3, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 3, 1, 0, 0, -1, -1, 0, -1, 0, 0, 1, 2, 3, 3, 2, 2, 3, 3, 1, 1, 2, 3, 2, 0, -1, 0, -1, 1, 1, 0, 2, 2, 1, 2, 1, -2, -2, -2, -2, -1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 2, 2, 2, 1, 2, 3, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -1, 0, 0, -1, 0, -1, 1, 0, 1, 0, 0, 0, 2, 2, 2, 2, 3, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, -1, 1, 0, 0, 1, 1, 1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, -1, -2, -3, -1, -1, -1, 0, 0, 0, 0, 1, 0, -1, -1, 1, 3, 3, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -2, -3, -2, -2, -2, 0, 0, -1, -1, 0, 0, -1, 0, 1, 0, 1, 2, 1, 0, 1, 0, 1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, -1, -2, -1, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 1, -1, -1, 0, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, 0, 1, 1, 0, 0, 2, 0, 1, 0, 1, 0, 1, 0, -1, 0, -1, -3, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, -2, 0, 0, 0, 1, 2, 0, 0, 0, 0, 2, 1, 2, 1, 1, 1, 0, 0, -1, -2, -3, -2, -1, -1, -1, -1, -1, 1, 1, 0, 0, 0, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 2, 1, -1, -1, -2, -2, 0, -1, -2, -2, -2, -2, 0, 1, 1, 0, 0, -1, 0, 0, 1, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 2, 1, 0, 0, -2, -3, 0, 0, 0, -1, 0, -3, -1, -1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 2, 1, 1, 0, 0, -2, -2, 0, 0, 0, -1, -2, -2, -2, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 2, 4, 3, 2, 3, 2, 3, 3, 3, 1, 2, 0, 0, 0, 1, 0, -1, -2, -2, 0, 0, 1, 0, 0, 0, 0, 1, 3, 2, 2, 1, 2, 0, 1, 3, 2, 4, 2, 3, 3, 2, 2, 0, 1, 0, 1, 1, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 2, 2, 2, 1, 0, 1, 0, 0, 0, 1, 2, 3, 4, 1, 2, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 1, 3, 1, 0, 0, 0, 0, 0, 1, 1, 2, 3, 1, 1, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 3, 3, 3, 2, 1, 1, 0, -2, -1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 3, 2, 0, 0, -1, 0, 1, 2, 2, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 1, 0, 0, 0, 2, 2, 1, 1, 2, 3, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 2, 2, 0, 1, 3, 2, 3, 2, 2, 1, 0, 0, -1, 1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 1, 1, 0, -1, 0, 2, 2, 1, 2, 3, 1, 2, 0, 1, 2, 1, 0, 0, 1, 1, -1, -2, -2, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 3, 2, 0, 0, 0, 0, 0, 0, 1, 1, 0, -2, -3, 0, 0, 0, 0, -2, -2, -2, -2, 0, 0, 1, 0, 0, -2, -1, 0, 0, 1, 2, 3, 2, 2, 0, 1, 0, 0, 0, 0, 0, -1, -1, -3, -3, 0, 0, -1, -4, -4, -4, -3, -1, 0, 0, 0, -1, -1, 0, 1, 1, 0, 1, 2, 2, 3, 1, 2, 1, -1, -1, 0, 0, 0, 0, -2, -2, -3, -2, -2, -1, -4, -6, -4, 0, 0, 0, 0, -1, 0, 0, 0, 2, 2, 1, 1, 2, 2, 2, 2, 2, 1, 1, 1, 0, 0, 0, -1, -1, -1, -1, 0, 0, -2, -2, -3, -1, 0, 0, 0, -1, -2, -1, 0, 0, 1, 1, 2, 2, 2, 3, 4, 3, 3, 2, 3, 2, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -3, -2, -1, -1, -1, -1, -1, 0, 0, 1, 1, 1, 0, 1, 2, 2, 2, 2, 2, 0, 0, 0, 0, 1, 2, 2, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 1, 2, 1, 0, 0, 1, 2, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, -1, 0, -1, -2, -1, -1, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -2, -1, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, -2, -1, 0, 1, 1, 1, 0, 0, 2, 1, 2, 2, 1, 2, 1, 1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 2, 1, 1, 1, 0, 0, -1, 0, -1, -2, -1, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 2, 1, 1, 0, 2, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, 1, 0, 1, 2, 1, 0, 0, 2, 1, 2, 1, 1, 3, 1, 0, 2, 0, 1, 1, 2, 1, 1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 1, 1, 2, 2, 1, 1, 1, 1, 1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 1, 1, 1, 1, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 2, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 1, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, -2, -2, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, -1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 1, 1, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 1, 0, 0, 1, 0, 1, 0, 0, 1, 2, 2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -3, -2, -2, -2, -1, 0, -1, -1, -1, 0, 0, 0, 2, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 3, 3, 1, 1, 1, 1, 0, 0, -1, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 3, 2, 3, 3, 3, 1, 1, 3, 5, 4, 3, 2, 1, 1, 2, 0, 0, -1, -2, -2, -2, -3, -2, -1, -1, -2, -2, -2, 0, 0, 1, 2, 2, 3, 3, 4, 2, 3, 1, 3, 3, 3, 1, 2, 0, 0, 0, -1, -2, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, -3, -1, 0, 0, 0, 1, 1, 2, 2, 2, 2, 1, 4, 4, 2, 2, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, -2, -2, -3, -2, -1, 0, -1, 0, 1, 2, 2, 1, 2, 0, 2, 3, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, -3, -3, -3, -3, -1, -2, 0, 1, 1, 0, 2, 1, 2, 5, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, -1, -1, 0, -1, -4, -4, -4, -4, -4, -4, -2, 0, 1, 1, 1, 1, 2, 4, 3, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 2, 0, 0, -1, -2, -6, -5, -5, -5, -5, -5, -3, 0, 0, 0, 2, 1, 3, 4, 3, 2, 0, 1, 1, 2, 2, 0, 1, 0, 0, 0, 2, 1, 0, -1, -2, -3, -4, -6, -6, -5, -6, -6, -4, 0, 0, 1, 2, 1, 2, 2, 1, 0, 0, 1, 2, 1, 2, 2, 2, 1, 0, 0, 2, 2, 1, -1, -1, -3, -5, -6, -5, -6, -6, -6, -6, -1, 0, 0, 2, 0, 2, 3, 1, 0, 1, 0, 0, 0, 2, 2, 0, 1, 2, 1, 3, 3, 2, 0, -1, -2, -4, -5, -4, -4, -4, -6, -5, -1, 1, 0, 2, 1, 1, 1, 1, 0, 0, 0, 0, 2, 1, 1, 0, 1, 1, 1, 3, 2, 2, 0, 0, -4, -4, -5, -4, -5, -5, -5, -5, -2, 0, 0, 2, 1, 2, 0, 0, 1, 1, -1, 0, 1, 0, 1, 0, 0, 1, 2, 3, 3, 3, 2, -1, -3, -4, -4, -5, -3, -5, -4, -4, -3, 0, 0, 2, 0, 2, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 3, 3, 3, 1, 0, -3, -3, -4, -3, -4, -4, -4, -4, -3, -1, 0, 3, 1, 3, 1, 0, 0, 0, 0, -1, 1, 0, 1, 1, 0, 1, 4, 4, 4, 5, 3, 0, -1, -3, -2, -3, -3, -3, -3, -5, -2, 0, 0, 2, 2, 2, 1, 0, 0, 0, -1, 0, 1, 1, 1, 1, 0, 2, 3, 5, 5, 6, 4, 0, -1, -1, -3, -2, -1, -3, -4, -3, -2, 0, 0, 2, 2, 2, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 4, 6, 6, 6, 4, 1, 0, -3, -4, -4, -2, -2, -3, -3, 0, 0, 0, 1, 0, 1, 1, -1, 0, 0, -2, -2, 0, 0, 1, 1, 2, 2, 4, 6, 7, 6, 4, 1, -1, -3, -4, -3, -1, -2, -2, -3, 0, 0, 0, 1, 2, 3, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 1, 3, 4, 6, 5, 4, 3, 1, -2, -2, -3, -3, -3, -2, -2, -3, 0, 0, 0, 2, 2, 2, 2, -1, 0, -2, -2, -3, -1, 0, 0, 0, 3, 2, 4, 4, 4, 3, 1, 0, -1, -3, -3, -3, -3, -2, -3, -3, -2, 0, 0, 2, 1, 1, 2, -1, 0, -2, -3, -2, 0, 0, 0, 1, 1, 3, 2, 4, 3, 3, 0, -1, -2, -3, -3, -5, -4, -3, -2, -3, -2, 0, -1, 1, 0, 3, 1, 0, -1, 0, -3, -2, -1, 0, 0, 0, 2, 3, 2, 2, 3, 1, 0, 0, -1, -4, -4, -5, -4, -4, -2, -4, -2, 0, 0, 2, 1, 1, 1, 0, -1, 0, -2, -2, 0, 0, 1, 1, 1, 2, 2, 2, 2, 2, 1, -1, -2, -4, -5, -5, -6, -4, -5, -5, -4, 0, 0, 1, 2, 1, 1, -1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 0, 2, 2, 0, 0, -2, -3, -5, -6, -6, -4, -5, -5, -4, -4, 0, 0, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 1, 1, 1, 0, -3, -3, -5, -5, -5, -6, -5, -4, -4, -3, -1, 1, 1, 1, 3, 2, 0, 0, 0, 0, 1, 2, 2, 1, 1, 1, 0, 2, 0, 0, 0, 0, -3, -6, -6, -7, -6, -5, -5, -5, -4, -2, -1, 0, 2, 0, 3, 3, 1, 2, 1, 1, 0, 1, 0, 3, 1, 0, 2, 2, 0, 0, -1, -2, -3, -6, -6, -6, -6, -5, -6, -4, -3, -2, 0, 1, 1, 1, 2, 5, 2, 2, 3, 1, 0, 1, 1, 1, 1, 0, 1, 0, 0, 1, 0, -1, -3, -4, -5, -6, -6, -5, -3, -3, -3, 0, 0, 1, 1, 2, 3, 4, 3, 4, 3, 2, 1, 1, 0, 3, 2, 1, 1, 0, 0, 0, -2, -2, -3, -4, -3, -4, -5, -2, -2, -2, -2, 0, 2, 2, 3, 1, 2, 5, 3, 2, 3, 1, 0, 1, 1, 2, 1, 0, -1, -1, -1, -1, -2, -2, -4, -4, -3, -2, -3, -2, -1, 0, 0, 2, 2, 1, 1, 0, 3, 4, 4, 2, 2, 0, 1, 0, 0, 0, 0, 0, -1, -3, -2, -2, -4, -3, -3, -2, -2, -2, 0, 0, 1, 2, 3, 4, 4, 2, 2, 2, 1, 3, 2, 2, 2, 1, 2, 0, 0, 0, 0, 0, 0, -2, -2, -2, -1, -2, -2, -1, -1, 0, 0, 0, 1, 2, 3, 4, 3, 1, 1, 0, 0, 1, 1, 2, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -2, -3, -2, -2, -2, -2, -2, -3, -3, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 1, 1, 0, 1, 0, 1, 1, 1, 0, -1, -1, 0, 0, -2, -2, -1, 0, 0, -3, -2, 0, -1, 0, 0, -1, -1, -2, -1, -1, -1, -2, 0, 0, -1, 0, 0, -1, 0, 0, 1, -1, 0, -1, -1, 0, -1, 0, 0, 1, 1, 0, -2, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 1, 1, 2, 1, 0, 0, 0, 1, 1, 1, 1, 1, 2, 0, -1, -1, 0, 0, 0, -2, -1, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 1, 1, 1, 0, 3, 1, 0, 1, 1, 0, 2, 0, 1, 2, 0, -1, -1, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 2, 3, 1, 0, 2, 1, 1, 0, 0, 2, 2, 1, 3, 4, 1, 0, -2, -1, 0, 0, -2, -1, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 2, 3, 1, 0, 3, 2, 1, 0, 0, 1, 4, 3, 2, 4, 0, 0, -1, -1, 0, 0, -2, -1, -1, 0, 1, 0, 1, 1, 1, 1, 0, 0, 2, 3, 2, 0, 2, 3, 1, 0, 0, 1, 4, 2, 3, 4, 1, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, 1, 1, 0, -1, 0, 3, 2, 2, 0, 2, 3, 1, 1, 0, 0, 1, 2, 2, 3, 3, 0, -1, 0, 0, 0, 0, -1, -3, -3, -2, 0, 0, 1, 1, 0, 0, 0, 2, 2, 1, 1, 2, 3, 3, 2, 0, 1, 2, 1, 0, 3, 1, 1, 0, -1, 0, 0, -1, -1, -2, -2, -2, -1, 0, 0, 1, 0, 0, 0, 1, 2, 1, 0, 2, 2, 3, 0, 0, 0, 1, 0, 0, 1, 2, 0, 0, -1, 0, 0, -1, 0, 0, -1, -3, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 1, 2, 3, 1, 0, 1, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -2, -2, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 3, 1, 0, 1, 0, 1, 0, 1, 1, -2, 0, 0, 0, -1, -2, 0, 0, -2, -1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, 1, 2, 1, 0, 0, 0, 0, 0, 2, 1, 0, 0, -1, 0, 0, -3, -1, -1, -2, -1, -2, -2, -1, -2, -2, 0, -2, -1, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 0, 2, 2, -1, 0, 0, 0, -1, -3, -2, 0, -2, -1, -3, -4, -1, -2, -2, -2, -1, -2, -1, 0, 0, 1, 1, 3, 2, 0, 0, 0, 0, 0, 1, 2, 0, 0, -1, 0, -1, -3, -2, 0, -1, 0, -1, -3, -1, -1, -1, -2, -1, -2, 0, 0, 1, 2, 1, 3, 1, 0, 0, 1, 1, 0, 1, 0, -1, 0, -1, 0, 0, -3, -1, 0, -1, 0, -2, -1, 0, 0, -1, -1, -2, -1, 0, 0, 1, 2, 1, 2, 1, 0, 1, 0, 0, 1, 3, 1, -2, 0, 0, -1, 0, -2, -1, -1, 0, 0, 0, -1, 1, 0, 1, 0, -1, 0, 0, 1, 2, 3, 1, 1, 1, 1, 3, 2, 2, 1, 3, 1, 0, 0, 0, 0, 1, -2, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, -1, -1, 0, 1, 2, 3, 0, 1, 1, 1, 2, 5, 2, 2, 3, 1, -1, -1, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 2, 3, 0, 2, 2, 0, 4, 3, 2, 4, 3, 1, -1, -2, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, -1, 0, -1, 0, 1, 3, 0, 2, 3, 0, 3, 3, 3, 5, 4, 0, -1, -2, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 2, 3, 2, 1, 2, 2, 2, 2, 2, 5, 4, 0, -2, -2, -1, 0, -2, -3, 0, -2, -1, -2, 1, 0, 0, 0, 0, 0, -1, 1, 0, 2, 3, 2, 1, 1, 2, 1, 2, 1, 3, 4, 4, 1, -2, -1, 0, 0, -1, -3, 0, -2, -2, -3, 0, 0, 0, -1, -1, 0, 0, 0, -1, 1, 1, 1, 1, 2, 1, 0, 2, 1, 2, 4, 4, 0, -3, -1, -1, 0, 0, -2, 0, 0, -2, -2, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 2, 2, 2, 0, 0, 1, 2, 1, 3, 3, 0, -1, -1, -1, 0, 0, -2, 0, 0, -2, -2, 0, 0, -2, -3, -2, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, -1, -2, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -3, -2, -1, -1, -1, -1, -1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, -3, 0, 0, 0, 1, -1, -1, 0, 0, 0, -1, -2, -2, -1, -2, 0, 0, -1, 0, 0, -1, -1, 0, -1, -2, 0, 0, 0, 0, -1, 0, 0, -2, 0, -1, 0, 1, 0, -2, 0, 0, 0, -1, -3, -2, -1, -1, -2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, -2, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, -1, -4, 0, 1, 0, 3, 2, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 5, 6, 4, 3, 2, 0, 0, 0, 2, 0, 0, 0, -2, -3, -4, -3, -4, -6, -4, -6, -5, -5, -4, -5, -3, -3, -2, -1, -1, 1, 2, 4, 6, 7, 4, 2, 1, 0, 0, 1, 1, 1, 0, 0, -1, -4, -3, -3, -3, -3, -5, -5, -7, -7, -6, -4, -3, -3, -3, -3, -2, 0, 0, 3, 6, 6, 4, 2, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -3, -5, -5, -4, -3, -2, -2, -3, -2, 0, 1, 2, 4, 5, 3, 1, 1, 1, 1, 1, 2, 1, 1, 1, 1, 0, 1, 0, 1, 0, 0, -1, -4, -3, -3, -2, -1, -1, -2, -2, -2, -1, 0, 2, 4, 5, 3, 1, 2, 2, 1, 2, 2, 2, 1, 2, 1, 3, 2, 1, 0, 0, 0, -1, -1, -2, -1, -1, -2, -2, -2, -3, -4, -1, 0, 3, 4, 4, 2, 1, 2, 2, 1, 1, 2, 2, 2, 1, 1, 2, 2, 1, 0, 0, 0, 0, -1, -1, -1, -1, -2, -2, -2, -4, -4, -2, 0, 3, 3, 3, 1, 1, 1, 1, 1, 0, 3, 3, 2, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -3, -2, -3, -4, -2, 0, 3, 2, 1, 0, 0, 1, 1, 1, 1, 2, 3, 2, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, -1, -1, -2, -1, -2, -1, -3, -2, -2, 0, 2, 3, 1, -2, -3, 0, 0, 0, 2, 2, 1, 1, 1, 0, 0, 1, 1, 0, 0, 1, 0, -1, -1, -2, -2, -1, -1, -1, -3, -3, -1, 0, 1, 1, 0, -3, -4, 0, 1, 0, 0, 0, 2, 2, 0, 1, 1, 1, 0, 0, 0, 1, 0, -1, -4, -4, -3, -2, -1, -1, -2, -2, 0, 1, 1, 1, 0, -4, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 0, -3, -3, -5, -3, -3, -1, -1, -2, -2, 0, 0, 1, 2, 0, -2, -1, -1, 0, 0, -2, 0, 0, 1, 1, 1, 1, 1, 0, 2, 2, 1, 0, -2, -4, -4, -3, -3, -1, -2, -2, -2, 0, 1, 3, 3, 0, 0, -1, -2, 0, -2, -1, 0, 0, 0, 2, 0, 1, 1, 1, 1, 2, 4, 1, 0, -2, -3, -4, -2, -3, -2, -1, -2, 0, 1, 3, 2, 2, 0, -1, -1, 0, -1, -1, 0, 0, 2, 2, 2, 1, 1, 1, 2, 4, 3, 3, 0, -1, -4, -4, -3, -3, -1, -1, -1, 1, 2, 4, 3, 3, 0, 0, 0, 0, -1, 0, 0, 1, 1, 2, 1, 1, 1, 0, 1, 4, 4, 3, 0, -1, -3, -4, -3, -1, -2, 0, -1, 0, 1, 3, 4, 2, 1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 1, 1, 3, 3, 3, 2, 1, -2, -3, -3, -2, -1, 0, 0, -1, 0, 1, 3, 4, 2, 0, -1, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 1, 3, 2, 3, 2, 1, -1, -3, -3, -3, -3, 0, -1, 0, 0, 0, 1, 2, 3, 2, 0, 0, -1, 0, 0, 0, 1, 1, 2, 2, 1, 1, 2, 2, 1, 2, 0, 0, -1, -2, -3, -2, -3, -2, 0, -1, 0, 0, 0, 2, 3, 2, 0, -1, -2, -1, -1, 0, 0, 1, 3, 2, 1, 1, 1, 1, 1, 3, 0, -1, -1, -2, -3, -1, -1, 0, -1, -2, -1, 0, 0, 2, 3, 1, -2, -2, -2, -1, 0, 0, 2, 2, 2, 1, 0, 0, 0, 2, 3, 1, 0, -1, -2, -2, -1, -1, -2, -2, -2, -2, -1, 0, 1, 2, 2, 1, -1, -1, -2, 0, 0, 2, 3, 3, 3, 0, 0, 0, 0, 2, 4, 3, 0, 0, 0, -1, -1, 0, -1, -2, -1, -3, -3, -1, 1, 1, 3, 2, 0, 0, 0, 0, 1, 2, 3, 3, 2, 0, 0, -1, 0, 2, 4, 1, 0, 0, -2, -3, -3, -2, -1, -2, -3, -4, -3, -2, 1, 1, 3, 2, 0, 0, 0, 0, 1, 2, 3, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, -1, -3, -4, -3, -2, -3, -1, -3, -3, -4, -2, 1, 2, 3, 3, 1, 1, 0, 2, 2, 1, 1, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, -2, -3, -3, -5, -3, -3, -3, -4, -5, -5, -3, 1, 2, 3, 3, 2, 1, 2, 2, 1, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -2, -3, -4, -2, -3, -3, -3, -4, -4, -2, 1, 1, 4, 4, 2, 2, 1, 1, 2, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -2, -3, -3, -2, -1, -1, -3, -4, -3, -1, 2, 3, 3, 4, 4, 1, 1, 0, 2, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, -4, -3, -4, -3, -2, -1, -1, -2, -2, 0, 1, 2, 5, 5, 4, 2, 2, 0, 1, 2, 0, 0, 0, -2, -2, -1, -2, -2, -1, -2, -3, -3, -4, -5, -5, -3, -2, -1, -1, -2, -1, 1, 1, 2, 4, 4, 4, 4, 3, 3, 1, 0, 0, -1, -1, 0, -1, -1, -3, -2, -3, -3, -4, -4, -6, -5, -4, -5, -3, -2, -1, -2, -2, 0, 1, 3, 5, 6, 5, 5, 4, 3, 2, 2, 0, 0, -1, -1, -1, -1, -2, -4, -4, -5, -5, -4, -5, -5, -3, -4, -4, -2, -1, -2, 0, 1, 3, 2, 5, 4, 4, 4, 5, 3, 1, 0, 0, 0, -1, -1, -1, 0, -3, -2, -3, -4, -4, -6, -5, -4, -3, -3, -3, -2, -1, -1, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, -1, -2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 1, 1, 2, 1, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -2, 0, 0, 0, -1, 0, 0, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 2, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 1, 1, 0, 2, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 1, 1, 1, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 2, 3, 1, 1, 0, 1, 0, 1, 0, 0, -1, -1, 0, -1, -1, 0, 0, 1, 1, 0, 2, 2, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 2, 1, 0, 1, 0, 0, 0, -1, 0, -2, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, -2, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -2, 0, 0, -1, 0, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 2, 0, 0, 1, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 2, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 2, 3, 3, 2, 2, 3, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 0, 2, 3, 2, 4, 5, 4, 4, 3, 4, 5, 2, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, -1, -1, -3, -2, -2, 0, 0, 1, 0, 0, 0, 1, 2, 2, 4, 4, 6, 5, 3, 5, 5, 2, 0, 0, -2, -1, -2, -1, -1, 0, 0, 0, 0, -1, -1, -3, 0, -1, -1, 0, 1, 0, -1, 0, 0, 2, 2, 4, 5, 3, 1, 3, 4, 1, 0, 0, -3, -2, 0, -1, -1, -1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 4, 1, 0, 0, -2, -3, -1, 0, -1, 0, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, 0, 1, 0, 0, 0, 3, 1, 0, -1, -2, -2, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -3, -2, -3, -1, -1, 0, 0, 1, 1, 0, 0, -3, -2, 0, 0, 0, 0, 0, -1, 0, 0, -2, -1, 0, -1, -1, 0, 0, -2, -1, -1, -3, -4, -3, -4, -3, -2, -2, 0, 1, 1, 0, -1, -2, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, -3, -3, -4, -5, -3, -4, -3, -2, 1, 1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -4, -4, -5, -3, -2, 0, 1, 1, -1, 0, -2, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -2, -3, -3, -2, -2, 0, 1, 0, -1, -1, -1, 0, 2, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 1, 0, 0, -1, -2, -4, -2, -1, -3, -3, -4, -1, 0, 2, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 2, 0, 0, 0, -4, -4, -3, -1, -2, -2, -3, -2, 0, 2, 1, 0, 0, -2, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, -2, -1, 0, 2, 1, 1, 0, -2, -4, -5, -2, -1, -1, -2, -3, -3, 0, 2, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 2, 1, 0, -1, -3, -4, -2, -1, -1, -3, -2, -4, -1, 0, 0, 0, 0, -2, 0, 1, 1, 0, 1, 1, 0, 0, -1, -1, -1, 0, 0, 1, 1, 2, 0, 0, -3, -2, -2, 0, -1, -1, -3, -2, -2, 1, 0, 0, 0, -1, 0, 0, 1, 3, 2, 0, 0, 0, -1, 0, -1, 0, 1, 2, 2, 2, 2, 0, -2, -2, 0, 0, -1, -1, -2, -4, 0, 1, 0, 0, 0, -2, -1, 0, 2, 2, 3, 0, 0, 0, 0, 0, -1, 0, 1, 1, 3, 2, 1, 1, -2, 0, 0, -1, 0, 0, -2, -2, -1, 0, 0, 0, 0, -2, -1, 0, 2, 3, 1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, -1, -1, 0, 1, 1, -1, 0, -2, -2, 1, 2, 3, 1, 0, -1, -2, 0, 0, 0, 1, 2, 0, 1, 0, -1, -2, -2, -1, -2, -1, 0, 0, -1, -1, 0, 1, 0, -1, 0, -1, -1, 0, 1, 2, 1, 1, 0, -2, -1, -1, 1, 1, 1, 1, 1, 0, 0, -2, -2, -1, -2, -1, -2, -1, -2, -2, 0, 1, 0, -1, 0, -2, 0, 1, 0, 1, 1, 1, 0, -1, -2, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -2, -2, -2, -2, -2, -2, -2, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, -1, -1, -2, -1, -2, -2, -3, -2, 0, 0, 1, 0, -1, -1, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -2, -2, -2, -2, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, 2, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, -1, -1, -1, -1, -3, -1, -3, -3, -2, -1, 0, 1, 1, 0, 0, -1, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 2, -1, -3, -3, -4, -3, -3, -2, -2, -2, -2, -1, 1, 1, 0, -1, 0, -1, -1, -1, -1, -1, 1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 2, 0, -2, -4, -4, -3, -2, -3, -2, -3, -3, -1, 1, 2, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, -1, -4, -4, -4, -2, -2, -2, -1, -3, -1, 1, 1, 0, 0, 0, -2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 1, 0, 0, 0, -2, -3, -3, -2, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 3, 2, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, -2, 0, 0, 0, 1, -1, 0, 1, 1, 2, 2, 2, 3, 3, 3, 4, 4, 4, 5, 4, 3, 4, 1, -1, 0, -1, -2, -1, 0, -1, 0, 0, -1, -2, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 1, 2, 1, 2, 2, 3, 4, 3, 3, 3, 0, 0, -2, 0, -1, 0, -1, 0, 0, 0, 2, 0, 0, 0, 2, 2, 1, 2, 1, 2, 0, 2, 1, 1, 1, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, -1, 0, 1, 0, 0, 0, 2, 3, 1, 0, 0, -1, 0, 1, 0, 0, 0, -1, -1, -2, -1, -2, 0, 0, -1, 0, -3, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 1, 3, 2, 1, 0, 0, 0, -1, -3, -4, -2, 1, -2, -1, -5, -1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -2, -1, 0, 0, 2, 5, 3, 1, 0, 1, 1, 0, -3, -3, -1, 0, -2, 0, -5, 0, -1, -1, -1, 0, 0, 1, 0, 1, -1, -1, -1, 0, -2, -1, -1, -1, 1, 1, 0, 0, 0, 0, 2, 2, 0, 0, 0, 1, -1, -1, -5, -2, 0, -1, -1, -1, -1, 0, -1, 0, -1, -1, -1, -1, -1, -1, -1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 3, -1, 0, -5, -1, 0, 0, -1, -1, -2, 0, -1, 0, 0, -2, -1, -2, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 1, 1, 2, 1, 1, 0, -1, -4, -2, 0, -1, 0, -1, -2, 0, -1, -1, -1, 0, -2, -3, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, -3, -2, -1, 0, -1, 0, -2, -1, -1, -1, -1, 0, -2, -3, -2, -1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, -3, 0, 0, -2, -1, 0, 0, 0, -2, -3, -1, -1, 0, 0, -1, 0, 0, 1, 4, 2, 1, 0, 0, -1, 0, 0, 3, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, 0, 0, 0, -2, -2, -1, 0, 0, 0, -1, 0, -1, 0, 2, 3, 3, 2, 3, 1, -1, 0, 2, 0, 0, -1, 0, 0, -3, 0, 0, -3, -2, -1, -1, 0, -1, -2, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 1, 2, 2, 1, 0, 0, 2, 2, 0, -1, 0, 0, -2, 0, 0, -1, -2, 0, 0, 0, -2, -2, 0, 1, 1, 0, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 2, 0, -1, -1, 0, -3, 0, 0, -1, -2, 0, 0, 0, -2, -1, 0, 3, 2, 1, 1, 0, 1, 2, 1, 0, -1, -1, -1, -1, -2, 0, 0, 1, 1, 0, 0, 0, -2, 0, 0, -1, -3, -1, -1, -1, -2, -2, -1, 2, 0, 0, 0, 1, 0, 1, 2, 0, -1, 0, -1, -1, 0, 0, -1, 0, 1, 0, 0, 0, -2, 0, 0, -1, -3, -1, 0, -1, -1, -1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, -1, -1, -1, -2, -1, 0, 0, 0, 1, -3, 0, 0, -2, -3, -3, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 0, -3, -3, -3, -2, -1, 0, 0, 0, -3, 0, 0, 0, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 3, 3, 1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, -2, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 3, 4, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -3, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 1, -1, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 1, 1, 0, 0, 1, 2, 0, 0, -1, 1, 0, 0, 1, 1, 1, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 1, 0, -2, 0, 0, 2, 0, -1, -1, -2, -2, -2, -1, 0, 0, 0, 0, 0, 1, 2, 3, 2, 1, -1, 0, 0, 0, 1, 3, 1, 0, 0, 1, 0, -2, 0, 0, 1, 0, 0, 0, -2, -2, -1, -2, 0, 2, 0, 0, 1, 0, 3, 4, 4, 2, -1, 1, 1, 0, 1, 2, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 2, 2, 0, -1, 0, 0, 2, 3, 3, 2, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 2, 2, 1, 0, -1, 0, 0, 0, 0, 2, 3, 0, 0, 0, 0, 1, 2, 3, 3, 0, -1, 1, 0, 0, 0, 0, 0, -4, 0, -1, -1, 0, 1, 1, 1, -1, 0, -1, -1, 0, 0, 3, 2, 0, 0, -1, 0, 2, 3, 3, 2, 0, -2, 0, 0, 0, 0, 0, -1, -3, -1, 0, -1, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 1, 1, 1, -1, -1, 0, 0, 1, 3, 0, -3, -2, -1, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, 0, 3, 2, 1, 2, 1, 0, 0, 2, 2, 2, 1, 0, 0, 0, 0, 1, -1, -3, -3, -2, -3, -2, -1, -1, -1, -5, -1, -1, 0, 2, 1, 2, 1, 2, 1, 2, 1, -1, 0, 2, 3, 3, 1, 2, 0, 1, 2, 1, 0, -1, -1, -2, -2, -2, 0, 0, -1, -5, -2, 0, -1, 0, 1, 1, 0, 1, 2, 1, 0, 0, 0, 1, 4, 2, 2, 4, 3, 4, 2, 2, 1, 0, -1, -1, -4, -2, -1, -2, 0, -3, -4, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 3, 4, 3, 5, 4, 2, 1, 0, 1, 0, -1, -2, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -2, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, -1, -1, -2, 0, 0, 0, -1, -1, 0, 0, -2, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -2, -1, -1, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 2, 2, 0, 1, 1, 1, 2, 1, 1, 0, 2, 3, 1, 1, 1, 1, 1, 1, 2, 0, 0, 2, 1, 0, 0, 2, 0, 0, 2, 2, 1, 1, 3, 3, 0, 0, 2, 2, 1, 0, 1, 0, 2, 5, 3, 1, 2, 2, 2, 2, 3, 1, 1, 4, 2, 0, 0, 3, 0, 0, 3, 2, 3, 3, 3, 2, 1, 0, 2, 2, 0, 0, -1, 0, 2, 4, 3, 2, 3, 0, 3, 2, 1, 1, 2, 5, 4, 0, 0, 3, 0, 0, 3, 2, 2, 3, 2, 4, 2, 2, 1, 3, 0, 0, -1, 0, 3, 3, 2, 4, 2, 0, 3, 4, 1, 1, 1, 5, 4, 2, -1, 1, 0, 0, 4, 1, 2, 3, 2, 4, 3, 0, 0, 2, 0, 0, 0, 1, 4, 2, 2, 6, 2, 0, 2, 3, 1, 2, 1, 4, 3, 0, -2, 0, 0, 0, 1, 0, 1, 4, 4, 6, 3, 0, 0, 0, 1, -1, 0, 1, 4, 2, 2, 5, 2, 0, 3, 3, 1, 4, 1, 2, 5, 1, -2, -2, 0, 1, 1, -3, 0, 3, 3, 5, 2, 2, 1, 1, 2, -1, -1, 0, 1, 0, 2, 4, 1, 1, 2, 1, 1, 3, 2, 3, 5, 2, -2, -1, 0, 0, 2, -3, 0, 1, 3, 4, 2, 1, 1, 0, 0, -1, -1, 0, 0, -2, 0, 3, 0, 2, 2, 0, 2, 5, 3, 2, 5, 2, 0, -1, 0, 1, 2, 0, 0, 1, 1, 4, 1, 0, 0, 1, 1, -1, -1, -1, -1, -2, -1, 2, 1, 2, 3, 0, 2, 5, 1, 3, 5, 3, 0, -1, 0, 0, 4, 2, 0, 0, 0, 1, 3, 0, -1, 0, -1, -2, -3, -1, 0, -3, -2, 1, 0, 2, 1, 0, 1, 5, 2, 3, 5, 4, 1, 0, 0, 0, 3, 2, 1, 0, 0, 0, 4, 1, 0, -1, -1, -3, -2, -1, 0, -2, -2, 1, 2, 2, 1, -1, 1, 3, 1, 3, 4, 4, 0, 3, 0, 0, 2, 1, 2, 1, 0, 0, 2, 0, 0, -1, -2, -3, -2, -4, -1, 0, 0, 0, 1, 4, 1, 0, 0, 4, 3, 2, 3, 3, 0, 4, 0, 0, 2, 2, 6, 3, 0, -1, 2, 0, 0, 0, -1, -3, -3, -3, -3, -1, 0, -1, 0, 2, 3, 0, 0, 2, 2, 0, 1, 4, 0, 4, 0, 0, 2, 2, 6, 4, -1, 0, 2, 0, 0, -2, -2, -3, -4, -3, -2, -2, 0, -3, 0, 3, 2, 0, 0, 2, 1, 0, 1, 1, -2, 4, 0, 0, 2, 3, 6, 4, 1, 1, 1, 0, 1, -3, -1, -1, -3, -3, -2, -3, -2, -3, -1, 1, 1, 0, 1, 1, 0, 0, 0, 1, -1, 2, 0, 0, 4, 2, 3, 4, 1, 2, 0, 0, 0, -4, -2, -3, -4, -4, -1, -2, -4, -4, 0, 1, 1, 0, 0, 0, 0, 0, 2, 1, -1, 3, 0, 0, 4, 0, 3, 4, 3, 2, 0, 0, -1, -4, -3, -3, -5, -4, -2, -1, -3, -3, -2, 0, 0, 1, 1, 0, 0, 0, 1, 2, -1, 2, 0, 0, 3, 0, 2, 2, 2, 4, 0, -2, -2, -4, -2, -3, -5, -5, -2, 0, 0, -2, -2, 0, 0, 1, 2, 1, 0, -1, 1, 2, -2, 1, 0, 0, 3, 0, 3, 2, 1, 3, 0, -1, -1, -4, -3, -3, -3, -2, -1, 0, 0, 0, -3, 0, 1, 1, 3, 1, 0, -1, 1, 2, -1, 1, -1, 0, 4, 1, 4, 3, 2, 2, 0, 0, 0, 0, -1, -1, -3, -2, -1, -1, 2, -1, -1, 0, 2, 2, 2, 2, 0, 0, 0, 0, -1, 0, 0, 1, 3, 0, 3, 3, 2, 1, 0, 0, 2, 1, 0, -1, -3, -3, -3, -1, 2, 0, -1, 2, 4, 2, 5, 5, 1, 2, 1, 1, 0, -1, 0, 0, 4, 1, 2, 3, 2, 0, 0, -1, 0, 1, 0, 0, -3, -4, -3, -1, 1, 0, -1, 4, 4, 3, 3, 3, 0, 2, 3, 0, 0, -2, 0, 1, 3, 0, 4, 2, 0, 1, 0, -2, 0, 0, 0, -1, 0, -2, -1, 0, 2, 0, 0, 2, 4, 3, 3, 2, 0, 3, 4, 1, 0, -2, 0, 0, 0, 0, 3, 2, 0, 1, 1, 0, -1, -1, -2, -1, 0, 1, 0, 0, 3, 0, 1, 3, 4, 3, 3, 0, 0, 5, 5, 2, -1, -2, 0, 0, -2, -2, 2, 1, 0, 0, 2, 0, 0, -1, -2, -2, 0, 3, 1, 2, 2, 0, 1, 4, 5, 4, 3, 1, 0, 4, 6, 3, -1, 0, 0, 0, -2, -1, 3, 1, -2, 1, 3, 4, 2, -1, -1, -1, 0, 2, 1, 1, 1, 1, 0, 2, 2, 2, 2, 1, 0, 2, 5, 1, -2, 0, 0, 0, 0, -1, 3, 0, -3, 0, 4, 3, 1, -2, 0, 0, 2, 2, 1, 3, 2, 0, 1, 2, 0, 0, 1, 2, 2, 3, 4, 1, -1, 0, 0, 0, 0, 0, 4, 3, 0, 0, 3, 2, 3, -1, -1, 0, 2, 1, 1, 5, 3, 0, 2, 2, 0, -1, 0, 0, 0, 3, 3, 1, -2, 1, 0, 0, 1, 0, 2, 2, 0, 0, 2, 1, 2, 0, 0, 0, 1, 2, 1, 4, 2, 1, 2, 2, 1, 0, 0, 0, 1, 1, 3, 0, -2, 1, 0, 0, 2, 0, 0, 2, 1, 0, 0, 0, 3, 2, 0, 0, 2, 1, 2, 4, 1, 2, 3, 1, 3, 2, 0, 1, 0, 0, 3, 1, -3, 1, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 1, 2, 2, 4, 4, 3, 4, 3, 3, 2, 2, 0, 0, 1, 0, 1, 1, -2, 2, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 1, 2, 1, 3, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 1, 3, 2, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -1, -3, -3, -3, -3, -2, -3, -1, -1, -2, 0, 0, 0, 1, 1, 1, 3, 4, 4, 2, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -2, -1, -1, -2, -3, -2, -4, -3, -3, -3, -2, 0, 0, 0, -1, 1, 0, 3, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -2, -3, -3, -2, -1, -1, -2, 0, -1, -2, 0, 0, 2, 3, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -2, -2, -1, -2, -1, -1, -1, -1, 1, 0, 2, 1, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, -1, -2, -1, 0, -2, -1, -1, -1, -2, 0, 0, 1, 2, 1, 1, 2, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -2, -1, -2, -2, -1, -2, 0, 0, 2, 2, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -2, -1, -1, -2, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, -1, -1, -2, -2, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, -2, -2, -1, -2, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, -2, -2, 0, -1, -1, 0, -2, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, -3, -2, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 0, -2, -2, -2, 0, -1, 0, 0, -1, -1, 1, 0, 1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 2, 1, 0, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 2, 1, 2, 1, 0, -1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 3, 2, 2, 2, 1, -1, 0, -2, 0, 0, 0, 0, 0, 1, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 2, 3, 2, 2, 3, 2, 1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 2, 0, 1, 2, 2, 1, 3, 2, 2, 1, -1, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 1, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 2, 3, 2, 1, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 1, 0, 1, 0, -1, -2, -1, -1, 0, 0, 2, 1, 1, 1, 0, 0, 1, 2, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 1, 0, 2, 1, 0, 0, 0, -1, 0, 0, 1, 2, 2, 1, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -1, 0, -1, 0, -2, -1, -2, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -2, -1, -2, -3, -2, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, -1, 0, -1, -2, -2, 0, 0, 1, 2, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, -1, -1, -3, -2, 0, 0, -1, -1, -1, 0, 0, 0, 2, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -2, -1, -1, -1, 0, -1, -1, 0, 0, 0, 2, 2, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, -2, -3, -2, -1, -1, 0, 0, 0, 0, 0, 0, 2, 3, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -2, -3, -3, -3, -3, -2, -1, 0, -1, -1, 0, 0, 2, 0, 3, 2, 3, 2, 2, 1, 1, 0, -1, -1, 0, -1, -1, -1, -1, -1, -2, -1, -2, -4, -4, -2, -2, -1, -2, -1, 0, -1, -1, 0, 1, 0, 3, 2, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, -2, -1, -2, -2, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 3, 1, 0, 1, 0, 0, -1, -2, 0, -1, -1, 0, 0, -2, -3, -1, -3, -3, -3, -4, -3, -3, -3, -2, -1, -1, -1, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -2, -2, 0, 0, 0, -1, -1, -3, -3, -3, -2, -2, -3, -2, 0, -1, -1, 0, 1, 1, 1, 1, 1, -1, 0, -1, -1, -1, -2, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -2, -3, -1, -2, -1, 0, -1, -1, -1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, -2, -2, -1, 0, -1, -1, 0, -1, 0, 0, 1, 2, 1, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 2, 1, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 2, 2, 0, 1, 2, 1, 1, 1, 1, 0, 1, 0, 0, 1, 3, 3, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 2, 1, 1, 0, 1, 1, 1, 2, 1, 0, 2, 1, 0, 0, 0, 4, 2, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 1, 2, 0, -1, 0, 1, 1, 1, 2, 1, 2, 1, 1, 0, 0, 3, 2, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 1, 1, 2, 2, 1, 1, 2, 3, 2, 2, 0, 1, 1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, -2, -2, -1, -1, 1, 1, 2, 1, 2, 2, 0, 2, 4, 3, 1, 2, 2, 1, 0, -1, 0, 0, 1, 0, 1, 2, 0, 0, 0, 0, 2, -1, 0, -2, -1, 0, 0, 1, 0, 0, 1, 2, 0, 2, 4, 3, 1, 2, 1, 2, 0, -1, -1, 0, 0, 1, 0, 1, 0, -1, 1, 2, 1, 0, -1, -1, -1, -2, 0, 0, 1, 2, 0, 1, 0, 2, 3, 3, 3, 2, 1, 2, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 1, 1, 1, 1, 2, 3, 2, 3, 3, 2, 1, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, -1, 0, 0, 1, 2, 2, 1, 2, 2, 3, 2, 3, 4, 3, 3, 2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, -1, -1, 1, 1, 0, 0, 0, 2, 3, 3, 3, 2, 2, 3, 2, 4, 2, 3, 3, 0, 0, -2, -1, -1, 0, 0, 0, 0, 1, 2, 1, 0, -1, -1, 0, 0, 0, 0, 1, 2, 2, 3, 2, 3, 2, 2, 3, 3, 2, 3, 2, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 2, 0, -1, 0, 0, 0, 1, 0, 0, 1, 2, 1, 1, 2, 3, 4, 3, 4, 1, 2, 2, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 2, 2, 2, 1, 3, 2, 3, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 2, 1, -1, 0, 0, 2, 0, -1, 0, 0, 0, 0, 0, 0, 1, 3, 2, 1, 2, 1, 1, 2, 3, 2, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 2, 3, 3, 2, 2, 1, 2, 3, 4, 1, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 1, 1, 0, 1, 3, 2, 3, 1, 2, 1, 3, 3, 4, 1, 0, 1, 0, 0, 2, 2, 2, 1, 0, -1, 0, 0, 2, 2, 0, 0, -1, 0, 1, 2, 2, 2, 3, 2, 2, 2, 0, 0, 1, 3, 3, 2, 0, 0, 1, 1, 0, 2, 2, 0, 1, 0, 0, 0, 2, 2, 0, 0, -1, 0, 0, 1, 0, 1, 1, 2, 2, 2, 0, 0, 1, 2, 2, 1, -1, 0, 0, 0, 0, 2, 2, 1, 2, 0, -2, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 1, 1, 1, 0, 0, -1, -1, 1, 1, 0, 0, -1, -1, 0, 1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 2, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 2, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 2, 3, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, 1, -1, -2, -1, 2, 2, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -1, -2, -1, -1, -2, -1, -1, -2, -1, -2, -1, 0, 0, -1, -1, 0, 1, 2, 1, 0, 1, 1, 0, -1, -1, 0, 0, -1, 0, -1, 0, -2, -1, -2, -3, -3, -3, -1, -1, -2, -1, -1, -1, -1, 0, -1, -1, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, -1, -1, -2, -2, -3, -3, -2, -3, -3, -3, -2, -3, -2, -2, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 2, 4, 2, 3, 2, 1, 0, 0, 0, 0, 0, 0, -1, -1, -2, -2, -2, -2, -2, -3, -2, -2, -3, -2, -1, 0, 1, 2, 2, 1, 1, 2, 2, 5, 4, 3, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, -1, -1, -1, -3, -4, -4, -4, -4, -2, -1, 0, 0, 0, 1, 2, 2, 1, 4, 4, 3, 2, 1, 1, 1, 2, 1, 1, 2, 1, 2, 2, 0, 1, 0, -1, -2, -2, -5, -5, -4, -2, -2, 0, 0, 0, 1, 0, 2, 1, 4, 3, 1, 0, 0, 0, 1, 0, 1, 0, 3, 1, 2, 1, 1, 0, -1, 0, 0, -3, -4, -4, -4, -3, -1, -2, -2, 0, 0, 0, 0, 2, 3, 3, 2, 2, 0, 0, 0, 1, 0, 1, 1, 2, 2, 2, 1, 0, 0, -1, 0, -2, -4, -3, -3, -4, -4, -4, -2, -2, -1, 0, 1, 0, 3, 3, 3, 0, 1, 0, 0, 1, 0, 1, 2, 1, 0, 1, 0, 1, -1, 0, -1, -3, -4, -3, -4, -5, -4, -4, -3, -3, -2, -1, 0, 1, 3, 3, 2, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -3, -4, -4, -3, -3, -3, -5, -4, -2, -3, -2, 0, 1, 4, 2, 0, 0, 0, 0, 0, 1, 3, 2, 2, 0, 0, 0, 1, 0, -1, -2, -1, -4, -5, -3, -4, -5, -3, -5, -5, -4, -2, -1, 0, 0, 3, 2, 0, 0, 0, 1, 0, 1, 1, 1, 2, 2, 1, 1, 2, 0, 0, 0, -1, -3, -4, -3, -3, -3, -3, -4, -4, -4, -1, -1, 0, 1, 3, 0, -1, -1, 0, 0, 1, 0, 1, 2, 3, 3, 3, 2, 3, 3, 0, 0, -1, -3, -3, -4, -3, -3, -4, -4, -5, -3, -1, -1, 0, 1, 2, 0, -1, -1, -1, -1, -1, 0, 1, 2, 0, 2, 3, 3, 2, 3, 2, 1, 0, -1, -4, -5, -5, -3, -4, -5, -5, -4, -2, -1, 1, 1, 2, 1, 0, 0, -1, -1, -1, -1, 0, 1, 1, 2, 3, 3, 5, 5, 4, 2, 0, -2, -4, -5, -5, -4, -4, -3, -5, -4, -2, -1, 0, 1, 4, 2, 0, 0, -1, -1, 0, 0, 1, 2, 3, 2, 4, 4, 5, 5, 5, 4, 2, 0, -2, -3, -5, -5, -2, -3, -5, -4, -3, -2, 1, 1, 3, 1, -1, -1, -2, -1, -1, 0, 0, 3, 2, 3, 4, 5, 6, 5, 5, 4, 3, 1, -1, -3, -4, -5, -4, -3, -4, -3, -3, -1, 1, 2, 3, 2, -1, 0, -1, 0, 0, 0, 2, 3, 3, 3, 5, 5, 7, 7, 5, 5, 3, 0, 0, -2, -4, -4, -2, -3, -4, -3, -3, -1, 1, 1, 2, 1, -1, -2, 0, 0, 0, 0, 2, 2, 3, 4, 5, 6, 7, 7, 7, 6, 4, 1, -1, -4, -4, -4, -2, -3, -3, -1, -2, 0, 0, 0, 2, 1, -1, -2, -2, -1, -1, 0, 0, 0, 3, 3, 4, 6, 6, 8, 6, 4, 1, 0, -3, -3, -5, -4, -1, -3, -2, -1, -1, -1, 1, 1, 3, 1, -1, -2, -3, -2, -1, 0, 0, 0, 2, 3, 4, 5, 6, 5, 4, 3, 1, -1, -2, -3, -5, -4, -2, -2, -3, -2, -2, 0, 1, 1, 1, 0, -2, -4, -3, -3, -2, 0, 0, 1, 2, 4, 4, 4, 5, 5, 4, 3, 1, -2, -3, -4, -5, -4, -4, -2, -4, -4, -1, -1, 0, 1, 2, 0, -1, -3, -3, -1, 0, 0, 1, 0, 2, 2, 3, 3, 3, 5, 5, 4, 0, -1, -2, -3, -4, -5, -3, -4, -5, -4, -3, -2, 1, 1, 3, 0, -2, -1, -2, -2, 0, 2, 3, 3, 3, 1, 3, 3, 3, 5, 3, 3, 1, -1, -3, -5, -4, -3, -5, -3, -5, -4, -3, -1, 0, 2, 3, 1, 0, -1, -1, -1, 0, 3, 2, 4, 3, 3, 3, 3, 3, 4, 3, 2, -1, -3, -3, -4, -5, -4, -4, -3, -4, -4, -3, -2, 0, 2, 3, 3, 1, 0, 0, 0, 1, 1, 2, 3, 2, 2, 2, 2, 1, 2, 2, 0, -2, -4, -5, -6, -5, -5, -4, -3, -4, -4, -3, 0, 0, 0, 3, 3, 0, 1, 1, 1, 1, 2, 1, 3, 3, 3, 3, 1, 1, 1, 0, 0, -1, -5, -5, -6, -6, -4, -4, -3, -5, -5, -4, -1, 1, 1, 3, 3, 2, 1, 0, 2, 1, 3, 3, 3, 1, 2, 1, 2, 0, 1, 0, 0, -2, -2, -6, -6, -6, -5, -5, -3, -5, -5, -3, 0, 0, 1, 3, 3, 1, 2, 0, 1, 0, 2, 3, 3, 0, 2, 2, 1, 0, 0, -1, 0, -2, -3, -5, -5, -6, -4, -4, -3, -3, -2, -1, 0, 0, 2, 4, 4, 2, 1, 2, 1, 0, 1, 1, 1, 2, 2, 1, 1, 0, 0, 0, -1, -1, -4, -4, -5, -4, -4, -2, -2, -1, -1, -1, 0, 1, 1, 4, 4, 2, 2, 3, 2, 2, 2, 1, 2, 2, 1, 0, 0, 0, 0, 0, -2, -2, -3, -4, -5, -5, -3, -3, -2, -1, 0, 0, 0, 2, 2, 5, 5, 4, 3, 3, 3, 3, 1, 1, 2, 1, 0, 0, 0, -1, -2, -2, -1, -2, -4, -3, -4, -3, -2, -3, -1, 0, 0, 1, 1, 3, 2, 4, 6, 3, 3, 3, 3, 2, 2, 0, 1, 0, 0, 0, 0, -3, -4, -2, -3, -3, -3, -3, -3, -3, -1, -2, -1, 0, 0, 1, 0, 3, 1, 3, 5, 4, 3, 4, 4, 2, 2, 0, 1, 1, 0, 0, 0, -2, -1, -1, -2, -3, -2, -4, -2, -2, -1, -2, 0, 0, 0, 1, 0, 2, 0, 0, 1, 2, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 2, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 2, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 1, 2, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 1, 0, 2, 1, 1, 0, 0, 1, 0, 0, 0, -1, 2, 0, 2, 0, 0, -1, 0, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, -1, -1, 2, 0, 1, -1, 0, 0, 0, 0, 2, 2, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 2, 0, 0, -1, 0, 1, 0, 1, 1, 1, 0, 1, 1, 1, 0, 0, 1, 0, 1, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, -1, 0, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 2, 1, 1, -2, -1, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, -2, -1, 0, 0, 2, 1, 2, 1, 0, 0, -1, 0, 1, -1, -1, -1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -3, 0, 0, 2, 1, 3, 1, 1, 0, -1, -2, 0, 0, -1, -2, -1, 0, 1, 2, 2, 0, 0, 1, 0, -1, 0, 1, 0, 0, 0, 0, 0, -2, 0, 0, 2, 2, 2, 1, 0, 1, 0, 0, 0, 0, -1, -1, -1, 1, 0, 0, 1, 0, 1, 2, 0, -1, 0, 0, 0, 0, 1, 0, 0, -3, 0, 1, 2, 2, 1, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 1, -1, 0, 3, 1, 0, 0, 1, 0, 1, 1, 0, 0, -2, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 1, 0, 0, 0, 2, 1, 0, 0, 2, 1, 1, 2, 0, 0, -1, 1, 2, 1, 1, 1, 1, 1, 1, 0, 0, 1, 1, -1, -2, 0, 0, 0, 0, 0, -1, -2, 1, 0, 0, 0, 1, 0, 1, 3, 0, 0, 0, 0, 2, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 0, 0, 3, 0, 1, 0, 1, 2, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, 0, -1, -3, 0, 0, -2, 0, 0, 1, -1, 0, 1, 0, 1, -1, 0, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 1, -1, 0, 0, 1, 0, -1, 1, 0, 1, 0, 0, 2, 2, 2, 2, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -2, -1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 2, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 3, 1, 2, 1, 3, 0, 0, 0, 1, -1, 0, 0, -1, 0, -1, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, 2, 0, 0, -1, 0, 2, 2, 3, 1, 2, 1, 1, 1, 0, 0, 1, 0, -1, 0, -1, -3, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, -2, 0, 2, 1, 1, 1, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -3, -1, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, 0, -2, 0, 1, 2, 0, 1, 2, 1, 1, 1, -1, 0, -1, -1, 1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, -1, 1, 2, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, 1, 0, 1, 0, 1, 2, 1, -1, 1, 1, 0, -2, 1, 3, 2, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 2, 0, -1, 2, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, -1, -2, -2, -1, 0, 0, 0, 1, 1, 1, 0, 0, 2, 0, 0, 0, 0, 1, 1, 0, 0, 1, 2, 0, 0, 1, 0, 0, 0, 0, 1, 1, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, 1, 0, 1, -1, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, -1, -2, -1, 1, 0, 1, 0, 0, -1, -1, 2, 0, 2, 0, 0, 1, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, -1, 0, -2, -1, 2, 1, 0, -1, 0, 1, 1, 1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 1, 2, 0, 0, -1, -1, -1, 3, 0, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 0, 2, 0, 1, 0, 1, 1, 1, 1, 1, -1, 0, 3, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 2, 1, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 0, 1, 2, 0, 2, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 1, 1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 0, 1, 1, 2, 1, 1, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 2, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 1, 1, 1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 1, 0, 1, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 3, 2, 0, -1, -1, 1, 1, 0, 0, 0, -1, 0, 0, 0, -3, -2, -1, -1, 0, 1, 1, 1, 1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 2, 0, 0, -2, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, -2, -3, -1, 0, 1, 1, 1, 1, 0, 1, -1, -1, 0, 0, 0, -2, -1, 0, 1, 0, 0, -2, -1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 1, 2, 2, 2, 1, 0, -2, -2, -1, -2, -1, -2, -2, -2, -1, 0, 0, -3, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 0, 0, 0, -1, -1, -2, -2, -4, -3, -3, -4, -1, 0, 0, -3, -3, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 3, 1, 0, 0, 0, -1, -3, -3, -4, -4, -4, -3, -3, 0, -1, -1, -3, -4, -1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, -3, -3, -3, -5, -3, -4, -3, -3, -2, 0, 0, -2, -2, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, -2, -3, -2, -4, -5, -3, -3, -4, -1, -1, 0, -2, -3, 0, 0, 1, 2, 1, 1, -1, 0, 0, 0, 0, 0, -1, -1, 2, 2, 3, 1, 0, -1, -1, -2, -3, -3, -3, -4, -2, 0, 0, 0, -3, -1, -1, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 3, 2, 2, 0, 0, -1, -1, -2, -3, -2, -3, -2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 2, 1, 1, 0, 1, 3, 4, 2, 2, 0, -1, 0, -1, -1, -1, -2, -1, -1, 0, 1, 0, -2, -2, 0, 2, 0, 2, 1, 1, 2, 1, 3, 3, 1, 0, 0, 3, 3, 3, 4, 1, -1, -3, -2, 0, -1, -1, -2, -1, 0, 1, 0, -1, -3, -1, 0, 1, 2, 2, 3, 3, 2, 3, 2, 3, 2, 1, 3, 3, 4, 4, 4, 1, -1, -2, -3, 0, -2, -1, -2, 0, -1, 1, 0, 0, -1, 0, 0, 0, 1, 1, 2, 2, 5, 3, 4, 2, 2, 1, 1, 2, 5, 5, 3, 0, -2, -4, -2, -2, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 2, 1, 3, 5, 4, 4, 4, 2, 2, 1, 2, 4, 4, 4, 3, 0, 0, -3, -2, -1, -1, -1, -3, -3, -2, 1, 0, 1, 0, 0, 0, 1, 3, 2, 3, 5, 4, 4, 3, 3, 1, 2, 3, 3, 5, 5, 4, 1, 0, -2, -1, -1, -2, -2, -3, -2, -2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 3, 4, 3, 2, 3, 2, 2, 3, 4, 5, 6, 4, 2, 2, 0, -2, -1, -1, -1, -1, -3, -4, -1, 0, 0, 0, 0, 0, 1, 2, 3, 3, 3, 3, 3, 1, 1, 3, 4, 3, 4, 5, 5, 4, 2, 0, -1, -2, -1, -1, -2, -1, -2, -3, -3, 0, 0, 1, 0, 0, 1, 1, 2, 3, 3, 4, 2, 1, 0, 2, 4, 3, 3, 5, 4, 2, 0, 0, -2, -2, -2, -2, -2, -2, -3, -2, -2, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 4, 2, 2, 1, 1, 3, 4, 3, 3, 4, 2, 0, 0, -2, -2, -3, -4, -3, -3, -4, -3, -3, -1, 0, 0, -1, 0, 0, 0, 1, 0, 2, 2, 1, 1, 1, 2, 3, 2, 2, 2, 3, 0, 1, 0, -1, -1, -2, -4, -4, -3, -3, -4, -2, 0, 0, 0, -1, 0, 0, 0, 1, 1, 2, 2, 1, 1, -1, 0, 0, 2, 1, 3, 3, 1, 1, 1, -1, 0, -2, -4, -4, -3, -3, -3, -3, -1, 0, 1, 0, -1, 0, 0, 0, 1, 1, 2, 1, 1, 0, 0, 1, 1, 1, 3, 1, 0, 0, 0, 0, -1, -1, -4, -4, -3, -4, -2, -3, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 2, 2, 3, 0, -1, 0, 0, 0, -2, -3, -2, -3, -2, -2, -2, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 2, 0, -1, 0, 0, 1, 1, 3, 3, 3, 0, -1, -2, -1, -2, -1, -2, -3, -2, -3, -1, -1, 0, 1, 0, -1, 0, 0, 0, -1, 0, 2, 1, 0, 0, 0, 0, 2, 1, 3, 4, 3, 1, 0, 0, -1, -2, -3, -3, -4, -4, -2, -2, -2, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 1, 1, 1, 1, 4, 2, 2, 0, 0, -1, -2, -3, -3, -2, -4, -4, -3, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 0, 1, 1, 0, 1, 4, 2, 2, 1, -1, -1, -2, -3, -2, -2, -3, -3, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 1, 1, 1, 2, 3, 3, 2, 1, 0, 0, -2, -1, 0, -2, -2, -1, -1, -1, 1, 1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 3, 4, 3, 3, 2, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, 2, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 1, 1, 1, 2, 3, 2, 1, 1, 1, 1, 1, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 2, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 2, 1, 0, 1, 0, 0, 1, 1, 1, 1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 2, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 1, 1, 1, 0, 0, 1, 1, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, -2, -1, -2, -1, -2, -2, -3, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 2, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -1, -2, -2, -1, -2, -1, -1, 0, 0, 1, 1, 0, 0, 2, 0, 0, 0, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, -2, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 2, 1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, 0, -1, 0, -1, -1, -2, -1, -1, 0, 0, -1, 0, 1, 0, 0, 2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -3, -3, -3, -2, -1, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -4, -3, -2, -3, -1, -2, -2, -2, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -2, -3, -2, -2, -3, -2, -1, -3, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 0, 0, -2, -2, -2, -2, -2, -3, -2, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, -1, -2, -4, -3, -3, -2, -3, -3, -1, -2, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, -3, -3, -2, -2, -2, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, -1, -2, -3, -2, -2, -3, -3, -2, -2, -1, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, 1, 1, 0, 1, 1, 1, 1, 0, -1, -2, -3, -3, -1, -2, -3, -2, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 3, 1, 1, 1, 0, -1, -3, -2, -3, -1, -1, -1, -1, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 3, 2, 3, 1, 0, -2, -2, -2, -3, -2, -2, -2, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 2, 2, 3, 1, 0, 0, -3, -2, -2, -2, -1, -1, -1, -1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 2, 2, 1, 2, 2, 0, -1, -3, -2, -2, -2, -1, -1, -1, -2, -1, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 0, 1, 0, 2, 2, 2, 2, 0, 0, -1, -3, -2, -3, -2, -3, -2, 0, -2, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 1, 0, 0, 2, 1, 1, 1, 1, -1, -1, -1, -2, -2, -2, -2, -2, -2, -1, 0, 0, 1, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, -2, -3, -3, -2, -3, -3, -3, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -2, -2, -2, -3, -3, -2, -2, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, -1, -2, -2, -3, -4, -2, -3, -2, -4, -2, -3, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -2, -1, -2, -3, -3, -3, -3, -3, -2, -2, -2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, -1, -2, -1, -2, -3, -3, -2, -2, -3, -2, -1, 0, 0, 0, 0, 2, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -2, -2, -2, -4, -3, -3, -3, -2, -2, -2, 0, 1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, -2, -2, -1, -2, -3, -3, -2, -3, -2, -1, -1, 0, 2, 0, 0, 3, 1, 1, 2, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, -1, -2, -2, -3, -2, -3, -2, -3, -1, -1, 0, 1, 2, 0, 1, 1, 1, 2, 1, 1, 2, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, -2, -3, -3, -2, -2, -1, -2, 0, -1, 0, 1, 1, 0, 1, 1, 1, 1, 2, 2, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, -2, -1, -1, -3, -2, -2, -2, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 3, 2, 2, 0, 0, 3, 3, 1, 3, 2, 2, 3, 4, 5, 5, 5, 5, 4, 2, 0, 2, 1, -1, 0, 0, -3, -1, 0, 0, -1, -1, 1, 3, 3, 1, -1, 0, 3, 2, 3, 3, 4, 3, 5, 6, 6, 6, 5, 8, 6, 1, 1, 0, 1, -1, 0, -1, -3, 0, 0, 1, -1, 0, 0, 1, 3, 0, -2, -1, 1, 0, 0, 3, 0, 0, 3, 4, 6, 5, 6, 8, 8, 2, 0, 1, 1, -1, 0, -2, -5, -1, 0, 0, 0, 1, 1, 2, 2, 0, -3, -3, 0, -2, 0, 0, -1, -1, 0, 3, 1, 2, 4, 8, 7, 3, -1, 1, 2, -1, -1, -2, -4, -1, 0, 1, 0, 0, 0, 1, 1, -1, -3, -4, -3, -3, -1, -2, -3, -3, -2, 0, -1, 0, 0, 4, 4, 3, 0, 0, 2, -1, 0, -3, -4, 0, 2, 2, 1, 0, 0, 0, -1, -3, -4, -3, -3, -4, -1, -2, -4, -3, -2, -1, -1, -1, -1, 0, 2, 2, 2, 0, 3, 0, 0, -3, -2, 0, 3, 2, 0, 0, -1, -1, -1, -4, -5, -4, -3, -4, -1, -1, -2, -3, -2, -2, -3, -3, -2, -2, 0, 0, 0, 0, 1, 0, 0, -3, -3, 0, 4, 2, 0, 0, -1, -2, -3, -2, -4, -3, -4, -2, -2, -1, -3, -2, 0, -2, -5, -5, -6, -5, -2, -1, 0, 0, 0, -2, 0, -2, -1, 0, 2, 1, 1, 1, 0, 0, -1, -2, -1, -1, -2, -2, -1, -1, -2, -1, 0, -1, -3, -4, -5, -5, -4, -1, 0, 0, 0, -1, 0, -2, -1, 0, 2, 2, 1, 2, 1, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 2, 1, 0, -2, -5, -5, -4, -1, 0, 0, 0, -4, -1, -3, 0, 3, 2, 0, 1, 0, 1, 0, 0, 0, -1, 0, -2, 0, 0, 0, -2, -1, 0, 0, -1, 0, -2, -5, -4, -2, 0, 0, -1, -3, 0, -2, 0, 2, 2, 1, 0, 0, 0, 0, -1, -1, -2, -1, -3, -2, 0, 0, -3, -1, -2, -2, -2, 0, 0, -5, -4, -3, 0, 1, 0, -3, 0, -2, 0, 2, 3, 0, 0, 0, 1, -2, -4, -4, -3, -2, -3, 0, 0, -1, -3, -1, -4, -5, -4, -2, -2, -4, -5, -4, 0, 1, 1, -1, 0, -2, 0, 3, 2, 0, 0, 0, -1, -3, -3, -5, -4, -2, -2, 0, 0, 0, -1, -1, -4, -5, -4, -2, 0, -4, -5, -4, -2, 0, 1, -2, -1, -2, -1, 2, 2, 1, 0, 0, -2, -2, -4, -5, -5, -4, -4, -2, 0, 0, -2, -3, -5, -7, -2, 0, 0, -2, -4, -6, -5, -1, 0, -2, 0, -3, -1, 2, 4, 1, 0, -1, -2, -4, -4, -6, -6, -4, -3, -2, 0, 0, -1, -2, -5, -5, -1, 1, 0, -3, -5, -6, -6, -2, -1, -2, 0, -1, 0, 1, 3, 1, 1, -1, -3, -5, -3, -4, -4, -3, -2, -1, 0, 2, -1, 0, -2, -3, -1, 1, 1, -1, -3, -5, -6, -3, 0, -3, -1, -1, 0, 1, 3, 3, 1, 0, -3, -4, -2, -3, -3, -2, -1, 0, 0, 2, 0, -1, -1, 0, 0, 0, 1, 0, -2, -5, -4, -2, 0, -2, 0, -1, -1, 1, 2, 6, 2, 1, -3, -5, -2, -3, -1, -1, 1, 0, 2, 1, 0, 0, -1, -1, 0, 0, 2, 0, -1, -3, -3, 0, 0, -1, 0, -1, -1, 0, 3, 5, 4, 0, 0, -4, -4, -2, -1, 0, 0, 1, 2, 0, 0, -1, -2, -2, -2, -1, 1, 1, 0, -3, -2, -1, 0, -1, 0, 0, 0, 3, 4, 3, 4, 1, 0, -2, -2, -3, -2, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 1, 0, -2, -2, -2, 0, 0, 0, -2, 1, 1, 2, 2, 2, 2, 1, -1, -4, -4, -2, -2, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -4, -3, -1, 0, 0, 0, 0, 0, 1, 0, 2, 1, 1, 0, -3, -3, -3, -2, -1, 0, 2, 1, 0, 0, 0, 0, 0, 1, 0, -1, -3, -3, -2, -2, -1, 0, 1, 0, 1, 0, 0, 0, 2, 3, 2, 0, -3, -2, -1, -2, -2, 0, 3, 0, 0, 0, 0, 0, 2, 2, 0, 0, -3, -2, -2, -2, -1, -1, 1, 0, 0, 0, 1, 1, 2, 5, 5, 2, -1, -1, -1, -2, -2, 0, 3, 1, -1, 0, -1, 0, 1, 2, 1, 0, -4, -4, -3, 0, 0, -1, 1, 0, 0, 0, 1, 0, 2, 6, 6, 1, -2, -2, -1, -3, -2, 0, 4, 2, 0, -2, -3, 0, 0, 0, 2, 0, -4, -4, -2, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 6, 5, 2, -1, -1, -1, -4, -4, -1, 3, 3, 0, -3, -3, -3, -1, 0, 0, -2, -4, -4, -2, 0, 0, -1, 0, -1, 0, 0, 0, 1, 4, 5, 6, 2, 0, 0, -2, -2, -5, -1, 1, 1, 0, -3, -3, -4, -2, 0, 2, 0, -5, -4, -3, 0, 0, -1, -1, -1, -1, -1, 0, 3, 4, 5, 4, 1, 0, 1, 0, -2, -3, -1, 0, 0, 0, 0, 0, -2, -1, 0, 3, 1, 0, -1, -2, 0, 0, -1, -1, -3, -2, 0, 1, 3, 5, 3, 3, 1, 0, 2, 2, 0, -1, -1, 1, 1, 2, 3, 3, 2, 4, 6, 6, 4, 4, 0, 0, 1, 0, -2, 0, -1, -5, -1, 0, 1, 3, 4, 2, 1, 0, 1, 1, 0, 0, 0, 0, 3, 4, 8, 8, 9, 9, 9, 9, 6, 6, 6, 3, 3, 3, -1, -1, 0, -1, 0, 0, 1, 1, 2, 1, 1, 0, 1, 0, 1, 0, 0, 1, 2, 5, 6, 6, 6, 6, 6, 7, 5, 6, 6, 4, 3, 2, 0, -1, 2, 5, 6, 5, 3, 3, 1, 1, 0, 0, 1, 0, -1, -2, -2, -2, -3, -2, -2, -1, -2, -1, -1, -2, -2, 0, 0, 0, 2, 1, 3, 2, 4, 8, 6, 7, 4, 3, 2, 1, 0, 1, 1, 0, 0, -1, -2, -2, -2, -3, -4, -2, -2, -3, -3, -3, -2, -1, -1, 0, 0, 0, 3, 1, 5, 9, 9, 6, 4, 2, 2, 1, 1, 2, 0, -1, -1, -2, -5, -4, -5, -6, -5, -3, -5, -4, -4, -4, -4, -3, 0, 0, 0, 2, 2, 4, 5, 9, 7, 5, 2, 0, 0, 1, 0, 2, 0, 0, 0, -1, -1, -1, -1, -2, -2, 0, -2, -4, -3, -4, -2, -1, -2, -1, -1, 0, 0, 1, 5, 7, 5, 4, 0, 1, 1, 0, 2, 1, 0, 3, 2, 0, 1, 0, 0, 0, 0, 0, 0, -2, -3, -2, -2, -3, -2, -2, -2, -2, 0, 1, 3, 5, 3, 1, 1, 1, 1, 1, 2, 2, 3, 3, 2, 0, 1, 2, 0, 1, 2, 0, -2, -2, -2, -2, -3, -4, -3, -3, -3, -3, 0, 1, 3, 5, 2, 1, 1, 1, 0, 1, 1, 3, 3, 2, 0, -1, 0, 0, 0, 0, 1, 0, 0, -3, -2, -3, -3, -3, -4, -2, -4, -3, 0, 0, 3, 4, 0, 0, 1, 1, 2, 1, 2, 2, 3, 1, 0, -2, -1, -1, 0, 0, 0, 0, 0, 0, -1, -3, -2, -4, -5, -3, -4, -4, 0, 2, 3, 2, 0, -2, -3, 0, 2, 2, 1, 1, 2, 0, 0, -3, -1, -2, -2, -2, -1, 0, 0, 0, -1, -2, -2, -3, -4, -3, -3, -2, 0, 1, 2, 1, -2, -4, -4, -2, 2, 0, 1, 0, 0, 0, -1, -2, -2, -1, -2, 0, 0, 0, 1, 0, -2, -3, -2, -2, -4, -3, -3, -2, 0, 2, 2, 0, -2, -6, -5, -2, 0, 1, 0, 0, -1, 0, -1, -2, -2, -1, -2, 0, 0, 1, 0, -1, -4, -3, -2, -2, -2, -2, -1, 0, 2, 3, 1, 0, -3, -5, -4, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, -2, -4, -5, -3, -1, -2, -2, 0, 0, 1, 3, 2, 0, -2, -4, -3, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, 0, 1, 0, 0, -1, -3, -4, -2, -2, -1, -1, 0, 0, 2, 5, 1, 3, 0, -1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -2, -2, 0, 0, 0, 1, 0, -4, -4, -3, -1, -1, -1, 0, 1, 5, 6, 2, 3, 2, 0, 0, 0, 0, 1, 2, 3, 3, 1, 0, -1, -2, -1, -2, 0, 1, 2, 2, 0, -3, -4, -4, -3, -2, 0, 0, 2, 4, 5, 3, 5, 2, 0, 0, 1, 3, 3, 2, 4, 2, 2, 1, 0, 0, 0, 0, 0, 3, 3, 2, 0, -2, -4, -2, -2, -1, 0, 1, 3, 4, 4, 4, 6, 3, 0, 0, 1, 3, 2, 3, 2, 2, 2, 0, -1, -1, 0, 0, 0, 2, 2, 1, 0, -2, -4, -2, -1, 0, 0, 2, 2, 3, 4, 3, 6, 2, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, -1, 1, 0, 1, 0, 0, 0, -2, -4, -3, -2, -1, -1, 1, 1, 1, 3, 4, 4, 3, 2, 0, -2, -2, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, -1, -3, -2, -3, -4, -2, -1, 0, 0, 1, 1, 5, 4, 3, 3, 0, -2, -3, -3, -2, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, -1, -2, -2, -2, -1, -2, -1, 0, 0, 1, 4, 3, 2, 2, -1, -3, -3, -2, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 1, 2, 2, 1, 0, 0, -1, -2, -2, -2, -1, 0, 0, 1, 3, 3, 3, 3, -1, -1, -3, -1, -1, 1, 0, 1, 0, 0, -2, -2, -2, 0, 2, 3, 3, 0, 0, 0, 0, -2, -3, -1, -1, -2, 0, 0, 3, 3, 2, 4, 0, -1, 0, -1, -1, 1, 2, 1, 2, 0, -1, -1, -2, 0, 1, 2, 2, 0, 0, 0, -2, -2, -3, -3, -2, -3, -2, 1, 2, 2, 3, 4, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, -1, -1, 0, 0, 0, 2, 1, -1, -2, -2, -3, -5, -4, -3, -4, -3, -2, 0, 1, 3, 3, 4, 1, 1, 1, 2, 1, 2, 2, 1, 0, -1, 0, 1, 1, 0, 2, 1, 0, -2, -2, -2, -4, -6, -4, -6, -5, -5, -4, 0, 1, 1, 2, 3, 3, 2, 2, 2, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -2, -4, -4, -6, -5, -5, -6, -4, -5, -1, 0, 2, 3, 4, 4, 3, 3, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, -3, -5, -7, -5, -4, -5, -5, -2, 0, 1, 3, 4, 6, 4, 2, 3, 2, 1, 2, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -4, -5, -7, -5, -3, -2, -1, 0, 0, 3, 4, 5, 6, 5, 5, 3, 2, 2, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -4, -6, -6, -4, -1, 0, 0, 0, 2, 4, 3, 4, 7, 5, 6, 6, 4, 4, 3, 2, 1, 0, 0, -1, 0, -2, -2, -3, -2, -3, -3, -5, -5, -6, -6, -2, -1, 0, 1, 2, 2, 4, 4, 5, 8, 8, 6, 6, 6, 3, 3, 2, 2, 0, -1, -1, 0, -2, -3, -3, -3, -4, -4, -5, -4, -4, -3, -2, -1, 0, 1, 2, 2, 5, 4, 2, 5, 5, 6, 4, 4, 4, 2, 2, 1, 0, 0, -2, 0, 0, -1, -2, -1, -1, -2, -2, -2, -2, -1, 0, -1, 0, 0, 0, 1, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 5, 4, 4, 4, 2, 1, 1, 1, 1, 0, 0, 0, -1, -2, -2, -3, -4, -3, -1, -1, -1, -1, 0, -1, -1, 0, 0, 2, 2, 3, 1, 3, 5, 6, 4, 4, 2, 1, 1, 2, 1, 0, 0, 0, -1, -2, -2, -2, -1, -3, -2, -1, -2, -3, -3, -3, -3, -2, -1, -1, 0, 1, 0, 5, 6, 7, 3, 2, 0, 0, 1, 1, 2, 1, 1, 0, -2, -1, -2, -1, -2, -1, -2, -3, -3, -3, -4, -3, -2, -1, -1, -2, 0, 1, 2, 4, 4, 4, 3, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -3, -2, -2, -3, -3, -1, -2, -2, -1, 0, 0, 4, 4, 3, 1, 1, 0, 0, 0, 1, 1, 1, 1, 2, 0, 2, 0, 0, 0, 0, 0, -1, -2, -1, -3, -2, -3, -2, -2, -3, -2, 0, 1, 4, 2, 1, 0, 1, 0, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, -1, -2, -2, -3, -3, -2, -3, 0, 0, 4, 3, 1, 0, 0, 1, 1, 1, 2, 2, 2, 1, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, -1, -2, -3, -3, -2, 0, 0, 2, 1, 1, 0, 0, 1, 1, 2, 2, 3, 1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -3, -2, -2, -3, -2, -1, 0, 2, 0, 0, -3, -1, 0, 1, 0, 2, 0, 1, 0, -1, -1, 0, -1, -1, 0, 1, 0, 1, 0, 0, -2, -2, -2, -3, -2, -2, -2, 0, 0, 2, 0, -3, -3, -2, -1, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 2, 1, 0, -2, -2, -2, -1, -1, -1, -2, -1, 0, 0, 2, 0, -3, -3, -2, 0, 1, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -2, -2, -2, -1, 0, -1, -2, 0, 1, 0, 2, 0, -2, -4, -3, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -3, -2, -2, -1, -1, 0, 0, 0, 2, 1, 1, 0, 0, -2, -2, -1, -1, -1, -1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 2, 1, 0, -3, -3, -1, 0, 0, 0, 0, 0, 2, 2, 2, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 2, -1, -2, -2, -2, -1, 0, -1, 1, 0, 2, 1, 2, 3, 3, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, -1, 0, -1, -1, 0, 2, 3, 2, 0, -1, -1, -1, -1, 0, 0, 1, 1, 3, 2, 3, 3, 1, 0, 0, 0, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 4, 2, 0, 0, -2, -1, 0, 0, 0, 0, 1, 3, 2, 3, 3, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 2, 2, 1, 0, 0, -1, -3, -3, -1, 0, 1, 1, 0, 2, 1, 4, 2, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -2, -1, -2, -3, 0, 0, 1, 0, 0, 3, 1, 2, 1, 0, -2, -3, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, -1, -2, -2, -2, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 3, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 2, 2, 1, 1, -1, -1, -1, -1, -1, 0, 1, 1, 0, -1, -2, -1, -1, 0, 2, 5, 2, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 0, -1, -1, -1, -1, 1, 1, 1, 2, 0, 0, -2, 0, 0, 2, 3, 2, 1, 2, 0, -1, 0, -1, 0, -1, 0, 0, 1, 0, 0, 3, 1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 2, 3, 2, 0, 0, 0, 0, -2, -3, -1, 0, -1, -1, 0, 0, 1, 2, 2, 1, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 1, 0, -2, -4, -2, -2, -1, -3, -2, -2, 0, 0, 3, 1, 1, 2, 0, 1, 2, 1, 1, 1, 0, 0, 1, 2, 1, 0, 2, 1, 0, 0, 0, 0, -2, -4, -3, -4, -2, -4, -3, -3, 0, 0, 1, 2, 3, 1, 2, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -3, -3, -3, -3, -2, -3, -4, -1, 0, 0, 3, 4, 3, 2, 2, 0, 2, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, -1, -2, -3, -4, -3, -2, 0, -1, -1, -1, 1, 1, 2, 4, 4, 3, 1, 1, 0, 2, 1, 1, 0, -1, 0, 0, -1, 0, 0, 1, 0, 1, -1, -3, -5, -3, -2, -1, 0, 0, -1, 0, 2, 0, 3, 4, 4, 3, 3, 2, 2, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -4, -3, -3, -2, -1, 0, 1, 1, 0, 3, 2, 4, 6, 5, 5, 4, 3, 2, 1, 1, 1, 0, -1, 0, 0, -2, -1, -2, -1, -1, -2, -4, -4, -3, -3, -3, 0, 0, 0, 0, 1, 3, 3, 2, 4, 5, 5, 5, 3, 4, 1, 0, 1, 0, -1, 0, -1, -2, -2, -2, -1, -2, -3, -2, -3, -2, -3, -2, -2, 0, 0, 0, 1, 2, 1, 1, 2, 3, 1, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 1, 1, 1, 0, 1, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 2, 1, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, -1, -2, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, -2, -3, -2, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 1, 0, 0, -2, 0, 0, -1, 0, -2, 0, 0, -2, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, -1, 0, 0, -1, -1, 0, -1, 1, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 2, 0, 0, -2, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 1, 2, 2, 2, 0, 0, 0, -2, 0, -2, -2, -1, 0, 0, 0, -1, -1, 0, 0, 0, -2, 0, 0, 0, 1, 2, 1, 1, 1, 0, 1, 2, 1, 2, 2, 2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -3, -1, 1, 2, 2, 2, 2, 2, 0, 0, 0, 1, 2, 1, 2, 1, 0, 0, 0, -2, -2, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 1, 2, 3, 3, 2, 2, 1, 0, 0, 1, 1, 1, 2, 2, 0, 0, 0, 0, -2, -2, -2, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 1, 3, 3, 4, 4, 3, 0, 0, 2, 3, 2, 0, 0, 0, 0, 0, -1, -1, -3, -1, 0, -1, -2, -1, -1, 0, 0, 1, 0, 0, -1, 0, 2, 1, 2, 2, 3, 2, 1, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, -1, -2, -2, 0, 0, -1, -1, 0, 1, 2, 1, 1, 0, 1, 0, 1, 2, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, -2, -2, 0, 0, -1, -2, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 2, 2, 2, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -2, -3, 0, -1, 0, -1, -1, -1, 1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -2, -3, -2, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 3, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 1, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 2, 2, 1, 1, 1, 0, 0, 1, 1, 0, 0, 2, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, 0, 1, 0, 0, 2, 2, 3, 2, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 2, 3, 1, 0, 0, 0, 1, 2, 2, 1, 2, 3, 1, -1, 0, -1, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 3, 1, 1, 0, 0, 0, 1, 1, 0, 3, 3, 1, 0, 0, -1, 0, -2, 0, 0, 0, -1, 0, 0, -2, -1, -2, -1, 0, 0, 1, 0, 1, 2, 2, 2, 1, 0, 1, 2, 1, 1, 3, 2, 0, 0, 0, 0, -2, -2, -2, -1, -1, -1, -1, 0, 0, -2, -2, -1, -1, 1, 0, 1, 1, 3, 3, 4, 3, 2, 1, 0, 1, 2, 3, 2, 0, 0, 0, 0, 0, -2, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 2, 3, 2, 3, 2, 2, 1, 0, 1, 1, 1, 0, 0, -1, -1, -1, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 3, 3, 2, 2, 1, 0, 1, 1, 2, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 3, 1, 1, 0, 1, 0, 1, 2, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -2, -1, 0, 1, 1, 0, 1, 3, 2, 2, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 2, 0, 2, 2, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, -1, -2, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 2, 1, 1, 2, 1, 0, 1, 0, 0, 0, -1, -2, 0, -1, -1, -2, -1, -3, -2, -1, -1, -2, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 0, 1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 2, 1, 0, 1, 2, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, -1, -1, -1, -2, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 2, 0, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, -2, -1, 0, 0, 0, 1, 0, 1, 0, 3, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 2, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 2, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 2, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, -1, 0, 0, 0, 0, 0, 3, 0, 1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -1, 1, 0, 0, 0, 1, 1, 2, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -2, -1, 0, 0, -1, 0, 0, 0, 1, 3, 0, 1, 1, 0, -1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 1, 2, 0, 1, 2, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, -2, -1, -1, 0, 0, 0, 1, 0, 1, 3, 0, 1, 1, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 1, 1, 0, 1, 3, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 1, 3, 0, 3, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, -1, 0, -1, 0, 1, 0, 1, 0, 0, -1, 0, -1, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, 0, 0, -1, -1, -1, 0, -1, -1, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 3, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -2, -2, -2, -1, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 3, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 2, 1, 0, 0, 0, 0, 2, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 1, 2, 0, 2, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 3, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 0, 1, 1, 1, 2, 3, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 1, 1, 0, 0, 1, 0, 0, 2, 1, 2, 1, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 2, 1, 2, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 2, 0, 0, 2, 2, 0, 0, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 3, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, 1, 1, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 0, 0, -1, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 1, 1, 1, 2, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 2, 0, -1, -2, -1, 1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 1, 0, 0, 0, 1, 1, 2, 1, 0, 0, -2, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 2, 2, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 1, 2, 1, 2, 1, 0, 0, -2, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 1, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, 1, 0, 1, 2, 0, 1, 0, 0, 1, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 2, 0, 1, 0, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 2, 0, 1, -1, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, -2, 0, 0, 0, 1, 1, 1, 0, 2, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 0, 0, -1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 2, 0, 0, 2, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, -1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 3, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, -1, -1, -1, -1, 0, 1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -2, -1, -2, -1, -1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, -2, -1, -3, 0, -1, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, -2, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 1, -1, 0, 0, 2, 1, 1, 1, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, -2, -1, 0, 1, 1, 0, 1, 0, 0, -1, 0, -1, 1, 1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, -1, -2, 0, 0, 1, 0, -3, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, -3, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 2, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, -2, -1, 0, 1, 0, 1, 0, 2, 1, 1, 1, 0, 0, 0, -1, 0, 0, 2, 3, 2, 2, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, -2, -3, 0, 0, 1, 0, 0, 2, 2, 2, 1, 1, 1, 1, 0, 0, -1, 2, 2, 2, 2, 2, 1, 0, 1, 0, 0, 1, 1, 1, 2, 0, -2, -3, -1, 0, 0, 0, 0, 2, 2, 3, 3, 1, 0, 2, 1, 0, 0, 2, 2, 1, 1, 3, 1, 0, 0, 0, 1, 0, 2, 1, 2, 1, -1, -2, 0, 0, 0, -1, -1, 0, 1, 3, 2, 2, 2, 1, 1, 0, 0, 2, 1, 2, 0, 2, 1, 0, 0, 0, 1, 1, 2, 1, 2, 2, -1, -2, -1, 0, 0, -1, -2, 0, 1, 3, 1, 1, 1, 1, 0, 0, 0, 1, 3, 1, 0, 3, 3, 2, 1, 0, 0, 2, 2, 2, 3, 1, 0, -2, 0, 0, 0, -1, 0, -3, -1, 2, 0, 1, 0, 1, 1, 0, 0, 2, 2, 2, 0, 1, 2, 2, 1, 0, 0, 2, 1, 3, 3, 2, 0, -1, 0, 0, 1, 0, 0, -2, -1, 0, 1, 0, 2, 0, 1, 0, 0, 1, 3, 1, 2, 2, 2, 4, 1, 0, 0, 1, 2, 2, 3, 3, 0, -1, -1, 1, 0, 0, 0, 0, -1, 0, 0, 1, 2, 2, 1, 1, 0, 0, 2, 1, 3, 2, 1, 2, 2, 0, 0, 0, 2, 2, 1, 2, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 1, 3, 2, 1, 3, 2, 2, 3, 3, 0, -1, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 2, 2, 1, 3, 1, 3, 2, 2, 4, 2, 1, 2, 2, 1, 0, 0, 0, 0, 1, 1, 0, -1, -1, 0, 1, 0, 1, 1, 1, 0, 0, 1, 0, 2, 2, 2, 2, 2, 3, 3, 3, 2, 2, 3, 3, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 2, 3, 2, 1, 2, 0, 2, 1, 0, -1, 0, -1, 0, 1, 2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 2, 1, -1, 1, 0, 0, 0, 0, 1, 2, 3, 2, 1, 1, 2, 2, 0, 0, 0, 0, -1, 2, 1, -1, -2, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, 0, 1, 2, 1, 1, 2, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, -1, -1, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 2, 2, 4, 3, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, -2, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 2, 1, 2, 1, 2, 2, 1, 2, 5, 3, 1, 0, 0, 0, 0, 2, 1, 0, 1, 0, -1, -3, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 1, 2, 1, 2, 0, 1, 0, 3, 3, 3, 0, 1, 2, 1, 1, 2, 2, 1, 3, 1, -2, -1, 0, 1, 2, -1, 0, 1, 0, 1, 2, 1, 2, 2, 2, 2, 2, 0, 0, 2, 4, 3, 0, 1, 1, 0, 2, 1, 2, 1, 2, 1, -1, -3, -1, 0, 0, -1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 0, 2, 2, 1, 0, 1, 1, 2, 3, 1, -1, -3, 0, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 2, 2, 0, 0, 1, 2, 3, 4, 3, -1, -4, 0, 0, 0, -2, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 2, 3, 1, 1, 0, 1, 3, 3, 2, -1, -2, 0, 0, 0, -2, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 2, 3, 3, -2, -3, -1, 0, -1, 0, 0, 0, -2, 0, 1, 2, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 2, 1, 0, 0, 0, 2, 3, 2, 2, -2, -2, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 2, 0, 0, 0, 0, 1, 1, 2, 1, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, -2, -3, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -3, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, 1, -2, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, -1, 0, -1, 0, 1, 0, 0, 2, 2, 1, 2, 1, 2, 2, 1, 2, 2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, 1, 1, 1, 1, 2, 0, 2, 2, 4, 2, 2, 2, 1, 1, 1, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 1, 0, 1, 2, 1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -2, -2, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, 0, 1, 0, 0, 0, -1, 0, -1, 0, -1, -2, -1, -1, -1, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, -2, 0, -1, 0, 0, 0, -1, -1, -2, -3, -2, -1, -2, -1, -1, -1, 0, 1, 0, 0, -1, 1, 0, 0, 0, -1, -1, 0, 0, -1, -2, -1, -2, 0, 0, -1, 0, -1, -1, -1, -4, -3, -3, -3, -2, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, -1, -1, 0, -1, -1, -2, -3, -4, -3, -4, -3, -3, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -3, -3, -4, -3, -3, -3, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, 0, -1, -2, -3, -2, -4, -4, -3, -1, -1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, -2, -3, -3, -3, -2, -2, -1, -1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, 0, 1, 1, 0, -1, 0, -2, -2, -2, -3, -2, -2, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, -2, -2, -3, -3, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, -2, 0, 0, -1, -2, -3, -2, -1, 0, 0, 1, 0, 0, 0, 1, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -1, -1, -2, -2, -3, -3, -1, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, -2, -2, -3, -1, 0, 0, 1, 0, 0, 0, 2, 2, 0, 0, 0, 0, -2, -1, -2, 0, 0, 0, 2, 1, 1, 0, -1, -1, -2, -1, 0, 0, -1, -2, -3, -2, -1, -1, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 2, 0, 0, -1, -1, -1, -2, -1, 0, -1, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 1, 1, 0, 0, -2, -1, -1, -2, -2, -3, -1, -2, -2, -1, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, -1, -1, -2, -2, -3, -3, -2, -3, -1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, -1, -1, -2, -1, 1, 0, 1, 0, 1, 0, 0, 0, -2, -1, -1, -2, -3, -3, -2, -3, -2, -2, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -3, -3, -2, -4, -4, -2, -2, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -2, -3, -3, -3, -2, -1, -1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -2, -1, -3, -3, -2, -2, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -2, -3, -3, -3, -1, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, -1, -1, -1, -2, -2, -3, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, -2, -2, -1, -1, -1, -2, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, 0, 0, -1, -2, -1, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 1, 1, 2, 2, 1, 3, 2, 3, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, -1, -1, 0, 1, 1, 1, 3, 2, 3, 2, 4, 3, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, -1, 4, 3, 2, 1, 0, 0, 0, 0, -1, -1, -2, -3, -5, -5, -3, -5, -3, -4, -1, 0, 0, 0, 0, 1, 3, 5, 5, 4, 4, 4, 5, 0, 4, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, -3, -4, -4, -3, -1, -2, -2, -1, -1, 0, 0, 1, 1, 3, 5, 4, 4, 3, 3, 5, -1, 3, 2, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 3, 3, 2, 1, 2, 3, 0, 4, 1, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -1, 0, 1, 2, 1, 0, 0, 1, 2, 3, 0, 3, 1, 0, 0, 0, 0, -2, -1, -2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, -2, -1, -2, 0, 0, -1, 0, -1, 0, 3, 2, 0, 3, 2, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -3, -2, -2, -3, -4, -3, -1, -1, 0, 1, 4, 0, 3, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, -4, -3, -4, -5, -3, -3, -1, -1, 3, 3, 0, 4, 1, -1, 0, 1, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -3, -4, -3, -3, -5, -3, -3, -2, 0, 2, 3, 0, 2, 0, 0, 0, 1, 0, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 1, 0, -2, -2, -1, -3, -3, -2, -4, -4, -4, -1, 0, 3, 3, 0, 1, 0, -2, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, -1, -2, -4, -3, -1, -4, -4, -4, -2, 0, 2, 3, 0, 1, -1, -1, 0, 1, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 1, 1, 1, -1, -1, -3, -3, -3, -2, -3, -3, -3, -1, 0, 3, 4, 0, 1, -1, -1, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 2, 1, 0, -1, -2, -4, -3, -2, -2, -3, -2, -1, 0, 4, 5, 0, 3, 1, -1, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 1, 3, 3, 3, 0, -1, -1, -3, -2, -2, -3, -2, -3, -1, 2, 3, 3, 0, 3, 0, -1, 0, 1, 0, 0, 1, 3, 3, 2, 0, 1, 0, 2, 2, 5, 3, 2, 0, -2, -4, -3, -1, -1, -1, -1, 0, 2, 2, 3, 1, 3, 1, 0, -1, 0, 0, 1, 0, 2, 1, 2, 1, 0, 1, 1, 3, 5, 4, 2, 0, -2, -2, -2, -1, -2, 0, 0, 0, 0, 3, 2, 0, 4, 0, -1, -2, 0, 1, 1, 0, 1, 0, 2, 1, 1, 1, 3, 3, 5, 5, 2, 1, -2, -4, -2, -1, -1, -1, 0, 1, 0, 3, 3, 0, 4, 0, -3, -2, -1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 4, 4, 5, 3, 0, 0, -3, -4, -2, -1, -1, 0, 1, 0, 0, 1, 3, 0, 4, 0, -3, -2, 0, -1, 0, -1, -1, 0, 0, 1, 0, 2, 3, 4, 4, 3, 0, -1, -5, -4, -2, -1, 0, 0, 0, 0, 0, 1, 3, 0, 2, 0, -2, -3, -1, -1, -1, 0, -2, 0, 0, 0, 1, 3, 1, 1, 1, 0, 0, -1, -4, -4, -4, -2, -2, 0, 0, 0, 1, 2, 2, 0, 2, 0, -2, -2, -1, -1, 0, 0, -2, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, -2, -3, -3, -2, -3, -3, -1, 0, 0, 0, 3, 3, 0, 3, 0, -2, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, -1, -3, -3, -2, -2, -3, -2, -3, -2, 0, 1, 3, 1, 2, 0, -2, -2, -2, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 2, 1, 1, 0, 0, -2, -4, -3, -4, -3, -3, -2, -2, 0, 2, 2, 0, 3, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, -1, -1, 0, 1, 0, 0, -1, -1, -3, -4, -4, -3, -3, -2, -3, -3, -1, 0, 0, 2, 0, 1, 0, -2, -1, -2, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, -1, -2, -3, -5, -6, -5, -4, -3, -3, -3, -1, 0, 0, 2, 0, 3, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, -2, -2, -5, -5, -5, -4, -3, -4, -4, -2, 0, 2, 4, 0, 3, 2, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, -1, -3, -4, -5, -6, -3, -2, -3, -3, -2, 1, 2, 3, 0, 3, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, -1, 0, -1, -1, -4, -4, -4, -5, -3, 0, -1, 0, 0, 2, 4, 3, 0, 4, 3, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -3, -4, -3, -3, -2, 0, 0, 0, 0, 1, 3, 4, 4, 0, 5, 2, 1, 1, 0, 0, 0, 1, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, -2, -2, -2, -1, 0, 1, 4, 3, 3, 4, 4, 5, 5, 0, 5, 3, 1, 0, 0, 1, 2, 1, 0, -2, -2, -1, -1, -3, -3, -3, -3, -2, -2, -2, -2, -1, 1, 3, 5, 5, 5, 5, 6, 7, 4, 0, 4, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -2, -2, -1, 0, 0, -1, 0, 0, 0, 3, 2, 2, 2, 4, 4, 4, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, -2, -2, 0, 0, 1, 0, 0, 2, 2, 3, 2, 0, 0, 2, 1, 2, 3, 3, 2, 3, 3, 2, 3, 3, 4, 3, 0, 0, 0, -1, -1, -2, -1, -2, 0, 2, 1, 1, 0, 2, 2, 3, 1, 1, 1, 3, 2, 3, 3, 2, 2, 2, 3, 3, 3, 4, 4, 3, 0, -2, -1, 0, -2, -2, -1, 0, 0, 1, 2, 0, 1, 2, 2, 2, 2, 0, 0, 2, 1, 1, 1, 0, 0, 1, 2, 1, 2, 2, 3, 1, 0, -3, -2, -2, -3, -1, -1, 0, 0, 2, 2, 0, 1, 0, 1, 2, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 1, 1, -1, -2, -2, -3, -3, -2, -1, 0, 1, 2, 1, 0, 0, 0, 0, 0, -1, -2, 0, -1, -2, 0, -2, -2, -2, 0, 0, -1, 0, 0, 0, 0, -1, -2, -1, -1, -3, -2, -1, -1, 1, 2, 2, 0, -1, 0, 0, 0, -1, -2, -1, -3, -3, -1, 0, -1, -1, -1, 0, -1, 0, -1, -1, 0, 0, -2, -2, -1, -2, -1, 0, 0, 1, 2, 3, 1, 0, 0, -1, -1, -2, -2, -1, -3, -3, -2, 0, -1, -2, 0, -1, -1, -2, -4, -1, -2, -1, 0, -2, -1, -1, -2, -1, 0, 1, 2, 2, 1, 0, -1, 0, -2, -3, -2, -2, -1, -2, -2, -1, 0, -1, 0, -1, -2, -2, -4, -4, -3, -2, -3, -1, -2, -1, 0, 0, 0, 1, 3, 3, 2, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -2, -3, -3, -1, -2, -1, -3, -2, 0, 0, 0, 2, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, -1, -3, -3, -1, 0, -2, -3, -3, 0, -1, 0, 3, 2, 1, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, -1, -3, -1, -2, -1, 0, -3, -5, -1, 0, 1, 2, 1, 0, 0, 1, 0, -1, -2, -1, -2, -1, -2, 0, 1, 0, 0, -1, 0, -2, 0, 0, 0, -1, -2, -1, -2, -1, -3, -3, -1, 0, 0, 1, 2, 0, 0, -1, 0, -1, -3, -3, -2, -3, -1, 0, 1, 0, -1, 0, -2, -2, -1, 0, 0, -1, -2, -3, -3, -1, -3, -3, -3, -1, 0, 1, 0, 1, 0, -1, 0, -3, -3, -3, -5, -1, -1, -1, 0, -1, -2, -2, -3, -3, -2, 0, 1, -2, -1, -2, -4, -2, -2, -3, -2, -1, 0, 1, 1, 0, 0, 0, -2, -2, -2, -4, -3, -2, -3, -2, 0, -1, -1, -2, -3, -4, -3, 0, 1, 0, -3, -3, -3, -3, -3, -3, -2, -2, 0, 0, 2, 1, 0, -1, -2, -3, -4, -3, -2, -2, -2, -1, 0, 0, 0, -2, -2, -4, -2, 0, 1, 0, -2, -1, -4, -4, -2, -3, -2, 0, 0, 0, 1, 1, 0, -2, -2, -4, -5, -5, -4, -2, -1, -1, 0, 0, 0, -1, -3, -2, 0, 0, 2, 0, -1, -2, -3, -4, -4, -3, -2, -1, 0, 1, 0, 2, 0, 0, -3, -4, -3, -3, -3, -3, -1, -1, 0, 1, -1, -2, -2, -1, 0, 0, 1, 0, -1, -1, -3, -4, -2, -3, -2, 0, 0, 1, 1, 2, 1, 0, -3, -4, -4, -3, -1, -2, 0, 0, 1, 0, -1, -1, -3, -2, 1, 0, 0, 0, -1, -1, -3, -2, -3, -3, -1, -1, 0, 1, 3, 3, 1, -1, -3, -4, -4, -1, -2, -3, 0, 0, 0, -1, 0, -2, -2, -1, 0, 0, -1, 0, -1, -2, -3, -2, -2, -3, -2, -2, 0, 2, 1, 2, 2, -1, -1, -3, -4, -2, -2, -2, -2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, -2, -2, -2, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -2, -2, -3, -4, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -2, -4, -3, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -3, -2, -3, -2, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -3, -3, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, -2, -3, -2, -2, 0, 0, 1, 0, 1, 0, 0, 1, 1, 1, 0, 0, -2, -3, -3, -2, -2, -2, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -2, -2, -2, -1, -2, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -2, -3, -3, -2, 0, -1, -1, -1, 0, 0, 1, 0, 2, 3, 2, 0, -2, -2, -1, -2, -2, 0, 1, 2, 0, -1, 0, 1, 0, 0, 0, 0, -2, -4, -2, -1, -1, -2, -1, -1, 0, 0, 1, 1, 3, 3, 1, 0, -2, 0, -1, -3, -3, 0, 1, 1, -1, 0, -1, 0, 0, 0, 0, -1, -2, -3, -3, -2, -2, -2, -1, -1, 0, 1, 0, 2, 3, 3, 3, 0, -2, 0, 0, -1, -3, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -1, -2, -1, -1, 0, 0, 0, 1, 3, 4, 2, 2, 0, -2, -1, 0, -2, -2, -1, 0, 0, 1, 0, 1, 2, 2, 0, 0, 0, 0, 0, -1, -2, -1, -1, -2, -1, -1, 0, 0, 2, 2, 2, 2, 0, 0, 0, 0, -2, -1, 0, 0, 0, 2, 3, 3, 4, 4, 2, 4, 2, 3, 1, 1, 0, 0, -1, -1, 0, 0, 0, 1, 2, 2, 2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 4, 5, 5, 5, 5, 3, 4, 4, 3, 2, 0, 0, 0, -2, -1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 2, 3, 3, 2, 3, 1, 1, 1, 2, 2, 0, 0, 0, 0,

    others => 0);
end iwght_package;
