library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    500, 500, 497, 498, 503, 503, 502, 507, 507, 497, 485, 495, 516, 532, 536, 537, 522, 507, 489, 477, 472, 473, 479, 482, 481, 491, 502, 516, 517, 510, 
    515, 516, 509, 502, 505, 502, 504, 507, 502, 464, 445, 469, 505, 527, 527, 517, 505, 473, 439, 412, 407, 426, 448, 464, 473, 483, 494, 510, 514, 509, 
    516, 518, 519, 515, 511, 507, 508, 510, 497, 409, 381, 402, 465, 494, 495, 497, 475, 414, 369, 320, 310, 322, 364, 395, 421, 456, 479, 492, 503, 505, 
    497, 497, 505, 514, 514, 515, 514, 517, 508, 434, 397, 370, 439, 479, 469, 449, 418, 369, 298, 235, 221, 244, 282, 313, 374, 415, 453, 466, 480, 490, 
    469, 476, 496, 507, 516, 519, 520, 523, 518, 457, 398, 378, 403, 411, 400, 407, 381, 313, 231, 187, 193, 215, 234, 275, 311, 368, 424, 448, 466, 480, 
    402, 409, 466, 497, 515, 526, 525, 520, 515, 492, 435, 379, 362, 355, 347, 345, 327, 280, 219, 183, 200, 235, 259, 273, 300, 354, 397, 429, 455, 470, 
    322, 334, 388, 443, 496, 520, 508, 480, 475, 451, 396, 332, 295, 293, 303, 304, 301, 293, 251, 215, 219, 263, 293, 295, 308, 334, 390, 424, 447, 464, 
    209, 228, 294, 358, 459, 506, 443, 348, 301, 293, 293, 262, 231, 255, 279, 295, 312, 319, 270, 240, 222, 249, 285, 306, 313, 321, 361, 416, 448, 464, 
    134, 135, 185, 295, 421, 491, 380, 247, 150, 168, 175, 191, 190, 233, 278, 296, 324, 328, 278, 226, 181, 227, 273, 290, 299, 306, 342, 393, 430, 459, 
    82, 98, 108, 245, 389, 475, 384, 218, 74, 82, 124, 148, 168, 217, 270, 279, 339, 312, 242, 182, 139, 211, 253, 286, 286, 280, 305, 354, 396, 437, 
    71, 74, 87, 221, 377, 471, 418, 231, 140, 124, 150, 132, 145, 184, 243, 259, 310, 272, 210, 133, 117, 203, 253, 286, 282, 285, 283, 312, 344, 409, 
    61, 66, 96, 214, 377, 467, 468, 320, 235, 166, 167, 121, 108, 145, 213, 241, 286, 231, 173, 98, 127, 212, 269, 297, 293, 282, 267, 278, 304, 379, 
    56, 68, 85, 193, 368, 457, 483, 382, 296, 195, 175, 107, 104, 126, 179, 215, 263, 214, 152, 101, 129, 201, 252, 276, 280, 268, 253, 255, 294, 369, 
    43, 58, 65, 176, 312, 408, 448, 383, 309, 173, 95, 50, 72, 138, 194, 223, 252, 225, 171, 113, 144, 222, 267, 278, 279, 257, 245, 270, 314, 384, 
    25, 36, 33, 140, 225, 324, 365, 387, 318, 190, 113, 84, 110, 189, 214, 239, 282, 256, 215, 162, 165, 195, 253, 279, 276, 262, 270, 312, 361, 424, 
    0, 6, 5, 96, 167, 237, 264, 324, 295, 250, 146, 148, 209, 234, 259, 257, 272, 296, 326, 256, 226, 245, 292, 318, 310, 290, 300, 344, 403, 442, 
    0, 0, 0, 51, 128, 169, 200, 242, 282, 291, 232, 240, 255, 248, 262, 245, 261, 295, 298, 291, 302, 290, 319, 347, 345, 333, 352, 385, 431, 451, 
    0, 0, 0, 23, 116, 150, 176, 184, 217, 274, 275, 306, 257, 219, 208, 211, 241, 275, 282, 305, 304, 326, 368, 346, 354, 350, 387, 410, 437, 459, 
    0, 0, 0, 16, 97, 122, 115, 128, 194, 279, 279, 287, 202, 157, 136, 161, 227, 293, 308, 318, 325, 362, 372, 340, 342, 352, 400, 424, 444, 460, 
    33, 0, 5, 35, 107, 116, 60, 14, 42, 153, 197, 167, 115, 64, 41, 100, 179, 262, 309, 314, 316, 313, 290, 266, 251, 281, 320, 343, 356, 365, 
    28, 0, 10, 41, 93, 72, 11, 0, 0, 31, 115, 113, 71, 33, 37, 91, 160, 236, 263, 270, 253, 234, 206, 175, 162, 168, 177, 199, 203, 204, 
    11, 0, 0, 16, 56, 27, 0, 0, 0, 8, 59, 92, 77, 69, 77, 93, 120, 173, 197, 185, 158, 136, 113, 91, 73, 64, 64, 71, 70, 72, 
    7, 0, 0, 17, 35, 0, 0, 0, 0, 0, 75, 103, 100, 105, 105, 110, 117, 128, 124, 106, 91, 80, 63, 43, 30, 21, 18, 23, 26, 22, 
    0, 14, 13, 24, 0, 0, 0, 0, 0, 64, 101, 110, 111, 117, 120, 113, 106, 102, 91, 74, 59, 50, 35, 16, 10, 8, 9, 7, 0, 0, 
    0, 29, 43, 50, 0, 0, 0, 0, 32, 88, 79, 84, 88, 94, 101, 104, 99, 92, 81, 60, 38, 21, 11, 9, 7, 12, 0, 0, 0, 0, 
    0, 21, 49, 60, 0, 0, 0, 0, 73, 84, 70, 71, 79, 94, 98, 97, 89, 79, 62, 45, 27, 9, 0, 0, 3, 1, 0, 0, 0, 0, 
    0, 3, 33, 52, 11, 0, 0, 16, 89, 76, 57, 62, 65, 81, 92, 92, 80, 63, 47, 32, 13, 2, 2, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 32, 33, 6, 38, 53, 109, 94, 73, 61, 55, 66, 70, 70, 59, 48, 35, 25, 23, 20, 17, 4, 0, 0, 0, 0, 0, 24, 
    0, 0, 3, 15, 43, 44, 73, 103, 116, 108, 98, 86, 77, 75, 73, 70, 52, 26, 13, 16, 26, 33, 28, 4, 0, 0, 0, 0, 3, 55, 
    0, 3, 15, 18, 45, 75, 94, 119, 126, 124, 117, 102, 103, 110, 111, 95, 62, 29, 14, 16, 29, 50, 41, 7, 0, 0, 0, 0, 6, 64, 
    
    -- channel=1
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 95, 87, 77, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    53, 57, 23, 0, 0, 0, 0, 0, 0, 0, 68, 129, 105, 64, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    145, 111, 80, 77, 52, 24, 0, 0, 0, 0, 5, 28, 9, 1, 0, 0, 0, 0, 0, 0, 10, 32, 44, 49, 36, 17, 1, 0, 0, 0, 
    200, 106, 67, 59, 79, 78, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 33, 41, 39, 22, 0, 0, 0, 0, 0, 
    187, 62, 0, 0, 23, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    147, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 27, 37, 47, 54, 53, 44, 
    55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 32, 33, 45, 69, 83, 90, 96, 98, 87, 71, 55, 
    183, 169, 154, 140, 127, 114, 107, 100, 91, 75, 54, 29, 19, 28, 41, 42, 42, 59, 81, 91, 98, 110, 122, 122, 112, 105, 103, 99, 90, 74, 
    318, 306, 274, 256, 258, 262, 267, 267, 263, 250, 218, 179, 148, 138, 135, 131, 131, 139, 151, 161, 166, 168, 162, 143, 118, 109, 118, 121, 110, 84, 
    400, 398, 351, 311, 311, 341, 369, 389, 400, 397, 362, 288, 232, 213, 218, 219, 218, 216, 219, 215, 202, 180, 150, 126, 120, 132, 139, 133, 120, 84, 
    441, 441, 392, 358, 346, 373, 407, 441, 465, 474, 451, 341, 228, 156, 164, 182, 186, 186, 186, 180, 169, 155, 153, 163, 163, 156, 150, 144, 116, 63, 
    462, 471, 439, 412, 401, 416, 441, 464, 482, 493, 483, 389, 269, 165, 138, 159, 169, 178, 186, 197, 213, 221, 214, 203, 195, 192, 175, 135, 88, 34, 
    456, 488, 485, 468, 464, 469, 478, 490, 499, 504, 501, 441, 337, 275, 256, 272, 278, 284, 293, 303, 303, 289, 271, 257, 240, 206, 157, 104, 55, 1, 
    429, 481, 505, 504, 503, 504, 505, 507, 509, 510, 509, 492, 439, 416, 419, 431, 433, 428, 415, 394, 369, 340, 306, 265, 220, 177, 137, 85, 30, 0, 
    402, 468, 508, 509, 508, 506, 507, 511, 512, 512, 511, 514, 508, 524, 555, 569, 554, 506, 450, 399, 353, 305, 256, 214, 184, 159, 125, 73, 17, 0, 
    384, 460, 501, 505, 503, 501, 503, 507, 509, 510, 506, 510, 517, 539, 559, 544, 507, 449, 388, 328, 279, 239, 209, 189, 169, 142, 105, 56, 4, 0, 
    374, 453, 482, 487, 486, 485, 487, 490, 492, 491, 483, 481, 481, 482, 475, 453, 419, 371, 316, 269, 234, 209, 194, 180, 157, 126, 88, 43, 0, 0, 
    366, 430, 450, 454, 453, 449, 448, 448, 447, 442, 435, 429, 422, 411, 394, 363, 328, 302, 277, 252, 224, 203, 188, 167, 142, 111, 76, 34, 0, 0, 
    
    -- channel=2
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 26, 71, 105, 112, 88, 48, 0, 0, 0, 0, 0, 0, 0, 
    0, 27, 28, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 45, 60, 98, 125, 118, 136, 142, 117, 65, 4, 0, 11, 0, 11, 
    62, 96, 106, 104, 88, 78, 77, 64, 63, 58, 45, 35, 24, 16, 20, 35, 73, 101, 124, 131, 144, 180, 171, 156, 99, 67, 76, 108, 114, 126, 
    149, 166, 165, 152, 150, 152, 149, 136, 136, 133, 118, 100, 74, 59, 57, 73, 93, 102, 110, 120, 123, 136, 151, 179, 127, 93, 107, 140, 174, 171, 
    189, 185, 168, 160, 160, 178, 182, 158, 151, 144, 130, 100, 69, 53, 53, 75, 93, 97, 104, 118, 100, 89, 69, 88, 126, 112, 133, 138, 187, 182, 
    168, 173, 161, 151, 141, 156, 149, 123, 95, 86, 92, 74, 44, 34, 55, 87, 102, 106, 111, 116, 87, 62, 21, 30, 99, 100, 132, 143, 174, 190, 
    141, 142, 139, 151, 145, 153, 149, 107, 59, 46, 40, 25, 8, 9, 33, 59, 77, 78, 78, 72, 51, 24, 0, 6, 69, 108, 128, 171, 188, 224, 
    111, 123, 142, 153, 150, 145, 103, 49, 13, 0, 0, 0, 0, 0, 0, 0, 2, 2, 14, 22, 24, 17, 3, 15, 52, 125, 159, 230, 237, 252, 
    70, 88, 101, 95, 79, 53, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 38, 56, 53, 47, 48, 51, 118, 169, 232, 266, 261, 
    33, 39, 40, 32, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 71, 96, 88, 76, 63, 52, 93, 130, 158, 192, 201, 
    0, 5, 22, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 77, 103, 94, 70, 61, 49, 68, 97, 131, 140, 131, 
    16, 30, 31, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 27, 55, 66, 56, 42, 41, 36, 56, 82, 103, 109, 116, 
    36, 31, 22, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 14, 20, 18, 23, 32, 54, 85, 117, 154, 173, 149, 
    19, 33, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 37, 31, 15, 0, 0, 5, 13, 39, 69, 101, 131, 172, 207, 222, 215, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 82, 117, 95, 58, 17, 14, 34, 56, 84, 113, 150, 191, 221, 239, 265, 272, 
    0, 0, 0, 0, 0, 0, 13, 24, 29, 4, 0, 0, 8, 62, 122, 159, 136, 106, 71, 68, 87, 104, 136, 178, 213, 237, 255, 278, 301, 318, 
    11, 0, 0, 0, 2, 37, 73, 87, 86, 56, 26, 0, 17, 76, 139, 176, 166, 139, 116, 121, 141, 170, 205, 224, 246, 264, 285, 305, 325, 359, 
    45, 2, 0, 0, 17, 58, 102, 112, 102, 79, 63, 54, 79, 123, 152, 164, 161, 157, 164, 186, 206, 217, 225, 243, 274, 291, 308, 326, 354, 377, 
    66, 32, 19, 21, 47, 85, 124, 139, 142, 138, 125, 120, 131, 148, 165, 179, 188, 200, 213, 224, 232, 249, 260, 275, 290, 308, 327, 343, 359, 370, 
    122, 104, 95, 102, 122, 148, 163, 168, 169, 172, 180, 191, 201, 205, 212, 223, 227, 227, 235, 251, 273, 285, 283, 293, 306, 325, 339, 347, 352, 359, 
    204, 196, 192, 198, 206, 213, 213, 219, 230, 243, 250, 253, 247, 242, 245, 249, 238, 241, 262, 281, 295, 302, 309, 317, 327, 341, 346, 345, 346, 357, 
    288, 289, 293, 293, 291, 290, 285, 282, 280, 282, 280, 274, 265, 264, 276, 281, 262, 256, 263, 291, 311, 323, 332, 336, 342, 346, 346, 344, 353, 374, 
    350, 354, 351, 343, 335, 329, 320, 308, 298, 292, 292, 292, 288, 290, 305, 305, 270, 257, 269, 308, 334, 340, 343, 349, 349, 348, 345, 347, 375, 405, 
    370, 369, 364, 352, 341, 335, 329, 320, 312, 308, 304, 301, 297, 304, 328, 332, 292, 274, 285, 329, 346, 346, 354, 355, 354, 349, 344, 361, 400, 440, 
    365, 360, 356, 347, 340, 335, 331, 325, 319, 317, 318, 325, 333, 351, 381, 383, 337, 308, 309, 344, 355, 359, 361, 360, 358, 350, 355, 385, 427, 475, 
    
    -- channel=3
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 47, 55, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 63, 115, 115, 81, 76, 77, 81, 86, 80, 77, 70, 68, 63, 54, 52, 69, 28, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 66, 129, 123, 111, 115, 115, 131, 133, 109, 89, 81, 72, 69, 60, 60, 76, 34, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 11, 90, 121, 99, 114, 130, 134, 151, 163, 133, 112, 85, 77, 81, 73, 80, 75, 60, 8, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 58, 138, 154, 99, 99, 90, 101, 120, 139, 113, 92, 68, 71, 76, 80, 86, 44, 59, 38, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 44, 135, 132, 83, 68, 55, 80, 87, 96, 80, 68, 54, 54, 73, 82, 85, 48, 54, 36, 10, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 53, 55, 45, 38, 37, 42, 39, 44, 41, 37, 31, 36, 58, 70, 70, 33, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 19, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 27, 85, 107, 79, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 36, 108, 149, 124, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 33, 128, 183, 170, 110, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 51, 161, 226, 215, 163, 110, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 131, 237, 286, 262, 225, 178, 135, 88, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 136, 265, 329, 319, 304, 273, 238, 208, 183, 158, 133, 92, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 13, 156, 293, 350, 342, 329, 314, 303, 289, 271, 252, 240, 226, 191, 151, 115, 73, 25, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 13, 137, 242, 309, 344, 349, 314, 262, 218, 216, 262, 279, 272, 252, 245, 231, 171, 93, 22, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 38, 97, 144, 182, 216, 194, 154, 103, 71, 104, 137, 170, 154, 154, 170, 148, 94, 18, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 67, 98, 86, 46, 2, 0, 11, 35, 45, 37, 44, 55, 46, 11, 0, 0, 0, 0, 0, 
    32, 0, 5, 18, 24, 30, 36, 41, 38, 46, 66, 89, 91, 71, 34, 0, 0, 0, 14, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    86, 60, 61, 71, 74, 80, 87, 90, 94, 98, 97, 97, 92, 84, 69, 54, 45, 41, 39, 40, 42, 37, 29, 24, 22, 22, 27, 35, 41, 64, 
    170, 144, 145, 150, 157, 172, 183, 192, 201, 203, 207, 208, 203, 192, 173, 165, 167, 172, 179, 179, 180, 179, 177, 170, 165, 164, 169, 180, 184, 184, 
    239, 225, 222, 219, 217, 226, 237, 248, 257, 265, 269, 266, 263, 261, 256, 254, 260, 271, 281, 284, 285, 283, 282, 282, 282, 281, 290, 295, 264, 241, 
    292, 289, 288, 289, 293, 302, 311, 323, 331, 337, 334, 333, 334, 334, 333, 332, 339, 347, 355, 360, 361, 360, 360, 359, 358, 356, 345, 312, 268, 255, 
    350, 352, 353, 353, 354, 356, 362, 366, 371, 375, 369, 363, 364, 368, 366, 365, 363, 366, 371, 373, 370, 370, 368, 367, 361, 331, 286, 259, 247, 243, 
    348, 351, 347, 348, 349, 353, 356, 358, 360, 350, 338, 333, 337, 342, 341, 338, 333, 337, 342, 352, 358, 365, 370, 360, 319, 267, 242, 234, 237, 280, 
    363, 368, 363, 359, 354, 357, 361, 366, 371, 363, 351, 336, 340, 347, 348, 346, 340, 340, 340, 348, 355, 366, 359, 321, 279, 248, 230, 241, 296, 352, 
    
    -- channel=4
    321, 344, 376, 378, 354, 317, 306, 325, 380, 414, 417, 374, 353, 360, 347, 336, 318, 318, 306, 291, 309, 318, 288, 262, 314, 356, 388, 356, 337, 339, 
    287, 323, 343, 351, 322, 298, 296, 326, 384, 423, 422, 373, 362, 370, 352, 330, 305, 309, 307, 294, 311, 314, 284, 250, 295, 331, 357, 320, 305, 320, 
    247, 300, 310, 329, 299, 290, 288, 330, 390, 442, 436, 393, 374, 367, 351, 328, 303, 304, 305, 294, 317, 314, 272, 225, 253, 289, 310, 270, 263, 276, 
    264, 301, 301, 317, 291, 293, 290, 342, 397, 447, 427, 389, 357, 347, 328, 301, 288, 301, 323, 313, 327, 309, 258, 197, 211, 237, 254, 227, 227, 252, 
    305, 320, 332, 310, 292, 297, 301, 367, 403, 430, 398, 359, 322, 312, 322, 319, 292, 309, 340, 330, 339, 301, 230, 168, 164, 186, 219, 197, 225, 266, 
    338, 328, 346, 311, 295, 299, 321, 392, 404, 399, 359, 313, 298, 327, 358, 364, 330, 324, 329, 334, 335, 278, 223, 154, 136, 154, 193, 174, 225, 275, 
    340, 322, 306, 262, 278, 303, 332, 383, 384, 369, 314, 277, 312, 359, 386, 383, 347, 320, 317, 305, 290, 252, 223, 152, 139, 143, 173, 159, 233, 308, 
    325, 301, 252, 200, 238, 295, 348, 366, 346, 319, 266, 280, 342, 383, 400, 372, 322, 276, 290, 275, 253, 258, 229, 173, 147, 143, 157, 161, 258, 342, 
    309, 278, 214, 150, 192, 261, 345, 366, 330, 281, 244, 272, 320, 363, 369, 323, 274, 262, 266, 240, 247, 273, 243, 214, 164, 142, 147, 164, 274, 367, 
    310, 281, 213, 134, 142, 221, 300, 327, 312, 262, 247, 278, 291, 292, 272, 238, 236, 255, 253, 241, 259, 259, 236, 221, 172, 141, 137, 162, 293, 393, 
    325, 305, 240, 151, 127, 167, 221, 267, 277, 254, 262, 295, 301, 282, 233, 211, 229, 246, 248, 259, 272, 283, 249, 207, 178, 159, 143, 172, 301, 386, 
    319, 309, 253, 179, 141, 134, 172, 227, 246, 268, 290, 303, 286, 264, 249, 243, 247, 253, 252, 264, 261, 277, 244, 213, 193, 162, 149, 187, 278, 347, 
    302, 295, 252, 211, 163, 140, 142, 201, 258, 300, 299, 304, 295, 277, 261, 262, 274, 281, 277, 269, 252, 246, 225, 230, 214, 187, 164, 188, 264, 330, 
    286, 290, 249, 221, 179, 157, 134, 160, 233, 305, 322, 315, 296, 283, 260, 256, 267, 273, 275, 276, 255, 225, 198, 199, 210, 205, 168, 203, 293, 327, 
    277, 278, 239, 202, 179, 154, 154, 164, 208, 265, 295, 312, 272, 250, 255, 255, 244, 244, 238, 240, 235, 229, 188, 159, 192, 196, 190, 222, 298, 323, 
    263, 260, 225, 205, 181, 167, 166, 171, 178, 216, 232, 274, 256, 233, 222, 219, 239, 248, 243, 243, 235, 213, 182, 184, 185, 198, 205, 235, 309, 344, 
    236, 227, 197, 213, 191, 208, 186, 205, 189, 188, 199, 221, 233, 232, 210, 206, 206, 197, 203, 211, 226, 232, 203, 190, 210, 261, 247, 264, 301, 282, 
    199, 214, 207, 236, 235, 245, 218, 213, 217, 192, 192, 183, 197, 203, 182, 195, 189, 181, 196, 213, 218, 226, 217, 215, 254, 266, 291, 299, 289, 241, 
    194, 218, 220, 266, 277, 262, 264, 237, 236, 224, 222, 216, 185, 172, 159, 155, 165, 166, 166, 184, 208, 216, 220, 230, 264, 263, 299, 276, 253, 221, 
    213, 230, 253, 277, 279, 267, 263, 245, 240, 252, 224, 228, 187, 135, 132, 132, 149, 161, 176, 190, 214, 221, 228, 235, 263, 274, 262, 227, 211, 171, 
    234, 263, 289, 266, 277, 274, 241, 232, 227, 243, 232, 204, 182, 135, 114, 119, 137, 145, 184, 202, 212, 216, 231, 240, 259, 263, 226, 201, 178, 153, 
    227, 225, 224, 226, 263, 266, 235, 216, 214, 219, 234, 199, 172, 141, 136, 128, 133, 155, 184, 201, 223, 221, 233, 252, 273, 265, 225, 187, 154, 168, 
    178, 166, 148, 162, 221, 240, 220, 207, 205, 206, 207, 199, 174, 151, 162, 148, 137, 151, 183, 189, 198, 202, 237, 261, 293, 296, 248, 192, 164, 182, 
    186, 142, 102, 110, 165, 211, 211, 207, 211, 212, 183, 158, 170, 179, 200, 194, 171, 160, 171, 172, 186, 194, 236, 260, 301, 321, 273, 227, 183, 205, 
    216, 194, 153, 123, 129, 162, 194, 211, 221, 220, 204, 177, 180, 225, 258, 262, 227, 189, 171, 174, 175, 191, 221, 260, 309, 339, 299, 262, 218, 233, 
    277, 294, 274, 204, 153, 142, 152, 184, 221, 218, 201, 204, 212, 234, 260, 283, 258, 215, 183, 167, 164, 207, 233, 266, 320, 350, 313, 281, 235, 259, 
    311, 356, 379, 311, 232, 159, 136, 142, 179, 218, 226, 226, 237, 237, 244, 252, 239, 224, 197, 179, 188, 202, 240, 302, 343, 343, 348, 271, 210, 252, 
    301, 359, 417, 389, 328, 222, 143, 114, 125, 165, 202, 218, 231, 236, 246, 246, 239, 223, 211, 190, 196, 224, 259, 313, 349, 359, 347, 259, 247, 237, 
    321, 360, 421, 410, 387, 314, 212, 140, 112, 113, 131, 164, 194, 199, 208, 235, 272, 266, 262, 257, 259, 261, 263, 284, 296, 294, 268, 246, 221, 205, 
    355, 364, 404, 397, 411, 381, 307, 215, 149, 119, 104, 107, 136, 152, 165, 197, 251, 284, 304, 278, 270, 250, 221, 214, 206, 215, 209, 201, 162, 178, 
    
    -- channel=5
    383, 411, 407, 416, 428, 431, 435, 427, 441, 449, 460, 464, 472, 467, 445, 431, 431, 449, 450, 446, 438, 436, 438, 434, 434, 432, 417, 413, 417, 427, 
    357, 377, 380, 413, 425, 423, 419, 417, 438, 441, 452, 463, 471, 470, 465, 460, 466, 474, 469, 458, 445, 439, 433, 426, 425, 417, 416, 422, 421, 417, 
    348, 355, 379, 411, 423, 422, 411, 417, 428, 426, 442, 459, 472, 475, 471, 464, 473, 476, 470, 462, 448, 445, 440, 430, 419, 413, 420, 426, 427, 424, 
    343, 347, 375, 399, 417, 420, 413, 413, 415, 422, 432, 444, 465, 474, 472, 471, 460, 457, 445, 438, 432, 434, 430, 432, 428, 422, 423, 425, 423, 415, 
    340, 340, 371, 382, 400, 412, 409, 406, 401, 412, 424, 435, 449, 463, 469, 473, 449, 429, 416, 416, 424, 434, 436, 442, 440, 441, 434, 428, 419, 409, 
    327, 348, 364, 371, 394, 398, 397, 396, 389, 406, 421, 436, 436, 450, 456, 453, 436, 422, 416, 426, 428, 442, 443, 448, 455, 454, 447, 433, 418, 411, 
    321, 360, 353, 374, 389, 394, 394, 388, 389, 414, 427, 433, 431, 448, 451, 450, 438, 428, 418, 430, 418, 440, 444, 449, 452, 446, 443, 430, 418, 412, 
    345, 350, 351, 371, 381, 397, 395, 393, 391, 407, 418, 418, 413, 420, 423, 426, 429, 435, 428, 434, 415, 421, 427, 439, 447, 444, 434, 421, 420, 412, 
    353, 350, 356, 360, 376, 388, 385, 389, 398, 413, 402, 381, 369, 360, 362, 375, 407, 432, 434, 423, 402, 402, 420, 431, 448, 441, 432, 423, 418, 410, 
    377, 385, 368, 367, 376, 378, 382, 392, 403, 399, 346, 300, 296, 298, 302, 322, 377, 409, 414, 403, 398, 412, 429, 434, 448, 437, 437, 432, 424, 417, 
    407, 377, 327, 332, 348, 354, 359, 380, 388, 377, 304, 249, 236, 268, 314, 337, 377, 390, 383, 373, 382, 408, 429, 452, 452, 451, 450, 438, 428, 421, 
    416, 369, 321, 323, 309, 310, 334, 365, 365, 341, 268, 224, 224, 261, 296, 313, 355, 347, 336, 344, 364, 412, 439, 449, 448, 455, 454, 444, 437, 429, 
    402, 363, 318, 293, 272, 285, 307, 320, 316, 294, 252, 252, 274, 284, 284, 262, 288, 270, 272, 306, 340, 396, 420, 435, 442, 447, 451, 444, 438, 435, 
    402, 365, 327, 279, 264, 282, 296, 292, 273, 245, 229, 266, 299, 282, 245, 216, 214, 208, 232, 257, 316, 377, 406, 431, 431, 425, 424, 426, 435, 438, 
    401, 386, 337, 283, 270, 294, 294, 277, 232, 215, 227, 281, 304, 276, 225, 190, 190, 196, 202, 228, 303, 363, 414, 436, 426, 409, 386, 392, 417, 437, 
    405, 370, 318, 273, 256, 295, 299, 265, 236, 239, 243, 273, 289, 293, 270, 233, 230, 234, 247, 275, 331, 386, 442, 455, 440, 404, 353, 361, 392, 430, 
    407, 371, 308, 256, 243, 293, 317, 275, 258, 236, 250, 275, 306, 327, 341, 321, 320, 319, 335, 359, 400, 439, 471, 470, 444, 393, 332, 320, 371, 417, 
    414, 375, 314, 239, 203, 254, 332, 306, 284, 251, 274, 285, 301, 305, 343, 338, 376, 390, 402, 427, 445, 467, 481, 465, 443, 386, 317, 274, 336, 402, 
    395, 370, 314, 228, 185, 230, 347, 368, 364, 315, 282, 298, 339, 349, 353, 335, 385, 437, 441, 448, 448, 458, 470, 462, 449, 384, 300, 236, 286, 371, 
    389, 380, 318, 235, 196, 243, 365, 416, 428, 407, 368, 366, 396, 393, 374, 372, 405, 452, 464, 465, 450, 441, 453, 451, 449, 396, 300, 213, 256, 352, 
    374, 370, 331, 268, 231, 280, 377, 429, 446, 430, 427, 429, 440, 425, 419, 429, 452, 481, 477, 472, 467, 463, 467, 459, 451, 410, 321, 234, 252, 345, 
    369, 370, 351, 297, 270, 302, 363, 425, 445, 433, 431, 431, 434, 444, 464, 473, 489, 505, 496, 485, 486, 487, 489, 482, 456, 430, 361, 287, 271, 349, 
    379, 375, 355, 325, 296, 288, 334, 402, 416, 434, 435, 433, 432, 442, 445, 466, 486, 492, 494, 490, 489, 487, 490, 480, 458, 456, 416, 359, 318, 345, 
    387, 385, 364, 347, 331, 315, 307, 344, 369, 405, 405, 417, 418, 421, 434, 454, 463, 476, 480, 482, 484, 487, 489, 477, 469, 471, 451, 429, 381, 359, 
    398, 380, 357, 350, 341, 341, 321, 349, 378, 407, 405, 399, 403, 409, 419, 430, 434, 446, 448, 453, 462, 462, 465, 463, 463, 463, 451, 428, 399, 383, 
    395, 392, 370, 359, 351, 361, 348, 352, 350, 372, 412, 401, 391, 387, 407, 423, 422, 418, 421, 433, 442, 439, 437, 433, 433, 445, 443, 414, 404, 380, 
    390, 386, 373, 367, 364, 390, 381, 375, 382, 375, 402, 391, 380, 378, 401, 409, 408, 406, 408, 416, 427, 424, 417, 413, 422, 431, 431, 418, 409, 390, 
    388, 370, 372, 369, 367, 386, 385, 373, 365, 383, 397, 386, 388, 387, 399, 406, 409, 410, 409, 421, 426, 416, 405, 402, 409, 414, 425, 419, 405, 399, 
    385, 368, 369, 363, 379, 387, 380, 376, 363, 364, 376, 390, 407, 408, 410, 416, 414, 417, 422, 429, 424, 413, 400, 398, 396, 405, 418, 427, 419, 391, 
    382, 367, 371, 384, 398, 394, 379, 382, 382, 384, 389, 400, 414, 421, 425, 431, 423, 425, 422, 415, 413, 404, 392, 391, 390, 396, 400, 407, 397, 384, 
    
    -- channel=6
    729, 748, 754, 762, 777, 789, 792, 791, 783, 773, 761, 751, 747, 744, 736, 728, 698, 636, 603, 618, 632, 627, 598, 555, 503, 482, 511, 559, 599, 615, 
    772, 772, 757, 758, 768, 779, 777, 771, 760, 749, 736, 726, 724, 721, 713, 704, 685, 658, 643, 646, 646, 631, 583, 524, 467, 469, 509, 568, 611, 624, 
    755, 742, 728, 733, 739, 753, 747, 738, 726, 715, 702, 696, 695, 693, 686, 677, 666, 656, 649, 630, 595, 573, 542, 503, 475, 483, 521, 574, 612, 623, 
    705, 700, 695, 702, 711, 721, 715, 706, 695, 683, 673, 669, 671, 671, 664, 656, 650, 649, 641, 585, 518, 471, 458, 482, 494, 497, 528, 565, 601, 608, 
    665, 659, 666, 677, 685, 688, 683, 679, 672, 661, 653, 651, 655, 655, 651, 645, 641, 644, 626, 548, 461, 391, 401, 456, 487, 514, 543, 573, 600, 603, 
    647, 652, 658, 662, 660, 661, 661, 662, 658, 651, 645, 642, 646, 645, 643, 634, 625, 624, 597, 517, 424, 372, 405, 462, 500, 541, 569, 591, 610, 616, 
    645, 648, 650, 649, 644, 645, 646, 650, 650, 647, 639, 626, 620, 611, 613, 608, 604, 602, 568, 496, 422, 406, 444, 494, 543, 580, 604, 616, 628, 630, 
    638, 646, 647, 647, 642, 642, 641, 644, 642, 633, 617, 594, 587, 580, 592, 593, 584, 570, 530, 462, 404, 412, 460, 520, 579, 616, 629, 630, 631, 628, 
    632, 644, 648, 649, 644, 644, 642, 640, 633, 618, 603, 564, 543, 524, 514, 483, 435, 387, 366, 333, 332, 375, 431, 494, 550, 592, 618, 624, 624, 620, 
    634, 644, 646, 646, 643, 643, 642, 637, 627, 601, 548, 452, 384, 336, 313, 289, 247, 203, 179, 125, 154, 259, 378, 475, 482, 514, 568, 608, 617, 613, 
    641, 644, 642, 642, 640, 639, 639, 630, 594, 521, 435, 345, 281, 239, 225, 212, 183, 158, 124, 43, 25, 120, 292, 440, 447, 455, 496, 563, 604, 609, 
    645, 642, 637, 637, 637, 636, 632, 593, 527, 456, 380, 284, 218, 203, 222, 232, 243, 245, 177, 48, 0, 0, 204, 386, 439, 425, 456, 508, 578, 602, 
    642, 639, 634, 634, 635, 630, 604, 543, 481, 402, 323, 263, 248, 270, 333, 367, 389, 354, 231, 63, 0, 0, 87, 285, 414, 430, 438, 472, 538, 584, 
    636, 637, 634, 626, 598, 574, 535, 491, 410, 353, 331, 318, 317, 344, 400, 404, 375, 273, 144, 0, 0, 0, 7, 188, 352, 429, 428, 424, 454, 521, 
    632, 635, 628, 603, 539, 488, 432, 380, 344, 361, 356, 335, 299, 258, 240, 197, 149, 77, 0, 0, 0, 0, 43, 192, 355, 426, 420, 351, 332, 414, 
    630, 631, 613, 575, 497, 423, 346, 306, 335, 348, 370, 362, 278, 167, 85, 13, 0, 0, 0, 0, 0, 0, 143, 291, 393, 391, 347, 258, 192, 290, 
    630, 617, 557, 492, 409, 350, 309, 303, 320, 356, 369, 356, 241, 107, 0, 0, 0, 0, 0, 0, 0, 21, 223, 343, 332, 290, 230, 150, 82, 211, 
    624, 547, 425, 362, 321, 327, 310, 320, 351, 408, 386, 349, 202, 43, 0, 0, 0, 0, 0, 0, 0, 0, 141, 222, 206, 151, 98, 55, 53, 197, 
    582, 421, 265, 184, 206, 286, 316, 356, 395, 443, 415, 352, 179, 18, 0, 0, 0, 0, 0, 0, 0, 0, 1, 36, 32, 3, 4, 30, 97, 234, 
    526, 347, 145, 52, 152, 258, 333, 387, 427, 461, 413, 330, 161, 13, 0, 0, 0, 11, 98, 170, 155, 60, 0, 0, 0, 0, 8, 83, 190, 310, 
    504, 350, 146, 85, 158, 233, 341, 400, 449, 432, 356, 268, 117, 0, 0, 0, 0, 105, 240, 323, 306, 203, 74, 0, 0, 0, 75, 182, 290, 405, 
    502, 359, 215, 164, 176, 226, 353, 418, 447, 389, 311, 208, 60, 0, 0, 0, 55, 197, 362, 393, 384, 325, 191, 66, 0, 45, 158, 268, 391, 465, 
    515, 397, 300, 199, 180, 221, 345, 414, 410, 331, 249, 132, 22, 0, 0, 0, 98, 250, 360, 356, 383, 392, 291, 163, 63, 93, 216, 350, 454, 478, 
    520, 411, 312, 196, 176, 225, 341, 391, 350, 260, 187, 102, 23, 0, 0, 0, 122, 263, 337, 335, 356, 392, 358, 239, 137, 147, 271, 410, 482, 486, 
    509, 404, 304, 199, 166, 198, 278, 298, 224, 128, 67, 15, 0, 0, 0, 0, 124, 251, 295, 269, 292, 360, 387, 306, 227, 230, 335, 447, 492, 492, 
    502, 404, 311, 213, 182, 210, 261, 273, 209, 139, 95, 59, 28, 9, 3, 47, 164, 252, 296, 274, 297, 348, 409, 380, 346, 343, 406, 474, 495, 490, 
    497, 431, 362, 284, 267, 286, 320, 318, 273, 234, 211, 199, 189, 182, 182, 210, 286, 309, 306, 265, 286, 349, 423, 437, 427, 432, 467, 488, 487, 475, 
    486, 443, 395, 357, 340, 348, 369, 373, 362, 352, 345, 340, 336, 338, 344, 361, 397, 397, 362, 300, 310, 385, 435, 476, 482, 486, 492, 489, 477, 461, 
    467, 434, 388, 353, 337, 345, 368, 385, 394, 391, 386, 390, 396, 404, 414, 429, 448, 439, 398, 370, 368, 399, 454, 488, 491, 490, 489, 483, 467, 453, 
    427, 380, 317, 271, 250, 256, 282, 304, 321, 319, 311, 317, 328, 342, 357, 377, 402, 410, 385, 353, 363, 410, 460, 473, 469, 469, 467, 460, 446, 438, 
    
    -- channel=7
    266, 273, 280, 284, 275, 271, 270, 285, 308, 323, 324, 317, 316, 313, 312, 317, 327, 334, 347, 353, 360, 369, 380, 392, 402, 407, 407, 409, 411, 417, 
    266, 271, 282, 285, 286, 298, 296, 314, 333, 347, 349, 338, 337, 344, 347, 342, 338, 343, 357, 369, 378, 382, 386, 391, 391, 389, 387, 387, 389, 393, 
    270, 273, 285, 288, 297, 316, 323, 356, 368, 386, 396, 387, 384, 386, 383, 374, 359, 353, 354, 363, 367, 369, 370, 371, 368, 363, 357, 357, 361, 369, 
    277, 278, 287, 296, 310, 331, 352, 381, 396, 423, 435, 433, 439, 445, 437, 411, 365, 338, 328, 335, 341, 342, 342, 342, 338, 335, 335, 343, 355, 369, 
    289, 289, 295, 311, 342, 371, 387, 402, 428, 457, 471, 479, 482, 483, 478, 451, 393, 336, 305, 304, 312, 313, 319, 324, 328, 331, 335, 348, 366, 383, 
    302, 301, 305, 325, 360, 397, 424, 446, 461, 482, 495, 504, 507, 511, 501, 477, 433, 370, 318, 292, 297, 312, 324, 327, 327, 328, 336, 355, 377, 397, 
    310, 304, 300, 299, 331, 395, 439, 470, 474, 476, 479, 485, 493, 501, 502, 496, 467, 425, 376, 340, 327, 331, 337, 337, 331, 330, 344, 366, 386, 400, 
    284, 266, 248, 233, 278, 359, 425, 481, 479, 463, 448, 438, 445, 463, 481, 501, 498, 475, 438, 405, 379, 369, 364, 349, 339, 336, 349, 366, 380, 393, 
    222, 200, 178, 161, 218, 313, 413, 479, 479, 451, 420, 393, 394, 421, 459, 491, 500, 497, 487, 470, 448, 422, 399, 365, 344, 341, 355, 369, 377, 385, 
    159, 136, 117, 103, 173, 291, 407, 463, 459, 435, 406, 382, 375, 401, 439, 474, 487, 495, 507, 505, 492, 464, 432, 393, 364, 354, 356, 360, 364, 370, 
    111, 101, 95, 92, 153, 277, 384, 437, 426, 408, 386, 373, 369, 400, 431, 448, 460, 473, 495, 508, 507, 487, 454, 417, 385, 364, 352, 350, 354, 362, 
    105, 105, 104, 106, 141, 249, 356, 421, 416, 394, 371, 365, 375, 404, 432, 432, 433, 438, 465, 488, 500, 495, 467, 436, 399, 375, 355, 345, 349, 359, 
    117, 118, 120, 121, 133, 197, 287, 362, 413, 415, 396, 390, 403, 420, 438, 424, 406, 404, 431, 461, 487, 496, 476, 446, 413, 384, 363, 347, 352, 364, 
    132, 132, 129, 124, 130, 164, 221, 284, 360, 398, 402, 399, 409, 434, 442, 415, 384, 374, 398, 438, 475, 495, 487, 452, 426, 397, 382, 362, 356, 365, 
    138, 131, 123, 121, 137, 172, 197, 242, 281, 334, 366, 380, 394, 428, 441, 414, 377, 358, 381, 422, 464, 489, 491, 458, 435, 407, 386, 369, 366, 380, 
    137, 128, 116, 101, 102, 150, 160, 177, 203, 260, 306, 315, 348, 392, 424, 410, 373, 354, 372, 410, 449, 475, 485, 464, 440, 415, 394, 388, 392, 417, 
    112, 88, 55, 22, 10, 63, 113, 141, 152, 157, 245, 258, 321, 362, 406, 412, 377, 358, 368, 397, 430, 455, 474, 466, 443, 425, 412, 418, 429, 453, 
    31, 0, 0, 0, 0, 0, 29, 80, 139, 128, 213, 240, 307, 348, 394, 410, 383, 361, 365, 384, 408, 434, 459, 467, 449, 440, 434, 448, 466, 488, 
    0, 0, 0, 0, 0, 0, 30, 92, 160, 168, 222, 255, 312, 360, 390, 405, 385, 364, 364, 377, 395, 424, 452, 468, 456, 447, 452, 473, 488, 494, 
    0, 0, 0, 0, 0, 74, 134, 179, 229, 242, 272, 316, 352, 382, 399, 406, 390, 373, 369, 378, 400, 429, 458, 474, 464, 447, 451, 468, 482, 486, 
    0, 0, 0, 0, 81, 179, 231, 279, 323, 335, 358, 386, 401, 414, 421, 420, 403, 392, 390, 395, 408, 428, 452, 468, 467, 446, 437, 448, 469, 484, 
    0, 0, 0, 41, 144, 226, 272, 323, 381, 421, 444, 436, 409, 408, 430, 449, 439, 425, 412, 401, 403, 420, 443, 464, 469, 448, 428, 433, 455, 481, 
    0, 5, 44, 110, 180, 223, 257, 305, 378, 452, 478, 447, 402, 388, 400, 429, 441, 431, 417, 397, 383, 385, 407, 446, 469, 465, 437, 425, 440, 468, 
    91, 130, 163, 189, 206, 221, 243, 283, 333, 388, 428, 425, 397, 379, 400, 423, 436, 428, 400, 362, 340, 350, 385, 424, 457, 472, 455, 432, 431, 451, 
    211, 224, 226, 229, 237, 254, 267, 288, 320, 357, 395, 416, 409, 394, 403, 415, 424, 417, 379, 335, 312, 329, 375, 419, 452, 465, 469, 447, 432, 439, 
    262, 261, 262, 271, 279, 292, 310, 333, 347, 358, 380, 404, 425, 422, 419, 425, 431, 427, 392, 347, 321, 337, 382, 417, 449, 470, 481, 469, 445, 438, 
    291, 297, 301, 311, 329, 352, 378, 402, 409, 403, 404, 415, 421, 428, 436, 452, 461, 453, 427, 392, 369, 371, 397, 426, 455, 478, 492, 491, 469, 450, 
    317, 331, 348, 369, 392, 416, 442, 464, 461, 436, 413, 412, 422, 442, 451, 478, 487, 478, 464, 445, 431, 424, 431, 447, 469, 491, 507, 506, 491, 470, 
    361, 386, 410, 432, 450, 469, 482, 494, 480, 451, 423, 414, 432, 454, 477, 503, 504, 496, 491, 486, 478, 472, 469, 474, 490, 509, 520, 516, 506, 490, 
    417, 444, 466, 484, 493, 497, 496, 501, 488, 463, 441, 426, 443, 465, 499, 518, 520, 515, 508, 504, 499, 497, 496, 501, 511, 521, 528, 524, 514, 503, 
    
    -- channel=8
    441, 447, 387, 318, 265, 247, 233, 217, 233, 257, 264, 257, 254, 249, 235, 214, 209, 248, 302, 314, 256, 201, 165, 179, 198, 202, 204, 207, 215, 225, 
    440, 451, 403, 329, 277, 246, 211, 166, 162, 193, 215, 211, 198, 191, 178, 155, 154, 197, 259, 272, 222, 156, 119, 143, 162, 172, 178, 184, 192, 202, 
    441, 448, 416, 345, 303, 264, 208, 130, 87, 123, 166, 192, 187, 171, 155, 137, 137, 173, 233, 236, 177, 101, 73, 94, 114, 131, 146, 157, 167, 179, 
    439, 441, 426, 364, 330, 286, 219, 116, 36, 56, 121, 176, 203, 195, 181, 164, 167, 186, 211, 186, 133, 70, 56, 64, 73, 83, 93, 102, 112, 126, 
    443, 441, 432, 372, 323, 274, 209, 104, 17, 12, 82, 169, 221, 228, 226, 209, 211, 207, 185, 123, 73, 39, 36, 30, 29, 28, 35, 43, 52, 62, 
    427, 442, 403, 317, 259, 229, 188, 101, 17, 0, 43, 128, 193, 230, 241, 232, 240, 216, 161, 86, 41, 23, 9, 0, 0, 0, 0, 0, 10, 8, 
    310, 346, 312, 247, 176, 164, 177, 124, 41, 0, 18, 75, 131, 179, 211, 225, 237, 215, 151, 71, 31, 11, 0, 0, 0, 0, 0, 1, 9, 0, 
    210, 229, 211, 147, 90, 130, 179, 146, 77, 14, 7, 33, 77, 125, 188, 217, 223, 207, 149, 76, 35, 4, 0, 0, 0, 0, 2, 45, 47, 3, 
    121, 137, 116, 72, 67, 131, 178, 158, 90, 24, 6, 20, 57, 112, 172, 197, 214, 197, 150, 96, 50, 12, 0, 0, 0, 0, 36, 87, 84, 33, 
    73, 79, 69, 53, 62, 121, 162, 149, 77, 21, 10, 29, 71, 133, 181, 196, 195, 183, 145, 102, 59, 18, 0, 0, 0, 0, 46, 101, 113, 76, 
    65, 69, 62, 58, 70, 113, 147, 133, 74, 34, 28, 45, 83, 143, 177, 171, 163, 148, 127, 95, 62, 19, 0, 0, 0, 0, 25, 86, 119, 104, 
    68, 76, 72, 86, 106, 122, 138, 122, 100, 83, 63, 69, 104, 137, 145, 128, 122, 108, 110, 86, 61, 24, 0, 0, 0, 0, 0, 49, 92, 93, 
    74, 86, 83, 119, 148, 144, 133, 87, 82, 77, 65, 67, 92, 135, 133, 100, 86, 93, 89, 65, 56, 22, 0, 0, 0, 0, 0, 3, 40, 55, 
    75, 89, 85, 128, 176, 161, 124, 60, 63, 65, 65, 59, 66, 95, 107, 98, 83, 95, 86, 75, 64, 45, 7, 0, 0, 0, 0, 0, 0, 9, 
    79, 100, 96, 124, 184, 167, 113, 34, 31, 40, 39, 42, 59, 82, 118, 119, 116, 120, 110, 103, 90, 121, 118, 59, 0, 0, 0, 0, 0, 0, 
    85, 115, 120, 121, 153, 141, 92, 17, 0, 0, 12, 28, 39, 62, 119, 145, 158, 160, 131, 113, 112, 151, 191, 180, 106, 34, 19, 17, 7, 0, 
    80, 117, 127, 110, 111, 106, 66, 16, 0, 0, 0, 0, 2, 29, 95, 173, 190, 196, 156, 137, 141, 170, 231, 234, 186, 132, 110, 98, 61, 11, 
    63, 102, 108, 88, 63, 55, 44, 20, 0, 0, 0, 0, 0, 0, 57, 145, 185, 197, 160, 138, 151, 179, 239, 249, 213, 180, 164, 154, 132, 79, 
    40, 80, 84, 63, 35, 30, 34, 21, 10, 0, 0, 0, 0, 0, 2, 69, 129, 151, 157, 146, 169, 198, 222, 215, 199, 185, 184, 187, 177, 143, 
    20, 53, 65, 50, 25, 17, 23, 25, 12, 18, 32, 23, 16, 3, 1, 27, 73, 106, 148, 162, 193, 210, 206, 183, 172, 167, 179, 196, 205, 197, 
    8, 34, 60, 50, 26, 6, 4, 10, 7, 20, 51, 66, 61, 32, 18, 16, 44, 95, 158, 194, 216, 207, 181, 156, 145, 153, 179, 206, 223, 234, 
    7, 26, 61, 56, 30, 0, 0, 0, 0, 12, 54, 75, 71, 52, 36, 29, 47, 109, 179, 218, 223, 191, 161, 134, 131, 147, 174, 206, 221, 239, 
    14, 30, 66, 62, 33, 0, 0, 0, 0, 40, 77, 82, 67, 54, 49, 50, 70, 129, 193, 230, 216, 184, 165, 143, 137, 140, 175, 202, 219, 243, 
    25, 45, 77, 76, 40, 0, 0, 0, 26, 105, 132, 117, 74, 58, 67, 76, 100, 150, 210, 229, 210, 187, 176, 163, 156, 159, 182, 199, 227, 245, 
    35, 63, 96, 104, 59, 0, 0, 0, 50, 144, 183, 159, 98, 81, 98, 114, 137, 183, 226, 229, 217, 202, 196, 192, 191, 198, 203, 208, 214, 222, 
    45, 82, 119, 133, 89, 19, 0, 0, 54, 139, 174, 161, 119, 117, 144, 164, 183, 225, 247, 246, 230, 217, 212, 219, 223, 234, 233, 216, 202, 212, 
    60, 98, 140, 163, 116, 34, 0, 0, 38, 104, 138, 140, 135, 159, 183, 199, 224, 262, 265, 263, 237, 224, 224, 234, 249, 260, 244, 215, 200, 203, 
    86, 114, 153, 184, 141, 52, 0, 0, 21, 66, 97, 122, 160, 191, 214, 230, 259, 287, 286, 277, 245, 235, 230, 240, 254, 258, 245, 221, 204, 206, 
    121, 135, 161, 195, 166, 78, 0, 0, 11, 42, 89, 151, 208, 237, 245, 251, 280, 295, 296, 275, 250, 239, 234, 237, 244, 251, 246, 229, 215, 214, 
    170, 177, 183, 217, 198, 117, 34, 4, 25, 63, 125, 196, 269, 300, 293, 288, 293, 297, 295, 274, 260, 247, 237, 235, 252, 258, 250, 234, 224, 219, 
    
    -- channel=9
    0, 0, 0, 0, 0, 0, 21, 51, 43, 25, 20, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 6, 20, 
    0, 0, 0, 0, 0, 0, 9, 44, 41, 13, 9, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 27, 63, 59, 29, 32, 27, 30, 29, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 40, 72, 54, 16, 12, 8, 10, 17, 18, 24, 22, 25, 48, 43, 6, 0, 0, 0, 0, 0, 25, 51, 19, 0, 
    0, 0, 0, 0, 0, 0, 40, 52, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 39, 21, 0, 0, 0, 0, 0, 53, 80, 57, 0, 
    0, 0, 0, 0, 0, 0, 26, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 77, 83, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 78, 96, 56, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 50, 29, 
    0, 0, 0, 0, 0, 0, 21, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 43, 63, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 45, 104, 94, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 17, 35, 48, 83, 83, 50, 0, 0, 0, 0, 20, 15, 0, 0, 0, 0, 22, 42, 27, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 45, 65, 72, 65, 76, 40, 14, 0, 0, 0, 13, 49, 55, 42, 16, 17, 51, 96, 117, 91, 45, 0, 0, 0, 0, 0, 0, 
    0, 24, 77, 119, 92, 73, 74, 46, 13, 36, 69, 76, 75, 84, 103, 100, 84, 66, 77, 117, 152, 158, 137, 114, 78, 45, 0, 0, 0, 0, 
    14, 75, 135, 167, 125, 97, 85, 51, 50, 52, 84, 115, 123, 140, 176, 204, 220, 222, 210, 210, 229, 240, 236, 200, 129, 75, 26, 0, 0, 0, 
    2, 91, 146, 172, 133, 132, 123, 110, 96, 100, 107, 117, 103, 132, 175, 205, 225, 229, 191, 175, 183, 203, 236, 201, 137, 59, 0, 0, 0, 0, 
    0, 85, 137, 161, 140, 176, 186, 180, 126, 123, 127, 110, 66, 93, 101, 132, 149, 142, 107, 92, 89, 113, 157, 125, 74, 33, 17, 4, 0, 0, 
    0, 49, 127, 164, 167, 209, 244, 238, 171, 149, 158, 160, 145, 128, 75, 89, 77, 78, 58, 31, 42, 76, 94, 50, 28, 32, 55, 55, 0, 0, 
    0, 44, 141, 199, 211, 233, 271, 267, 207, 186, 200, 212, 194, 178, 131, 73, 19, 32, 41, 34, 35, 47, 51, 31, 42, 61, 102, 113, 9, 0, 
    0, 30, 120, 207, 236, 250, 269, 285, 270, 260, 234, 219, 199, 202, 175, 145, 122, 116, 117, 112, 123, 115, 114, 112, 101, 106, 112, 110, 18, 0, 
    0, 26, 117, 200, 231, 245, 256, 288, 311, 314, 262, 217, 145, 161, 201, 201, 144, 107, 105, 112, 125, 94, 72, 109, 138, 136, 106, 94, 18, 0, 
    0, 27, 135, 215, 229, 195, 211, 259, 312, 347, 319, 279, 193, 199, 231, 258, 207, 149, 113, 115, 126, 88, 80, 142, 178, 209, 172, 126, 41, 0, 
    0, 28, 157, 248, 246, 163, 150, 201, 275, 346, 349, 318, 269, 265, 288, 311, 264, 194, 136, 114, 98, 73, 98, 158, 220, 254, 222, 190, 87, 0, 
    0, 0, 114, 212, 210, 142, 114, 140, 240, 322, 359, 367, 351, 338, 346, 349, 282, 163, 76, 8, 0, 0, 59, 161, 277, 306, 279, 234, 99, 0, 
    0, 0, 28, 116, 150, 98, 95, 117, 206, 280, 347, 386, 396, 388, 372, 361, 317, 210, 102, 0, 0, 0, 80, 191, 305, 338, 294, 227, 77, 0, 
    0, 0, 0, 22, 71, 70, 107, 118, 182, 246, 319, 373, 394, 384, 363, 337, 294, 204, 103, 14, 0, 0, 79, 211, 332, 352, 291, 205, 56, 0, 
    0, 0, 0, 0, 44, 78, 132, 134, 176, 220, 296, 361, 384, 375, 356, 334, 296, 218, 137, 79, 41, 16, 102, 233, 356, 358, 287, 195, 47, 0, 
    0, 0, 0, 0, 49, 98, 152, 169, 189, 220, 284, 341, 362, 356, 337, 312, 279, 243, 202, 158, 110, 68, 130, 241, 355, 356, 291, 198, 48, 0, 
    0, 0, 0, 0, 28, 113, 175, 206, 211, 235, 279, 318, 329, 324, 312, 301, 282, 256, 226, 191, 154, 117, 156, 253, 337, 348, 289, 177, 31, 0, 
    0, 0, 0, 0, 0, 97, 188, 246, 244, 248, 269, 289, 284, 277, 271, 264, 247, 225, 201, 178, 161, 145, 165, 229, 289, 305, 243, 127, 0, 0, 
    
    
    others => 0);
end gold_package;
