library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 7, 1, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=1
    55, 56, 57, 59, 57, 54, 58, 62, 58, 47, 37, 38, 44, 51, 53, 
    54, 60, 60, 60, 59, 47, 55, 46, 33, 19, 15, 15, 18, 35, 50, 
    35, 34, 58, 61, 59, 45, 26, 21, 18, 9, 17, 16, 15, 17, 35, 
    32, 15, 55, 57, 47, 35, 30, 21, 10, 10, 16, 12, 10, 11, 21, 
    23, 17, 51, 50, 43, 32, 23, 16, 9, 0, 22, 22, 14, 17, 11, 
    7, 3, 47, 30, 0, 14, 19, 26, 19, 0, 17, 14, 13, 16, 15, 
    11, 0, 23, 54, 15, 9, 20, 17, 24, 0, 14, 13, 6, 10, 21, 
    3, 10, 15, 35, 31, 18, 18, 6, 20, 13, 11, 14, 7, 14, 32, 
    2, 0, 5, 2, 19, 4, 15, 13, 15, 18, 14, 11, 6, 26, 46, 
    2, 1, 10, 0, 20, 11, 8, 21, 12, 16, 9, 7, 10, 31, 42, 
    0, 1, 9, 0, 18, 21, 0, 0, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=2
    25, 25, 26, 26, 25, 21, 27, 27, 23, 19, 16, 19, 21, 23, 25, 
    26, 24, 27, 26, 27, 21, 17, 16, 12, 6, 3, 0, 4, 21, 25, 
    10, 26, 26, 26, 26, 9, 5, 0, 10, 14, 10, 15, 11, 11, 25, 
    3, 15, 24, 24, 13, 10, 12, 13, 14, 16, 8, 8, 10, 12, 22, 
    8, 16, 21, 22, 20, 6, 0, 6, 8, 12, 4, 8, 13, 17, 8, 
    0, 6, 20, 3, 0, 2, 6, 9, 9, 20, 0, 3, 13, 14, 14, 
    0, 0, 10, 21, 11, 6, 7, 6, 10, 13, 0, 3, 6, 12, 16, 
    0, 1, 0, 13, 19, 19, 2, 5, 14, 16, 5, 0, 11, 14, 24, 
    0, 0, 0, 12, 1, 0, 1, 5, 15, 0, 3, 6, 10, 25, 29, 
    0, 0, 0, 0, 5, 7, 6, 9, 0, 16, 10, 11, 21, 25, 18, 
    0, 0, 0, 11, 12, 9, 12, 4, 7, 0, 2, 10, 0, 0, 0, 
    0, 0, 9, 5, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 6, 5, 0, 0, 0, 4, 0, 0, 
    
    -- channel=3
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 11, 5, 0, 0, 0, 0, 
    0, 7, 0, 0, 0, 0, 0, 0, 3, 16, 0, 4, 0, 1, 0, 
    0, 10, 0, 0, 0, 0, 0, 0, 2, 16, 1, 0, 2, 0, 7, 
    13, 8, 0, 0, 14, 0, 0, 0, 0, 32, 0, 0, 7, 0, 0, 
    9, 8, 0, 0, 9, 5, 0, 0, 0, 31, 0, 1, 9, 9, 0, 
    12, 0, 6, 0, 4, 13, 0, 0, 0, 15, 0, 1, 12, 2, 0, 
    10, 16, 3, 4, 1, 5, 0, 5, 4, 0, 13, 0, 7, 0, 0, 
    8, 17, 0, 26, 2, 2, 5, 0, 14, 0, 0, 5, 7, 0, 0, 
    25, 14, 0, 38, 0, 14, 22, 4, 0, 5, 25, 26, 32, 28, 25, 
    56, 20, 1, 33, 10, 25, 40, 37, 34, 36, 38, 42, 43, 46, 43, 
    48, 53, 28, 20, 9, 35, 35, 35, 37, 41, 45, 47, 45, 45, 49, 
    48, 47, 65, 0, 25, 39, 35, 38, 39, 43, 49, 49, 46, 59, 49, 
    44, 49, 48, 36, 38, 44, 38, 33, 38, 41, 44, 45, 50, 50, 37, 
    
    -- channel=4
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=5
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 13, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 0, 0, 2, 
    0, 15, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 
    0, 16, 0, 0, 43, 0, 0, 0, 0, 54, 0, 0, 0, 0, 0, 
    0, 10, 0, 0, 29, 9, 9, 0, 0, 62, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 45, 0, 0, 0, 38, 0, 0, 0, 0, 0, 
    0, 20, 0, 10, 0, 3, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    11, 18, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    45, 12, 0, 55, 0, 0, 36, 14, 0, 0, 0, 0, 6, 7, 0, 
    60, 34, 0, 72, 3, 0, 13, 9, 0, 4, 9, 13, 13, 16, 9, 
    10, 49, 31, 38, 0, 5, 6, 6, 5, 8, 14, 15, 19, 18, 18, 
    7, 15, 66, 10, 0, 11, 1, 6, 10, 13, 17, 20, 13, 26, 26, 
    5, 18, 20, 18, 2, 17, 15, 7, 12, 11, 8, 12, 27, 18, 0, 
    
    -- channel=6
    2, 0, 1, 4, 3, 0, 2, 3, 3, 4, 5, 0, 2, 6, 8, 
    1, 0, 0, 5, 0, 0, 22, 4, 16, 0, 6, 3, 0, 0, 4, 
    9, 0, 1, 4, 0, 0, 26, 10, 0, 0, 8, 7, 20, 0, 0, 
    51, 0, 3, 0, 6, 0, 1, 18, 4, 0, 26, 0, 18, 15, 0, 
    57, 0, 32, 0, 0, 16, 25, 24, 9, 0, 1, 36, 0, 22, 0, 
    48, 0, 42, 4, 0, 16, 17, 19, 28, 0, 36, 43, 0, 13, 18, 
    50, 0, 9, 30, 0, 0, 0, 25, 34, 0, 44, 25, 0, 0, 17, 
    34, 4, 27, 17, 0, 0, 50, 0, 23, 0, 22, 26, 0, 0, 11, 
    27, 0, 64, 0, 19, 0, 9, 0, 0, 9, 0, 36, 0, 0, 0, 
    0, 0, 56, 0, 27, 11, 0, 0, 8, 5, 34, 3, 0, 0, 8, 
    0, 0, 49, 0, 56, 19, 0, 3, 46, 22, 0, 0, 0, 0, 6, 
    0, 0, 21, 0, 52, 32, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 75, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 18, 18, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 
    
    -- channel=7
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=8
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=9
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 14, 8, 9, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 8, 9, 0, 1, 2, 4, 0, 0, 
    27, 7, 0, 0, 0, 9, 1, 3, 4, 1, 4, 8, 3, 6, 0, 
    35, 7, 0, 0, 0, 0, 0, 3, 7, 3, 12, 5, 3, 9, 7, 
    33, 20, 0, 0, 0, 0, 1, 6, 6, 10, 13, 9, 9, 10, 4, 
    32, 20, 12, 0, 0, 0, 8, 0, 0, 0, 6, 7, 7, 1, 0, 
    35, 30, 30, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    19, 29, 25, 25, 9, 3, 1, 16, 12, 0, 2, 6, 1, 0, 0, 
    20, 23, 25, 19, 45, 37, 34, 23, 25, 23, 33, 46, 47, 32, 32, 
    53, 31, 28, 29, 42, 41, 46, 46, 52, 59, 65, 69, 74, 76, 75, 
    89, 51, 28, 30, 42, 62, 64, 61, 64, 69, 76, 78, 77, 79, 84, 
    91, 78, 50, 31, 55, 66, 68, 64, 67, 72, 82, 80, 84, 89, 89, 
    91, 83, 76, 46, 62, 62, 63, 63, 70, 75, 79, 77, 83, 95, 87, 
    
    -- channel=10
    31, 33, 31, 28, 29, 28, 33, 35, 31, 30, 27, 31, 23, 19, 21, 
    28, 31, 34, 30, 33, 19, 8, 31, 31, 15, 0, 0, 17, 30, 21, 
    26, 54, 32, 31, 36, 69, 11, 6, 0, 16, 0, 0, 0, 12, 31, 
    0, 18, 26, 36, 23, 21, 0, 0, 0, 42, 0, 2, 0, 0, 43, 
    0, 0, 0, 46, 0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 6, 
    0, 12, 0, 26, 84, 8, 0, 0, 0, 57, 0, 0, 5, 0, 0, 
    0, 0, 16, 8, 57, 22, 18, 0, 0, 62, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 24, 57, 0, 14, 0, 51, 0, 0, 7, 5, 0, 
    0, 4, 0, 19, 0, 28, 0, 0, 4, 0, 35, 0, 8, 12, 16, 
    8, 3, 0, 16, 0, 0, 7, 0, 0, 23, 0, 0, 1, 26, 21, 
    44, 0, 0, 41, 0, 0, 15, 13, 0, 0, 0, 0, 0, 5, 0, 
    44, 26, 0, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 26, 23, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 47, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=11
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 3, 19, 14, 7, 0, 0, 
    10, 0, 0, 0, 0, 0, 1, 15, 13, 2, 10, 9, 15, 13, 0, 
    30, 0, 0, 0, 0, 0, 8, 16, 11, 4, 9, 15, 10, 14, 0, 
    40, 12, 0, 0, 1, 11, 9, 9, 11, 3, 16, 20, 10, 14, 14, 
    44, 9, 0, 0, 0, 7, 7, 13, 15, 0, 21, 20, 12, 16, 13, 
    42, 18, 15, 0, 0, 5, 12, 7, 16, 0, 16, 18, 14, 8, 0, 
    37, 25, 40, 8, 13, 0, 10, 11, 8, 0, 13, 11, 8, 0, 0, 
    26, 25, 34, 9, 28, 10, 7, 12, 17, 11, 8, 15, 5, 0, 0, 
    18, 23, 28, 19, 34, 36, 23, 25, 33, 18, 34, 38, 32, 23, 30, 
    38, 31, 31, 2, 36, 56, 41, 44, 53, 49, 53, 53, 59, 57, 63, 
    67, 40, 33, 18, 59, 53, 51, 50, 52, 56, 59, 62, 59, 62, 66, 
    74, 61, 41, 31, 56, 51, 54, 53, 54, 58, 61, 65, 65, 74, 65, 
    71, 66, 56, 39, 52, 55, 55, 53, 53, 56, 62, 60, 63, 68, 70, 
    
    -- channel=12
    19, 15, 17, 17, 18, 11, 21, 27, 20, 10, 6, 8, 8, 13, 14, 
    19, 18, 18, 19, 16, 0, 7, 10, 1, 0, 0, 0, 0, 9, 11, 
    2, 24, 22, 22, 22, 4, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 17, 19, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=13
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    11, 4, 0, 0, 13, 0, 0, 0, 0, 1, 0, 3, 3, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 5, 4, 0, 0, 0, 0, 6, 0, 0, 
    4, 6, 0, 1, 0, 7, 0, 0, 5, 0, 0, 9, 5, 0, 0, 
    7, 7, 0, 3, 1, 2, 4, 0, 0, 5, 6, 7, 0, 0, 0, 
    8, 2, 0, 9, 0, 0, 1, 15, 12, 3, 10, 9, 14, 17, 13, 
    45, 27, 8, 0, 4, 41, 31, 32, 33, 29, 32, 33, 35, 35, 36, 
    39, 40, 31, 0, 41, 30, 28, 29, 30, 32, 36, 35, 36, 39, 40, 
    46, 38, 42, 20, 30, 32, 28, 29, 32, 35, 38, 43, 42, 44, 42, 
    41, 42, 32, 42, 33, 38, 40, 34, 28, 30, 33, 40, 36, 33, 41, 
    
    -- channel=14
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 14, 0, 0, 
    2, 0, 0, 0, 0, 24, 0, 13, 0, 0, 0, 0, 0, 19, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 
    0, 0, 0, 40, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 11, 0, 0, 0, 15, 24, 0, 13, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    50, 0, 0, 0, 0, 0, 41, 33, 0, 0, 0, 0, 0, 0, 0, 
    0, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 19, 20, 11, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 2, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 0, 
    1, 13, 0, 0, 18, 0, 0, 0, 0, 10, 0, 0, 1, 0, 0, 
    0, 24, 0, 0, 28, 0, 15, 0, 0, 35, 0, 0, 0, 0, 0, 
    0, 23, 0, 0, 4, 18, 11, 3, 0, 37, 0, 0, 0, 7, 0, 
    8, 26, 0, 0, 0, 24, 0, 1, 0, 13, 7, 0, 3, 0, 0, 
    22, 33, 0, 21, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    30, 26, 8, 29, 0, 0, 10, 18, 0, 0, 0, 0, 3, 0, 0, 
    50, 21, 5, 51, 38, 5, 36, 28, 9, 3, 11, 26, 26, 19, 12, 
    38, 47, 15, 53, 12, 17, 24, 23, 27, 30, 36, 39, 45, 41, 40, 
    42, 33, 40, 36, 6, 36, 33, 33, 32, 36, 43, 45, 43, 46, 55, 
    46, 43, 36, 45, 28, 36, 35, 32, 38, 41, 45, 45, 47, 57, 47, 
    45, 50, 42, 24, 24, 34, 36, 37, 42, 45, 38, 41, 57, 53, 38, 
    
    -- channel=16
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 16, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 12, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 0, 8, 1, 0, 0, 10, 0, 0, 0, 0, 4, 0, 0, 
    5, 2, 0, 30, 28, 25, 11, 2, 0, 0, 12, 21, 14, 0, 0, 
    19, 8, 16, 19, 0, 0, 0, 3, 14, 19, 27, 27, 34, 34, 33, 
    38, 17, 11, 0, 0, 27, 27, 25, 26, 31, 36, 40, 36, 33, 46, 
    41, 35, 18, 0, 11, 30, 29, 29, 29, 33, 32, 35, 35, 46, 31, 
    40, 41, 24, 16, 14, 22, 25, 30, 35, 37, 35, 36, 50, 49, 41, 
    
    -- channel=17
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 3, 0, 0, 
    7, 11, 0, 0, 0, 11, 18, 10, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 12, 39, 11, 0, 0, 0, 0, 0, 10, 0, 0, 0, 
    0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 12, 14, 4, 0, 5, 1, 0, 0, 0, 
    0, 0, 1, 0, 0, 25, 6, 0, 0, 0, 17, 29, 10, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 20, 18, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 
    15, 9, 0, 0, 32, 61, 28, 27, 12, 0, 0, 0, 0, 0, 0, 
    0, 13, 0, 0, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 30, 10, 0, 0, 0, 0, 0, 0, 1, 0, 0, 9, 
    0, 0, 0, 23, 9, 10, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=18
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 5, 0, 0, 0, 0, 2, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 7, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 23, 14, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 7, 9, 13, 13, 13, 11, 10, 9, 
    13, 0, 0, 0, 0, 10, 10, 14, 17, 18, 16, 11, 3, 4, 4, 
    11, 16, 0, 0, 0, 10, 11, 15, 13, 12, 13, 9, 13, 11, 0, 
    8, 17, 11, 0, 17, 16, 7, 8, 8, 8, 11, 16, 5, 0, 12, 
    
    -- channel=19
    5, 7, 7, 5, 7, 7, 6, 8, 11, 12, 14, 12, 10, 9, 10, 
    7, 7, 8, 5, 6, 0, 10, 14, 24, 13, 6, 11, 14, 7, 6, 
    17, 6, 6, 7, 7, 10, 21, 22, 12, 0, 0, 0, 5, 7, 3, 
    6, 0, 0, 9, 14, 11, 0, 5, 2, 0, 2, 7, 10, 8, 3, 
    0, 0, 1, 7, 0, 1, 4, 8, 8, 5, 0, 5, 1, 3, 14, 
    6, 0, 0, 29, 0, 12, 0, 2, 3, 0, 0, 11, 0, 3, 5, 
    5, 0, 2, 14, 3, 0, 0, 0, 1, 0, 2, 6, 5, 0, 0, 
    3, 0, 2, 0, 1, 0, 3, 6, 0, 0, 2, 7, 2, 0, 0, 
    0, 0, 7, 0, 9, 14, 6, 2, 0, 14, 2, 17, 9, 0, 0, 
    0, 0, 0, 0, 0, 14, 4, 0, 2, 6, 15, 14, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 15, 3, 0, 0, 0, 6, 
    0, 0, 0, 0, 6, 15, 10, 10, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=20
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=21
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=22
    18, 14, 15, 17, 18, 11, 18, 20, 18, 13, 8, 6, 6, 17, 18, 
    17, 14, 17, 17, 14, 0, 19, 10, 3, 0, 0, 1, 4, 3, 13, 
    13, 0, 16, 17, 20, 10, 0, 1, 0, 0, 0, 0, 3, 11, 0, 
    0, 0, 14, 14, 8, 0, 0, 4, 0, 0, 0, 3, 0, 13, 0, 
    0, 0, 18, 0, 0, 0, 0, 0, 5, 0, 0, 3, 0, 1, 23, 
    0, 0, 12, 32, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 8, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 9, 
    0, 0, 2, 0, 10, 0, 0, 0, 0, 4, 0, 6, 1, 0, 16, 
    0, 0, 0, 0, 0, 10, 0, 0, 17, 0, 0, 0, 0, 2, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=23
    4, 7, 2, 6, 5, 3, 6, 4, 3, 8, 7, 2, 4, 6, 6, 
    2, 3, 1, 8, 0, 20, 17, 9, 13, 5, 27, 19, 3, 0, 7, 
    22, 0, 4, 6, 2, 23, 32, 13, 0, 6, 48, 32, 41, 0, 4, 
    71, 0, 13, 0, 19, 0, 38, 23, 25, 0, 61, 26, 37, 20, 0, 
    71, 31, 30, 0, 55, 24, 62, 41, 35, 0, 47, 47, 24, 37, 0, 
    47, 56, 38, 0, 30, 29, 79, 45, 61, 0, 73, 50, 17, 31, 18, 
    36, 96, 19, 41, 0, 10, 76, 52, 67, 0, 79, 45, 18, 19, 35, 
    45, 86, 22, 43, 0, 26, 79, 42, 46, 1, 62, 53, 9, 28, 20, 
    72, 63, 72, 29, 23, 23, 42, 41, 8, 43, 26, 44, 4, 11, 8, 
    68, 59, 102, 14, 60, 0, 1, 73, 25, 29, 45, 8, 0, 4, 15, 
    46, 55, 100, 0, 114, 48, 25, 71, 67, 35, 16, 16, 22, 30, 36, 
    32, 43, 61, 33, 143, 68, 43, 43, 46, 36, 41, 41, 46, 48, 52, 
    62, 20, 0, 111, 94, 43, 45, 41, 42, 39, 41, 45, 53, 48, 48, 
    68, 45, 0, 144, 54, 40, 51, 42, 38, 42, 49, 54, 54, 42, 78, 
    73, 51, 44, 68, 46, 35, 42, 42, 40, 51, 57, 42, 34, 81, 79, 
    
    -- channel=24
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 3, 0, 0, 0, 0, 3, 
    25, 9, 0, 0, 5, 0, 0, 0, 0, 3, 5, 2, 3, 0, 0, 
    24, 6, 0, 0, 0, 0, 0, 0, 0, 7, 3, 3, 5, 0, 2, 
    21, 5, 5, 0, 0, 0, 10, 4, 0, 3, 0, 5, 6, 7, 0, 
    18, 18, 18, 0, 0, 8, 0, 0, 0, 0, 0, 4, 10, 0, 0, 
    12, 20, 6, 13, 6, 8, 0, 0, 20, 0, 0, 0, 0, 0, 0, 
    10, 16, 11, 16, 0, 6, 13, 13, 8, 4, 13, 13, 22, 11, 5, 
    53, 24, 10, 9, 23, 38, 41, 40, 34, 33, 37, 42, 45, 47, 47, 
    55, 53, 27, 15, 34, 38, 39, 39, 39, 41, 44, 48, 48, 47, 50, 
    56, 49, 59, 15, 29, 42, 39, 41, 41, 45, 51, 53, 50, 56, 62, 
    57, 53, 50, 40, 40, 45, 42, 39, 39, 44, 49, 49, 47, 55, 50, 
    
    -- channel=25
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 15, 0, 0, 0, 4, 0, 0, 
    19, 13, 0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 4, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 14, 47, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 11, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 16, 11, 15, 0, 6, 0, 0, 0, 6, 0, 
    0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 23, 17, 8, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 13, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 21, 0, 0, 0, 0, 0, 0, 0, 
    44, 13, 0, 0, 33, 25, 18, 16, 2, 0, 0, 0, 0, 0, 0, 
    0, 34, 0, 13, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 38, 28, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 20, 
    0, 0, 1, 22, 3, 11, 10, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=26
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 9, 3, 0, 0, 11, 20, 14, 9, 2, 0, 
    0, 5, 0, 0, 0, 17, 0, 6, 12, 41, 40, 32, 21, 13, 3, 
    15, 21, 1, 0, 0, 11, 25, 24, 22, 48, 25, 26, 14, 7, 16, 
    41, 57, 9, 27, 54, 51, 35, 19, 15, 33, 42, 23, 24, 13, 13, 
    51, 59, 10, 0, 47, 40, 34, 30, 14, 57, 45, 20, 32, 24, 15, 
    51, 51, 16, 0, 38, 40, 58, 34, 24, 66, 38, 22, 25, 31, 25, 
    54, 58, 39, 15, 36, 73, 43, 32, 20, 49, 31, 21, 31, 33, 12, 
    63, 74, 31, 41, 21, 34, 22, 24, 37, 21, 26, 10, 17, 17, 10, 
    60, 71, 36, 57, 41, 27, 39, 48, 38, 23, 13, 12, 30, 20, 6, 
    68, 66, 40, 83, 61, 60, 73, 64, 39, 23, 31, 40, 50, 47, 37, 
    85, 71, 64, 99, 64, 35, 46, 45, 43, 49, 54, 58, 61, 64, 61, 
    66, 73, 72, 81, 39, 53, 54, 51, 51, 54, 62, 67, 68, 68, 75, 
    67, 61, 88, 59, 45, 59, 54, 53, 55, 60, 65, 66, 63, 75, 73, 
    67, 64, 58, 58, 47, 53, 57, 55, 60, 63, 62, 62, 77, 82, 60, 
    
    -- channel=27
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 3, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 15, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=28
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 5, 4, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 9, 1, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 5, 0, 1, 0, 4, 5, 0, 
    3, 14, 0, 0, 24, 0, 0, 0, 4, 0, 0, 4, 7, 5, 0, 
    1, 13, 0, 0, 0, 0, 6, 0, 10, 2, 8, 4, 5, 9, 0, 
    0, 22, 0, 0, 0, 0, 0, 2, 9, 0, 6, 8, 8, 0, 0, 
    8, 18, 1, 13, 0, 6, 8, 3, 5, 0, 11, 4, 7, 0, 0, 
    15, 13, 18, 16, 10, 0, 0, 10, 0, 0, 6, 14, 7, 0, 0, 
    33, 8, 20, 9, 4, 0, 0, 17, 15, 11, 26, 23, 23, 28, 28, 
    50, 31, 17, 0, 25, 51, 47, 47, 49, 43, 47, 48, 54, 50, 53, 
    55, 41, 19, 11, 44, 44, 44, 43, 46, 48, 53, 51, 50, 54, 58, 
    65, 54, 26, 48, 42, 44, 45, 44, 46, 49, 53, 60, 60, 61, 59, 
    58, 60, 47, 64, 46, 50, 50, 45, 43, 48, 52, 54, 54, 57, 62, 
    
    -- channel=29
    3, 5, 6, 7, 6, 6, 8, 8, 8, 5, 4, 4, 6, 7, 5, 
    7, 9, 8, 7, 5, 8, 14, 12, 0, 0, 0, 0, 0, 0, 6, 
    8, 0, 6, 7, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 6, 7, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 13, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=30
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 5, 0, 0, 1, 0, 0, 0, 0, 4, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 7, 0, 0, 0, 0, 3, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 2, 5, 0, 
    3, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 1, 16, 0, 0, 1, 12, 0, 0, 0, 0, 0, 0, 0, 
    9, 3, 2, 21, 20, 14, 1, 0, 0, 8, 22, 25, 16, 8, 8, 
    11, 5, 7, 10, 0, 5, 18, 17, 20, 25, 28, 31, 37, 33, 32, 
    36, 14, 8, 0, 1, 28, 28, 27, 28, 32, 36, 37, 31, 32, 43, 
    38, 35, 10, 0, 18, 30, 31, 29, 29, 32, 34, 33, 37, 42, 28, 
    38, 38, 30, 16, 23, 23, 21, 27, 33, 37, 34, 36, 45, 43, 36, 
    
    -- channel=31
    8, 7, 7, 9, 7, 3, 9, 5, 3, 3, 2, 0, 4, 7, 5, 
    3, 2, 4, 10, 4, 17, 24, 5, 4, 0, 18, 8, 0, 0, 5, 
    10, 0, 6, 8, 3, 0, 34, 2, 0, 0, 48, 37, 30, 0, 0, 
    53, 0, 10, 0, 14, 0, 30, 31, 21, 0, 64, 21, 32, 13, 0, 
    84, 13, 42, 0, 57, 53, 66, 48, 23, 0, 44, 53, 16, 28, 0, 
    85, 47, 61, 20, 8, 63, 81, 45, 45, 0, 89, 61, 8, 29, 20, 
    90, 69, 23, 36, 0, 26, 62, 68, 54, 0, 88, 48, 12, 14, 37, 
    91, 77, 41, 29, 0, 17, 103, 40, 47, 0, 69, 49, 3, 24, 29, 
    103, 64, 102, 16, 45, 17, 37, 29, 7, 26, 6, 46, 0, 9, 11, 
    80, 68, 108, 0, 61, 28, 14, 56, 37, 32, 37, 0, 0, 0, 12, 
    21, 66, 98, 0, 138, 60, 31, 72, 76, 28, 4, 11, 12, 9, 21, 
    0, 48, 79, 24, 131, 71, 24, 27, 36, 25, 28, 29, 36, 37, 43, 
    52, 2, 27, 92, 114, 37, 36, 31, 30, 28, 30, 36, 42, 40, 44, 
    59, 33, 0, 114, 57, 32, 44, 31, 29, 34, 38, 39, 44, 35, 59, 
    69, 39, 33, 25, 32, 21, 31, 38, 34, 43, 46, 34, 30, 69, 68, 
    
    -- channel=32
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=33
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 2, 0, 5, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 23, 14, 0, 0, 0, 0, 8, 0, 0, 
    44, 0, 0, 0, 3, 0, 3, 0, 0, 0, 18, 0, 17, 2, 0, 
    38, 0, 5, 0, 0, 0, 13, 12, 5, 0, 2, 18, 0, 15, 0, 
    11, 0, 12, 0, 0, 0, 18, 13, 28, 0, 9, 26, 0, 6, 4, 
    13, 0, 0, 32, 0, 0, 0, 10, 28, 0, 30, 17, 0, 0, 0, 
    3, 10, 0, 16, 0, 0, 15, 0, 15, 0, 18, 23, 0, 0, 0, 
    6, 0, 31, 0, 0, 0, 15, 3, 0, 16, 0, 23, 0, 0, 0, 
    0, 0, 44, 0, 4, 0, 0, 8, 0, 0, 19, 2, 0, 0, 0, 
    0, 0, 42, 0, 36, 0, 0, 0, 11, 16, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 40, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 25, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    
    -- channel=34
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 
    0, 18, 0, 0, 0, 11, 14, 11, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 24, 16, 0, 0, 0, 0, 0, 14, 0, 0, 0, 
    4, 0, 10, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 21, 13, 5, 0, 6, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 33, 6, 0, 0, 0, 0, 31, 6, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 18, 28, 9, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 15, 11, 0, 0, 0, 0, 0, 1, 
    14, 16, 0, 0, 29, 56, 22, 22, 11, 0, 0, 0, 0, 0, 0, 
    0, 8, 9, 0, 59, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    3, 0, 0, 32, 14, 0, 0, 0, 0, 0, 0, 4, 6, 0, 9, 
    0, 0, 0, 30, 10, 8, 12, 2, 0, 0, 0, 0, 0, 0, 5, 
    
    -- channel=35
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 11, 0, 0, 
    7, 7, 0, 0, 0, 35, 17, 28, 0, 0, 0, 0, 0, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 10, 4, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 12, 
    23, 0, 0, 26, 25, 16, 0, 0, 0, 0, 2, 14, 0, 0, 0, 
    9, 0, 16, 0, 2, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 17, 19, 0, 0, 3, 11, 0, 0, 0, 
    0, 0, 8, 0, 0, 45, 14, 0, 0, 18, 21, 29, 10, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 6, 11, 19, 7, 0, 0, 0, 
    0, 0, 10, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 6, 
    34, 0, 0, 0, 59, 59, 42, 39, 13, 0, 0, 0, 0, 0, 0, 
    0, 29, 0, 0, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 22, 15, 5, 0, 0, 0, 0, 0, 0, 5, 2, 0, 18, 
    0, 0, 9, 39, 16, 11, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=36
    17, 19, 19, 18, 18, 18, 22, 24, 18, 11, 8, 10, 12, 16, 14, 
    18, 23, 21, 20, 18, 9, 16, 15, 8, 0, 0, 0, 0, 8, 12, 
    5, 10, 21, 22, 21, 9, 2, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 18, 20, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 10, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=37
    0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    4, 3, 2, 1, 2, 31, 17, 0, 0, 0, 21, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 9, 9, 8, 15, 0, 0, 
    24, 25, 5, 0, 0, 0, 23, 16, 5, 0, 1, 0, 0, 3, 0, 
    34, 48, 18, 4, 62, 59, 6, 8, 0, 3, 21, 25, 6, 16, 0, 
    8, 0, 17, 0, 0, 0, 18, 18, 20, 14, 4, 0, 0, 9, 29, 
    26, 0, 0, 0, 0, 9, 0, 15, 4, 0, 0, 10, 4, 10, 20, 
    25, 3, 34, 12, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 0, 21, 0, 21, 0, 0, 5, 6, 4, 0, 0, 0, 0, 19, 
    0, 0, 10, 4, 3, 2, 3, 34, 15, 0, 0, 0, 16, 15, 0, 
    0, 0, 0, 24, 95, 71, 7, 0, 0, 7, 19, 34, 11, 0, 0, 
    0, 0, 17, 22, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 5, 7, 12, 0, 0, 14, 
    0, 2, 0, 0, 0, 1, 10, 2, 0, 1, 0, 0, 0, 5, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 12, 15, 6, 1, 23, 21, 7, 
    
    -- channel=38
    34, 31, 33, 33, 34, 30, 35, 36, 34, 31, 29, 29, 28, 32, 31, 
    36, 31, 32, 33, 31, 24, 32, 32, 23, 18, 16, 23, 28, 30, 31, 
    32, 30, 35, 34, 36, 20, 27, 20, 21, 8, 10, 10, 17, 31, 27, 
    10, 33, 35, 33, 32, 18, 13, 17, 19, 14, 12, 19, 16, 29, 27, 
    0, 14, 32, 17, 0, 7, 7, 16, 19, 19, 7, 16, 15, 16, 34, 
    11, 11, 31, 38, 7, 9, 5, 9, 15, 16, 10, 15, 14, 12, 20, 
    10, 8, 32, 22, 11, 16, 0, 10, 8, 9, 8, 16, 18, 14, 20, 
    12, 0, 24, 16, 14, 3, 6, 15, 14, 15, 12, 16, 15, 18, 24, 
    2, 0, 19, 12, 28, 12, 16, 16, 15, 18, 21, 17, 21, 22, 31, 
    1, 2, 6, 4, 12, 21, 9, 0, 25, 18, 14, 15, 19, 28, 30, 
    0, 4, 3, 1, 0, 7, 5, 0, 6, 9, 11, 9, 10, 11, 12, 
    4, 0, 0, 0, 1, 11, 8, 7, 8, 5, 5, 2, 1, 4, 3, 
    6, 12, 7, 1, 0, 3, 3, 5, 5, 5, 1, 1, 1, 0, 0, 
    0, 5, 14, 0, 5, 2, 4, 5, 3, 2, 2, 1, 0, 1, 3, 
    0, 1, 11, 0, 9, 9, 5, 3, 1, 0, 2, 2, 0, 0, 0, 
    
    -- channel=39
    44, 44, 44, 45, 46, 42, 47, 50, 45, 39, 35, 36, 36, 38, 37, 
    44, 45, 46, 47, 45, 39, 43, 43, 32, 19, 10, 17, 27, 34, 38, 
    37, 42, 48, 47, 48, 47, 26, 20, 8, 7, 0, 0, 4, 20, 33, 
    8, 28, 47, 47, 43, 29, 15, 2, 1, 10, 6, 5, 0, 1, 28, 
    0, 16, 40, 36, 21, 15, 10, 2, 2, 6, 9, 2, 3, 0, 16, 
    0, 13, 35, 26, 18, 9, 8, 5, 0, 9, 9, 1, 5, 0, 0, 
    0, 9, 31, 31, 21, 14, 16, 7, 1, 13, 4, 0, 2, 0, 2, 
    0, 3, 11, 28, 15, 17, 11, 10, 3, 18, 4, 2, 1, 7, 16, 
    0, 3, 0, 10, 12, 13, 9, 6, 9, 25, 12, 4, 3, 15, 32, 
    2, 2, 0, 4, 3, 7, 9, 4, 7, 10, 4, 0, 5, 30, 37, 
    7, 5, 0, 3, 0, 0, 1, 3, 0, 0, 0, 0, 0, 11, 9, 
    0, 0, 0, 16, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=40
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 12, 0, 0, 4, 15, 27, 16, 5, 0, 0, 
    9, 0, 0, 0, 0, 3, 21, 13, 10, 18, 37, 30, 28, 2, 1, 
    44, 0, 0, 0, 6, 5, 29, 22, 24, 5, 42, 20, 31, 18, 0, 
    57, 28, 9, 0, 44, 17, 40, 31, 25, 0, 37, 32, 23, 27, 0, 
    46, 50, 17, 0, 33, 27, 54, 32, 38, 0, 50, 38, 21, 28, 18, 
    43, 63, 15, 13, 4, 25, 53, 42, 43, 7, 56, 36, 22, 26, 27, 
    48, 66, 23, 27, 0, 30, 52, 31, 37, 7, 47, 38, 18, 23, 13, 
    64, 57, 56, 34, 21, 19, 34, 34, 20, 21, 26, 30, 12, 12, 0, 
    62, 54, 72, 26, 45, 9, 18, 54, 22, 25, 30, 15, 10, 0, 4, 
    54, 51, 69, 21, 87, 44, 34, 58, 55, 33, 32, 34, 39, 45, 50, 
    46, 55, 56, 39, 93, 69, 49, 50, 56, 49, 52, 54, 59, 58, 62, 
    69, 38, 35, 78, 81, 53, 51, 50, 52, 53, 57, 60, 61, 62, 68, 
    76, 58, 20, 103, 62, 51, 57, 50, 50, 55, 61, 65, 66, 66, 74, 
    75, 63, 54, 63, 53, 50, 54, 53, 52, 60, 62, 57, 58, 80, 76, 
    
    -- channel=41
    36, 35, 35, 37, 37, 34, 37, 42, 40, 33, 29, 28, 30, 34, 35, 
    36, 38, 35, 38, 35, 16, 41, 34, 27, 11, 6, 13, 18, 25, 33, 
    29, 25, 39, 40, 37, 23, 31, 26, 13, 0, 1, 3, 5, 15, 19, 
    25, 0, 36, 37, 34, 22, 8, 9, 1, 0, 11, 4, 10, 11, 4, 
    14, 0, 39, 17, 0, 3, 12, 12, 6, 0, 4, 14, 1, 9, 9, 
    15, 0, 42, 23, 0, 11, 4, 13, 11, 0, 12, 21, 0, 5, 8, 
    18, 0, 29, 40, 0, 0, 0, 10, 14, 0, 16, 13, 0, 0, 10, 
    7, 0, 14, 24, 0, 0, 19, 3, 17, 0, 6, 16, 0, 1, 21, 
    0, 0, 18, 0, 18, 5, 14, 1, 0, 13, 6, 22, 2, 5, 18, 
    0, 0, 12, 0, 12, 11, 0, 0, 8, 11, 14, 5, 0, 8, 33, 
    0, 0, 12, 0, 0, 0, 0, 0, 7, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=42
    63, 73, 67, 68, 65, 68, 69, 72, 68, 61, 54, 54, 57, 55, 53, 
    62, 71, 69, 71, 68, 90, 60, 68, 55, 44, 32, 27, 35, 47, 53, 
    61, 55, 68, 72, 69, 98, 63, 34, 18, 46, 50, 36, 24, 17, 52, 
    36, 21, 63, 71, 72, 51, 58, 25, 25, 46, 62, 41, 32, 8, 32, 
    48, 54, 57, 59, 96, 55, 71, 40, 28, 24, 63, 35, 31, 16, 3, 
    47, 86, 64, 65, 127, 83, 92, 47, 30, 46, 77, 42, 34, 26, 5, 
    44, 91, 56, 69, 70, 81, 106, 61, 45, 65, 72, 36, 26, 35, 27, 
    64, 91, 23, 56, 40, 103, 80, 64, 47, 70, 75, 42, 31, 44, 41, 
    87, 91, 45, 65, 43, 61, 58, 53, 35, 51, 66, 37, 23, 43, 53, 
    106, 91, 69, 53, 56, 24, 47, 74, 32, 58, 31, 5, 16, 51, 60, 
    98, 88, 72, 75, 83, 35, 63, 88, 44, 13, 0, 0, 9, 27, 24, 
    49, 82, 67, 115, 123, 49, 35, 33, 19, 9, 8, 11, 13, 14, 14, 
    1, 35, 64, 137, 56, 14, 11, 9, 7, 4, 6, 10, 16, 16, 17, 
    7, 3, 38, 119, 25, 13, 11, 8, 9, 10, 11, 16, 10, 13, 24, 
    10, 9, 10, 43, 8, 12, 16, 12, 13, 16, 11, 6, 16, 28, 3, 
    
    -- channel=43
    5, 4, 7, 2, 3, 5, 4, 4, 3, 2, 2, 7, 4, 0, 0, 
    4, 4, 8, 1, 9, 0, 0, 0, 4, 9, 0, 0, 5, 9, 0, 
    0, 25, 4, 2, 10, 10, 0, 0, 7, 23, 0, 0, 0, 9, 9, 
    0, 31, 0, 8, 0, 14, 0, 0, 0, 39, 0, 0, 0, 0, 34, 
    0, 0, 0, 47, 0, 0, 0, 0, 0, 53, 0, 0, 0, 0, 17, 
    0, 0, 0, 22, 33, 1, 0, 0, 0, 84, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 39, 23, 0, 0, 0, 66, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 30, 27, 0, 0, 0, 40, 0, 0, 10, 0, 0, 
    0, 0, 0, 5, 0, 11, 0, 0, 6, 0, 6, 0, 13, 6, 5, 
    0, 0, 0, 25, 0, 5, 17, 0, 0, 0, 0, 0, 13, 11, 0, 
    17, 0, 0, 62, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 9, 0, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 23, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    
    -- channel=44
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 0, 0, 0, 1, 5, 0, 0, 0, 0, 9, 6, 0, 0, 0, 
    21, 6, 0, 0, 0, 0, 1, 0, 0, 0, 12, 0, 0, 0, 0, 
    20, 4, 0, 0, 0, 0, 15, 4, 0, 0, 4, 3, 0, 0, 0, 
    21, 13, 22, 0, 0, 3, 0, 0, 0, 0, 1, 6, 0, 0, 0, 
    12, 13, 18, 0, 11, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 
    4, 12, 17, 0, 0, 2, 8, 23, 17, 0, 1, 4, 10, 15, 21, 
    35, 23, 11, 0, 51, 48, 32, 33, 31, 27, 28, 30, 32, 31, 34, 
    39, 32, 10, 23, 50, 26, 27, 25, 25, 26, 27, 30, 34, 36, 31, 
    44, 35, 29, 38, 30, 25, 26, 27, 27, 30, 35, 40, 39, 37, 52, 
    44, 38, 35, 33, 31, 31, 32, 27, 24, 26, 34, 31, 24, 38, 42, 
    
    -- channel=45
    0, 5, 1, 5, 4, 2, 2, 5, 3, 0, 3, 0, 6, 6, 7, 
    4, 2, 0, 6, 0, 9, 12, 3, 9, 1, 13, 2, 0, 0, 7, 
    5, 0, 3, 7, 0, 0, 29, 7, 0, 0, 7, 14, 19, 0, 0, 
    55, 0, 3, 0, 11, 0, 11, 9, 6, 0, 36, 0, 24, 11, 0, 
    61, 0, 21, 0, 26, 0, 28, 24, 11, 0, 10, 29, 2, 28, 0, 
    20, 0, 36, 0, 0, 7, 41, 21, 39, 0, 29, 39, 0, 16, 17, 
    26, 17, 9, 35, 0, 0, 8, 31, 41, 0, 46, 25, 0, 0, 15, 
    17, 31, 7, 30, 0, 0, 43, 2, 32, 0, 31, 27, 0, 0, 18, 
    25, 0, 48, 0, 0, 0, 18, 4, 0, 6, 0, 34, 0, 0, 0, 
    10, 0, 67, 0, 20, 0, 0, 22, 0, 1, 34, 3, 0, 0, 7, 
    0, 0, 58, 0, 82, 6, 0, 9, 47, 23, 0, 0, 0, 0, 5, 
    0, 0, 27, 0, 40, 34, 0, 0, 7, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 56, 21, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 29, 
    
    -- channel=46
    0, 6, 8, 10, 8, 7, 6, 6, 9, 0, 0, 0, 4, 6, 8, 
    9, 10, 9, 9, 11, 49, 13, 2, 0, 2, 20, 0, 0, 0, 7, 
    0, 0, 5, 8, 5, 0, 0, 0, 0, 17, 15, 17, 17, 0, 0, 
    30, 8, 5, 9, 13, 5, 34, 17, 9, 0, 14, 0, 0, 0, 0, 
    40, 42, 12, 14, 88, 49, 15, 13, 0, 0, 25, 23, 13, 22, 0, 
    0, 6, 10, 0, 0, 0, 37, 21, 27, 17, 10, 0, 0, 16, 21, 
    7, 13, 0, 17, 0, 18, 12, 20, 19, 5, 4, 9, 1, 15, 16, 
    13, 26, 9, 19, 11, 12, 0, 0, 0, 0, 6, 0, 0, 0, 2, 
    20, 9, 9, 9, 8, 0, 0, 17, 6, 0, 0, 0, 0, 5, 21, 
    2, 5, 24, 5, 8, 0, 5, 51, 0, 0, 0, 0, 12, 15, 2, 
    0, 5, 8, 31, 108, 61, 22, 0, 8, 8, 13, 32, 8, 0, 0, 
    0, 0, 23, 38, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 1, 
    3, 0, 0, 4, 0, 3, 2, 0, 1, 6, 8, 11, 2, 0, 15, 
    1, 0, 0, 0, 0, 2, 9, 1, 2, 4, 0, 0, 0, 8, 0, 
    6, 2, 0, 0, 0, 0, 0, 3, 15, 15, 4, 0, 25, 25, 8, 
    
    -- channel=47
    0, 5, 2, 3, 0, 4, 2, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 2, 3, 2, 26, 4, 1, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 2, 3, 0, 10, 5, 0, 0, 9, 18, 9, 0, 0, 0, 
    5, 0, 3, 2, 6, 0, 14, 0, 0, 4, 24, 2, 0, 0, 0, 
    28, 28, 9, 2, 52, 29, 30, 8, 0, 0, 26, 8, 0, 0, 0, 
    28, 47, 19, 1, 45, 37, 46, 13, 1, 10, 38, 10, 0, 0, 0, 
    31, 48, 10, 1, 9, 34, 48, 29, 11, 20, 35, 8, 0, 5, 3, 
    44, 52, 10, 9, 0, 42, 37, 17, 10, 17, 32, 8, 0, 7, 5, 
    57, 53, 27, 27, 8, 12, 16, 12, 8, 6, 8, 0, 0, 4, 3, 
    57, 52, 39, 22, 22, 0, 15, 37, 8, 7, 0, 0, 0, 3, 2, 
    47, 50, 38, 41, 73, 24, 32, 44, 22, 0, 0, 0, 1, 3, 1, 
    15, 45, 43, 66, 64, 20, 8, 6, 5, 0, 2, 4, 10, 11, 10, 
    9, 11, 39, 74, 26, 7, 5, 3, 1, 2, 6, 10, 13, 11, 19, 
    13, 6, 14, 61, 10, 7, 8, 3, 4, 7, 8, 10, 9, 14, 17, 
    15, 10, 8, 9, 0, 0, 4, 7, 9, 13, 9, 6, 18, 28, 11, 
    
    -- channel=48
    45, 44, 42, 43, 42, 42, 45, 46, 41, 41, 40, 41, 37, 35, 33, 
    41, 41, 43, 44, 43, 38, 39, 41, 41, 31, 19, 24, 35, 40, 35, 
    40, 54, 46, 44, 47, 74, 46, 33, 18, 34, 35, 25, 15, 30, 38, 
    11, 25, 45, 45, 40, 38, 28, 18, 22, 50, 40, 35, 25, 10, 36, 
    26, 34, 43, 44, 35, 30, 44, 24, 23, 34, 40, 20, 21, 6, 19, 
    51, 66, 48, 51, 98, 67, 48, 28, 10, 41, 56, 35, 30, 17, 2, 
    45, 59, 57, 34, 53, 57, 70, 42, 24, 57, 54, 27, 26, 27, 20, 
    54, 56, 29, 36, 35, 72, 63, 57, 36, 58, 54, 33, 30, 41, 34, 
    62, 71, 38, 47, 38, 65, 47, 32, 33, 44, 56, 35, 29, 32, 32, 
    79, 73, 42, 47, 41, 29, 42, 36, 35, 48, 29, 11, 14, 36, 43, 
    80, 71, 51, 58, 27, 15, 49, 70, 33, 15, 5, 1, 16, 42, 37, 
    76, 81, 53, 84, 102, 66, 53, 51, 32, 24, 24, 27, 27, 29, 28, 
    24, 64, 74, 99, 61, 24, 22, 23, 21, 20, 21, 23, 30, 32, 29, 
    26, 24, 73, 90, 34, 26, 21, 21, 22, 23, 28, 35, 29, 29, 46, 
    27, 23, 33, 59, 29, 33, 33, 24, 21, 24, 25, 25, 26, 31, 19, 
    
    -- channel=49
    35, 36, 40, 42, 41, 40, 41, 40, 40, 31, 21, 24, 34, 35, 32, 
    41, 43, 42, 42, 45, 80, 56, 35, 8, 30, 47, 30, 14, 23, 35, 
    15, 13, 40, 41, 37, 15, 16, 12, 24, 46, 46, 44, 33, 8, 27, 
    54, 43, 45, 44, 43, 43, 62, 36, 25, 22, 44, 18, 16, 7, 13, 
    78, 86, 56, 63, 134, 93, 57, 35, 10, 26, 70, 48, 34, 32, 2, 
    47, 60, 58, 0, 1, 38, 74, 57, 40, 50, 58, 27, 28, 36, 35, 
    63, 52, 28, 38, 19, 59, 66, 59, 44, 44, 51, 38, 26, 39, 40, 
    66, 80, 58, 62, 41, 62, 42, 17, 30, 31, 38, 29, 21, 23, 30, 
    75, 72, 44, 46, 41, 1, 30, 39, 46, 35, 6, 0, 0, 27, 45, 
    56, 63, 59, 47, 53, 26, 50, 87, 36, 9, 3, 6, 34, 50, 43, 
    51, 67, 52, 89, 144, 102, 59, 46, 43, 33, 37, 46, 36, 31, 28, 
    5, 40, 80, 99, 29, 0, 0, 0, 10, 19, 23, 22, 29, 30, 29, 
    30, 2, 51, 67, 14, 27, 24, 21, 23, 26, 33, 40, 31, 27, 51, 
    29, 23, 9, 33, 22, 30, 33, 24, 22, 28, 22, 18, 22, 37, 8, 
    32, 22, 9, 6, 7, 3, 10, 26, 36, 42, 29, 26, 55, 58, 31, 
    
    -- channel=50
    2, 3, 3, 3, 1, 3, 6, 1, 0, 11, 16, 13, 8, 4, 0, 
    1, 4, 4, 5, 2, 1, 13, 17, 16, 0, 4, 2, 1, 9, 7, 
    19, 15, 3, 0, 0, 0, 0, 0, 0, 2, 9, 4, 12, 8, 8, 
    7, 2, 9, 1, 6, 0, 10, 13, 9, 11, 3, 4, 0, 4, 8, 
    12, 28, 18, 4, 45, 33, 6, 0, 1, 0, 0, 12, 1, 8, 7, 
    4, 12, 17, 0, 0, 2, 2, 0, 2, 8, 18, 0, 4, 6, 7, 
    0, 14, 9, 2, 0, 0, 26, 9, 7, 10, 1, 0, 0, 0, 10, 
    6, 1, 15, 14, 8, 40, 16, 0, 0, 0, 0, 0, 1, 12, 0, 
    5, 10, 4, 9, 9, 0, 0, 0, 7, 0, 0, 0, 0, 0, 9, 
    0, 2, 5, 0, 22, 14, 0, 13, 8, 20, 12, 0, 23, 22, 13, 
    5, 6, 0, 0, 31, 42, 55, 38, 36, 4, 0, 21, 20, 17, 14, 
    16, 14, 17, 24, 14, 0, 0, 0, 0, 4, 8, 3, 0, 0, 2, 
    10, 7, 0, 24, 0, 2, 7, 2, 0, 1, 1, 6, 14, 8, 1, 
    2, 7, 16, 14, 0, 1, 1, 3, 5, 5, 1, 1, 0, 3, 19, 
    7, 1, 2, 0, 0, 0, 8, 7, 8, 0, 1, 0, 0, 8, 7, 
    
    -- channel=51
    23, 20, 22, 24, 25, 19, 25, 26, 24, 19, 13, 11, 17, 24, 26, 
    24, 24, 23, 25, 21, 16, 29, 17, 17, 4, 15, 13, 6, 13, 23, 
    12, 7, 25, 26, 25, 2, 18, 12, 7, 0, 1, 0, 19, 5, 12, 
    34, 0, 28, 21, 22, 8, 14, 9, 6, 0, 9, 2, 9, 13, 0, 
    16, 0, 32, 0, 7, 7, 7, 9, 7, 0, 5, 18, 4, 17, 3, 
    0, 0, 27, 15, 0, 0, 10, 11, 24, 0, 4, 8, 0, 8, 15, 
    0, 3, 6, 34, 0, 0, 0, 7, 16, 0, 9, 10, 2, 0, 12, 
    0, 0, 8, 25, 1, 0, 0, 0, 7, 0, 3, 11, 0, 0, 10, 
    0, 0, 12, 0, 11, 0, 5, 6, 0, 25, 0, 5, 0, 6, 20, 
    0, 0, 14, 0, 2, 0, 0, 11, 0, 0, 8, 3, 0, 8, 17, 
    0, 0, 12, 0, 24, 7, 0, 0, 0, 10, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=52
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 3, 0, 0, 
    19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 2, 0, 0, 
    15, 0, 0, 0, 1, 0, 2, 3, 1, 0, 0, 5, 0, 9, 0, 
    0, 0, 0, 0, 0, 0, 10, 5, 19, 0, 0, 1, 0, 3, 0, 
    0, 7, 0, 0, 0, 0, 0, 0, 16, 0, 4, 2, 0, 0, 0, 
    0, 10, 0, 0, 0, 0, 5, 0, 1, 0, 3, 5, 0, 0, 0, 
    1, 0, 6, 0, 0, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 23, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 17, 0, 34, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 1, 5, 5, 7, 
    9, 0, 0, 0, 16, 4, 5, 3, 5, 5, 6, 5, 4, 2, 5, 
    14, 0, 0, 18, 6, 3, 9, 5, 3, 5, 6, 4, 8, 3, 7, 
    18, 9, 0, 0, 3, 0, 0, 5, 6, 10, 11, 6, 4, 22, 21, 
    
    -- channel=53
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 
    0, 11, 0, 0, 38, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 
    0, 8, 0, 0, 11, 4, 0, 0, 0, 29, 0, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 4, 0, 5, 0, 20, 0, 0, 0, 0, 0, 
    6, 20, 0, 3, 0, 18, 1, 0, 0, 0, 6, 0, 3, 0, 0, 
    18, 22, 0, 26, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 16, 0, 34, 0, 0, 0, 3, 0, 0, 0, 0, 5, 10, 0, 
    53, 30, 0, 34, 20, 32, 40, 39, 20, 15, 17, 24, 26, 28, 23, 
    25, 48, 35, 26, 12, 17, 16, 18, 19, 20, 24, 24, 24, 27, 30, 
    28, 26, 55, 19, 9, 23, 17, 18, 19, 22, 30, 33, 31, 35, 34, 
    24, 29, 34, 42, 21, 29, 23, 16, 18, 24, 24, 29, 32, 29, 17, 
    
    -- channel=54
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 19, 0, 6, 0, 11, 8, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 19, 9, 0, 0, 13, 6, 32, 0, 0, 
    77, 0, 0, 0, 10, 0, 13, 9, 2, 0, 32, 0, 18, 13, 0, 
    56, 0, 24, 0, 11, 4, 35, 23, 16, 0, 13, 37, 0, 30, 0, 
    20, 0, 27, 0, 0, 0, 33, 28, 53, 0, 37, 36, 0, 14, 13, 
    11, 37, 0, 36, 0, 0, 18, 19, 54, 0, 48, 27, 0, 0, 16, 
    4, 32, 16, 27, 0, 0, 45, 0, 18, 0, 20, 34, 0, 0, 1, 
    18, 0, 51, 0, 0, 0, 13, 8, 0, 28, 0, 33, 0, 0, 0, 
    0, 0, 71, 0, 31, 0, 0, 29, 2, 0, 34, 0, 0, 0, 6, 
    0, 0, 68, 0, 72, 23, 0, 8, 42, 28, 0, 0, 0, 0, 6, 
    0, 0, 13, 0, 82, 22, 0, 0, 3, 0, 0, 0, 0, 0, 2, 
    14, 0, 0, 17, 68, 0, 3, 0, 1, 0, 0, 0, 0, 0, 0, 
    18, 0, 0, 64, 12, 0, 9, 0, 0, 0, 0, 0, 2, 0, 13, 
    24, 0, 0, 13, 6, 0, 0, 0, 0, 0, 10, 0, 0, 21, 41, 
    
    -- channel=55
    23, 23, 22, 24, 24, 20, 20, 25, 27, 23, 20, 16, 17, 20, 25, 
    22, 20, 20, 24, 21, 19, 19, 21, 17, 12, 10, 9, 12, 16, 22, 
    28, 14, 24, 25, 23, 18, 31, 18, 12, 0, 12, 12, 13, 8, 13, 
    28, 0, 19, 22, 26, 12, 12, 13, 10, 0, 22, 9, 20, 18, 0, 
    21, 0, 21, 0, 2, 0, 13, 20, 16, 0, 7, 17, 10, 18, 1, 
    16, 6, 25, 17, 7, 11, 20, 14, 21, 0, 19, 26, 6, 13, 10, 
    15, 10, 17, 32, 0, 3, 11, 16, 22, 0, 24, 19, 7, 6, 15, 
    11, 9, 6, 15, 0, 0, 27, 14, 25, 0, 24, 23, 4, 7, 20, 
    15, 0, 28, 3, 12, 5, 19, 15, 3, 5, 17, 28, 8, 13, 15, 
    16, 4, 30, 0, 16, 8, 0, 5, 7, 22, 22, 9, 0, 1, 20, 
    0, 2, 26, 0, 17, 1, 0, 8, 21, 9, 4, 0, 0, 1, 10, 
    0, 0, 8, 0, 29, 30, 5, 7, 14, 5, 2, 0, 0, 0, 2, 
    3, 0, 0, 7, 45, 3, 1, 2, 3, 1, 0, 0, 0, 0, 0, 
    7, 0, 0, 34, 19, 0, 4, 1, 0, 0, 0, 2, 3, 0, 3, 
    6, 0, 0, 8, 9, 4, 5, 4, 0, 0, 3, 0, 0, 0, 10, 
    
    -- channel=56
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 8, 6, 0, 
    13, 26, 0, 0, 0, 24, 11, 10, 0, 0, 0, 0, 0, 11, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 48, 9, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 17, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 15, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 32, 0, 0, 0, 0, 19, 25, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 22, 7, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 20, 7, 0, 0, 0, 0, 10, 10, 
    46, 20, 0, 0, 31, 52, 28, 26, 13, 0, 0, 0, 0, 0, 0, 
    0, 33, 10, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 34, 32, 5, 0, 0, 0, 0, 0, 0, 5, 0, 0, 15, 
    0, 0, 1, 36, 8, 14, 15, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=57
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=58
    27, 26, 30, 26, 27, 26, 28, 31, 29, 23, 25, 30, 27, 22, 21, 
    29, 27, 31, 25, 32, 11, 15, 24, 24, 22, 0, 0, 17, 31, 21, 
    8, 50, 30, 28, 30, 8, 13, 9, 17, 9, 0, 0, 0, 18, 26, 
    0, 28, 22, 33, 15, 32, 0, 0, 0, 26, 0, 0, 0, 0, 38, 
    0, 0, 9, 66, 0, 0, 0, 0, 0, 51, 0, 0, 0, 0, 19, 
    0, 0, 9, 22, 20, 24, 0, 0, 0, 55, 0, 0, 1, 0, 0, 
    4, 0, 27, 0, 15, 26, 0, 0, 0, 25, 0, 0, 0, 1, 0, 
    0, 0, 2, 0, 25, 7, 0, 0, 0, 11, 0, 0, 8, 0, 11, 
    0, 0, 0, 10, 1, 13, 0, 0, 17, 0, 2, 0, 9, 13, 16, 
    0, 0, 0, 4, 0, 20, 28, 0, 0, 11, 0, 7, 12, 20, 21, 
    0, 0, 0, 37, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=59
    29, 33, 29, 29, 29, 29, 31, 34, 30, 23, 23, 26, 26, 27, 27, 
    28, 33, 28, 30, 26, 25, 20, 30, 24, 14, 1, 10, 20, 24, 25, 
    29, 29, 31, 33, 29, 35, 34, 21, 4, 0, 0, 0, 0, 11, 27, 
    6, 3, 27, 29, 30, 13, 3, 0, 0, 0, 12, 5, 11, 9, 14, 
    0, 0, 19, 0, 0, 0, 9, 8, 11, 0, 0, 0, 2, 2, 5, 
    0, 4, 24, 25, 36, 10, 13, 0, 8, 0, 1, 11, 0, 0, 0, 
    0, 8, 25, 34, 8, 3, 2, 3, 6, 0, 7, 5, 1, 0, 0, 
    0, 1, 0, 14, 0, 0, 11, 13, 14, 1, 12, 11, 0, 4, 18, 
    0, 0, 0, 4, 1, 15, 17, 8, 0, 12, 17, 22, 13, 17, 16, 
    4, 0, 7, 0, 0, 0, 0, 0, 0, 15, 14, 3, 0, 8, 19, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 15, 2, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=60
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 0, 0, 0, 14, 21, 11, 12, 1, 0, 
    10, 0, 0, 0, 0, 0, 11, 6, 8, 21, 14, 13, 5, 0, 0, 
    21, 29, 0, 0, 27, 19, 22, 6, 8, 2, 21, 10, 7, 3, 0, 
    25, 37, 0, 0, 37, 20, 22, 12, 7, 16, 28, 9, 13, 8, 0, 
    17, 46, 5, 0, 18, 14, 44, 15, 17, 32, 26, 9, 8, 11, 7, 
    26, 40, 16, 5, 9, 46, 25, 21, 7, 20, 19, 11, 13, 14, 0, 
    37, 48, 18, 25, 3, 19, 11, 12, 13, 10, 19, 5, 1, 0, 0, 
    36, 43, 28, 30, 30, 2, 10, 31, 15, 15, 9, 3, 11, 3, 0, 
    48, 40, 31, 30, 37, 32, 45, 50, 29, 11, 13, 20, 32, 35, 29, 
    63, 46, 35, 58, 67, 30, 35, 33, 31, 30, 34, 36, 37, 41, 39, 
    44, 49, 32, 68, 29, 32, 34, 31, 30, 32, 37, 40, 45, 44, 43, 
    45, 41, 51, 60, 27, 34, 32, 33, 34, 37, 41, 45, 41, 45, 56, 
    44, 42, 40, 47, 30, 34, 37, 32, 35, 37, 39, 36, 41, 54, 43, 
    
    -- channel=61
    46, 47, 47, 49, 48, 46, 48, 54, 50, 39, 32, 31, 38, 45, 46, 
    46, 50, 50, 50, 49, 27, 50, 36, 35, 15, 11, 11, 15, 29, 40, 
    24, 28, 48, 52, 49, 36, 32, 28, 16, 0, 12, 13, 13, 13, 24, 
    36, 0, 43, 48, 36, 31, 19, 18, 4, 0, 16, 11, 14, 10, 11, 
    36, 0, 45, 41, 20, 22, 23, 16, 6, 0, 19, 24, 7, 16, 5, 
    22, 0, 45, 23, 0, 27, 18, 28, 15, 0, 17, 24, 7, 13, 14, 
    28, 0, 28, 47, 4, 0, 12, 16, 26, 0, 25, 16, 4, 4, 17, 
    13, 9, 21, 28, 23, 0, 19, 7, 24, 0, 16, 19, 3, 5, 32, 
    8, 0, 15, 0, 10, 15, 23, 4, 10, 15, 10, 19, 3, 19, 31, 
    1, 0, 18, 0, 21, 8, 8, 10, 7, 11, 14, 11, 1, 14, 38, 
    0, 0, 19, 0, 15, 10, 0, 0, 10, 3, 0, 0, 0, 0, 0, 
    0, 0, 20, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=62
    34, 41, 38, 37, 35, 39, 41, 41, 36, 34, 33, 34, 33, 32, 27, 
    34, 42, 39, 40, 36, 43, 38, 44, 37, 18, 12, 13, 20, 28, 29, 
    37, 33, 39, 40, 37, 44, 34, 12, 4, 10, 14, 6, 8, 9, 30, 
    14, 5, 38, 39, 42, 21, 23, 6, 4, 13, 25, 15, 7, 1, 16, 
    14, 20, 36, 24, 48, 31, 34, 14, 6, 0, 22, 14, 4, 0, 2, 
    15, 34, 41, 36, 55, 43, 41, 14, 6, 8, 35, 15, 6, 2, 0, 
    12, 41, 35, 37, 25, 33, 48, 25, 15, 17, 30, 10, 2, 5, 6, 
    26, 33, 12, 28, 12, 45, 33, 26, 14, 20, 29, 11, 5, 15, 14, 
    33, 34, 18, 27, 19, 24, 21, 15, 9, 21, 26, 12, 1, 13, 28, 
    36, 30, 26, 12, 26, 9, 13, 27, 10, 27, 12, 0, 4, 27, 33, 
    34, 34, 26, 12, 32, 11, 27, 40, 20, 0, 0, 0, 0, 4, 5, 
    4, 28, 23, 41, 55, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 16, 59, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=63
    2, 0, 4, 0, 0, 4, 4, 0, 0, 0, 0, 2, 1, 0, 0, 
    4, 6, 6, 0, 6, 21, 0, 0, 0, 4, 0, 0, 7, 6, 0, 
    0, 14, 5, 0, 8, 11, 0, 0, 3, 42, 0, 0, 0, 12, 14, 
    0, 66, 3, 7, 0, 5, 0, 0, 0, 52, 0, 0, 0, 0, 42, 
    0, 49, 0, 35, 2, 5, 0, 0, 0, 59, 0, 0, 1, 0, 27, 
    0, 13, 0, 15, 36, 0, 0, 0, 0, 129, 0, 0, 9, 0, 0, 
    0, 0, 0, 0, 55, 36, 0, 0, 0, 111, 0, 0, 5, 11, 0, 
    0, 0, 0, 0, 35, 59, 0, 0, 0, 74, 0, 0, 15, 8, 0, 
    0, 2, 0, 19, 0, 0, 0, 0, 14, 0, 12, 0, 14, 13, 17, 
    0, 1, 0, 46, 0, 0, 15, 0, 2, 0, 0, 0, 32, 37, 0, 
    45, 0, 0, 108, 0, 0, 46, 0, 0, 0, 3, 15, 15, 6, 0, 
    48, 13, 0, 97, 0, 0, 0, 0, 0, 0, 0, 3, 1, 3, 0, 
    0, 47, 40, 5, 0, 0, 0, 0, 0, 2, 5, 7, 1, 0, 6, 
    0, 2, 90, 0, 0, 2, 0, 0, 1, 3, 1, 0, 0, 20, 0, 
    0, 0, 9, 0, 0, 7, 0, 0, 6, 1, 0, 0, 27, 0, 0, 
    
    -- channel=64
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=65
    1, 1, 1, 1, 1, 1, 1, 1, 2, 0, 0, 1, 1, 1, 1, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 5, 1, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 1, 3, 0, 0, 0, 0, 0, 0, 0, 
    12, 7, 0, 0, 0, 0, 0, 0, 0, 0, 4, 9, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 14, 13, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 8, 7, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 9, 14, 14, 9, 5, 0, 4, 0, 0, 3, 12, 5, 0, 3, 
    20, 3, 2, 8, 10, 9, 0, 26, 32, 24, 5, 0, 9, 7, 2, 
    23, 12, 10, 10, 11, 11, 6, 20, 15, 8, 18, 16, 10, 5, 1, 
    24, 20, 17, 15, 15, 14, 6, 9, 24, 24, 17, 11, 10, 7, 1, 
    
    -- channel=66
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 13, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    13, 7, 0, 0, 0, 10, 16, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 7, 11, 6, 0, 0, 0, 6, 10, 10, 12, 7, 4, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 
    22, 25, 27, 21, 19, 18, 20, 0, 0, 0, 5, 12, 16, 3, 6, 
    16, 15, 9, 12, 19, 20, 12, 14, 15, 12, 1, 0, 5, 9, 5, 
    16, 21, 19, 19, 21, 21, 10, 0, 0, 0, 9, 15, 8, 7, 4, 
    17, 24, 24, 23, 22, 21, 11, 0, 12, 22, 13, 10, 11, 8, 3, 
    
    -- channel=67
    16, 16, 16, 16, 16, 16, 16, 15, 16, 17, 17, 16, 16, 16, 16, 
    16, 17, 17, 17, 17, 17, 17, 16, 18, 16, 24, 21, 17, 17, 17, 
    15, 16, 17, 16, 17, 17, 18, 18, 22, 17, 29, 20, 16, 17, 17, 
    24, 21, 18, 16, 16, 12, 22, 11, 21, 22, 26, 40, 19, 20, 18, 
    38, 37, 25, 15, 17, 10, 23, 14, 21, 20, 21, 23, 26, 30, 20, 
    12, 16, 23, 17, 18, 17, 16, 16, 18, 16, 20, 18, 13, 40, 23, 
    33, 36, 27, 15, 14, 14, 37, 43, 46, 20, 16, 14, 12, 16, 28, 
    22, 29, 18, 34, 19, 9, 20, 19, 24, 25, 29, 29, 31, 27, 35, 
    53, 13, 11, 16, 22, 20, 26, 6, 16, 19, 17, 17, 21, 26, 25, 
    34, 28, 37, 37, 38, 37, 36, 38, 37, 29, 36, 27, 30, 25, 24, 
    25, 28, 29, 28, 28, 30, 33, 31, 29, 27, 27, 26, 30, 23, 19, 
    0, 15, 0, 0, 2, 9, 17, 27, 29, 27, 23, 20, 6, 7, 17, 
    0, 11, 3, 0, 0, 3, 29, 0, 0, 0, 0, 0, 7, 13, 23, 
    0, 1, 1, 0, 1, 1, 2, 0, 0, 0, 0, 7, 9, 18, 24, 
    0, 0, 2, 1, 1, 3, 7, 0, 0, 1, 4, 8, 12, 17, 24, 
    
    -- channel=68
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=69
    25, 26, 26, 26, 27, 27, 27, 26, 26, 27, 28, 27, 27, 26, 27, 
    25, 27, 27, 26, 27, 26, 27, 26, 25, 19, 39, 33, 26, 27, 27, 
    27, 27, 27, 26, 27, 26, 28, 22, 24, 11, 41, 45, 26, 27, 28, 
    31, 27, 29, 27, 27, 19, 36, 9, 14, 9, 11, 43, 29, 29, 29, 
    30, 37, 48, 28, 27, 16, 33, 22, 29, 24, 30, 31, 30, 48, 33, 
    9, 20, 39, 24, 32, 27, 44, 43, 44, 21, 6, 7, 0, 45, 36, 
    28, 42, 32, 21, 17, 0, 5, 13, 38, 33, 32, 29, 32, 35, 44, 
    16, 19, 2, 45, 19, 0, 20, 22, 25, 9, 0, 0, 7, 9, 26, 
    48, 28, 9, 29, 39, 31, 38, 9, 20, 26, 30, 25, 32, 31, 18, 
    66, 30, 37, 34, 32, 27, 20, 14, 22, 2, 19, 3, 9, 12, 18, 
    0, 6, 0, 7, 14, 22, 24, 22, 17, 9, 7, 8, 9, 3, 14, 
    0, 2, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 10, 1, 12, 
    0, 0, 0, 0, 0, 0, 58, 0, 0, 0, 0, 0, 0, 9, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 12, 28, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 14, 27, 
    
    -- channel=70
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 14, 0, 0, 
    0, 0, 0, 0, 2, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 0, 5, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 1, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 0, 16, 23, 12, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 
    33, 0, 0, 14, 10, 2, 0, 10, 12, 14, 10, 0, 0, 0, 0, 
    64, 4, 0, 7, 4, 3, 0, 0, 25, 2, 0, 0, 0, 0, 0, 
    56, 10, 4, 4, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=71
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=72
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=73
    31, 31, 31, 31, 30, 30, 31, 30, 29, 31, 32, 30, 30, 31, 31, 
    31, 31, 31, 31, 31, 30, 30, 30, 31, 34, 28, 28, 31, 31, 31, 
    29, 30, 30, 30, 30, 30, 32, 34, 34, 34, 34, 29, 31, 30, 31, 
    37, 37, 32, 29, 30, 30, 27, 33, 46, 52, 52, 44, 35, 34, 33, 
    30, 25, 22, 27, 30, 30, 34, 32, 40, 41, 44, 37, 27, 26, 33, 
    51, 52, 40, 24, 23, 27, 22, 24, 32, 42, 45, 48, 50, 45, 37, 
    29, 27, 23, 30, 44, 46, 44, 41, 39, 34, 31, 26, 21, 30, 29, 
    29, 40, 28, 22, 29, 43, 51, 48, 31, 31, 37, 37, 41, 41, 47, 
    28, 40, 40, 40, 43, 40, 35, 36, 44, 49, 45, 46, 42, 39, 34, 
    48, 39, 46, 46, 49, 49, 54, 52, 50, 50, 51, 44, 45, 41, 36, 
    19, 21, 25, 22, 18, 24, 34, 38, 38, 38, 39, 39, 42, 34, 28, 
    4, 8, 10, 12, 7, 8, 34, 56, 47, 44, 39, 32, 25, 16, 22, 
    7, 3, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 19, 26, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 13, 19, 29, 
    3, 0, 2, 2, 1, 3, 0, 0, 0, 0, 7, 11, 15, 23, 31, 
    
    -- channel=74
    6, 8, 8, 8, 9, 9, 9, 8, 9, 8, 9, 9, 9, 8, 9, 
    7, 9, 9, 9, 9, 9, 9, 8, 9, 4, 33, 19, 8, 9, 9, 
    11, 11, 10, 8, 9, 8, 12, 6, 17, 1, 30, 36, 9, 10, 10, 
    9, 5, 10, 10, 9, 2, 27, 0, 0, 0, 0, 9, 8, 9, 9, 
    40, 52, 45, 14, 12, 0, 10, 3, 1, 0, 12, 26, 36, 55, 15, 
    0, 0, 6, 20, 32, 35, 60, 54, 42, 0, 0, 0, 0, 8, 15, 
    39, 56, 40, 9, 0, 0, 0, 0, 7, 15, 25, 31, 41, 33, 48, 
    13, 0, 0, 45, 9, 0, 0, 0, 21, 4, 0, 0, 0, 0, 0, 
    26, 0, 0, 0, 11, 13, 29, 0, 0, 0, 7, 3, 21, 26, 14, 
    42, 30, 32, 27, 22, 15, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 12, 2, 17, 30, 39, 29, 24, 14, 3, 0, 0, 0, 0, 0, 
    0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 8, 0, 0, 0, 74, 14, 0, 5, 18, 19, 0, 3, 11, 
    0, 0, 0, 0, 0, 0, 9, 32, 30, 17, 0, 0, 2, 9, 18, 
    0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 4, 2, 6, 6, 13, 
    
    -- channel=75
    28, 27, 27, 27, 27, 27, 27, 27, 26, 28, 28, 27, 27, 27, 27, 
    28, 27, 27, 27, 27, 27, 27, 26, 27, 30, 26, 28, 27, 27, 27, 
    27, 26, 26, 27, 27, 27, 27, 29, 33, 38, 28, 23, 27, 27, 27, 
    33, 31, 28, 26, 26, 26, 27, 31, 38, 38, 36, 30, 30, 29, 28, 
    35, 35, 28, 25, 27, 26, 23, 29, 31, 39, 38, 34, 33, 29, 29, 
    38, 32, 16, 27, 27, 34, 30, 30, 28, 33, 42, 38, 33, 29, 29, 
    36, 29, 36, 32, 27, 47, 31, 31, 36, 31, 33, 32, 31, 23, 30, 
    24, 31, 22, 15, 32, 45, 34, 25, 26, 32, 37, 36, 31, 35, 36, 
    27, 20, 36, 25, 28, 32, 37, 48, 39, 41, 41, 40, 37, 32, 36, 
    14, 41, 42, 46, 45, 46, 45, 46, 43, 50, 41, 44, 42, 37, 29, 
    26, 25, 32, 31, 29, 33, 42, 42, 42, 41, 41, 38, 35, 34, 22, 
    18, 14, 17, 15, 13, 16, 19, 37, 35, 35, 31, 32, 17, 14, 19, 
    13, 9, 4, 10, 12, 9, 0, 0, 0, 0, 0, 0, 17, 13, 20, 
    21, 8, 6, 8, 8, 8, 0, 0, 0, 0, 1, 5, 11, 19, 22, 
    19, 7, 8, 9, 8, 8, 0, 0, 0, 0, 5, 14, 16, 19, 23, 
    
    -- channel=76
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=77
    3, 3, 3, 3, 4, 4, 4, 3, 3, 4, 5, 4, 3, 3, 3, 
    4, 4, 4, 3, 4, 4, 4, 3, 3, 4, 16, 7, 3, 4, 3, 
    5, 4, 4, 4, 3, 3, 7, 3, 19, 22, 18, 16, 3, 4, 4, 
    7, 5, 5, 3, 3, 0, 11, 6, 7, 5, 1, 5, 7, 6, 5, 
    35, 39, 19, 5, 4, 5, 0, 4, 3, 9, 17, 26, 30, 34, 9, 
    1, 0, 0, 10, 13, 25, 36, 32, 26, 10, 8, 0, 0, 0, 9, 
    38, 39, 29, 16, 0, 14, 15, 8, 2, 10, 19, 25, 28, 21, 30, 
    30, 0, 12, 8, 17, 0, 0, 0, 19, 19, 12, 8, 4, 3, 3, 
    11, 3, 0, 0, 5, 11, 20, 25, 16, 20, 25, 22, 29, 31, 29, 
    11, 39, 40, 41, 37, 36, 29, 26, 24, 25, 26, 29, 24, 20, 16, 
    21, 25, 25, 32, 36, 41, 46, 44, 40, 36, 33, 27, 21, 10, 8, 
    7, 15, 1, 0, 2, 7, 2, 0, 1, 2, 0, 0, 0, 8, 2, 
    0, 3, 7, 3, 4, 0, 15, 0, 0, 0, 0, 4, 0, 0, 3, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 4, 8, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 4, 7, 
    
    -- channel=78
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    58, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    49, 42, 0, 0, 0, 0, 19, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 21, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 3, 21, 15, 12, 1, 0, 4, 4, 0, 13, 0, 0, 0, 0, 
    77, 60, 76, 77, 78, 68, 51, 35, 24, 23, 15, 6, 0, 0, 0, 
    0, 10, 0, 0, 7, 18, 0, 0, 5, 0, 0, 0, 0, 0, 0, 
    7, 39, 35, 12, 8, 15, 79, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 16, 9, 11, 11, 36, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 4, 5, 5, 29, 3, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=79
    35, 35, 35, 35, 35, 36, 36, 35, 35, 35, 38, 36, 35, 35, 36, 
    35, 35, 35, 35, 35, 35, 35, 35, 34, 30, 41, 38, 35, 35, 36, 
    35, 35, 36, 35, 36, 35, 36, 31, 28, 29, 32, 47, 35, 36, 36, 
    39, 38, 36, 35, 36, 33, 38, 31, 39, 37, 38, 38, 37, 37, 37, 
    18, 23, 50, 34, 35, 34, 36, 35, 40, 38, 35, 30, 23, 38, 40, 
    42, 48, 35, 19, 37, 12, 33, 36, 43, 44, 36, 36, 34, 45, 39, 
    23, 26, 31, 43, 36, 1, 21, 31, 36, 33, 29, 26, 31, 31, 36, 
    25, 44, 7, 30, 36, 37, 45, 25, 24, 24, 19, 23, 25, 33, 32, 
    49, 41, 40, 42, 44, 38, 38, 36, 42, 36, 49, 38, 37, 30, 29, 
    46, 37, 41, 41, 44, 42, 42, 35, 36, 31, 31, 28, 29, 27, 30, 
    0, 12, 3, 7, 7, 16, 27, 30, 30, 25, 25, 26, 32, 23, 23, 
    0, 0, 6, 0, 0, 0, 52, 13, 18, 22, 25, 22, 19, 17, 21, 
    0, 0, 0, 0, 0, 0, 6, 10, 5, 0, 0, 2, 6, 16, 27, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 7, 8, 15, 28, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 4, 11, 18, 29, 
    
    -- channel=80
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 7, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 5, 3, 0, 0, 7, 6, 6, 6, 
    4, 5, 5, 6, 6, 5, 6, 0, 0, 4, 6, 6, 6, 6, 6, 
    10, 8, 7, 5, 6, 0, 4, 7, 20, 27, 27, 20, 8, 7, 7, 
    0, 0, 3, 3, 4, 10, 10, 10, 14, 12, 3, 0, 0, 0, 8, 
    42, 38, 15, 0, 0, 0, 0, 0, 0, 10, 24, 33, 29, 23, 10, 
    0, 0, 0, 11, 12, 0, 8, 17, 24, 8, 0, 0, 0, 0, 0, 
    15, 24, 0, 0, 10, 36, 45, 10, 0, 0, 0, 11, 16, 25, 19, 
    33, 32, 31, 25, 14, 3, 0, 11, 21, 18, 20, 12, 2, 0, 0, 
    11, 0, 0, 0, 0, 4, 8, 9, 12, 11, 9, 11, 16, 14, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 10, 16, 19, 12, 
    0, 2, 7, 2, 0, 0, 32, 35, 30, 31, 34, 33, 14, 2, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 3, 7, 
    
    -- channel=81
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 17, 11, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    62, 53, 6, 0, 0, 0, 0, 0, 0, 0, 6, 33, 47, 25, 0, 
    0, 0, 0, 9, 11, 38, 50, 39, 16, 0, 0, 0, 0, 0, 0, 
    70, 64, 32, 0, 0, 8, 0, 0, 0, 0, 17, 36, 32, 27, 27, 
    2, 0, 0, 3, 0, 0, 0, 0, 30, 26, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 9, 3, 0, 0, 0, 0, 20, 35, 31, 
    0, 51, 48, 49, 42, 32, 20, 13, 10, 12, 13, 17, 0, 0, 0, 
    43, 44, 50, 64, 71, 74, 70, 63, 54, 47, 35, 19, 0, 0, 0, 
    8, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 8, 24, 18, 4, 0, 11, 20, 0, 7, 31, 31, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 16, 34, 15, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=82
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    36, 34, 30, 27, 21, 14, 7, 1, 1, 7, 11, 11, 7, 0, 0, 
    35, 31, 15, 33, 48, 50, 33, 32, 37, 33, 21, 0, 0, 0, 0, 
    39, 50, 38, 39, 49, 51, 12, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 51, 49, 49, 52, 51, 34, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 44, 47, 49, 49, 50, 42, 14, 10, 0, 0, 0, 0, 0, 0, 
    
    -- channel=83
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 13, 0, 0, 0, 11, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 4, 7, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 7, 7, 7, 3, 2, 2, 0, 4, 2, 2, 0, 0, 0, 
    24, 24, 26, 27, 25, 26, 23, 22, 17, 20, 16, 12, 3, 0, 0, 
    15, 4, 3, 12, 18, 19, 0, 0, 3, 2, 0, 0, 0, 6, 0, 
    15, 19, 25, 27, 19, 19, 6, 22, 25, 30, 37, 32, 7, 0, 0, 
    7, 17, 21, 22, 19, 18, 25, 79, 97, 60, 17, 0, 0, 0, 0, 
    3, 9, 11, 11, 13, 14, 19, 42, 20, 0, 0, 0, 0, 0, 0, 
    
    -- channel=84
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 10, 11, 0, 0, 23, 10, 4, 0, 0, 0, 0, 0, 
    25, 11, 0, 6, 11, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28, 12, 10, 10, 11, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 17, 15, 15, 14, 13, 16, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=85
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=86
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 8, 7, 9, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 9, 0, 15, 19, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 22, 13, 13, 17, 18, 7, 0, 2, 8, 7, 0, 0, 0, 0, 
    17, 19, 18, 16, 18, 17, 22, 0, 1, 0, 0, 0, 0, 0, 0, 
    13, 20, 18, 18, 17, 15, 19, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=87
    82, 80, 80, 80, 80, 81, 80, 81, 79, 82, 81, 81, 81, 80, 80, 
    82, 81, 81, 81, 80, 81, 80, 82, 83, 103, 65, 71, 81, 81, 81, 
    80, 79, 80, 82, 79, 84, 77, 95, 83, 87, 50, 56, 83, 80, 81, 
    77, 82, 81, 81, 81, 105, 61, 97, 71, 80, 67, 49, 85, 83, 83, 
    62, 45, 62, 77, 80, 96, 68, 86, 76, 89, 92, 82, 73, 37, 81, 
    60, 54, 79, 71, 76, 79, 63, 64, 61, 98, 80, 70, 84, 33, 78, 
    55, 33, 57, 49, 107, 77, 28, 24, 28, 83, 82, 77, 67, 75, 46, 
    0, 39, 47, 27, 72, 73, 51, 90, 70, 69, 64, 50, 42, 51, 48, 
    0, 83, 57, 56, 68, 90, 82, 88, 61, 66, 66, 76, 62, 63, 62, 
    26, 59, 59, 62, 62, 65, 76, 62, 60, 58, 55, 54, 39, 38, 37, 
    20, 11, 27, 21, 18, 17, 31, 32, 40, 38, 32, 26, 23, 35, 30, 
    11, 0, 23, 17, 0, 0, 0, 38, 25, 19, 13, 22, 31, 33, 24, 
    18, 0, 0, 4, 0, 0, 0, 23, 14, 22, 23, 17, 15, 24, 31, 
    58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 32, 27, 40, 
    53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 34, 31, 35, 44, 
    
    -- channel=88
    18, 18, 18, 18, 18, 18, 18, 18, 17, 19, 20, 18, 18, 18, 18, 
    19, 19, 19, 19, 19, 19, 19, 18, 18, 22, 22, 20, 19, 19, 19, 
    19, 19, 19, 18, 19, 18, 20, 20, 27, 25, 29, 20, 19, 18, 19, 
    21, 21, 20, 18, 18, 17, 20, 18, 20, 22, 22, 29, 20, 19, 19, 
    43, 40, 20, 18, 19, 13, 17, 16, 21, 25, 30, 33, 36, 29, 20, 
    13, 14, 23, 23, 21, 29, 29, 27, 24, 19, 19, 16, 14, 23, 22, 
    44, 41, 31, 13, 14, 29, 28, 29, 29, 25, 28, 30, 24, 28, 30, 
    23, 16, 28, 25, 20, 8, 12, 26, 30, 28, 28, 22, 22, 18, 27, 
    23, 14, 6, 11, 22, 24, 27, 18, 23, 27, 25, 30, 32, 36, 33, 
    32, 43, 48, 49, 48, 44, 43, 43, 40, 39, 42, 36, 33, 29, 27, 
    34, 32, 41, 44, 44, 45, 50, 49, 46, 44, 40, 36, 34, 26, 19, 
    2, 11, 0, 3, 5, 10, 4, 25, 27, 27, 24, 21, 16, 15, 10, 
    0, 6, 6, 2, 0, 0, 34, 9, 5, 5, 8, 7, 2, 5, 10, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 3, 8, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 8, 14, 
    
    -- channel=89
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 16, 6, 18, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    48, 44, 8, 0, 0, 0, 0, 0, 0, 0, 20, 36, 46, 22, 0, 
    0, 0, 0, 16, 17, 58, 69, 56, 25, 0, 0, 0, 0, 0, 0, 
    64, 56, 31, 0, 0, 0, 0, 0, 0, 8, 34, 48, 44, 42, 31, 
    0, 0, 0, 10, 0, 0, 0, 0, 22, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 22, 8, 0, 14, 14, 26, 40, 39, 21, 
    41, 57, 54, 52, 41, 29, 14, 3, 10, 3, 17, 11, 2, 5, 0, 
    30, 28, 40, 56, 68, 73, 73, 66, 55, 45, 31, 16, 0, 0, 0, 
    4, 9, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 9, 25, 11, 0, 0, 54, 43, 29, 35, 45, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 23, 48, 42, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=90
    89, 89, 89, 89, 90, 90, 90, 89, 89, 89, 91, 89, 90, 89, 90, 
    89, 90, 90, 89, 89, 89, 89, 89, 87, 77, 81, 88, 89, 89, 90, 
    89, 89, 89, 89, 90, 89, 91, 83, 79, 72, 84, 90, 90, 90, 91, 
    92, 92, 92, 90, 90, 80, 86, 80, 83, 83, 81, 98, 93, 92, 92, 
    59, 69, 84, 88, 90, 86, 92, 89, 93, 91, 88, 76, 68, 85, 92, 
    87, 90, 96, 78, 79, 78, 77, 81, 90, 86, 82, 84, 73, 91, 96, 
    51, 61, 71, 76, 81, 36, 46, 58, 86, 91, 85, 75, 75, 75, 82, 
    45, 58, 52, 69, 76, 74, 92, 85, 65, 56, 51, 53, 62, 70, 83, 
    64, 94, 80, 92, 97, 89, 89, 77, 83, 86, 83, 79, 73, 68, 60, 
    81, 64, 69, 69, 70, 71, 69, 63, 66, 54, 60, 49, 53, 55, 58, 
    11, 16, 18, 19, 22, 29, 38, 42, 41, 37, 37, 39, 47, 48, 55, 
    0, 23, 14, 5, 0, 2, 30, 35, 32, 33, 39, 49, 50, 42, 55, 
    0, 0, 0, 0, 0, 0, 44, 19, 22, 22, 18, 18, 30, 50, 66, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 38, 43, 54, 72, 
    3, 0, 0, 0, 0, 0, 0, 0, 6, 31, 38, 41, 49, 60, 75, 
    
    -- channel=91
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 26, 19, 20, 19, 18, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 15, 0, 2, 14, 24, 28, 0, 10, 9, 5, 0, 0, 0, 0, 
    1, 19, 23, 17, 16, 20, 36, 0, 4, 4, 5, 11, 0, 0, 0, 
    0, 18, 21, 18, 18, 19, 20, 46, 47, 31, 8, 0, 0, 0, 0, 
    0, 9, 14, 13, 16, 17, 15, 30, 12, 0, 0, 0, 0, 0, 0, 
    
    -- channel=92
    11, 11, 11, 11, 11, 11, 11, 11, 10, 12, 13, 11, 11, 11, 11, 
    12, 12, 12, 12, 12, 12, 12, 12, 12, 19, 27, 17, 12, 12, 12, 
    11, 12, 12, 12, 12, 11, 13, 13, 26, 33, 18, 19, 12, 12, 12, 
    19, 15, 14, 11, 11, 14, 17, 18, 20, 21, 19, 13, 16, 15, 14, 
    42, 40, 29, 11, 12, 19, 8, 16, 12, 16, 20, 27, 30, 32, 17, 
    7, 2, 7, 11, 17, 17, 24, 23, 24, 27, 25, 15, 13, 7, 17, 
    41, 41, 36, 17, 20, 23, 36, 32, 16, 14, 16, 18, 23, 19, 27, 
    31, 11, 13, 17, 32, 15, 0, 3, 27, 36, 34, 30, 23, 24, 10, 
    3, 19, 5, 0, 10, 20, 25, 28, 14, 17, 24, 21, 26, 31, 38, 
    11, 40, 44, 47, 46, 48, 49, 44, 43, 38, 40, 42, 34, 27, 23, 
    28, 36, 35, 37, 36, 39, 47, 45, 45, 42, 41, 36, 35, 21, 13, 
    8, 9, 5, 2, 5, 7, 28, 18, 27, 26, 19, 7, 0, 9, 9, 
    0, 4, 9, 8, 7, 4, 0, 0, 0, 0, 0, 6, 4, 3, 9, 
    4, 4, 2, 5, 4, 4, 0, 0, 0, 0, 0, 0, 3, 8, 14, 
    10, 0, 2, 4, 3, 4, 0, 0, 0, 0, 0, 6, 7, 8, 13, 
    
    -- channel=93
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 11, 8, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 6, 41, 33, 8, 4, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 1, 5, 10, 0, 0, 0, 0, 0, 0, 
    
    -- channel=94
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 1, 1, 1, 1, 
    1, 1, 1, 1, 2, 2, 1, 1, 1, 0, 1, 3, 2, 2, 2, 
    0, 0, 1, 2, 2, 0, 1, 0, 0, 1, 0, 0, 1, 1, 1, 
    7, 5, 3, 1, 1, 0, 1, 5, 17, 23, 27, 17, 3, 3, 3, 
    0, 0, 0, 0, 0, 3, 7, 4, 8, 2, 0, 0, 0, 0, 2, 
    20, 22, 7, 0, 0, 0, 0, 0, 0, 9, 21, 24, 26, 20, 4, 
    0, 0, 0, 5, 9, 15, 30, 40, 24, 0, 0, 0, 0, 0, 0, 
    15, 24, 7, 4, 9, 23, 25, 3, 0, 9, 21, 25, 27, 27, 16, 
    32, 12, 12, 11, 4, 0, 0, 0, 5, 0, 0, 0, 0, 0, 3, 
    4, 0, 1, 3, 8, 10, 19, 21, 18, 18, 15, 15, 15, 12, 11, 
    4, 8, 7, 0, 0, 0, 0, 0, 3, 5, 10, 15, 25, 19, 9, 
    0, 1, 4, 5, 4, 5, 43, 52, 47, 45, 42, 24, 1, 0, 8, 
    2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 5, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 5, 0, 2, 4, 
    0, 3, 3, 4, 4, 5, 0, 0, 11, 5, 0, 0, 0, 3, 6, 
    
    -- channel=95
    101, 98, 98, 98, 98, 98, 98, 99, 97, 99, 98, 98, 98, 98, 98, 
    101, 98, 98, 98, 98, 98, 97, 98, 98, 107, 69, 84, 99, 98, 98, 
    99, 97, 98, 99, 98, 101, 95, 106, 89, 90, 53, 68, 100, 98, 98, 
    89, 98, 96, 98, 100, 112, 75, 112, 89, 92, 79, 57, 99, 98, 99, 
    50, 43, 64, 95, 98, 105, 80, 100, 94, 108, 102, 86, 72, 47, 95, 
    86, 80, 77, 84, 85, 88, 69, 74, 75, 105, 96, 89, 96, 43, 89, 
    45, 26, 56, 73, 99, 98, 16, 20, 37, 94, 96, 90, 77, 77, 56, 
    0, 38, 53, 20, 76, 100, 76, 96, 68, 65, 61, 47, 42, 55, 59, 
    0, 74, 81, 70, 80, 97, 86, 107, 82, 81, 80, 84, 67, 61, 61, 
    10, 61, 56, 61, 62, 63, 67, 59, 51, 64, 45, 51, 36, 37, 36, 
    3, 0, 9, 5, 2, 5, 20, 24, 31, 30, 24, 19, 21, 37, 32, 
    4, 0, 23, 12, 0, 0, 0, 39, 19, 18, 19, 34, 40, 39, 27, 
    8, 0, 0, 0, 0, 0, 0, 62, 57, 52, 35, 16, 20, 24, 33, 
    51, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 9, 30, 29, 40, 
    48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 32, 30, 38, 48, 
    
    -- channel=96
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=97
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 
    0, 0, 0, 0, 0, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 18, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 
    12, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 4, 10, 6, 0, 0, 23, 13, 7, 0, 0, 0, 0, 0, 
    22, 0, 0, 12, 6, 1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    48, 2, 0, 4, 2, 1, 0, 0, 5, 5, 0, 0, 0, 0, 0, 
    43, 8, 4, 5, 4, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=98
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 18, 14, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    49, 46, 3, 0, 0, 0, 0, 0, 0, 0, 8, 33, 41, 33, 0, 
    0, 0, 0, 9, 6, 39, 53, 44, 31, 0, 0, 0, 0, 0, 0, 
    56, 60, 24, 0, 0, 10, 0, 0, 0, 0, 19, 37, 36, 31, 31, 
    23, 0, 3, 0, 1, 0, 0, 0, 27, 22, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 8, 17, 0, 0, 3, 8, 26, 38, 31, 
    0, 49, 44, 44, 37, 30, 20, 10, 6, 9, 12, 18, 0, 0, 0, 
    29, 29, 31, 46, 55, 62, 58, 55, 48, 43, 31, 18, 1, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 1, 17, 15, 4, 0, 2, 23, 3, 6, 28, 28, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 16, 8, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=99
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 11, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 6, 29, 14, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    80, 64, 0, 0, 0, 0, 0, 0, 0, 0, 13, 41, 56, 27, 0, 
    0, 0, 0, 24, 9, 52, 43, 32, 16, 0, 0, 0, 0, 0, 0, 
    75, 77, 31, 0, 0, 26, 12, 0, 0, 0, 20, 37, 24, 33, 31, 
    5, 0, 21, 17, 0, 0, 0, 0, 47, 41, 22, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 10, 0, 0, 0, 0, 0, 17, 43, 36, 
    0, 50, 53, 53, 47, 38, 29, 24, 21, 15, 24, 20, 1, 0, 0, 
    62, 48, 63, 70, 76, 76, 68, 60, 49, 48, 34, 20, 1, 0, 0, 
    3, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 28, 17, 3, 0, 21, 0, 0, 0, 35, 35, 0, 0, 0, 
    0, 0, 1, 1, 0, 0, 9, 17, 42, 17, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=100
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 23, 23, 18, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 14, 64, 48, 12, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=101
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 25, 39, 50, 21, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 11, 1, 11, 0, 0, 0, 0, 0, 0, 
    68, 71, 12, 0, 0, 0, 0, 0, 0, 0, 33, 58, 64, 39, 0, 
    0, 0, 0, 0, 9, 10, 6, 33, 33, 0, 0, 0, 0, 0, 0, 
    0, 51, 0, 0, 0, 69, 87, 14, 0, 0, 0, 17, 30, 39, 29, 
    49, 16, 55, 37, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 3, 
    0, 0, 16, 23, 7, 0, 47, 96, 58, 58, 65, 57, 12, 0, 13, 
    25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 13, 11, 
    23, 3, 0, 0, 1, 1, 0, 0, 0, 0, 28, 31, 2, 2, 0, 
    5, 24, 18, 15, 16, 16, 11, 0, 32, 41, 10, 0, 3, 7, 4, 
    
    -- channel=102
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    13, 9, 1, 0, 0, 0, 0, 0, 0, 0, 0, 4, 8, 0, 0, 
    0, 0, 0, 3, 1, 6, 3, 1, 0, 0, 0, 0, 0, 5, 0, 
    12, 7, 4, 0, 0, 10, 9, 7, 7, 0, 0, 3, 0, 0, 1, 
    2, 12, 11, 7, 0, 0, 0, 2, 4, 3, 6, 6, 4, 0, 6, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 4, 6, 4, 
    22, 17, 17, 17, 18, 13, 7, 5, 5, 5, 6, 6, 2, 7, 7, 
    23, 17, 11, 17, 21, 20, 0, 5, 5, 5, 3, 5, 6, 5, 7, 
    25, 30, 22, 21, 24, 25, 14, 0, 0, 2, 9, 8, 13, 8, 8, 
    23, 25, 24, 22, 24, 24, 30, 3, 0, 2, 10, 13, 11, 12, 6, 
    21, 26, 25, 25, 24, 24, 30, 8, 10, 15, 14, 15, 12, 10, 6, 
    
    -- channel=103
    9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 10, 9, 9, 9, 
    9, 9, 9, 9, 9, 9, 9, 10, 10, 7, 7, 9, 9, 9, 9, 
    9, 9, 9, 9, 9, 9, 9, 9, 6, 0, 5, 8, 9, 9, 9, 
    7, 8, 10, 10, 9, 9, 8, 4, 0, 0, 0, 6, 9, 9, 10, 
    3, 6, 9, 10, 10, 8, 10, 7, 4, 1, 1, 3, 6, 7, 9, 
    0, 0, 10, 9, 10, 6, 7, 6, 6, 3, 0, 0, 0, 2, 8, 
    0, 0, 3, 1, 4, 0, 0, 0, 1, 6, 3, 3, 2, 5, 5, 
    0, 0, 0, 7, 1, 0, 0, 2, 4, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 3, 5, 6, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 3, 0, 4, 5, 
    0, 0, 0, 0, 0, 0, 1, 22, 17, 15, 7, 8, 7, 5, 6, 
    0, 0, 0, 0, 0, 0, 0, 15, 10, 8, 9, 7, 6, 6, 6, 
    
    -- channel=104
    72, 71, 71, 71, 71, 71, 71, 71, 70, 72, 72, 71, 71, 71, 71, 
    72, 71, 71, 72, 71, 71, 71, 72, 73, 79, 66, 68, 71, 71, 72, 
    71, 70, 71, 72, 71, 73, 71, 77, 73, 77, 52, 61, 73, 71, 72, 
    74, 75, 73, 71, 71, 81, 63, 80, 71, 73, 67, 58, 77, 75, 74, 
    60, 55, 68, 68, 71, 80, 64, 75, 70, 78, 77, 72, 65, 55, 75, 
    61, 57, 62, 60, 69, 64, 60, 62, 65, 86, 79, 69, 70, 48, 72, 
    53, 43, 61, 61, 81, 66, 40, 44, 46, 69, 68, 64, 62, 61, 55, 
    13, 46, 41, 36, 70, 72, 56, 65, 61, 65, 62, 55, 50, 58, 54, 
    0, 67, 60, 55, 64, 77, 76, 82, 63, 62, 66, 66, 59, 59, 62, 
    27, 58, 59, 62, 63, 66, 71, 62, 59, 59, 53, 54, 45, 43, 41, 
    18, 19, 23, 21, 19, 22, 33, 36, 41, 38, 37, 33, 36, 38, 33, 
    11, 0, 19, 11, 1, 0, 16, 36, 30, 27, 23, 25, 20, 30, 34, 
    10, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 12, 23, 30, 42, 
    35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 16, 33, 36, 49, 
    36, 3, 2, 1, 0, 0, 0, 0, 0, 1, 24, 36, 37, 42, 52, 
    
    -- channel=105
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 3, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 1, 7, 12, 9, 4, 0, 1, 0, 0, 0, 6, 1, 0, 0, 
    26, 7, 6, 9, 7, 6, 1, 19, 27, 18, 4, 0, 0, 0, 0, 
    30, 11, 7, 8, 7, 6, 1, 12, 8, 0, 0, 0, 0, 0, 0, 
    
    -- channel=106
    129, 129, 129, 129, 129, 129, 129, 130, 129, 129, 129, 128, 129, 129, 129, 
    130, 130, 130, 130, 129, 129, 129, 129, 129, 125, 121, 128, 129, 129, 130, 
    130, 130, 131, 130, 130, 131, 127, 128, 114, 100, 94, 121, 130, 130, 131, 
    122, 124, 128, 131, 132, 134, 124, 121, 94, 86, 78, 100, 127, 128, 129, 
    93, 98, 130, 130, 131, 127, 118, 126, 119, 122, 114, 108, 107, 111, 129, 
    68, 75, 110, 115, 128, 111, 115, 118, 119, 121, 93, 81, 74, 87, 125, 
    81, 86, 105, 99, 107, 37, 28, 48, 86, 123, 120, 114, 113, 109, 109, 
    13, 54, 54, 94, 110, 79, 74, 93, 100, 90, 67, 57, 55, 67, 74, 
    16, 98, 77, 92, 111, 120, 123, 102, 79, 78, 86, 82, 80, 83, 82, 
    60, 85, 86, 87, 86, 85, 78, 64, 68, 52, 53, 45, 37, 39, 53, 
    7, 19, 21, 23, 30, 38, 45, 41, 42, 34, 26, 23, 28, 38, 51, 
    0, 0, 6, 0, 0, 0, 5, 0, 0, 0, 9, 30, 46, 54, 57, 
    0, 0, 2, 0, 0, 0, 29, 103, 91, 83, 70, 60, 47, 51, 70, 
    0, 0, 0, 0, 0, 0, 0, 91, 77, 45, 29, 37, 52, 59, 80, 
    4, 0, 0, 0, 0, 0, 0, 27, 17, 29, 52, 50, 55, 64, 82, 
    
    -- channel=107
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 10, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 7, 0, 0, 0, 
    0, 15, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 
    0, 0, 0, 0, 0, 0, 5, 4, 7, 0, 0, 0, 0, 20, 0, 
    2, 28, 2, 0, 0, 0, 3, 9, 18, 0, 0, 0, 0, 0, 18, 
    37, 1, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    91, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    37, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 17, 1, 11, 17, 24, 13, 11, 1, 0, 0, 3, 6, 0, 5, 
    0, 31, 0, 0, 0, 14, 31, 0, 0, 0, 0, 0, 1, 0, 9, 
    0, 15, 12, 0, 0, 6, 94, 1, 4, 0, 6, 9, 4, 8, 11, 
    0, 2, 7, 3, 3, 4, 47, 29, 25, 27, 15, 12, 0, 7, 8, 
    0, 0, 0, 0, 0, 2, 16, 25, 19, 21, 0, 0, 1, 2, 4, 
    
    -- channel=108
    19, 18, 18, 18, 18, 18, 18, 18, 17, 18, 19, 18, 18, 18, 18, 
    19, 18, 18, 18, 18, 18, 18, 17, 19, 31, 21, 18, 18, 18, 18, 
    20, 19, 18, 18, 18, 19, 19, 26, 33, 30, 22, 17, 19, 18, 18, 
    21, 20, 19, 18, 18, 23, 16, 21, 14, 13, 8, 10, 21, 20, 19, 
    44, 37, 18, 19, 19, 16, 11, 17, 17, 26, 36, 40, 41, 24, 20, 
    3, 1, 11, 26, 24, 45, 41, 37, 29, 23, 14, 6, 7, 3, 19, 
    47, 39, 32, 13, 19, 31, 10, 0, 6, 25, 35, 39, 32, 33, 29, 
    3, 0, 13, 9, 15, 2, 0, 21, 30, 28, 21, 10, 5, 4, 13, 
    0, 7, 1, 5, 19, 28, 32, 33, 20, 30, 28, 35, 37, 37, 33, 
    20, 49, 51, 53, 50, 46, 43, 35, 34, 35, 33, 32, 22, 20, 15, 
    20, 15, 28, 31, 33, 37, 46, 46, 42, 38, 31, 24, 14, 9, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    
    -- channel=109
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 16, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 14, 0, 21, 5, 11, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 16, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 16, 15, 8, 29, 0, 0, 
    0, 0, 0, 0, 16, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 29, 0, 0, 0, 7, 12, 1, 0, 0, 0, 
    0, 0, 6, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 10, 0, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 22, 19, 6, 0, 0, 14, 1, 0, 0, 0, 0, 0, 0, 
    21, 0, 0, 11, 7, 0, 0, 20, 12, 6, 0, 0, 0, 0, 0, 
    61, 1, 0, 4, 1, 0, 0, 0, 5, 5, 0, 0, 0, 0, 0, 
    56, 8, 2, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=110
    12, 11, 11, 11, 11, 11, 11, 11, 11, 11, 10, 11, 11, 11, 11, 
    10, 10, 10, 10, 9, 10, 9, 10, 8, 0, 0, 2, 10, 10, 10, 
    6, 7, 10, 10, 11, 11, 6, 0, 0, 0, 0, 0, 9, 10, 10, 
    8, 9, 8, 10, 10, 7, 0, 16, 34, 43, 44, 17, 8, 9, 9, 
    0, 0, 0, 5, 7, 17, 19, 17, 22, 15, 0, 0, 0, 0, 6, 
    78, 78, 21, 0, 0, 0, 0, 0, 0, 12, 39, 61, 64, 36, 7, 
    0, 0, 0, 16, 27, 0, 0, 11, 23, 3, 0, 0, 0, 0, 0, 
    0, 53, 0, 0, 2, 76, 89, 18, 0, 0, 0, 8, 18, 37, 25, 
    35, 41, 67, 50, 18, 0, 0, 6, 29, 11, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 7, 
    0, 0, 29, 22, 2, 0, 55, 66, 37, 38, 50, 55, 21, 0, 15, 
    14, 0, 0, 0, 0, 0, 0, 4, 27, 12, 0, 0, 8, 17, 16, 
    22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 29, 8, 7, 8, 
    6, 17, 13, 9, 10, 10, 0, 0, 26, 37, 18, 4, 10, 14, 13, 
    
    -- channel=111
    82, 81, 81, 81, 81, 81, 81, 82, 81, 81, 82, 81, 81, 81, 81, 
    82, 82, 82, 82, 81, 81, 81, 82, 80, 74, 69, 78, 82, 81, 82, 
    81, 81, 82, 82, 82, 82, 80, 78, 63, 57, 50, 72, 82, 82, 82, 
    78, 80, 81, 82, 83, 81, 73, 76, 66, 64, 60, 65, 81, 81, 82, 
    38, 43, 75, 80, 82, 80, 74, 80, 78, 79, 68, 57, 51, 58, 82, 
    57, 63, 70, 63, 71, 53, 53, 59, 67, 78, 67, 62, 59, 58, 79, 
    29, 31, 51, 62, 67, 24, 11, 30, 55, 74, 67, 58, 56, 54, 56, 
    0, 34, 25, 42, 65, 64, 61, 58, 49, 46, 37, 33, 33, 45, 48, 
    5, 63, 59, 62, 71, 74, 70, 63, 53, 48, 53, 47, 41, 39, 41, 
    22, 39, 40, 44, 45, 47, 46, 38, 36, 30, 25, 22, 17, 18, 26, 
    0, 0, 0, 0, 0, 0, 3, 5, 8, 5, 1, 1, 11, 19, 23, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 8, 19, 20, 21, 26, 
    0, 0, 0, 0, 0, 0, 0, 49, 44, 33, 16, 9, 11, 19, 35, 
    0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 6, 17, 24, 41, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 15, 20, 30, 45, 
    
    -- channel=112
    99, 99, 99, 99, 99, 100, 100, 100, 99, 99, 99, 100, 99, 99, 100, 
    101, 100, 100, 100, 100, 100, 101, 100, 100, 100, 105, 102, 100, 100, 101, 
    102, 101, 101, 101, 100, 100, 101, 100, 103, 86, 88, 103, 101, 101, 102, 
    98, 99, 103, 101, 101, 100, 102, 90, 71, 62, 57, 86, 102, 102, 103, 
    110, 113, 110, 103, 102, 94, 92, 95, 91, 93, 99, 107, 110, 112, 105, 
    37, 44, 85, 101, 105, 107, 114, 112, 110, 95, 69, 53, 42, 69, 102, 
    96, 104, 101, 77, 76, 41, 41, 49, 70, 97, 103, 104, 100, 100, 107, 
    28, 31, 59, 86, 88, 41, 39, 73, 97, 87, 64, 50, 48, 49, 62, 
    17, 65, 44, 61, 85, 100, 106, 81, 60, 65, 69, 70, 79, 90, 84, 
    59, 89, 92, 92, 90, 86, 76, 64, 66, 52, 56, 48, 38, 42, 51, 
    32, 37, 39, 45, 53, 60, 59, 59, 55, 45, 38, 33, 32, 31, 43, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 28, 43, 47, 
    0, 0, 11, 0, 0, 0, 52, 46, 26, 27, 42, 48, 33, 41, 59, 
    0, 0, 0, 0, 0, 0, 3, 17, 18, 21, 10, 24, 44, 53, 71, 
    7, 0, 0, 0, 0, 0, 0, 12, 0, 14, 36, 46, 49, 56, 72, 
    
    -- channel=113
    92, 92, 92, 92, 91, 91, 92, 91, 91, 91, 91, 92, 92, 92, 92, 
    91, 91, 91, 91, 90, 91, 90, 91, 88, 62, 55, 83, 91, 91, 91, 
    86, 88, 91, 92, 92, 91, 88, 76, 48, 54, 49, 68, 91, 91, 92, 
    91, 94, 92, 91, 92, 80, 74, 91, 97, 105, 107, 98, 92, 93, 93, 
    0, 0, 60, 85, 89, 99, 97, 98, 98, 89, 55, 23, 7, 37, 88, 
    126, 126, 94, 53, 55, 17, 4, 19, 47, 87, 108, 121, 114, 96, 89, 
    0, 0, 24, 78, 89, 41, 30, 68, 90, 76, 46, 21, 26, 22, 29, 
    8, 77, 36, 32, 74, 127, 139, 76, 22, 30, 45, 62, 74, 94, 84, 
    68, 108, 119, 112, 89, 71, 57, 67, 80, 59, 58, 44, 18, 6, 17, 
    13, 0, 0, 0, 1, 15, 26, 29, 28, 27, 14, 15, 26, 28, 34, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 44, 43, 
    0, 0, 23, 13, 0, 0, 49, 77, 49, 50, 63, 69, 37, 35, 58, 
    12, 0, 0, 0, 0, 0, 0, 9, 25, 15, 0, 0, 42, 55, 68, 
    22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 56, 46, 51, 64, 
    22, 11, 5, 1, 1, 3, 0, 5, 42, 56, 47, 43, 52, 62, 72, 
    
    -- channel=114
    8, 8, 8, 8, 8, 8, 8, 8, 6, 8, 9, 9, 8, 8, 8, 
    7, 6, 6, 6, 6, 6, 6, 5, 6, 8, 0, 0, 6, 5, 6, 
    8, 7, 5, 5, 6, 7, 7, 9, 0, 1, 20, 9, 7, 6, 6, 
    6, 8, 8, 6, 7, 7, 0, 0, 2, 2, 0, 1, 9, 8, 7, 
    0, 0, 0, 6, 5, 5, 11, 9, 12, 16, 26, 6, 0, 0, 6, 
    46, 43, 24, 9, 6, 33, 31, 29, 18, 0, 0, 13, 13, 11, 9, 
    0, 0, 0, 8, 20, 0, 0, 0, 0, 24, 29, 23, 23, 19, 0, 
    0, 7, 0, 0, 0, 11, 38, 32, 0, 0, 0, 0, 0, 0, 16, 
    0, 39, 44, 52, 38, 22, 19, 36, 43, 54, 47, 49, 35, 4, 0, 
    51, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 12, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    5, 8, 21, 11, 2, 0, 0, 0, 0, 0, 0, 8, 33, 0, 0, 
    4, 0, 0, 0, 0, 0, 1, 10, 21, 23, 9, 0, 0, 7, 6, 
    10, 0, 0, 0, 0, 0, 7, 16, 6, 0, 0, 19, 3, 2, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 11, 2, 5, 6, 6, 
    
    -- channel=115
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 9, 18, 15, 3, 0, 25, 11, 7, 1, 0, 0, 0, 0, 
    29, 9, 0, 9, 14, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 16, 13, 15, 15, 15, 0, 0, 0, 3, 8, 2, 0, 0, 0, 
    29, 24, 21, 20, 19, 19, 13, 12, 15, 5, 0, 0, 0, 0, 0, 
    
    -- channel=116
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 5, 15, 0, 0, 
    0, 0, 0, 0, 7, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 13, 4, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 11, 12, 3, 0, 6, 24, 14, 11, 9, 7, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 
    23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 5, 3, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=117
    27, 28, 28, 28, 28, 28, 28, 27, 28, 28, 29, 28, 28, 28, 28, 
    29, 29, 29, 29, 29, 29, 30, 29, 29, 27, 44, 36, 29, 29, 30, 
    28, 29, 30, 29, 29, 28, 31, 28, 36, 25, 32, 38, 30, 29, 30, 
    33, 31, 31, 29, 29, 25, 38, 22, 20, 18, 22, 41, 31, 31, 31, 
    65, 63, 46, 30, 31, 23, 29, 24, 27, 24, 27, 40, 46, 54, 34, 
    0, 0, 27, 29, 33, 23, 33, 32, 37, 31, 20, 7, 1, 31, 35, 
    52, 64, 44, 20, 15, 8, 36, 46, 38, 25, 24, 27, 25, 31, 47, 
    21, 11, 23, 49, 36, 0, 0, 15, 45, 46, 36, 28, 26, 19, 21, 
    27, 7, 0, 0, 19, 28, 33, 3, 2, 4, 9, 9, 21, 40, 40, 
    24, 41, 50, 50, 52, 48, 42, 40, 38, 24, 33, 23, 18, 14, 22, 
    25, 36, 33, 37, 39, 42, 41, 37, 32, 28, 25, 22, 25, 13, 15, 
    0, 0, 0, 0, 0, 0, 5, 0, 11, 8, 4, 0, 0, 10, 13, 
    0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 0, 17, 1, 5, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 12, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 5, 11, 23, 
    
    -- channel=118
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 9, 0, 13, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 18, 0, 19, 0, 12, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 9, 7, 4, 31, 0, 0, 
    0, 0, 0, 0, 32, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 0, 0, 11, 0, 22, 0, 2, 12, 0, 0, 0, 0, 
    0, 11, 0, 0, 0, 1, 0, 12, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 4, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 0, 12, 24, 9, 0, 0, 32, 9, 0, 0, 0, 0, 0, 0, 
    37, 0, 0, 9, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    73, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    62, 10, 4, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=119
    4, 3, 3, 3, 3, 3, 3, 3, 4, 4, 3, 3, 3, 3, 3, 
    4, 3, 3, 4, 3, 4, 3, 4, 5, 13, 2, 1, 3, 3, 3, 
    4, 3, 3, 4, 2, 5, 3, 11, 12, 18, 0, 0, 4, 4, 3, 
    2, 3, 4, 3, 2, 12, 2, 14, 3, 1, 0, 0, 5, 5, 4, 
    14, 10, 3, 3, 4, 10, 0, 5, 0, 9, 12, 14, 16, 0, 4, 
    0, 0, 0, 7, 12, 17, 14, 12, 3, 11, 9, 0, 1, 0, 0, 
    13, 1, 11, 5, 7, 27, 0, 0, 0, 2, 10, 15, 14, 8, 2, 
    0, 0, 4, 0, 9, 10, 0, 0, 9, 12, 10, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 10, 21, 3, 2, 5, 8, 6, 8, 12, 
    0, 7, 2, 2, 2, 2, 1, 0, 0, 6, 0, 7, 0, 0, 0, 
    12, 7, 8, 10, 10, 8, 7, 3, 5, 4, 4, 0, 0, 0, 0, 
    18, 0, 10, 10, 8, 3, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    17, 5, 6, 14, 12, 7, 0, 0, 0, 0, 0, 5, 8, 0, 0, 
    33, 9, 7, 10, 9, 9, 0, 0, 0, 2, 3, 0, 6, 4, 0, 
    36, 15, 13, 12, 10, 9, 0, 0, 4, 0, 4, 13, 8, 4, 1, 
    
    -- channel=120
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 12, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 21, 13, 13, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    62, 61, 11, 0, 0, 0, 0, 0, 0, 0, 14, 41, 53, 39, 0, 
    0, 0, 0, 14, 15, 59, 74, 61, 34, 0, 0, 0, 0, 0, 0, 
    75, 75, 40, 0, 0, 0, 0, 0, 0, 0, 29, 48, 48, 40, 41, 
    15, 0, 0, 5, 0, 0, 0, 0, 31, 17, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 20, 14, 0, 5, 8, 16, 37, 46, 32, 
    15, 62, 59, 58, 48, 37, 21, 8, 10, 6, 16, 16, 1, 1, 0, 
    33, 34, 40, 60, 72, 79, 77, 72, 60, 51, 37, 19, 0, 0, 0, 
    6, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 24, 15, 2, 0, 31, 14, 0, 3, 31, 25, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 9, 9, 31, 11, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=121
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=122
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 
    0, 0, 0, 0, 0, 0, 8, 7, 8, 0, 0, 0, 0, 0, 0, 
    0, 18, 1, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    31, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 3, 9, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    1, 20, 0, 0, 0, 9, 11, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 10, 12, 5, 6, 6, 48, 20, 13, 8, 11, 18, 8, 0, 0, 
    0, 4, 8, 6, 6, 6, 47, 49, 48, 39, 17, 1, 0, 1, 0, 
    0, 0, 0, 0, 2, 2, 16, 25, 19, 9, 0, 0, 0, 0, 0, 
    
    -- channel=123
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 11, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 11, 0, 0, 
    0, 0, 0, 0, 2, 0, 5, 1, 0, 0, 0, 0, 0, 0, 0, 
    22, 16, 7, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 12, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 9, 7, 8, 6, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 21, 21, 25, 26, 23, 20, 14, 12, 11, 5, 0, 0, 0, 0, 
    8, 0, 0, 0, 3, 2, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 7, 24, 19, 10, 6, 6, 48, 33, 29, 32, 30, 3, 0, 0, 
    8, 6, 9, 9, 7, 6, 23, 83, 68, 41, 3, 0, 0, 0, 0, 
    8, 0, 0, 1, 2, 0, 9, 37, 6, 0, 0, 0, 0, 0, 0, 
    
    -- channel=124
    57, 57, 57, 57, 57, 57, 57, 57, 56, 58, 58, 57, 57, 57, 57, 
    57, 57, 57, 57, 57, 57, 57, 57, 57, 60, 55, 57, 57, 57, 58, 
    57, 58, 57, 57, 57, 58, 58, 60, 57, 51, 55, 57, 58, 57, 58, 
    60, 59, 58, 57, 58, 58, 53, 52, 47, 48, 44, 56, 60, 59, 59, 
    47, 49, 56, 56, 58, 57, 56, 57, 57, 60, 64, 57, 53, 52, 59, 
    45, 47, 63, 54, 55, 63, 60, 60, 60, 56, 46, 45, 42, 49, 61, 
    46, 47, 52, 43, 59, 19, 23, 24, 46, 63, 62, 57, 55, 57, 54, 
    17, 28, 28, 41, 46, 35, 44, 58, 49, 41, 33, 30, 32, 37, 46, 
    11, 63, 45, 56, 64, 64, 65, 55, 50, 58, 56, 58, 54, 50, 43, 
    58, 54, 58, 59, 57, 57, 55, 47, 50, 39, 45, 37, 35, 35, 35, 
    7, 10, 17, 18, 20, 26, 37, 39, 37, 34, 29, 26, 25, 26, 29, 
    0, 0, 1, 0, 0, 0, 1, 8, 9, 8, 10, 21, 30, 22, 26, 
    0, 0, 0, 0, 0, 0, 13, 15, 15, 18, 19, 10, 10, 23, 33, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 20, 25, 39, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 18, 18, 22, 29, 40, 
    
    -- channel=125
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 8, 12, 11, 4, 0, 5, 0, 0, 0, 0, 0, 2, 0, 
    19, 0, 7, 17, 12, 8, 0, 35, 37, 31, 18, 18, 11, 0, 0, 
    25, 11, 9, 12, 10, 10, 3, 42, 58, 37, 21, 3, 3, 0, 0, 
    31, 16, 12, 11, 12, 11, 3, 23, 27, 8, 6, 4, 0, 0, 0, 
    
    -- channel=126
    50, 50, 50, 50, 50, 51, 51, 51, 50, 50, 50, 50, 50, 50, 50, 
    51, 51, 51, 51, 50, 50, 50, 51, 50, 52, 44, 49, 51, 50, 50, 
    51, 52, 51, 50, 51, 52, 49, 51, 41, 33, 33, 45, 50, 50, 51, 
    44, 46, 48, 51, 53, 55, 44, 42, 26, 21, 17, 28, 47, 47, 48, 
    27, 29, 46, 52, 51, 47, 43, 47, 43, 44, 43, 38, 39, 34, 47, 
    18, 24, 42, 48, 50, 49, 48, 48, 44, 39, 22, 20, 21, 26, 45, 
    29, 29, 38, 32, 38, 2, 0, 0, 23, 49, 50, 48, 45, 43, 38, 
    0, 8, 11, 30, 30, 18, 17, 35, 35, 28, 15, 8, 6, 12, 19, 
    0, 34, 28, 38, 46, 48, 46, 38, 25, 28, 30, 30, 29, 25, 23, 
    24, 34, 32, 35, 33, 30, 26, 18, 20, 14, 12, 9, 4, 7, 13, 
    0, 0, 0, 1, 4, 7, 13, 14, 13, 10, 2, 0, 0, 6, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 23, 17, 13, 
    0, 0, 0, 0, 0, 0, 14, 83, 78, 69, 53, 28, 14, 11, 15, 
    0, 0, 0, 0, 0, 0, 16, 113, 91, 39, 11, 11, 12, 11, 18, 
    0, 0, 0, 0, 0, 0, 0, 27, 9, 9, 16, 9, 10, 12, 19, 
    
    -- channel=127
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 21, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 16, 0, 0, 0, 4, 47, 0, 0, 0, 
    0, 5, 27, 0, 0, 0, 19, 0, 6, 0, 0, 0, 0, 22, 3, 
    4, 24, 22, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 67, 7, 
    0, 7, 1, 5, 0, 0, 12, 37, 64, 0, 0, 0, 0, 0, 12, 
    26, 51, 0, 50, 0, 0, 35, 0, 0, 0, 0, 0, 14, 13, 30, 
    142, 3, 6, 25, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 13, 
    0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 10, 19, 
    0, 37, 0, 0, 0, 13, 50, 0, 8, 12, 25, 28, 14, 0, 24, 
    0, 16, 3, 0, 0, 4, 117, 0, 0, 0, 0, 0, 8, 22, 34, 
    0, 1, 5, 0, 0, 2, 62, 13, 0, 0, 17, 33, 7, 21, 28, 
    0, 0, 2, 1, 3, 4, 29, 9, 14, 44, 13, 0, 13, 19, 26, 
    
    -- channel=128
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=129
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 3, 4, 2, 1, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 1, 9, 6, 10, 2, 0, 0, 0, 0, 0, 1, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 5, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 10, 11, 11, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 15, 14, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 4, 2, 0, 4, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 1, 3, 
    3, 2, 1, 0, 2, 2, 0, 1, 0, 2, 0, 0, 1, 1, 6, 
    
    -- channel=130
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 5, 11, 8, 0, 0, 
    3, 9, 8, 1, 0, 0, 0, 0, 5, 7, 11, 17, 0, 13, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 1, 0, 1, 
    1, 3, 10, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 6, 0, 0, 1, 3, 
    0, 5, 2, 0, 0, 0, 3, 2, 3, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 5, 8, 11, 
    1, 0, 0, 0, 0, 0, 7, 11, 3, 0, 8, 6, 6, 10, 11, 
    7, 5, 8, 9, 2, 0, 3, 11, 10, 5, 10, 12, 10, 12, 14, 
    3, 4, 10, 14, 15, 12, 6, 8, 16, 11, 11, 11, 13, 14, 15, 
    15, 15, 13, 12, 14, 16, 15, 14, 13, 9, 13, 12, 15, 15, 15, 
    
    -- channel=131
    27, 38, 35, 31, 27, 24, 22, 16, 24, 21, 16, 19, 19, 19, 20, 
    24, 32, 30, 22, 20, 19, 19, 17, 21, 16, 27, 20, 16, 16, 20, 
    16, 26, 23, 14, 15, 14, 12, 19, 21, 1, 38, 19, 11, 12, 18, 
    7, 19, 12, 6, 3, 9, 5, 10, 22, 21, 40, 42, 26, 7, 9, 
    17, 20, 19, 22, 14, 17, 19, 16, 17, 19, 23, 14, 16, 6, 22, 
    26, 23, 13, 22, 23, 27, 29, 23, 22, 20, 25, 11, 2, 3, 7, 
    30, 23, 22, 35, 37, 30, 35, 29, 32, 29, 28, 15, 0, 12, 0, 
    29, 23, 24, 32, 32, 33, 31, 29, 25, 15, 20, 14, 10, 0, 10, 
    34, 27, 42, 37, 35, 33, 33, 28, 28, 7, 19, 16, 16, 11, 6, 
    32, 37, 32, 34, 34, 32, 26, 22, 20, 20, 20, 15, 12, 9, 14, 
    34, 36, 34, 24, 31, 30, 23, 22, 37, 24, 17, 15, 13, 11, 10, 
    43, 34, 27, 30, 31, 39, 12, 12, 22, 21, 18, 15, 16, 14, 7, 
    32, 24, 17, 19, 24, 25, 19, 19, 17, 17, 15, 18, 8, 13, 11, 
    21, 20, 18, 18, 16, 16, 20, 17, 19, 13, 13, 13, 12, 13, 11, 
    9, 12, 16, 17, 17, 16, 17, 10, 24, 7, 13, 11, 13, 13, 3, 
    
    -- channel=132
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=133
    19, 28, 41, 34, 35, 29, 33, 26, 36, 34, 27, 32, 24, 31, 30, 
    17, 25, 40, 25, 34, 24, 31, 33, 32, 19, 31, 36, 22, 32, 30, 
    14, 18, 35, 18, 30, 20, 22, 31, 33, 0, 49, 43, 20, 30, 33, 
    11, 11, 29, 24, 21, 21, 14, 12, 11, 0, 16, 18, 48, 30, 28, 
    12, 9, 11, 25, 17, 22, 17, 9, 0, 3, 8, 0, 18, 3, 8, 
    6, 1, 0, 1, 6, 2, 15, 1, 5, 1, 10, 17, 0, 24, 0, 
    15, 0, 0, 20, 21, 6, 11, 1, 3, 7, 26, 23, 0, 5, 0, 
    7, 2, 9, 22, 25, 24, 23, 19, 25, 6, 22, 17, 6, 0, 0, 
    18, 20, 29, 32, 28, 27, 23, 12, 16, 0, 15, 11, 8, 0, 15, 
    0, 20, 29, 23, 17, 18, 20, 18, 19, 19, 16, 9, 8, 0, 0, 
    28, 20, 20, 14, 29, 30, 7, 0, 12, 25, 13, 0, 0, 0, 0, 
    39, 18, 5, 0, 3, 32, 4, 0, 6, 0, 0, 0, 0, 0, 0, 
    26, 16, 7, 7, 8, 4, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 
    
    -- channel=134
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 46, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 12, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 7, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 6, 0, 0, 0, 0, 33, 0, 39, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 59, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 54, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 4, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 12, 0, 
    0, 0, 0, 1, 0, 0, 8, 13, 0, 0, 0, 6, 7, 6, 3, 
    0, 0, 7, 0, 0, 0, 11, 10, 0, 0, 4, 2, 3, 3, 9, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 3, 0, 13, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 2, 3, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 4, 0, 30, 0, 2, 0, 0, 18, 
    
    -- channel=135
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=136
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=137
    62, 60, 59, 57, 50, 45, 40, 37, 38, 36, 35, 34, 37, 36, 35, 
    52, 49, 45, 42, 36, 35, 31, 31, 35, 36, 23, 30, 33, 30, 31, 
    41, 39, 33, 29, 25, 27, 25, 23, 24, 33, 24, 27, 26, 20, 25, 
    26, 24, 15, 9, 10, 14, 16, 26, 35, 21, 37, 18, 2, 8, 6, 
    12, 19, 10, 7, 1, 6, 15, 25, 36, 42, 42, 22, 25, 8, 7, 
    34, 35, 36, 32, 39, 41, 49, 47, 42, 40, 37, 33, 27, 0, 28, 
    46, 39, 33, 46, 46, 56, 59, 60, 59, 51, 36, 20, 9, 8, 14, 
    55, 50, 55, 65, 63, 64, 62, 59, 48, 37, 17, 10, 17, 27, 18, 
    54, 50, 48, 58, 61, 60, 55, 46, 40, 34, 31, 27, 26, 21, 11, 
    56, 57, 64, 58, 55, 55, 50, 42, 37, 34, 33, 28, 25, 16, 13, 
    58, 63, 57, 50, 46, 45, 47, 35, 32, 31, 29, 23, 22, 20, 17, 
    52, 55, 54, 45, 46, 43, 34, 36, 35, 28, 29, 28, 23, 23, 13, 
    41, 42, 35, 38, 36, 28, 26, 31, 29, 26, 23, 24, 21, 19, 19, 
    24, 21, 24, 24, 25, 25, 26, 24, 25, 32, 20, 20, 19, 20, 17, 
    14, 18, 21, 22, 24, 26, 27, 18, 22, 24, 19, 17, 20, 19, 12, 
    
    -- channel=138
    0, 0, 0, 0, 0, 0, 7, 1, 13, 11, 8, 13, 0, 8, 8, 
    0, 0, 12, 0, 11, 3, 15, 17, 13, 0, 31, 21, 2, 14, 12, 
    0, 0, 18, 1, 18, 6, 10, 29, 30, 0, 47, 38, 8, 23, 22, 
    2, 1, 27, 29, 24, 20, 12, 0, 7, 4, 7, 34, 80, 39, 40, 
    29, 19, 27, 44, 43, 45, 34, 12, 0, 0, 0, 0, 2, 2, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 22, 3, 0, 0, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 3, 0, 0, 6, 4, 9, 
    0, 0, 0, 0, 13, 15, 0, 0, 3, 18, 11, 2, 0, 0, 0, 
    13, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 4, 2, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 
    
    -- channel=139
    50, 47, 44, 44, 40, 37, 33, 31, 29, 32, 30, 29, 33, 29, 31, 
    43, 42, 34, 38, 29, 31, 28, 27, 28, 30, 30, 26, 31, 26, 28, 
    36, 36, 26, 28, 21, 26, 23, 21, 27, 30, 31, 23, 27, 20, 24, 
    27, 31, 18, 16, 12, 18, 18, 26, 27, 35, 26, 28, 23, 14, 12, 
    24, 24, 20, 15, 15, 16, 24, 31, 41, 36, 34, 34, 10, 8, 19, 
    30, 34, 28, 26, 29, 36, 39, 43, 36, 37, 33, 21, 22, 4, 25, 
    33, 38, 34, 33, 39, 46, 46, 47, 44, 39, 28, 16, 20, 11, 30, 
    44, 40, 43, 43, 45, 47, 49, 47, 41, 33, 19, 18, 21, 28, 21, 
    51, 37, 43, 49, 51, 48, 45, 42, 37, 33, 22, 22, 26, 30, 10, 
    49, 51, 42, 43, 48, 47, 42, 37, 33, 30, 29, 30, 25, 24, 22, 
    46, 49, 49, 46, 38, 38, 40, 36, 35, 30, 28, 29, 31, 26, 20, 
    37, 46, 44, 42, 40, 36, 38, 34, 28, 31, 32, 26, 30, 25, 22, 
    35, 39, 38, 36, 30, 30, 34, 32, 29, 26, 32, 25, 25, 23, 22, 
    26, 28, 28, 28, 26, 25, 26, 28, 29, 26, 24, 24, 24, 22, 22, 
    19, 19, 22, 23, 26, 26, 26, 22, 20, 31, 21, 23, 23, 22, 16, 
    
    -- channel=140
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=141
    20, 24, 19, 18, 14, 14, 9, 6, 8, 8, 9, 6, 7, 4, 7, 
    16, 20, 15, 12, 9, 8, 6, 8, 7, 2, 24, 5, 5, 4, 7, 
    12, 18, 11, 6, 1, 5, 0, 12, 17, 4, 22, 17, 6, 4, 6, 
    10, 14, 5, 7, 0, 2, 3, 0, 13, 31, 16, 27, 32, 8, 11, 
    25, 17, 19, 16, 17, 16, 21, 20, 22, 16, 20, 16, 0, 0, 9, 
    14, 14, 8, 15, 1, 9, 14, 23, 19, 16, 16, 0, 0, 0, 0, 
    15, 17, 21, 16, 21, 17, 16, 15, 7, 8, 4, 3, 3, 2, 11, 
    18, 11, 8, 8, 15, 18, 21, 19, 24, 14, 18, 6, 2, 0, 0, 
    26, 29, 31, 26, 26, 30, 29, 23, 15, 7, 0, 0, 7, 6, 9, 
    24, 17, 17, 23, 28, 20, 17, 19, 27, 16, 10, 8, 14, 17, 17, 
    32, 25, 24, 26, 28, 32, 15, 23, 22, 17, 21, 23, 18, 18, 7, 
    26, 28, 20, 26, 19, 18, 25, 19, 15, 19, 18, 20, 13, 13, 12, 
    26, 29, 33, 26, 23, 25, 21, 16, 19, 21, 18, 16, 13, 12, 10, 
    19, 23, 20, 19, 17, 18, 18, 17, 18, 7, 15, 10, 13, 10, 9, 
    9, 9, 11, 11, 12, 11, 13, 13, 16, 16, 9, 10, 11, 11, 3, 
    
    -- channel=142
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 21, 15, 62, 109, 0, 0, 0, 
    12, 18, 28, 36, 16, 14, 0, 0, 0, 0, 0, 0, 0, 0, 39, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 9, 26, 0, 0, 0, 0, 0, 3, 
    7, 0, 0, 4, 0, 11, 0, 0, 0, 2, 0, 0, 5, 5, 0, 
    4, 0, 0, 0, 14, 25, 0, 0, 2, 4, 0, 5, 0, 2, 0, 
    37, 27, 12, 5, 0, 3, 12, 8, 0, 0, 0, 5, 0, 1, 1, 
    0, 4, 6, 6, 0, 0, 0, 1, 14, 0, 5, 1, 3, 0, 9, 
    
    -- channel=143
    48, 41, 56, 47, 51, 42, 43, 42, 42, 42, 34, 40, 35, 43, 37, 
    40, 33, 46, 36, 43, 33, 39, 43, 37, 30, 28, 40, 32, 40, 36, 
    33, 21, 36, 29, 33, 29, 32, 25, 30, 20, 32, 38, 30, 33, 34, 
    26, 17, 27, 27, 21, 25, 20, 26, 14, 10, 16, 0, 28, 25, 15, 
    14, 11, 10, 11, 10, 12, 18, 19, 23, 25, 24, 17, 13, 18, 1, 
    25, 14, 21, 19, 30, 20, 36, 27, 25, 25, 25, 37, 8, 26, 0, 
    28, 18, 15, 32, 34, 38, 39, 36, 35, 31, 30, 21, 14, 0, 0, 
    35, 36, 45, 50, 50, 49, 47, 41, 40, 21, 19, 18, 18, 5, 17, 
    35, 33, 40, 51, 45, 43, 38, 31, 26, 27, 26, 22, 22, 16, 10, 
    31, 44, 47, 38, 42, 39, 36, 27, 26, 32, 28, 22, 14, 5, 5, 
    52, 42, 39, 33, 33, 42, 28, 9, 15, 25, 18, 11, 7, 3, 2, 
    41, 36, 32, 19, 26, 31, 21, 21, 18, 12, 7, 9, 2, 2, 0, 
    28, 26, 22, 22, 17, 10, 12, 13, 9, 10, 4, 4, 1, 1, 1, 
    4, 3, 5, 7, 7, 6, 7, 4, 11, 2, 3, 1, 0, 2, 1, 
    0, 0, 1, 1, 3, 5, 5, 0, 10, 0, 2, 0, 1, 3, 0, 
    
    -- channel=144
    30, 26, 30, 25, 23, 17, 14, 12, 12, 12, 6, 8, 9, 11, 11, 
    21, 16, 19, 14, 13, 7, 5, 8, 8, 0, 0, 6, 5, 7, 5, 
    13, 8, 9, 5, 4, 1, 1, 0, 0, 0, 3, 1, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 14, 13, 20, 5, 0, 0, 
    14, 16, 11, 11, 17, 15, 16, 17, 15, 16, 27, 30, 0, 5, 0, 
    18, 6, 7, 11, 16, 21, 30, 33, 32, 29, 20, 0, 2, 0, 0, 
    31, 31, 41, 41, 36, 31, 31, 24, 19, 2, 0, 0, 0, 0, 17, 
    21, 9, 14, 25, 24, 16, 12, 15, 19, 20, 18, 3, 2, 2, 0, 
    26, 38, 31, 18, 20, 29, 24, 9, 3, 10, 8, 2, 0, 0, 0, 
    26, 28, 23, 16, 9, 11, 6, 0, 4, 3, 0, 0, 0, 0, 0, 
    22, 19, 14, 11, 18, 19, 8, 6, 2, 1, 0, 0, 0, 0, 0, 
    14, 6, 7, 5, 0, 0, 4, 7, 0, 0, 2, 1, 0, 1, 1, 
    0, 0, 0, 4, 2, 0, 0, 0, 11, 6, 0, 0, 0, 3, 2, 
    0, 0, 1, 2, 5, 7, 4, 0, 0, 0, 0, 0, 1, 3, 0, 
    
    -- channel=145
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 14, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 6, 5, 13, 5, 2, 0, 0, 0, 
    3, 1, 2, 7, 0, 0, 0, 0, 32, 48, 22, 61, 47, 12, 17, 
    46, 36, 38, 38, 46, 42, 37, 25, 7, 0, 0, 0, 0, 2, 30, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 18, 2, 0, 0, 0, 
    0, 16, 9, 0, 0, 8, 9, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 17, 30, 26, 
    0, 0, 0, 5, 15, 12, 5, 20, 3, 7, 24, 28, 17, 10, 6, 
    0, 0, 3, 8, 0, 0, 13, 2, 1, 9, 11, 12, 4, 5, 6, 
    2, 19, 25, 14, 21, 26, 10, 0, 9, 16, 6, 1, 7, 0, 0, 
    22, 24, 13, 4, 3, 8, 10, 7, 0, 0, 4, 1, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 2, 7, 0, 0, 0, 0, 3, 
    
    -- channel=146
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 9, 
    0, 0, 0, 4, 3, 0, 0, 0, 0, 0, 0, 9, 16, 22, 28, 
    0, 0, 0, 0, 1, 6, 5, 2, 4, 10, 16, 18, 19, 30, 31, 
    27, 27, 25, 22, 15, 15, 19, 20, 19, 13, 24, 26, 30, 32, 30, 
    31, 33, 32, 31, 27, 23, 22, 23, 19, 18, 29, 31, 33, 31, 31, 
    
    -- channel=147
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 12, 12, 18, 0, 0, 0, 
    13, 16, 13, 12, 14, 13, 11, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 2, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 21, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 11, 
    0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 1, 4, 2, 3, 5, 
    0, 0, 0, 2, 0, 0, 0, 0, 1, 0, 0, 2, 3, 7, 10, 
    0, 0, 0, 1, 4, 5, 3, 0, 2, 4, 1, 2, 8, 9, 8, 
    12, 11, 6, 2, 1, 3, 6, 2, 0, 0, 7, 9, 8, 7, 6, 
    9, 9, 5, 5, 1, 0, 1, 3, 6, 5, 9, 12, 8, 6, 11, 
    
    -- channel=148
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 8, 
    
    -- channel=149
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=150
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 2, 2, 
    6, 3, 1, 1, 1, 0, 0, 0, 0, 5, 0, 4, 2, 3, 5, 
    5, 4, 3, 2, 0, 1, 2, 5, 0, 3, 3, 3, 5, 1, 14, 
    
    -- channel=151
    96, 44, 75, 81, 85, 77, 82, 97, 75, 85, 82, 80, 83, 90, 73, 
    95, 42, 68, 80, 84, 77, 83, 87, 74, 115, 35, 72, 84, 91, 68, 
    92, 35, 59, 77, 82, 74, 94, 66, 56, 133, 10, 59, 87, 83, 65, 
    81, 25, 57, 55, 74, 62, 82, 80, 74, 68, 34, 28, 25, 69, 44, 
    44, 30, 44, 33, 43, 41, 44, 77, 51, 52, 36, 18, 17, 75, 27, 
    22, 17, 54, 18, 44, 39, 48, 60, 43, 47, 6, 44, 82, 53, 52, 
    36, 36, 41, 18, 42, 59, 60, 56, 54, 56, 29, 54, 84, 37, 51, 
    43, 46, 41, 46, 59, 67, 73, 74, 66, 85, 33, 40, 54, 71, 38, 
    54, 54, 33, 59, 73, 74, 72, 68, 50, 73, 34, 50, 55, 54, 52, 
    54, 34, 55, 65, 60, 61, 64, 67, 44, 59, 56, 69, 61, 56, 28, 
    45, 61, 62, 65, 51, 49, 88, 54, 6, 53, 59, 58, 44, 31, 33, 
    28, 55, 82, 44, 37, 31, 70, 43, 32, 43, 43, 36, 32, 22, 20, 
    24, 48, 56, 37, 39, 37, 33, 32, 32, 33, 28, 15, 31, 13, 12, 
    21, 19, 21, 15, 21, 22, 22, 28, 6, 40, 19, 16, 15, 11, 14, 
    12, 6, 11, 11, 14, 16, 20, 24, 0, 42, 13, 12, 10, 8, 28, 
    
    -- channel=152
    36, 42, 37, 38, 33, 32, 25, 21, 24, 24, 24, 20, 23, 21, 23, 
    32, 35, 31, 29, 23, 24, 22, 18, 22, 22, 28, 19, 22, 19, 23, 
    25, 32, 24, 19, 14, 17, 15, 23, 24, 17, 28, 22, 19, 15, 19, 
    18, 26, 18, 14, 9, 12, 10, 9, 27, 29, 35, 44, 20, 12, 17, 
    24, 22, 22, 21, 18, 18, 21, 22, 24, 24, 26, 18, 16, 8, 17, 
    20, 20, 16, 19, 12, 21, 25, 30, 25, 20, 23, 4, 7, 0, 13, 
    29, 26, 26, 28, 34, 29, 34, 30, 26, 25, 23, 18, 1, 20, 11, 
    31, 23, 19, 29, 33, 35, 36, 37, 34, 29, 22, 11, 11, 4, 0, 
    41, 37, 44, 40, 43, 42, 40, 31, 27, 12, 12, 15, 17, 15, 13, 
    39, 31, 34, 42, 38, 32, 30, 30, 26, 22, 22, 20, 20, 19, 18, 
    37, 40, 40, 35, 38, 33, 29, 31, 32, 23, 25, 24, 17, 15, 11, 
    37, 38, 34, 35, 29, 34, 26, 20, 23, 22, 19, 18, 17, 15, 11, 
    33, 34, 31, 28, 30, 29, 21, 20, 20, 20, 17, 18, 13, 13, 10, 
    26, 24, 20, 19, 17, 16, 19, 19, 13, 17, 15, 13, 12, 12, 12, 
    8, 9, 11, 12, 12, 12, 14, 14, 16, 16, 12, 12, 12, 12, 8, 
    
    -- channel=153
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 14, 9, 2, 19, 14, 0, 0, 0, 
    7, 3, 20, 14, 6, 0, 0, 0, 27, 19, 9, 47, 51, 27, 24, 
    41, 29, 31, 42, 44, 43, 31, 23, 1, 0, 0, 0, 0, 0, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 13, 17, 2, 0, 0, 0, 
    11, 19, 6, 0, 6, 12, 3, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 1, 0, 0, 0, 15, 15, 0, 0, 6, 22, 25, 19, 
    0, 0, 0, 13, 30, 11, 0, 0, 0, 20, 27, 19, 12, 5, 13, 
    4, 0, 0, 0, 0, 5, 22, 5, 1, 4, 12, 4, 0, 4, 0, 
    19, 30, 31, 21, 18, 15, 2, 1, 15, 9, 0, 4, 4, 0, 0, 
    16, 15, 7, 5, 8, 10, 5, 1, 0, 0, 2, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 6, 6, 0, 0, 0, 0, 0, 6, 
    
    -- channel=154
    86, 88, 99, 99, 98, 95, 95, 91, 95, 96, 93, 94, 93, 94, 95, 
    83, 82, 95, 90, 91, 86, 86, 89, 92, 78, 79, 94, 90, 92, 92, 
    78, 77, 87, 81, 84, 79, 77, 80, 84, 57, 77, 91, 82, 83, 88, 
    67, 64, 71, 70, 71, 73, 73, 63, 51, 37, 44, 40, 63, 70, 72, 
    39, 38, 39, 45, 42, 48, 52, 54, 49, 51, 50, 47, 61, 40, 37, 
    44, 50, 46, 46, 54, 56, 63, 58, 53, 50, 62, 73, 43, 54, 41, 
    55, 42, 41, 53, 65, 64, 70, 66, 66, 67, 71, 69, 53, 54, 14, 
    65, 61, 70, 83, 86, 87, 87, 80, 77, 57, 53, 56, 58, 31, 32, 
    65, 61, 68, 81, 84, 80, 74, 67, 70, 59, 65, 63, 60, 53, 57, 
    56, 70, 80, 74, 70, 76, 76, 69, 65, 67, 66, 60, 51, 35, 29, 
    70, 75, 72, 64, 67, 69, 57, 39, 49, 61, 52, 40, 32, 27, 22, 
    68, 67, 56, 45, 49, 67, 55, 44, 43, 41, 37, 30, 24, 20, 11, 
    57, 55, 49, 43, 39, 35, 33, 38, 34, 29, 24, 27, 18, 16, 14, 
    20, 19, 22, 26, 28, 27, 26, 24, 31, 29, 19, 17, 15, 17, 15, 
    12, 14, 17, 19, 22, 25, 26, 18, 30, 18, 16, 13, 15, 17, 6, 
    
    -- channel=155
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 
    7, 6, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 2, 
    4, 6, 3, 2, 0, 0, 0, 0, 9, 0, 5, 5, 4, 3, 0, 
    
    -- channel=156
    38, 25, 33, 28, 26, 19, 18, 20, 16, 16, 13, 14, 13, 17, 12, 
    32, 19, 25, 18, 19, 13, 16, 20, 14, 20, 19, 13, 10, 15, 9, 
    24, 12, 15, 11, 12, 11, 15, 15, 13, 26, 18, 14, 11, 13, 9, 
    16, 2, 3, 4, 3, 4, 11, 8, 21, 47, 30, 29, 35, 9, 1, 
    28, 18, 25, 18, 18, 16, 22, 34, 31, 26, 28, 14, 0, 8, 8, 
    28, 17, 19, 20, 24, 21, 28, 34, 26, 28, 15, 4, 0, 23, 4, 
    28, 23, 30, 27, 36, 35, 38, 35, 29, 27, 8, 5, 17, 0, 6, 
    30, 25, 25, 21, 28, 31, 34, 28, 31, 23, 19, 11, 8, 13, 11, 
    36, 35, 38, 40, 37, 39, 41, 38, 24, 22, 4, 7, 15, 10, 9, 
    41, 33, 30, 35, 42, 33, 25, 22, 24, 25, 17, 17, 17, 21, 18, 
    42, 39, 36, 34, 32, 38, 35, 34, 22, 26, 24, 29, 24, 22, 16, 
    38, 39, 42, 39, 36, 27, 31, 21, 20, 28, 25, 28, 24, 20, 19, 
    29, 30, 36, 27, 29, 33, 30, 22, 22, 27, 25, 17, 21, 19, 17, 
    26, 29, 26, 23, 20, 21, 25, 26, 22, 15, 21, 17, 19, 17, 15, 
    15, 15, 18, 19, 20, 18, 19, 18, 16, 23, 17, 17, 17, 17, 13, 
    
    -- channel=157
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=158
    21, 21, 21, 16, 13, 8, 6, 5, 6, 3, 0, 2, 4, 5, 4, 
    14, 13, 12, 6, 5, 3, 0, 2, 3, 0, 0, 2, 0, 0, 1, 
    6, 6, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 14, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 11, 14, 10, 2, 0, 0, 
    21, 14, 9, 16, 23, 19, 19, 14, 13, 15, 22, 17, 6, 0, 1, 
    19, 12, 12, 22, 22, 26, 32, 34, 35, 29, 14, 0, 0, 0, 0, 
    27, 27, 30, 31, 26, 24, 22, 16, 10, 0, 0, 0, 0, 11, 28, 
    15, 10, 19, 21, 16, 13, 15, 17, 15, 12, 13, 5, 5, 0, 0, 
    31, 29, 24, 19, 22, 22, 13, 0, 0, 8, 7, 0, 0, 0, 0, 
    22, 26, 18, 9, 4, 9, 11, 11, 12, 0, 0, 0, 0, 1, 0, 
    22, 18, 19, 20, 25, 15, 0, 3, 8, 5, 0, 7, 7, 5, 3, 
    9, 1, 0, 3, 5, 5, 8, 6, 1, 4, 6, 4, 3, 7, 8, 
    6, 4, 6, 6, 2, 2, 7, 7, 12, 8, 6, 6, 7, 9, 7, 
    5, 7, 9, 10, 10, 9, 7, 3, 5, 5, 7, 6, 7, 8, 0, 
    
    -- channel=159
    101, 66, 83, 97, 100, 99, 99, 108, 89, 102, 103, 99, 107, 103, 97, 
    99, 66, 77, 100, 94, 97, 94, 94, 91, 115, 58, 88, 109, 102, 95, 
    99, 63, 72, 97, 89, 92, 96, 71, 74, 129, 20, 75, 107, 92, 86, 
    90, 60, 70, 74, 84, 78, 88, 86, 69, 52, 17, 17, 15, 72, 64, 
    35, 31, 31, 22, 37, 37, 45, 64, 56, 48, 32, 35, 26, 65, 29, 
    11, 24, 48, 19, 34, 39, 46, 58, 41, 41, 23, 53, 93, 24, 62, 
    24, 39, 34, 14, 36, 62, 56, 60, 54, 53, 39, 63, 86, 43, 76, 
    46, 52, 49, 56, 67, 75, 81, 84, 71, 83, 31, 44, 64, 87, 33, 
    55, 49, 35, 63, 79, 76, 70, 67, 55, 78, 40, 57, 62, 67, 46, 
    55, 35, 55, 64, 62, 64, 68, 70, 53, 59, 61, 71, 60, 51, 25, 
    45, 60, 63, 66, 46, 48, 78, 49, 11, 42, 55, 50, 36, 24, 17, 
    12, 54, 69, 38, 29, 21, 66, 47, 28, 32, 33, 23, 18, 10, 7, 
    16, 45, 48, 35, 28, 22, 25, 24, 22, 19, 18, 7, 19, 1, 0, 
    5, 5, 7, 4, 10, 9, 8, 13, 1, 27, 6, 4, 3, 0, 1, 
    0, 0, 0, 0, 0, 4, 6, 10, 0, 35, 0, 0, 0, 0, 8, 
    
    -- channel=160
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=161
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 26, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 33, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 9, 17, 0, 0, 0, 4, 1, 0, 0, 
    0, 0, 10, 5, 0, 0, 0, 0, 0, 0, 0, 3, 4, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 8, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 12, 
    
    -- channel=162
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 9, 6, 15, 0, 11, 0, 0, 0, 
    8, 2, 0, 10, 2, 0, 1, 0, 28, 44, 12, 38, 40, 13, 21, 
    39, 29, 28, 28, 36, 34, 34, 27, 11, 0, 3, 0, 0, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 35, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 8, 18, 0, 0, 0, 0, 
    0, 23, 6, 0, 0, 12, 12, 1, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 1, 0, 0, 2, 23, 0, 0, 0, 18, 27, 22, 
    2, 0, 0, 8, 15, 19, 2, 20, 0, 4, 25, 26, 15, 14, 4, 
    0, 3, 2, 8, 0, 0, 20, 10, 3, 7, 11, 18, 1, 5, 7, 
    3, 20, 30, 17, 20, 22, 9, 0, 11, 17, 5, 3, 10, 1, 0, 
    15, 20, 11, 4, 5, 11, 10, 6, 0, 0, 7, 1, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 4, 11, 0, 1, 0, 0, 3, 
    
    -- channel=163
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 22, 0, 0, 0, 0, 
    0, 7, 0, 0, 0, 0, 0, 21, 11, 22, 8, 9, 4, 0, 0, 
    5, 6, 4, 5, 4, 0, 2, 0, 52, 58, 45, 89, 39, 12, 27, 
    47, 44, 48, 50, 51, 49, 41, 30, 4, 0, 2, 0, 0, 5, 41, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 4, 11, 0, 3, 0, 0, 0, 0, 0, 0, 4, 0, 23, 27, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 24, 7, 0, 0, 0, 
    3, 24, 14, 0, 3, 14, 17, 5, 0, 0, 0, 0, 0, 0, 14, 
    0, 0, 0, 10, 0, 0, 0, 4, 16, 0, 0, 3, 24, 35, 29, 
    0, 0, 0, 7, 20, 9, 13, 34, 12, 11, 30, 33, 18, 12, 11, 
    0, 6, 10, 19, 0, 0, 12, 0, 7, 15, 15, 17, 8, 8, 8, 
    4, 19, 21, 12, 27, 34, 11, 0, 14, 18, 5, 4, 10, 2, 0, 
    29, 28, 14, 5, 3, 11, 15, 11, 0, 0, 6, 4, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 4, 11, 1, 1, 0, 0, 11, 
    
    -- channel=164
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=165
    5, 8, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 13, 0, 0, 
    6, 16, 7, 6, 26, 18, 3, 0, 0, 7, 34, 56, 47, 0, 11, 
    2, 0, 0, 0, 0, 14, 22, 38, 51, 40, 29, 0, 0, 0, 0, 
    24, 36, 48, 49, 25, 16, 11, 3, 0, 0, 0, 0, 0, 29, 64, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 22, 35, 6, 0, 0, 0, 
    11, 28, 11, 0, 0, 13, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 10, 0, 0, 0, 1, 1, 
    0, 0, 1, 2, 3, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=166
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 0, 0, 0, 0, 0, 1, 4, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 1, 0, 11, 0, 0, 0, 0, 
    0, 10, 4, 1, 0, 1, 0, 6, 11, 6, 16, 26, 8, 3, 5, 
    10, 16, 12, 14, 12, 10, 7, 1, 3, 5, 7, 9, 9, 11, 22, 
    7, 10, 6, 7, 3, 6, 1, 2, 6, 6, 6, 0, 15, 0, 8, 
    5, 13, 6, 7, 2, 0, 0, 0, 2, 2, 10, 5, 0, 13, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 11, 8, 3, 7, 9, 
    4, 1, 1, 0, 0, 0, 2, 3, 4, 0, 5, 4, 4, 9, 3, 
    0, 0, 0, 0, 0, 1, 1, 5, 5, 1, 3, 4, 9, 13, 16, 
    0, 0, 1, 2, 4, 1, 6, 10, 17, 8, 8, 10, 15, 14, 18, 
    4, 2, 4, 8, 6, 8, 2, 8, 13, 13, 15, 14, 17, 19, 18, 
    8, 7, 5, 10, 13, 14, 12, 14, 15, 15, 17, 18, 15, 17, 17, 
    19, 18, 17, 17, 17, 17, 16, 18, 13, 16, 16, 18, 18, 17, 19, 
    19, 19, 19, 19, 17, 17, 17, 19, 17, 16, 17, 17, 18, 17, 21, 
    
    -- channel=167
    0, 0, 0, 0, 0, 0, 4, 4, 6, 6, 7, 7, 6, 7, 6, 
    0, 0, 0, 0, 4, 4, 7, 8, 7, 7, 7, 10, 8, 9, 9, 
    0, 0, 5, 6, 11, 8, 9, 11, 9, 2, 3, 10, 10, 12, 10, 
    2, 0, 9, 11, 14, 11, 11, 4, 3, 0, 0, 7, 9, 15, 15, 
    1, 0, 7, 10, 13, 11, 7, 1, 0, 0, 0, 0, 5, 12, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 5, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=168
    85, 57, 76, 77, 78, 72, 75, 81, 70, 76, 72, 73, 75, 78, 69, 
    82, 54, 68, 73, 74, 69, 72, 76, 69, 85, 51, 68, 74, 76, 66, 
    76, 46, 59, 68, 69, 66, 74, 58, 58, 92, 35, 60, 74, 70, 62, 
    64, 36, 48, 49, 57, 55, 64, 65, 58, 62, 39, 34, 41, 56, 41, 
    42, 34, 41, 33, 39, 39, 46, 65, 54, 48, 41, 33, 21, 53, 30, 
    35, 32, 47, 31, 48, 46, 53, 57, 46, 50, 31, 46, 56, 44, 39, 
    41, 41, 43, 35, 52, 63, 63, 61, 60, 58, 39, 47, 63, 25, 43, 
    51, 52, 51, 53, 63, 69, 73, 70, 64, 64, 37, 41, 49, 56, 40, 
    56, 52, 49, 66, 70, 71, 71, 68, 54, 64, 39, 47, 51, 49, 40, 
    58, 50, 57, 62, 67, 65, 63, 59, 49, 58, 53, 57, 49, 46, 31, 
    58, 63, 63, 61, 51, 58, 72, 51, 29, 50, 51, 51, 43, 34, 27, 
    42, 59, 70, 49, 46, 41, 58, 43, 37, 44, 42, 38, 33, 25, 21, 
    35, 47, 50, 39, 39, 39, 38, 36, 34, 35, 33, 22, 29, 19, 18, 
    23, 25, 27, 24, 26, 27, 29, 32, 24, 33, 23, 20, 20, 18, 18, 
    16, 15, 19, 20, 24, 24, 25, 24, 12, 36, 17, 17, 17, 16, 18, 
    
    -- channel=169
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 5, 22, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 1, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 5, 
    
    -- channel=170
    88, 68, 103, 108, 119, 115, 126, 130, 125, 134, 127, 134, 126, 135, 127, 
    96, 74, 110, 112, 126, 118, 130, 134, 125, 130, 105, 134, 129, 139, 129, 
    101, 72, 110, 115, 128, 118, 126, 116, 117, 112, 86, 123, 129, 135, 130, 
    103, 73, 112, 120, 126, 119, 118, 102, 80, 68, 44, 60, 108, 122, 114, 
    70, 55, 71, 78, 90, 91, 87, 84, 48, 37, 30, 31, 47, 91, 69, 
    23, 20, 38, 26, 45, 38, 49, 43, 34, 35, 27, 68, 65, 95, 37, 
    30, 28, 32, 31, 56, 53, 50, 39, 38, 45, 60, 97, 98, 64, 38, 
    33, 37, 41, 48, 64, 71, 74, 71, 77, 74, 71, 89, 87, 47, 37, 
    49, 52, 59, 76, 78, 75, 72, 69, 65, 66, 57, 76, 78, 71, 79, 
    33, 38, 54, 63, 63, 62, 67, 71, 64, 79, 78, 82, 69, 57, 42, 
    51, 53, 58, 57, 60, 69, 69, 38, 31, 70, 67, 55, 35, 20, 19, 
    42, 53, 53, 28, 28, 48, 60, 33, 30, 39, 29, 19, 14, 4, 0, 
    33, 45, 45, 28, 29, 33, 27, 20, 20, 20, 11, 5, 7, 0, 0, 
    9, 9, 6, 4, 8, 9, 10, 9, 5, 5, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 7, 5, 0, 0, 0, 0, 0, 
    
    -- channel=171
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 
    0, 5, 1, 0, 0, 0, 0, 0, 3, 0, 41, 8, 0, 0, 0, 
    0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 8, 14, 36, 0, 10, 
    0, 8, 0, 16, 5, 10, 4, 0, 0, 0, 0, 0, 14, 0, 10, 
    2, 2, 0, 3, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 
    0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 3, 0, 0, 0, 
    0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 3, 0, 0, 18, 0, 0, 0, 0, 0, 0, 
    19, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 
    
    -- channel=172
    32, 27, 26, 30, 27, 26, 23, 22, 19, 23, 24, 19, 22, 20, 20, 
    28, 23, 21, 25, 19, 22, 21, 19, 19, 31, 21, 17, 23, 20, 19, 
    24, 21, 15, 17, 13, 17, 18, 21, 21, 32, 15, 22, 22, 16, 17, 
    22, 17, 16, 13, 11, 11, 12, 15, 34, 32, 21, 34, 21, 17, 15, 
    25, 22, 21, 20, 22, 22, 25, 29, 23, 19, 17, 2, 0, 5, 15, 
    4, 7, 11, 3, 3, 11, 20, 26, 16, 10, 0, 0, 4, 0, 11, 
    14, 17, 17, 12, 19, 21, 19, 15, 9, 9, 4, 10, 8, 10, 21, 
    16, 9, 8, 13, 21, 25, 27, 31, 29, 29, 12, 7, 10, 8, 0, 
    34, 32, 26, 31, 38, 39, 33, 22, 15, 8, 0, 8, 14, 14, 8, 
    22, 16, 23, 32, 26, 21, 21, 28, 24, 16, 16, 21, 23, 21, 14, 
    25, 29, 30, 33, 32, 25, 29, 24, 12, 21, 26, 23, 17, 9, 8, 
    17, 28, 30, 23, 14, 17, 29, 17, 13, 15, 17, 11, 8, 6, 2, 
    20, 31, 29, 23, 21, 18, 13, 10, 15, 12, 9, 4, 7, 1, 0, 
    12, 11, 8, 6, 7, 8, 8, 8, 0, 7, 4, 3, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 4, 0, 11, 0, 0, 0, 0, 1, 
    
    -- channel=173
    14, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 
    14, 0, 0, 1, 0, 0, 4, 0, 0, 60, 0, 0, 6, 0, 0, 
    14, 0, 0, 0, 0, 0, 8, 7, 4, 21, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 11, 12, 2, 0, 0, 0, 13, 0, 
    0, 0, 11, 0, 0, 0, 0, 9, 0, 4, 0, 0, 33, 0, 20, 
    0, 0, 3, 0, 0, 7, 0, 9, 2, 0, 0, 0, 38, 0, 50, 
    0, 4, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 61, 14, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 28, 0, 0, 0, 6, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 11, 0, 
    0, 0, 0, 1, 0, 0, 18, 15, 0, 0, 0, 10, 8, 7, 1, 
    0, 0, 17, 2, 0, 0, 14, 9, 0, 0, 0, 7, 5, 2, 10, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 1, 6, 0, 13, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 8, 2, 0, 3, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 4, 0, 28, 0, 1, 0, 0, 14, 
    
    -- channel=174
    19, 6, 15, 10, 13, 8, 11, 16, 10, 10, 2, 12, 12, 15, 10, 
    11, 0, 6, 7, 9, 4, 3, 7, 7, 0, 0, 6, 7, 9, 5, 
    10, 0, 2, 9, 10, 6, 5, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 1, 4, 14, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 20, 8, 0, 0, 
    8, 12, 17, 4, 29, 16, 12, 0, 2, 13, 26, 63, 40, 12, 9, 
    4, 0, 0, 0, 0, 16, 21, 32, 43, 35, 22, 0, 13, 0, 0, 
    24, 38, 56, 51, 33, 25, 21, 10, 0, 0, 0, 0, 1, 24, 58, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 34, 35, 12, 0, 6, 0, 
    6, 31, 20, 0, 0, 17, 16, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 8, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 3, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=175
    64, 49, 72, 75, 81, 78, 83, 85, 79, 86, 81, 85, 83, 87, 83, 
    64, 49, 71, 74, 79, 75, 79, 82, 79, 77, 59, 83, 83, 86, 82, 
    64, 45, 66, 72, 75, 71, 73, 61, 65, 65, 40, 70, 79, 78, 78, 
    58, 42, 60, 66, 68, 67, 65, 57, 35, 24, 12, 11, 42, 62, 57, 
    20, 14, 19, 21, 29, 31, 34, 36, 22, 15, 11, 15, 19, 41, 19, 
    5, 5, 16, 8, 24, 18, 27, 23, 15, 16, 18, 47, 40, 40, 13, 
    12, 10, 9, 12, 30, 36, 35, 33, 31, 33, 38, 52, 53, 20, 9, 
    24, 27, 33, 39, 49, 52, 53, 49, 47, 40, 29, 41, 45, 29, 19, 
    28, 24, 30, 49, 51, 47, 44, 42, 38, 42, 34, 40, 42, 38, 31, 
    23, 26, 37, 39, 40, 42, 43, 39, 32, 43, 44, 43, 28, 16, 4, 
    31, 35, 36, 32, 27, 37, 38, 13, 7, 30, 26, 17, 4, 0, 0, 
    18, 31, 30, 10, 12, 21, 28, 12, 7, 9, 1, 0, 0, 0, 0, 
    8, 16, 14, 5, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=176
    70, 68, 85, 90, 94, 94, 99, 98, 99, 104, 104, 104, 100, 102, 101, 
    77, 73, 92, 92, 98, 96, 100, 102, 100, 102, 103, 105, 102, 106, 103, 
    80, 73, 93, 92, 98, 93, 95, 100, 103, 84, 86, 109, 104, 105, 103, 
    80, 69, 89, 95, 96, 91, 88, 74, 83, 74, 63, 90, 107, 100, 103, 
    73, 65, 75, 83, 88, 90, 86, 77, 46, 35, 37, 26, 45, 67, 71, 
    24, 26, 30, 31, 32, 35, 42, 42, 38, 34, 30, 39, 40, 64, 30, 
    32, 35, 35, 38, 56, 46, 43, 33, 30, 36, 53, 81, 66, 60, 38, 
    29, 26, 21, 31, 50, 58, 62, 63, 70, 67, 74, 74, 68, 32, 12, 
    48, 59, 64, 68, 70, 76, 76, 66, 59, 44, 42, 59, 65, 56, 69, 
    34, 30, 47, 63, 62, 55, 58, 65, 69, 68, 65, 65, 65, 59, 50, 
    52, 52, 55, 55, 65, 71, 62, 48, 46, 66, 68, 60, 41, 29, 23, 
    50, 56, 51, 40, 32, 51, 54, 34, 39, 44, 37, 33, 20, 15, 8, 
    42, 52, 49, 36, 44, 47, 33, 27, 31, 33, 20, 17, 14, 6, 1, 
    25, 25, 19, 17, 19, 23, 25, 22, 12, 11, 13, 8, 5, 2, 2, 
    3, 2, 5, 6, 7, 6, 11, 13, 21, 14, 5, 3, 2, 3, 2, 
    
    -- channel=177
    78, 67, 83, 84, 88, 86, 90, 93, 89, 92, 84, 93, 95, 96, 94, 
    75, 63, 79, 81, 85, 79, 78, 83, 87, 64, 51, 89, 91, 90, 88, 
    73, 58, 74, 82, 83, 78, 75, 52, 61, 52, 35, 61, 77, 77, 80, 
    54, 47, 50, 55, 66, 68, 74, 64, 6, 0, 0, 0, 0, 45, 42, 
    0, 0, 0, 0, 0, 0, 10, 22, 30, 32, 24, 57, 50, 40, 2, 
    35, 45, 42, 41, 63, 58, 47, 39, 37, 46, 68, 104, 74, 57, 43, 
    33, 23, 22, 27, 43, 60, 68, 76, 84, 78, 70, 57, 70, 36, 2, 
    61, 73, 88, 90, 82, 79, 77, 62, 49, 32, 17, 44, 58, 60, 85, 
    30, 13, 28, 51, 50, 37, 37, 52, 63, 80, 79, 64, 54, 52, 38, 
    49, 65, 60, 41, 49, 68, 65, 40, 28, 53, 57, 46, 18, 2, 0, 
    37, 52, 45, 30, 13, 28, 36, 13, 21, 25, 10, 7, 6, 8, 0, 
    25, 36, 31, 20, 35, 34, 24, 22, 17, 17, 9, 4, 8, 0, 0, 
    12, 4, 2, 1, 0, 0, 11, 18, 1, 0, 8, 5, 1, 1, 5, 
    0, 0, 0, 1, 3, 0, 0, 3, 23, 21, 1, 0, 1, 5, 5, 
    1, 3, 6, 8, 14, 16, 9, 0, 0, 9, 0, 0, 2, 5, 0, 
    
    -- channel=178
    10, 4, 5, 7, 7, 7, 9, 8, 6, 10, 10, 5, 6, 7, 6, 
    4, 3, 3, 6, 5, 4, 5, 5, 6, 7, 0, 6, 6, 7, 3, 
    6, 3, 4, 3, 6, 3, 6, 2, 3, 0, 1, 16, 7, 2, 4, 
    13, 6, 19, 10, 10, 4, 7, 18, 0, 0, 0, 0, 0, 18, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 13, 6, 6, 23, 0, 0, 
    0, 13, 18, 0, 2, 5, 15, 11, 11, 7, 5, 28, 13, 1, 7, 
    11, 1, 0, 0, 0, 0, 0, 0, 0, 1, 12, 4, 3, 21, 0, 
    12, 11, 25, 32, 24, 17, 16, 18, 14, 11, 0, 0, 3, 0, 0, 
    15, 6, 0, 2, 14, 8, 0, 0, 0, 10, 20, 10, 2, 12, 13, 
    0, 17, 27, 3, 0, 5, 20, 25, 11, 4, 6, 13, 13, 0, 0, 
    4, 5, 9, 17, 14, 0, 0, 0, 0, 13, 5, 0, 1, 0, 11, 
    0, 0, 0, 0, 0, 9, 20, 20, 1, 0, 6, 0, 0, 0, 0, 
    13, 17, 11, 14, 0, 0, 0, 9, 9, 0, 0, 3, 1, 0, 1, 
    0, 0, 0, 0, 8, 4, 0, 0, 0, 14, 0, 0, 0, 1, 2, 
    0, 0, 0, 0, 0, 6, 6, 5, 0, 0, 2, 0, 1, 1, 6, 
    
    -- channel=179
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 3, 3, 3, 4, 
    5, 5, 4, 4, 2, 2, 1, 3, 0, 8, 3, 3, 3, 2, 16, 
    
    -- channel=180
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 2, 0, 0, 11, 0, 5, 
    0, 0, 0, 0, 0, 1, 4, 5, 5, 4, 0, 0, 4, 0, 3, 
    0, 3, 3, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 10, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 4, 
    
    -- channel=181
    27, 35, 41, 39, 38, 35, 33, 29, 35, 33, 31, 33, 29, 32, 32, 
    28, 32, 40, 31, 35, 30, 32, 32, 33, 29, 45, 35, 29, 32, 34, 
    23, 27, 35, 25, 29, 25, 25, 35, 36, 13, 42, 36, 27, 31, 33, 
    15, 17, 19, 21, 18, 21, 17, 8, 31, 38, 45, 59, 48, 21, 27, 
    28, 26, 33, 35, 30, 31, 31, 22, 10, 8, 13, 0, 7, 17, 25, 
    12, 2, 0, 12, 9, 9, 13, 12, 11, 7, 10, 0, 0, 12, 0, 
    15, 11, 13, 25, 34, 22, 25, 17, 14, 14, 19, 24, 0, 4, 0, 
    11, 5, 0, 8, 19, 24, 24, 22, 26, 17, 32, 21, 12, 0, 0, 
    21, 29, 45, 37, 32, 36, 41, 33, 24, 0, 5, 12, 17, 4, 12, 
    25, 14, 19, 34, 37, 24, 17, 15, 22, 23, 19, 12, 13, 13, 15, 
    31, 29, 26, 18, 29, 37, 23, 25, 30, 22, 21, 21, 6, 1, 0, 
    37, 31, 25, 27, 22, 27, 7, 0, 14, 17, 6, 9, 1, 0, 0, 
    20, 17, 14, 9, 22, 28, 12, 4, 5, 12, 0, 0, 0, 0, 0, 
    15, 14, 7, 3, 0, 2, 9, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 
    
    -- channel=182
    16, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 31, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 0, 8, 0, 0, 73, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 9, 10, 16, 20, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 15, 3, 6, 0, 0, 0, 17, 0, 
    0, 0, 16, 0, 0, 0, 0, 11, 0, 2, 0, 0, 46, 0, 38, 
    0, 0, 6, 0, 0, 1, 1, 7, 4, 1, 0, 0, 32, 0, 35, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 26, 0, 0, 0, 52, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 6, 6, 13, 0, 
    0, 0, 0, 3, 0, 0, 27, 18, 0, 0, 0, 11, 7, 5, 6, 
    0, 0, 27, 2, 0, 0, 17, 2, 0, 0, 6, 5, 8, 2, 10, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 3, 0, 15, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 22, 0, 1, 2, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 6, 0, 31, 0, 0, 0, 0, 24, 
    
    -- channel=183
    6, 0, 0, 0, 0, 0, 1, 7, 0, 3, 3, 2, 4, 3, 0, 
    9, 0, 0, 4, 3, 4, 5, 5, 0, 16, 1, 0, 6, 4, 0, 
    11, 0, 0, 8, 5, 8, 11, 4, 5, 31, 0, 0, 12, 8, 1, 
    11, 1, 0, 3, 6, 6, 10, 14, 13, 24, 0, 8, 5, 8, 3, 
    14, 9, 13, 6, 12, 9, 11, 17, 14, 7, 1, 5, 0, 15, 11, 
    0, 0, 7, 0, 0, 1, 0, 8, 4, 7, 0, 0, 15, 1, 14, 
    0, 5, 8, 0, 0, 2, 0, 0, 0, 0, 0, 0, 19, 2, 34, 
    0, 0, 0, 0, 0, 0, 1, 4, 3, 15, 2, 4, 7, 20, 4, 
    3, 0, 0, 0, 1, 5, 8, 10, 2, 11, 0, 0, 5, 12, 4, 
    4, 0, 0, 0, 5, 2, 2, 8, 5, 5, 2, 10, 13, 20, 13, 
    0, 0, 3, 8, 2, 3, 14, 15, 0, 6, 13, 21, 19, 16, 11, 
    0, 4, 12, 8, 2, 0, 15, 10, 4, 12, 17, 13, 13, 10, 14, 
    0, 8, 15, 8, 8, 13, 14, 10, 11, 12, 16, 6, 14, 10, 9, 
    9, 13, 13, 10, 10, 10, 10, 13, 6, 9, 10, 8, 11, 7, 9, 
    10, 7, 8, 7, 9, 8, 9, 12, 0, 21, 5, 9, 8, 6, 13, 
    
    -- channel=184
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 13, 11, 3, 17, 16, 0, 0, 0, 
    4, 2, 8, 11, 1, 0, 0, 0, 32, 42, 18, 57, 64, 22, 26, 
    51, 38, 41, 48, 53, 51, 44, 31, 6, 0, 0, 0, 0, 0, 29, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 21, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 8, 23, 4, 0, 0, 0, 
    4, 23, 9, 0, 0, 13, 9, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 7, 23, 0, 0, 0, 22, 31, 26, 
    0, 0, 0, 10, 26, 19, 0, 12, 1, 15, 30, 29, 18, 13, 8, 
    0, 0, 0, 2, 0, 0, 22, 6, 2, 8, 14, 13, 1, 5, 4, 
    13, 27, 34, 20, 22, 23, 8, 0, 15, 16, 4, 3, 7, 0, 0, 
    17, 22, 11, 6, 8, 12, 9, 5, 0, 0, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 7, 2, 0, 0, 0, 0, 2, 
    
    -- channel=185
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=186
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 
    0, 4, 0, 0, 0, 0, 0, 0, 1, 0, 25, 4, 0, 0, 0, 
    0, 14, 0, 5, 0, 0, 0, 0, 0, 0, 0, 2, 32, 0, 14, 
    1, 9, 0, 7, 7, 9, 8, 0, 0, 0, 0, 4, 1, 0, 9, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 
    
    -- channel=187
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 
    0, 0, 1, 6, 4, 0, 0, 0, 7, 24, 3, 21, 17, 8, 2, 
    20, 10, 20, 17, 24, 18, 11, 8, 0, 0, 0, 0, 0, 20, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 3, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 14, 11, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 3, 10, 2, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 2, 0, 0, 2, 0, 0, 
    6, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 6, 
    
    -- channel=188
    59, 49, 63, 63, 63, 59, 62, 61, 60, 63, 60, 60, 58, 62, 59, 
    56, 45, 59, 56, 59, 54, 58, 60, 59, 62, 45, 60, 57, 62, 56, 
    52, 40, 52, 49, 55, 50, 55, 54, 52, 50, 44, 58, 54, 55, 55, 
    48, 32, 49, 46, 49, 45, 49, 45, 43, 31, 29, 30, 46, 51, 43, 
    33, 27, 31, 35, 35, 38, 38, 45, 30, 32, 29, 17, 29, 30, 25, 
    21, 23, 29, 20, 32, 31, 40, 39, 31, 28, 22, 37, 25, 37, 22, 
    34, 24, 25, 29, 40, 39, 42, 36, 35, 36, 36, 43, 37, 33, 6, 
    37, 33, 39, 47, 53, 54, 55, 52, 51, 44, 32, 35, 36, 15, 8, 
    46, 44, 41, 54, 59, 56, 49, 41, 40, 35, 34, 37, 37, 32, 38, 
    32, 41, 51, 50, 42, 45, 48, 48, 40, 42, 42, 43, 38, 27, 18, 
    43, 48, 48, 46, 47, 44, 44, 25, 21, 44, 38, 29, 21, 14, 15, 
    41, 42, 42, 26, 27, 41, 42, 26, 24, 25, 24, 16, 13, 9, 3, 
    35, 38, 36, 28, 25, 22, 18, 20, 21, 17, 11, 12, 10, 4, 3, 
    11, 9, 9, 10, 14, 13, 12, 11, 8, 16, 8, 7, 4, 4, 3, 
    1, 1, 3, 4, 6, 8, 10, 8, 10, 9, 6, 3, 3, 4, 3, 
    
    -- channel=189
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 3, 8, 0, 0, 2, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 1, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 7, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 23, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 1, 0, 0, 7, 
    
    -- channel=190
    22, 12, 28, 33, 40, 41, 47, 49, 45, 51, 49, 50, 47, 51, 48, 
    27, 17, 33, 39, 44, 44, 51, 51, 46, 53, 36, 52, 51, 55, 50, 
    33, 20, 37, 42, 47, 44, 50, 44, 42, 43, 26, 47, 51, 53, 51, 
    41, 28, 53, 55, 56, 50, 46, 41, 31, 16, 6, 17, 41, 55, 50, 
    26, 20, 25, 32, 40, 40, 34, 29, 8, 3, 0, 1, 14, 36, 28, 
    0, 0, 7, 0, 7, 2, 9, 6, 0, 0, 0, 20, 26, 35, 9, 
    0, 0, 0, 0, 7, 6, 2, 0, 0, 0, 15, 38, 40, 29, 14, 
    0, 1, 5, 8, 15, 15, 14, 17, 21, 25, 22, 34, 34, 15, 3, 
    11, 11, 7, 17, 20, 18, 11, 9, 12, 16, 17, 27, 27, 27, 30, 
    0, 0, 10, 13, 5, 7, 15, 22, 16, 22, 26, 31, 25, 19, 10, 
    2, 4, 9, 13, 14, 12, 17, 1, 0, 21, 20, 12, 4, 0, 2, 
    0, 4, 7, 0, 0, 6, 18, 4, 0, 1, 0, 0, 0, 0, 0, 
    0, 8, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=191
    0, 15, 16, 1, 2, 0, 2, 0, 10, 1, 0, 2, 0, 0, 2, 
    0, 12, 18, 0, 4, 0, 0, 0, 5, 0, 14, 11, 0, 0, 5, 
    0, 6, 18, 0, 4, 0, 0, 1, 8, 0, 57, 13, 0, 0, 9, 
    0, 5, 10, 0, 0, 0, 0, 0, 0, 0, 12, 7, 31, 0, 6, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 6, 31, 0, 3, 
    17, 13, 0, 9, 10, 5, 7, 0, 0, 0, 32, 29, 0, 18, 0, 
    16, 0, 0, 29, 15, 0, 0, 0, 6, 8, 42, 10, 0, 0, 0, 
    3, 3, 13, 24, 12, 5, 0, 0, 0, 0, 13, 9, 0, 0, 9, 
    0, 0, 20, 9, 0, 0, 0, 0, 8, 0, 29, 5, 0, 0, 0, 
    0, 27, 15, 0, 0, 4, 2, 0, 0, 0, 1, 0, 0, 0, 0, 
    12, 0, 0, 0, 5, 6, 0, 0, 28, 8, 0, 0, 0, 0, 0, 
    42, 0, 0, 0, 2, 39, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 10, 0, 0, 0, 0, 1, 1, 
    0, 4, 3, 4, 3, 3, 2, 0, 30, 0, 1, 0, 0, 4, 0, 
    
    -- channel=192
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=193
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 3, 5, 6, 5, 7, 6, 5, 5, 0, 0, 0, 
    0, 0, 0, 16, 11, 13, 18, 15, 13, 16, 12, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 15, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 16, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 4, 5, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 18, 17, 5, 12, 17, 21, 12, 11, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 2, 6, 8, 7, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 1, 5, 3, 3, 4, 8, 9, 9, 10, 9, 7, 10, 
    16, 9, 9, 10, 11, 11, 13, 14, 15, 15, 16, 15, 8, 13, 7, 
    
    -- channel=194
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 10, 11, 0, 0, 0, 0, 8, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 8, 0, 7, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 7, 14, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 4, 6, 12, 16, 17, 16, 9, 8, 10, 9, 8, 8, 7, 3, 
    0, 0, 0, 3, 5, 3, 6, 8, 11, 12, 13, 14, 13, 12, 18, 
    10, 12, 12, 12, 13, 12, 12, 14, 12, 13, 15, 17, 18, 23, 17, 
    
    -- channel=195
    31, 26, 21, 19, 24, 22, 21, 23, 22, 24, 22, 22, 24, 21, 20, 
    36, 33, 23, 0, 5, 0, 0, 0, 0, 0, 1, 4, 22, 21, 22, 
    35, 34, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 23, 22, 
    34, 33, 13, 0, 6, 7, 0, 3, 9, 0, 6, 5, 23, 26, 27, 
    29, 33, 25, 16, 21, 22, 24, 22, 22, 18, 20, 28, 20, 26, 27, 
    26, 27, 22, 19, 23, 21, 22, 20, 19, 21, 20, 27, 25, 24, 27, 
    27, 20, 21, 35, 23, 21, 25, 25, 23, 22, 23, 22, 24, 24, 26, 
    29, 25, 10, 0, 21, 31, 19, 19, 23, 21, 23, 23, 24, 24, 28, 
    28, 22, 20, 12, 0, 10, 26, 28, 13, 12, 21, 24, 25, 25, 27, 
    26, 21, 21, 16, 0, 10, 7, 3, 13, 25, 36, 18, 11, 15, 22, 
    27, 21, 22, 6, 2, 0, 21, 26, 5, 9, 11, 18, 34, 26, 29, 
    21, 12, 13, 13, 14, 2, 6, 19, 22, 17, 21, 17, 26, 30, 27, 
    14, 10, 9, 6, 5, 4, 7, 13, 9, 10, 9, 12, 11, 9, 12, 
    13, 12, 10, 9, 7, 9, 9, 7, 5, 4, 5, 4, 5, 7, 18, 
    2, 3, 5, 6, 3, 6, 5, 5, 4, 5, 4, 3, 9, 22, 12, 
    
    -- channel=196
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=197
    33, 29, 5, 12, 21, 17, 13, 14, 12, 15, 16, 14, 18, 24, 23, 
    35, 36, 19, 0, 17, 18, 9, 15, 13, 16, 15, 18, 31, 26, 25, 
    34, 33, 26, 0, 0, 1, 0, 3, 1, 1, 3, 9, 31, 27, 28, 
    29, 32, 12, 0, 5, 3, 0, 6, 5, 0, 7, 9, 20, 28, 29, 
    24, 32, 23, 13, 16, 17, 15, 19, 18, 13, 18, 28, 22, 27, 27, 
    28, 27, 26, 24, 17, 18, 21, 20, 16, 18, 20, 28, 26, 25, 27, 
    31, 2, 0, 27, 44, 35, 28, 27, 24, 23, 27, 25, 27, 28, 29, 
    37, 27, 7, 0, 0, 45, 47, 30, 24, 22, 24, 24, 25, 24, 27, 
    38, 30, 26, 14, 0, 0, 21, 37, 40, 33, 31, 24, 24, 25, 27, 
    37, 29, 27, 19, 0, 0, 0, 0, 0, 6, 33, 39, 41, 34, 28, 
    39, 26, 27, 2, 0, 0, 0, 3, 0, 0, 0, 0, 23, 21, 27, 
    43, 33, 32, 32, 34, 12, 23, 40, 27, 17, 28, 20, 31, 28, 28, 
    1, 0, 0, 0, 0, 0, 0, 12, 5, 9, 9, 13, 14, 11, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=198
    0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 25, 6, 0, 11, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 7, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 11, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 48, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 100, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 101, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 19, 51, 0, 0, 5, 25, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 3, 1, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 1, 0, 0, 0, 1, 0, 2, 0, 0, 0, 6, 
    
    -- channel=199
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=200
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=201
    39, 49, 47, 32, 33, 38, 35, 34, 36, 35, 35, 34, 34, 36, 38, 
    47, 53, 46, 4, 0, 0, 0, 0, 0, 0, 0, 4, 36, 37, 40, 
    45, 54, 40, 0, 0, 0, 0, 0, 0, 1, 1, 5, 29, 41, 42, 
    48, 53, 31, 0, 6, 8, 3, 3, 10, 0, 1, 11, 17, 42, 44, 
    48, 52, 48, 40, 36, 36, 37, 33, 37, 32, 32, 33, 43, 45, 48, 
    43, 47, 44, 41, 49, 48, 47, 46, 47, 48, 44, 49, 45, 44, 46, 
    40, 49, 39, 16, 20, 39, 45, 45, 45, 44, 43, 44, 44, 43, 44, 
    40, 46, 36, 38, 29, 12, 24, 37, 41, 40, 41, 43, 44, 45, 49, 
    37, 39, 40, 33, 29, 8, 10, 3, 10, 26, 38, 44, 44, 44, 47, 
    33, 35, 38, 31, 16, 3, 0, 3, 11, 9, 5, 2, 13, 31, 42, 
    32, 37, 39, 36, 26, 44, 27, 18, 37, 31, 35, 33, 28, 39, 38, 
    19, 21, 19, 16, 17, 13, 22, 30, 30, 33, 35, 35, 43, 38, 38, 
    22, 23, 24, 22, 20, 20, 22, 23, 22, 19, 19, 19, 18, 18, 17, 
    6, 4, 3, 3, 1, 2, 4, 3, 1, 3, 2, 3, 4, 7, 18, 
    3, 5, 5, 4, 3, 5, 7, 5, 6, 6, 5, 2, 13, 25, 27, 
    
    -- channel=202
    15, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    11, 2, 0, 0, 22, 25, 19, 25, 20, 24, 23, 24, 10, 2, 3, 
    11, 0, 0, 0, 0, 1, 0, 9, 0, 0, 0, 1, 23, 0, 2, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 16, 3, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 3, 10, 0, 0, 0, 
    2, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 34, 59, 14, 0, 0, 0, 0, 0, 0, 0, 1, 4, 
    15, 0, 0, 0, 0, 61, 51, 8, 0, 0, 0, 0, 0, 0, 0, 
    17, 4, 0, 0, 0, 3, 32, 67, 60, 29, 12, 0, 0, 0, 0, 
    20, 6, 3, 0, 0, 3, 7, 0, 3, 21, 64, 73, 60, 26, 3, 
    23, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    54, 42, 46, 49, 53, 32, 25, 36, 29, 12, 19, 10, 12, 17, 21, 
    0, 0, 0, 0, 0, 0, 0, 4, 3, 10, 11, 16, 18, 14, 20, 
    0, 8, 5, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=203
    29, 36, 38, 29, 27, 30, 29, 29, 29, 29, 29, 29, 30, 29, 30, 
    35, 41, 42, 8, 12, 9, 8, 9, 9, 12, 10, 12, 30, 32, 33, 
    34, 42, 42, 12, 1, 4, 0, 0, 5, 6, 9, 15, 16, 34, 34, 
    36, 42, 26, 8, 10, 10, 11, 5, 12, 7, 3, 9, 18, 35, 37, 
    36, 41, 42, 31, 31, 32, 33, 30, 32, 29, 26, 31, 33, 37, 39, 
    33, 41, 38, 37, 38, 39, 36, 35, 37, 37, 35, 35, 38, 36, 38, 
    30, 37, 35, 24, 31, 32, 37, 38, 38, 37, 36, 37, 36, 36, 37, 
    30, 37, 38, 30, 22, 20, 25, 31, 35, 36, 35, 36, 37, 37, 39, 
    27, 33, 33, 30, 39, 10, 8, 21, 25, 27, 31, 36, 36, 37, 39, 
    24, 30, 33, 34, 32, 12, 11, 10, 8, 13, 22, 25, 24, 28, 35, 
    25, 32, 33, 26, 36, 23, 16, 20, 21, 25, 21, 19, 22, 23, 32, 
    23, 28, 28, 27, 26, 34, 27, 22, 33, 42, 31, 39, 31, 38, 39, 
    23, 25, 26, 22, 21, 22, 23, 21, 25, 25, 24, 24, 25, 24, 22, 
    17, 14, 16, 14, 12, 13, 14, 13, 13, 11, 11, 11, 10, 10, 21, 
    13, 11, 11, 11, 11, 11, 12, 10, 11, 12, 12, 9, 10, 29, 13, 
    
    -- channel=204
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=205
    12, 13, 10, 3, 9, 4, 3, 6, 3, 4, 3, 5, 7, 3, 5, 
    14, 20, 17, 0, 0, 4, 1, 0, 0, 1, 0, 5, 9, 10, 8, 
    16, 19, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 10, 9, 
    13, 19, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 13, 
    9, 16, 18, 5, 8, 10, 13, 9, 9, 11, 6, 14, 2, 13, 13, 
    10, 14, 24, 19, 7, 7, 6, 5, 5, 7, 8, 5, 13, 11, 11, 
    9, 7, 0, 18, 36, 20, 11, 10, 10, 10, 12, 12, 13, 13, 14, 
    10, 12, 11, 0, 0, 26, 27, 13, 10, 10, 10, 10, 11, 11, 12, 
    9, 10, 9, 9, 0, 0, 7, 29, 31, 21, 17, 9, 10, 13, 14, 
    7, 7, 9, 5, 8, 7, 5, 0, 0, 10, 31, 36, 33, 22, 13, 
    8, 8, 9, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    24, 27, 30, 31, 32, 35, 24, 20, 29, 25, 24, 24, 19, 27, 26, 
    5, 8, 7, 7, 6, 9, 9, 12, 15, 19, 19, 21, 23, 21, 21, 
    7, 8, 9, 8, 5, 6, 5, 4, 4, 2, 2, 2, 2, 2, 5, 
    0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 10, 
    
    -- channel=206
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 81, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 38, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 67, 57, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 22, 0, 0, 25, 83, 99, 25, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 14, 
    30, 31, 23, 19, 16, 18, 14, 10, 1, 1, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    
    -- channel=207
    43, 50, 34, 29, 35, 37, 33, 31, 32, 32, 33, 32, 35, 39, 39, 
    46, 50, 42, 5, 18, 18, 14, 19, 17, 20, 20, 20, 46, 40, 41, 
    44, 48, 41, 9, 23, 25, 16, 23, 28, 29, 31, 30, 45, 42, 43, 
    44, 48, 30, 17, 20, 23, 16, 24, 22, 17, 20, 29, 28, 42, 41, 
    46, 47, 43, 37, 36, 33, 34, 34, 36, 32, 34, 38, 46, 42, 44, 
    45, 39, 33, 54, 43, 44, 45, 45, 45, 43, 42, 45, 43, 42, 43, 
    45, 38, 14, 0, 38, 52, 45, 45, 44, 42, 42, 43, 43, 42, 43, 
    47, 46, 37, 28, 0, 22, 47, 47, 41, 40, 40, 42, 43, 42, 44, 
    46, 42, 40, 35, 0, 4, 3, 9, 30, 43, 47, 43, 42, 41, 44, 
    45, 38, 40, 33, 0, 0, 1, 3, 0, 0, 3, 17, 36, 45, 46, 
    45, 41, 40, 35, 22, 12, 7, 20, 29, 1, 23, 4, 29, 33, 36, 
    29, 29, 26, 25, 25, 22, 29, 40, 33, 37, 37, 40, 41, 38, 39, 
    14, 21, 19, 17, 15, 15, 17, 19, 18, 16, 17, 16, 18, 17, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 
    
    -- channel=208
    10, 22, 16, 8, 8, 11, 8, 10, 9, 9, 9, 8, 12, 14, 12, 
    14, 22, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 12, 12, 
    14, 20, 19, 0, 2, 0, 0, 0, 0, 1, 1, 0, 5, 15, 14, 
    15, 21, 17, 0, 0, 6, 1, 0, 0, 0, 0, 0, 0, 14, 13, 
    17, 21, 23, 14, 7, 6, 8, 10, 8, 8, 7, 14, 15, 16, 16, 
    16, 17, 10, 22, 27, 26, 26, 26, 26, 25, 24, 18, 16, 15, 17, 
    12, 16, 3, 0, 0, 13, 18, 19, 19, 18, 17, 16, 15, 14, 13, 
    12, 19, 27, 22, 0, 0, 3, 12, 13, 13, 15, 16, 17, 17, 17, 
    12, 14, 14, 17, 0, 0, 0, 0, 0, 1, 12, 17, 16, 15, 16, 
    9, 10, 11, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 14, 
    7, 13, 12, 13, 32, 21, 15, 30, 29, 23, 27, 16, 25, 15, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 8, 3, 0, 2, 
    0, 9, 10, 9, 7, 8, 8, 5, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 
    
    -- channel=209
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 12, 24, 25, 19, 21, 21, 17, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 36, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 36, 22, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 26, 60, 48, 17, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 31, 9, 4, 0, 4, 44, 73, 73, 44, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 43, 51, 55, 58, 48, 17, 19, 38, 24, 15, 12, 10, 29, 26, 
    0, 0, 0, 0, 0, 0, 0, 1, 17, 22, 26, 30, 34, 37, 39, 
    24, 27, 25, 19, 15, 14, 11, 9, 5, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    
    -- channel=210
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 14, 6, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 6, 6, 8, 9, 14, 13, 11, 10, 13, 15, 14, 15, 15, 8, 
    10, 13, 14, 14, 13, 16, 12, 12, 12, 14, 13, 13, 13, 0, 0, 
    
    -- channel=211
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 16, 17, 15, 17, 16, 14, 13, 13, 12, 0, 0, 0, 
    0, 0, 0, 17, 14, 18, 19, 22, 13, 8, 10, 8, 0, 0, 0, 
    0, 0, 0, 40, 25, 22, 22, 27, 29, 27, 28, 19, 19, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 11, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 8, 17, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 14, 15, 10, 9, 15, 24, 22, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 3, 4, 6, 0, 0, 5, 8, 2, 2, 0, 5, 9, 6, 
    3, 3, 1, 0, 0, 0, 1, 5, 6, 6, 8, 8, 9, 10, 16, 
    19, 18, 16, 14, 12, 14, 12, 11, 8, 9, 8, 7, 9, 8, 0, 
    13, 10, 9, 8, 8, 6, 6, 4, 4, 3, 3, 4, 3, 0, 0, 
    
    -- channel=212
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 27, 13, 0, 0, 2, 0, 12, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=213
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=214
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 6, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    8, 3, 2, 4, 6, 5, 4, 5, 4, 6, 6, 4, 4, 0, 0, 
    8, 4, 1, 3, 3, 0, 3, 1, 2, 3, 7, 8, 0, 0, 9, 
    
    -- channel=215
    42, 69, 78, 61, 51, 67, 69, 59, 63, 62, 66, 64, 55, 66, 69, 
    48, 67, 80, 67, 37, 38, 48, 36, 45, 45, 48, 33, 61, 71, 70, 
    48, 68, 80, 40, 50, 30, 33, 20, 37, 47, 37, 32, 52, 74, 70, 
    52, 66, 89, 29, 39, 40, 43, 34, 40, 54, 42, 55, 24, 72, 70, 
    67, 67, 73, 83, 59, 58, 57, 57, 63, 65, 57, 47, 67, 73, 71, 
    71, 77, 67, 67, 70, 66, 64, 69, 71, 70, 66, 66, 74, 73, 70, 
    67, 89, 83, 36, 31, 61, 71, 75, 76, 77, 71, 74, 74, 74, 71, 
    64, 79, 85, 96, 38, 11, 39, 70, 76, 76, 71, 74, 74, 74, 71, 
    65, 75, 79, 85, 113, 17, 11, 24, 40, 58, 58, 74, 75, 74, 71, 
    64, 73, 76, 94, 116, 9, 7, 14, 20, 32, 9, 35, 40, 55, 66, 
    58, 74, 75, 103, 58, 72, 23, 0, 57, 40, 35, 34, 6, 47, 61, 
    45, 62, 62, 59, 55, 67, 44, 36, 61, 56, 53, 54, 55, 57, 57, 
    29, 36, 38, 36, 33, 31, 27, 26, 42, 34, 36, 33, 35, 41, 33, 
    21, 22, 25, 18, 22, 16, 16, 15, 20, 17, 12, 13, 12, 11, 3, 
    15, 14, 15, 11, 14, 9, 16, 10, 18, 15, 15, 14, 4, 20, 50, 
    
    -- channel=216
    20, 28, 30, 25, 21, 24, 21, 22, 22, 23, 22, 22, 22, 21, 21, 
    30, 35, 32, 20, 24, 26, 23, 24, 23, 22, 22, 21, 25, 26, 26, 
    30, 35, 42, 8, 0, 0, 0, 0, 0, 0, 0, 5, 18, 26, 28, 
    31, 35, 24, 2, 10, 15, 4, 8, 15, 11, 10, 10, 21, 30, 31, 
    28, 34, 32, 25, 25, 25, 28, 26, 27, 24, 22, 26, 24, 31, 31, 
    24, 33, 35, 24, 25, 24, 25, 24, 24, 24, 23, 29, 30, 30, 30, 
    22, 27, 25, 42, 31, 29, 32, 32, 30, 30, 30, 29, 30, 31, 31, 
    24, 29, 16, 0, 25, 35, 25, 27, 30, 28, 28, 28, 29, 30, 31, 
    24, 26, 26, 20, 9, 8, 25, 34, 26, 24, 29, 30, 30, 31, 32, 
    20, 24, 25, 27, 12, 9, 5, 2, 11, 27, 41, 32, 24, 24, 29, 
    20, 27, 27, 15, 1, 0, 6, 4, 0, 8, 0, 6, 10, 22, 29, 
    25, 31, 30, 31, 32, 23, 20, 27, 36, 28, 33, 27, 36, 42, 39, 
    13, 17, 17, 13, 11, 11, 15, 23, 24, 25, 26, 28, 29, 29, 27, 
    14, 16, 15, 11, 7, 8, 9, 7, 3, 2, 2, 1, 2, 0, 0, 
    1, 2, 2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 5, 12, 
    
    -- channel=217
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 23, 39, 33, 34, 35, 33, 31, 20, 0, 0, 0, 
    0, 0, 3, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 45, 54, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 56, 35, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 30, 70, 62, 29, 2, 0, 0, 0, 0, 
    0, 0, 0, 8, 3, 12, 7, 0, 2, 34, 72, 83, 59, 19, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    57, 63, 68, 72, 74, 59, 45, 44, 47, 34, 34, 26, 27, 36, 34, 
    0, 0, 0, 1, 3, 4, 7, 19, 26, 32, 35, 39, 42, 43, 42, 
    10, 16, 15, 9, 6, 5, 4, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    
    -- channel=218
    77, 87, 74, 66, 71, 74, 70, 72, 71, 72, 72, 72, 77, 84, 86, 
    82, 90, 83, 44, 48, 52, 49, 49, 50, 53, 54, 60, 82, 85, 86, 
    81, 87, 82, 47, 47, 50, 41, 50, 55, 55, 57, 59, 80, 86, 87, 
    80, 87, 66, 34, 50, 55, 48, 48, 52, 44, 47, 53, 66, 85, 88, 
    80, 86, 84, 73, 68, 68, 68, 70, 71, 68, 68, 79, 84, 86, 88, 
    84, 85, 80, 80, 85, 83, 85, 85, 84, 84, 84, 87, 85, 85, 88, 
    84, 73, 47, 55, 68, 81, 86, 88, 87, 85, 86, 86, 86, 86, 86, 
    88, 90, 83, 50, 42, 59, 77, 84, 84, 82, 83, 84, 85, 85, 87, 
    89, 89, 88, 84, 27, 25, 35, 51, 65, 73, 82, 85, 85, 85, 86, 
    86, 86, 86, 77, 19, 17, 19, 22, 25, 23, 39, 52, 67, 78, 84, 
    84, 85, 87, 71, 52, 34, 30, 53, 57, 44, 43, 37, 64, 74, 81, 
    70, 68, 65, 62, 62, 56, 60, 67, 66, 62, 70, 67, 72, 69, 71, 
    43, 44, 45, 43, 41, 39, 41, 46, 41, 40, 39, 40, 41, 38, 36, 
    17, 18, 18, 17, 14, 14, 15, 16, 15, 13, 14, 14, 14, 17, 34, 
    13, 15, 15, 15, 13, 16, 17, 18, 17, 17, 16, 14, 24, 42, 37, 
    
    -- channel=219
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 1, 0, 0, 8, 13, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 4, 3, 1, 0, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=220
    23, 28, 22, 17, 18, 21, 20, 20, 17, 19, 20, 19, 18, 15, 14, 
    28, 31, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 19, 17, 
    28, 31, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 20, 18, 
    27, 33, 24, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 24, 22, 
    26, 30, 29, 20, 22, 22, 24, 19, 22, 21, 18, 22, 15, 24, 23, 
    27, 25, 24, 30, 20, 19, 17, 17, 18, 19, 17, 16, 25, 23, 23, 
    24, 29, 19, 19, 31, 25, 23, 23, 22, 21, 21, 22, 22, 23, 23, 
    25, 25, 24, 4, 0, 20, 24, 20, 21, 22, 20, 22, 22, 23, 24, 
    23, 20, 18, 21, 4, 6, 6, 23, 22, 18, 22, 21, 22, 23, 24, 
    21, 17, 19, 15, 18, 10, 8, 3, 3, 19, 27, 27, 22, 20, 21, 
    22, 18, 19, 27, 13, 0, 10, 8, 0, 0, 4, 3, 10, 7, 19, 
    20, 19, 21, 21, 21, 28, 13, 13, 30, 28, 23, 26, 23, 33, 32, 
    11, 14, 12, 10, 7, 9, 8, 9, 16, 16, 17, 18, 19, 20, 17, 
    10, 14, 16, 12, 10, 11, 11, 9, 9, 6, 7, 6, 6, 9, 11, 
    1, 5, 7, 5, 5, 5, 3, 3, 4, 4, 2, 2, 8, 11, 13, 
    
    -- channel=221
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 5, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 13, 0, 0, 3, 6, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=222
    12, 18, 16, 13, 10, 15, 14, 14, 15, 15, 14, 12, 13, 10, 9, 
    17, 17, 16, 3, 0, 0, 0, 0, 0, 0, 0, 0, 4, 8, 8, 
    14, 18, 14, 0, 0, 1, 2, 0, 5, 8, 4, 3, 6, 8, 10, 
    16, 19, 9, 0, 1, 4, 0, 9, 2, 0, 0, 6, 7, 9, 9, 
    17, 19, 15, 12, 12, 11, 13, 12, 10, 8, 11, 11, 17, 13, 13, 
    14, 10, 2, 15, 20, 20, 18, 17, 17, 16, 16, 16, 14, 14, 16, 
    12, 24, 20, 0, 0, 7, 15, 15, 13, 12, 11, 10, 11, 10, 10, 
    11, 15, 11, 20, 8, 0, 0, 7, 10, 10, 11, 12, 13, 13, 15, 
    9, 9, 8, 7, 0, 0, 0, 0, 0, 0, 8, 13, 13, 12, 13, 
    7, 7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    8, 9, 9, 14, 27, 37, 37, 32, 30, 29, 36, 34, 29, 21, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 4, 1, 
    4, 6, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 6, 4, 3, 4, 4, 0, 0, 4, 9, 0, 
    
    -- channel=223
    44, 77, 93, 71, 62, 74, 76, 69, 74, 71, 74, 73, 69, 79, 86, 
    49, 75, 91, 87, 49, 63, 72, 62, 73, 71, 71, 62, 78, 88, 87, 
    48, 74, 93, 90, 72, 56, 64, 52, 69, 73, 70, 72, 71, 88, 87, 
    54, 71, 91, 55, 50, 51, 61, 48, 54, 61, 46, 55, 42, 81, 84, 
    70, 72, 86, 91, 68, 67, 68, 68, 73, 75, 64, 58, 85, 87, 87, 
    72, 84, 82, 80, 85, 83, 82, 87, 89, 85, 82, 81, 88, 88, 86, 
    69, 97, 85, 28, 38, 76, 86, 91, 93, 94, 87, 90, 87, 87, 85, 
    66, 90, 100, 113, 43, 8, 50, 87, 91, 90, 85, 88, 87, 88, 85, 
    66, 89, 95, 97, 135, 8, 2, 17, 50, 74, 75, 90, 89, 88, 87, 
    64, 86, 91, 105, 129, 0, 0, 12, 11, 13, 0, 33, 52, 72, 84, 
    59, 89, 90, 105, 81, 82, 11, 0, 64, 56, 35, 33, 1, 57, 70, 
    44, 72, 70, 66, 62, 75, 55, 45, 65, 70, 59, 67, 61, 63, 64, 
    32, 43, 44, 41, 38, 37, 33, 30, 46, 37, 38, 36, 38, 43, 34, 
    17, 11, 15, 9, 10, 4, 5, 5, 8, 6, 1, 3, 2, 0, 0, 
    16, 7, 4, 1, 5, 2, 9, 3, 9, 7, 6, 4, 0, 10, 29, 
    
    -- channel=224
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=225
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 15, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 74, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 20, 18, 42, 12, 0, 0, 18, 4, 16, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 2, 4, 0, 4, 3, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 
    
    -- channel=226
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 22, 20, 15, 18, 17, 19, 18, 0, 0, 0, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 18, 45, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 25, 29, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 13, 44, 48, 23, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 39, 8, 2, 0, 0, 26, 50, 60, 49, 19, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    33, 43, 50, 52, 55, 53, 27, 23, 37, 24, 19, 17, 14, 25, 24, 
    0, 0, 0, 0, 0, 0, 0, 2, 14, 19, 23, 24, 28, 30, 33, 
    18, 19, 18, 13, 11, 10, 7, 6, 3, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    
    -- channel=227
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 24, 10, 21, 26, 17, 19, 16, 19, 19, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 0, 0, 1, 0, 1, 8, 13, 9, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 6, 2, 0, 2, 3, 0, 0, 0, 0, 0, 
    0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 66, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 19, 42, 14, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 45, 67, 38, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 36, 21, 3, 0, 19, 67, 88, 67, 30, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 40, 46, 50, 55, 34, 6, 17, 39, 13, 16, 3, 17, 34, 28, 
    0, 0, 0, 0, 0, 0, 0, 3, 16, 20, 24, 30, 32, 35, 43, 
    37, 37, 32, 25, 23, 22, 18, 15, 9, 8, 5, 1, 3, 1, 0, 
    6, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    
    -- channel=228
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 6, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 0, 0, 0, 3, 0, 4, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=229
    0, 0, 13, 2, 0, 3, 4, 4, 10, 6, 5, 2, 6, 9, 2, 
    0, 0, 2, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 12, 10, 4, 14, 18, 12, 11, 0, 0, 0, 
    0, 0, 2, 22, 3, 6, 13, 11, 5, 0, 0, 6, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 
    0, 0, 0, 0, 26, 25, 23, 20, 22, 20, 19, 11, 0, 0, 1, 
    0, 18, 28, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 
    0, 0, 17, 82, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 34, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 80, 124, 73, 69, 98, 87, 101, 85, 54, 32, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 
    0, 0, 0, 0, 0, 10, 16, 14, 16, 17, 11, 3, 13, 30, 0, 
    
    -- channel=230
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 12, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 16, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 17, 20, 14, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 18, 16, 14, 18, 20, 20, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 10, 4, 0, 4, 5, 10, 5, 0, 0, 
    0, 2, 4, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 3, 4, 5, 8, 7, 6, 6, 6, 8, 8, 8, 8, 8, 10, 
    19, 18, 18, 20, 22, 20, 20, 20, 21, 21, 21, 21, 20, 20, 17, 
    19, 19, 18, 20, 20, 17, 18, 19, 18, 20, 21, 22, 17, 21, 22, 
    
    -- channel=231
    0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 1, 3, 3, 4, 3, 
    0, 0, 0, 2, 0, 0, 2, 3, 3, 0, 4, 1, 0, 0, 1, 
    0, 0, 0, 1, 8, 9, 14, 10, 10, 11, 9, 7, 5, 0, 0, 
    0, 0, 0, 3, 1, 3, 1, 5, 0, 2, 4, 2, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 2, 0, 0, 5, 6, 0, 0, 0, 0, 0, 0, 0, 
    5, 2, 1, 3, 0, 0, 0, 0, 3, 4, 3, 2, 0, 0, 0, 
    3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 1, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 6, 
    
    -- channel=232
    52, 67, 68, 55, 50, 62, 62, 57, 59, 59, 61, 60, 57, 62, 65, 
    56, 68, 72, 32, 22, 21, 25, 21, 24, 27, 29, 25, 58, 65, 65, 
    56, 69, 70, 23, 29, 24, 18, 15, 29, 34, 31, 28, 47, 67, 67, 
    57, 68, 61, 15, 28, 28, 30, 22, 27, 31, 27, 39, 29, 67, 67, 
    65, 67, 71, 66, 56, 55, 57, 53, 58, 58, 54, 53, 62, 68, 68, 
    68, 69, 62, 68, 66, 64, 62, 64, 65, 66, 63, 62, 69, 69, 68, 
    66, 76, 64, 31, 42, 61, 66, 69, 69, 68, 66, 68, 68, 68, 67, 
    66, 73, 77, 71, 26, 23, 46, 65, 67, 68, 66, 68, 68, 68, 68, 
    65, 70, 70, 72, 71, 17, 14, 28, 41, 54, 58, 67, 68, 68, 68, 
    62, 67, 69, 74, 72, 10, 13, 16, 18, 25, 19, 36, 44, 55, 63, 
    60, 66, 68, 78, 58, 51, 26, 18, 50, 38, 37, 34, 26, 46, 58, 
    44, 51, 52, 50, 48, 57, 41, 37, 55, 55, 49, 54, 50, 54, 56, 
    31, 34, 35, 32, 30, 29, 26, 24, 34, 29, 30, 28, 30, 31, 27, 
    21, 20, 23, 19, 20, 17, 17, 17, 20, 17, 15, 16, 15, 17, 28, 
    16, 15, 16, 15, 16, 15, 17, 15, 19, 18, 16, 15, 17, 39, 39, 
    
    -- channel=233
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 34, 2, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 3, 5, 5, 8, 6, 4, 4, 5, 7, 5, 5, 3, 1, 0, 
    12, 4, 3, 2, 5, 2, 2, 2, 4, 4, 5, 4, 0, 0, 0, 
    
    -- channel=234
    89, 96, 83, 86, 93, 94, 95, 91, 91, 93, 96, 95, 95, 105, 108, 
    86, 96, 98, 91, 110, 116, 115, 114, 119, 120, 118, 108, 116, 112, 111, 
    85, 93, 101, 98, 100, 97, 93, 101, 100, 102, 101, 101, 114, 110, 111, 
    83, 92, 98, 90, 96, 92, 90, 95, 97, 103, 103, 103, 99, 107, 109, 
    91, 92, 93, 94, 86, 85, 85, 90, 92, 89, 88, 96, 102, 105, 105, 
    102, 97, 90, 99, 88, 86, 91, 95, 92, 89, 91, 96, 105, 105, 106, 
    107, 90, 66, 75, 100, 106, 107, 109, 108, 106, 106, 106, 105, 107, 109, 
    111, 110, 101, 64, 34, 79, 108, 114, 111, 109, 105, 105, 105, 103, 103, 
    114, 116, 115, 112, 52, 31, 51, 89, 106, 109, 106, 107, 106, 105, 105, 
    116, 117, 117, 120, 62, 17, 26, 31, 35, 51, 67, 98, 106, 106, 107, 
    116, 113, 115, 108, 60, 22, 14, 34, 51, 21, 25, 19, 52, 80, 101, 
    103, 105, 105, 104, 102, 94, 74, 83, 97, 84, 84, 83, 84, 92, 93, 
    48, 50, 45, 41, 39, 37, 35, 44, 51, 50, 50, 52, 56, 57, 53, 
    33, 36, 36, 28, 26, 23, 21, 22, 22, 14, 13, 13, 12, 10, 10, 
    16, 13, 13, 13, 12, 13, 13, 13, 14, 12, 10, 11, 6, 16, 24, 
    
    -- channel=235
    10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 8, 5, 0, 6, 0, 4, 0, 9, 0, 0, 0, 
    6, 0, 0, 0, 0, 7, 0, 16, 4, 0, 7, 14, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 19, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 39, 26, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 27, 29, 20, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 9, 3, 7, 5, 38, 24, 20, 4, 0, 
    4, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 24, 0, 0, 
    16, 0, 0, 1, 6, 0, 1, 20, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 6, 0, 1, 1, 5, 5, 1, 6, 
    0, 3, 0, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    
    -- channel=236
    13, 26, 26, 19, 16, 19, 17, 16, 16, 16, 17, 18, 16, 18, 20, 
    18, 29, 27, 17, 5, 12, 13, 15, 16, 13, 17, 16, 15, 22, 23, 
    17, 29, 30, 19, 0, 0, 4, 0, 3, 4, 2, 9, 16, 22, 24, 
    17, 28, 19, 0, 0, 3, 0, 0, 1, 3, 0, 0, 7, 23, 26, 
    18, 27, 26, 26, 23, 25, 23, 22, 25, 22, 19, 17, 24, 25, 27, 
    16, 30, 35, 21, 18, 19, 18, 19, 20, 18, 17, 22, 25, 23, 25, 
    15, 22, 16, 28, 31, 24, 25, 26, 25, 25, 24, 26, 26, 27, 27, 
    15, 26, 16, 0, 11, 22, 25, 23, 26, 25, 22, 24, 24, 24, 27, 
    14, 22, 22, 18, 24, 0, 8, 28, 30, 27, 24, 25, 26, 26, 27, 
    12, 21, 22, 29, 31, 0, 0, 0, 0, 17, 30, 35, 29, 24, 25, 
    13, 24, 23, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 19, 
    28, 40, 40, 40, 41, 38, 26, 28, 40, 38, 33, 33, 34, 41, 40, 
    6, 11, 10, 8, 6, 7, 7, 12, 19, 18, 20, 21, 22, 23, 22, 
    4, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    
    -- channel=237
    0, 0, 17, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 26, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 8, 14, 0, 10, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 23, 9, 0, 0, 4, 0, 0, 12, 0, 6, 0, 0, 0, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    0, 29, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 22, 68, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 92, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 101, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 40, 44, 59, 2, 0, 24, 28, 15, 12, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 1, 4, 3, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    10, 0, 1, 0, 2, 0, 2, 0, 4, 2, 1, 0, 0, 0, 1, 
    
    -- channel=238
    10, 12, 12, 7, 5, 7, 9, 7, 11, 8, 9, 6, 12, 20, 15, 
    6, 4, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 4, 8, 
    3, 5, 0, 9, 24, 28, 21, 26, 33, 35, 30, 26, 7, 8, 8, 
    9, 6, 3, 9, 3, 3, 11, 2, 0, 0, 0, 4, 0, 1, 2, 
    17, 7, 10, 10, 0, 0, 0, 0, 0, 0, 0, 3, 16, 9, 7, 
    17, 7, 0, 17, 35, 34, 33, 32, 33, 32, 30, 19, 6, 8, 10, 
    13, 20, 11, 0, 0, 0, 9, 11, 13, 13, 9, 9, 6, 2, 1, 
    11, 13, 36, 87, 0, 0, 0, 3, 6, 5, 8, 9, 11, 10, 8, 
    10, 11, 11, 17, 32, 0, 0, 0, 0, 0, 0, 12, 8, 5, 7, 
    10, 7, 8, 1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 7, 
    5, 6, 6, 20, 77, 99, 45, 54, 93, 64, 86, 56, 45, 27, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 7, 11, 11, 11, 12, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 
    0, 0, 0, 0, 0, 9, 13, 11, 13, 14, 9, 5, 11, 31, 0, 
    
    -- channel=239
    49, 63, 57, 53, 55, 59, 58, 56, 57, 58, 60, 58, 60, 68, 69, 
    50, 62, 68, 55, 52, 59, 57, 58, 62, 61, 63, 57, 71, 71, 71, 
    50, 61, 65, 57, 53, 50, 48, 51, 55, 56, 55, 56, 66, 70, 71, 
    51, 61, 65, 45, 48, 48, 47, 47, 50, 53, 49, 54, 51, 67, 70, 
    58, 60, 62, 59, 49, 49, 50, 53, 54, 52, 49, 56, 66, 69, 69, 
    63, 62, 53, 65, 62, 61, 64, 66, 65, 62, 62, 64, 68, 69, 70, 
    65, 65, 41, 21, 43, 65, 70, 73, 72, 70, 68, 69, 68, 69, 69, 
    67, 74, 70, 53, 8, 23, 55, 72, 72, 70, 67, 68, 68, 68, 67, 
    69, 75, 74, 72, 35, 0, 3, 23, 44, 58, 66, 71, 69, 68, 68, 
    69, 74, 74, 73, 31, 0, 0, 0, 0, 0, 5, 28, 45, 60, 69, 
    66, 73, 73, 71, 48, 26, 5, 18, 41, 19, 22, 13, 28, 51, 62, 
    41, 49, 46, 43, 41, 39, 31, 38, 47, 45, 43, 46, 46, 49, 51, 
    16, 21, 19, 15, 11, 9, 9, 11, 15, 11, 11, 10, 12, 13, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=240
    67, 75, 68, 68, 68, 74, 73, 72, 70, 73, 74, 73, 74, 77, 82, 
    70, 81, 77, 64, 73, 77, 78, 77, 79, 80, 78, 77, 81, 86, 86, 
    70, 78, 87, 55, 49, 43, 46, 46, 47, 50, 52, 57, 77, 85, 88, 
    66, 76, 69, 51, 55, 58, 52, 57, 62, 63, 62, 65, 70, 87, 87, 
    67, 75, 74, 68, 69, 70, 70, 70, 72, 71, 71, 75, 76, 82, 84, 
    75, 76, 82, 73, 61, 61, 63, 65, 63, 64, 65, 74, 83, 84, 83, 
    81, 66, 54, 84, 95, 85, 82, 83, 82, 80, 81, 82, 84, 86, 87, 
    85, 84, 69, 23, 34, 83, 95, 88, 86, 83, 82, 81, 81, 80, 82, 
    87, 89, 89, 82, 27, 30, 61, 96, 98, 88, 84, 81, 82, 83, 83, 
    87, 90, 90, 90, 46, 23, 25, 23, 37, 63, 89, 103, 97, 88, 82, 
    87, 88, 89, 75, 21, 0, 3, 15, 12, 4, 0, 6, 32, 59, 79, 
    92, 97, 99, 99, 101, 84, 63, 76, 89, 71, 74, 68, 74, 84, 84, 
    36, 35, 30, 29, 28, 27, 26, 38, 45, 46, 48, 52, 55, 55, 53, 
    38, 42, 39, 34, 32, 28, 26, 26, 24, 19, 18, 16, 16, 14, 17, 
    15, 15, 15, 15, 15, 12, 10, 13, 13, 10, 11, 11, 12, 21, 44, 
    
    -- channel=241
    62, 77, 76, 61, 62, 72, 72, 72, 75, 73, 73, 72, 80, 86, 84, 
    61, 68, 78, 53, 32, 20, 23, 24, 26, 27, 28, 38, 70, 76, 80, 
    58, 67, 64, 49, 68, 70, 62, 67, 77, 78, 76, 70, 62, 80, 80, 
    63, 68, 67, 71, 64, 69, 72, 65, 63, 60, 59, 66, 66, 73, 74, 
    72, 68, 75, 68, 53, 49, 54, 58, 54, 57, 57, 68, 81, 76, 76, 
    76, 67, 43, 74, 94, 92, 93, 93, 93, 91, 91, 80, 74, 78, 79, 
    77, 83, 61, 0, 0, 56, 77, 80, 82, 79, 75, 75, 73, 71, 71, 
    77, 83, 105, 119, 33, 0, 25, 70, 75, 74, 76, 76, 78, 78, 76, 
    77, 82, 83, 92, 63, 13, 0, 0, 0, 34, 61, 79, 76, 73, 73, 
    76, 79, 81, 67, 24, 0, 7, 19, 7, 0, 0, 0, 0, 44, 71, 
    70, 79, 79, 88, 129, 119, 75, 100, 127, 110, 109, 93, 90, 86, 70, 
    6, 2, 0, 0, 0, 2, 15, 10, 9, 21, 25, 34, 28, 17, 21, 
    33, 36, 39, 35, 32, 30, 27, 14, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 7, 8, 8, 9, 9, 16, 54, 
    14, 12, 13, 13, 14, 23, 26, 27, 29, 29, 22, 18, 33, 57, 9, 
    
    -- channel=242
    3, 11, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 9, 
    2, 6, 11, 3, 0, 0, 0, 0, 0, 0, 0, 0, 4, 6, 7, 
    1, 4, 9, 14, 20, 23, 24, 18, 28, 30, 28, 30, 8, 11, 9, 
    3, 4, 7, 6, 0, 0, 6, 3, 0, 0, 0, 0, 0, 4, 3, 
    3, 2, 7, 13, 1, 0, 0, 0, 3, 0, 0, 0, 16, 6, 5, 
    3, 17, 16, 5, 17, 20, 20, 19, 21, 20, 19, 14, 3, 1, 1, 
    1, 0, 0, 0, 1, 6, 2, 4, 6, 9, 8, 10, 9, 7, 4, 
    2, 4, 15, 28, 5, 0, 10, 4, 3, 4, 6, 6, 7, 6, 5, 
    3, 6, 7, 7, 17, 0, 0, 0, 11, 16, 4, 4, 4, 4, 4, 
    3, 6, 6, 16, 0, 0, 0, 4, 0, 0, 0, 0, 17, 15, 6, 
    0, 5, 3, 0, 0, 9, 0, 0, 23, 0, 5, 0, 0, 3, 0, 
    21, 27, 23, 20, 18, 25, 47, 31, 7, 23, 23, 27, 19, 0, 7, 
    5, 9, 16, 21, 23, 22, 25, 18, 10, 8, 7, 3, 2, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 14, 16, 
    
    -- channel=243
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 23, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 43, 19, 0, 15, 17, 19, 21, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 1, 1, 3, 7, 5, 6, 6, 8, 1, 
    8, 6, 6, 6, 8, 6, 10, 8, 11, 10, 10, 9, 6, 1, 9, 
    
    -- channel=244
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 11, 29, 1, 0, 11, 9, 9, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=245
    26, 29, 21, 21, 28, 27, 26, 27, 25, 28, 27, 26, 25, 21, 25, 
    32, 38, 25, 5, 15, 16, 16, 16, 13, 14, 17, 20, 29, 29, 29, 
    33, 36, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 29, 30, 
    30, 35, 19, 0, 10, 14, 4, 9, 18, 13, 17, 14, 30, 32, 34, 
    27, 35, 28, 19, 26, 27, 28, 26, 25, 24, 26, 30, 23, 30, 33, 
    28, 25, 27, 25, 16, 14, 16, 16, 14, 15, 16, 26, 33, 33, 33, 
    30, 26, 22, 46, 40, 34, 33, 32, 29, 26, 29, 28, 30, 32, 34, 
    34, 32, 9, 0, 4, 43, 37, 32, 31, 29, 29, 28, 29, 29, 32, 
    34, 30, 29, 21, 0, 3, 33, 47, 32, 26, 32, 29, 31, 31, 32, 
    32, 29, 30, 21, 0, 0, 0, 0, 10, 37, 57, 42, 30, 27, 30, 
    33, 31, 32, 20, 0, 0, 3, 5, 0, 0, 0, 0, 14, 21, 35, 
    26, 27, 27, 28, 32, 12, 1, 22, 33, 15, 22, 13, 27, 38, 35, 
    0, 2, 0, 0, 0, 0, 0, 5, 9, 11, 13, 18, 20, 19, 24, 
    9, 17, 13, 9, 3, 3, 3, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    
    -- channel=246
    0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 19, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 25, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 13, 62, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 106, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 107, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 38, 26, 72, 8, 0, 23, 35, 10, 23, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 3, 0, 4, 2, 3, 1, 0, 0, 16, 
    
    -- channel=247
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 1, 0, 0, 3, 0, 0, 0, 0, 0, 
    1, 3, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 11, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 7, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 4, 36, 2, 0, 8, 8, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 44, 4, 4, 3, 1, 10, 7, 15, 9, 0, 0, 
    0, 0, 0, 7, 6, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 8, 13, 14, 13, 24, 6, 0, 4, 6, 0, 0, 0, 0, 0, 
    4, 0, 2, 3, 5, 6, 2, 0, 9, 9, 9, 9, 11, 11, 11, 
    16, 10, 14, 13, 15, 12, 11, 12, 15, 14, 13, 12, 10, 10, 14, 
    17, 10, 9, 9, 11, 8, 8, 7, 9, 9, 10, 13, 8, 17, 13, 
    
    -- channel=248
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 20, 17, 14, 16, 17, 16, 13, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 38, 60, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 50, 37, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 25, 71, 64, 27, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 15, 13, 7, 0, 0, 36, 78, 88, 63, 19, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    52, 60, 68, 71, 75, 66, 39, 37, 49, 33, 30, 24, 21, 35, 35, 
    0, 0, 0, 0, 0, 0, 0, 7, 18, 25, 28, 32, 36, 37, 40, 
    18, 21, 20, 15, 12, 11, 8, 6, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    
    -- channel=249
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=250
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 0, 9, 2, 2, 3, 14, 0, 0, 0, 
    0, 0, 0, 13, 0, 5, 4, 15, 2, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 15, 1, 1, 0, 2, 2, 0, 1, 0, 11, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 18, 18, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 16, 19, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 10, 5, 0, 0, 20, 19, 20, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 1, 0, 0, 
    3, 0, 1, 3, 6, 0, 4, 8, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 3, 0, 0, 0, 1, 0, 0, 1, 0, 1, 4, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 
    
    -- channel=251
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 19, 23, 28, 28, 27, 28, 25, 23, 12, 0, 0, 0, 
    0, 0, 0, 20, 16, 10, 19, 14, 7, 7, 7, 4, 0, 0, 0, 
    0, 0, 3, 20, 10, 6, 10, 11, 10, 22, 16, 12, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 5, 12, 22, 13, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 27, 8, 9, 6, 7, 25, 27, 24, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 10, 13, 15, 15, 14, 0, 0, 10, 1, 0, 0, 0, 6, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 6, 8, 9, 11, 14, 13, 
    13, 18, 19, 14, 13, 12, 10, 9, 8, 5, 5, 4, 4, 0, 0, 
    4, 5, 4, 3, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=252
    48, 59, 48, 42, 47, 49, 47, 45, 45, 45, 47, 47, 48, 55, 54, 
    50, 59, 56, 36, 35, 39, 36, 35, 37, 39, 40, 38, 55, 57, 57, 
    49, 56, 54, 33, 35, 32, 27, 29, 35, 37, 32, 33, 53, 58, 57, 
    50, 56, 58, 25, 38, 36, 33, 36, 38, 38, 39, 41, 40, 57, 58, 
    51, 55, 56, 53, 45, 46, 44, 46, 49, 46, 45, 51, 54, 57, 57, 
    53, 58, 55, 51, 53, 52, 54, 55, 53, 53, 53, 54, 56, 55, 56, 
    53, 46, 30, 39, 49, 54, 56, 58, 57, 56, 56, 57, 57, 58, 58, 
    55, 58, 53, 28, 23, 40, 52, 55, 57, 56, 55, 55, 56, 56, 57, 
    56, 57, 57, 55, 22, 12, 20, 38, 47, 51, 54, 57, 57, 56, 56, 
    55, 56, 57, 57, 21, 9, 8, 9, 12, 18, 29, 43, 47, 52, 55, 
    54, 57, 57, 51, 22, 12, 7, 16, 27, 11, 14, 10, 29, 42, 52, 
    52, 55, 53, 52, 51, 47, 44, 49, 55, 50, 53, 52, 55, 56, 56, 
    23, 28, 28, 26, 23, 21, 23, 27, 27, 26, 26, 26, 27, 27, 26, 
    5, 10, 9, 6, 5, 3, 4, 3, 4, 1, 1, 2, 2, 3, 1, 
    0, 2, 3, 2, 0, 0, 2, 0, 1, 0, 1, 1, 1, 11, 20, 
    
    -- channel=253
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 15, 12, 14, 17, 14, 16, 13, 14, 12, 0, 0, 0, 
    0, 0, 0, 25, 17, 17, 23, 20, 16, 15, 12, 3, 0, 0, 0, 
    0, 0, 0, 12, 12, 11, 11, 8, 9, 12, 12, 10, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 10, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 36, 8, 3, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 21, 15, 5, 2, 5, 21, 3, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 4, 7, 7, 9, 7, 6, 7, 8, 9, 8, 7, 7, 7, 0, 
    20, 8, 8, 6, 10, 7, 10, 9, 11, 10, 11, 8, 5, 0, 0, 
    
    -- channel=254
    27, 35, 30, 36, 36, 37, 36, 34, 34, 35, 37, 36, 37, 44, 42, 
    23, 29, 37, 62, 67, 70, 68, 69, 73, 71, 69, 58, 49, 45, 44, 
    22, 26, 40, 70, 67, 65, 69, 70, 66, 67, 65, 63, 50, 42, 43, 
    24, 27, 48, 68, 56, 52, 56, 59, 58, 64, 59, 60, 47, 39, 40, 
    27, 27, 30, 40, 34, 34, 30, 37, 38, 35, 35, 35, 44, 38, 37, 
    31, 33, 31, 34, 30, 31, 35, 38, 36, 32, 33, 36, 38, 37, 36, 
    34, 27, 19, 25, 38, 40, 40, 42, 41, 40, 40, 40, 39, 41, 41, 
    35, 38, 35, 26, 12, 29, 43, 44, 44, 43, 40, 39, 39, 38, 36, 
    38, 42, 43, 42, 27, 9, 15, 34, 45, 46, 42, 43, 40, 38, 37, 
    41, 45, 45, 52, 30, 4, 8, 12, 10, 14, 22, 40, 42, 42, 41, 
    40, 46, 44, 41, 18, 5, 0, 2, 16, 0, 1, 0, 11, 28, 37, 
    41, 51, 48, 48, 46, 41, 35, 40, 44, 42, 39, 40, 40, 43, 43, 
    14, 20, 18, 15, 13, 12, 12, 15, 18, 16, 16, 16, 17, 20, 16, 
    4, 8, 7, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=255
    25, 4, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 6, 7, 0, 
    26, 9, 0, 0, 17, 0, 0, 2, 0, 0, 0, 2, 9, 0, 0, 
    23, 7, 0, 0, 0, 8, 0, 10, 0, 1, 2, 12, 14, 0, 0, 
    18, 7, 0, 0, 1, 0, 0, 8, 1, 0, 6, 0, 28, 0, 0, 
    6, 8, 0, 0, 0, 0, 0, 1, 0, 0, 1, 17, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 5, 0, 0, 0, 3, 10, 0, 0, 2, 
    12, 0, 0, 14, 14, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 0, 0, 0, 0, 42, 19, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 1, 0, 0, 0, 15, 31, 20, 4, 0, 3, 0, 0, 0, 0, 
    20, 1, 0, 0, 0, 0, 10, 5, 10, 0, 23, 5, 4, 1, 1, 
    22, 0, 0, 0, 0, 0, 16, 56, 3, 0, 15, 3, 68, 26, 11, 
    10, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 25, 
    0, 0, 0, 3, 0, 7, 1, 7, 0, 1, 0, 0, 10, 28, 0, 
    
    -- channel=256
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=257
    18, 24, 17, 13, 20, 12, 20, 17, 20, 16, 20, 12, 32, 10, 16, 
    20, 23, 21, 13, 22, 10, 13, 13, 20, 18, 23, 8, 36, 22, 18, 
    7, 7, 15, 13, 19, 17, 26, 21, 11, 15, 14, 14, 27, 17, 23, 
    19, 12, 22, 13, 22, 22, 25, 21, 10, 23, 24, 18, 21, 19, 15, 
    21, 7, 20, 24, 13, 26, 30, 21, 30, 25, 26, 25, 26, 12, 22, 
    20, 4, 17, 26, 23, 25, 35, 23, 27, 28, 31, 23, 27, 12, 29, 
    23, 11, 12, 19, 31, 25, 29, 23, 23, 23, 22, 20, 28, 16, 32, 
    15, 10, 8, 15, 19, 30, 15, 29, 29, 29, 25, 17, 21, 16, 19, 
    19, 20, 16, 14, 14, 15, 24, 23, 19, 17, 29, 18, 24, 17, 19, 
    14, 12, 11, 6, 8, 18, 15, 15, 23, 19, 19, 24, 18, 12, 19, 
    15, 13, 26, 16, 20, 9, 15, 20, 14, 20, 15, 23, 28, 22, 14, 
    26, 33, 43, 23, 17, 18, 13, 20, 17, 22, 18, 24, 28, 18, 18, 
    5, 10, 33, 43, 28, 20, 18, 17, 8, 18, 23, 23, 26, 17, 17, 
    16, 6, 6, 31, 46, 32, 26, 27, 19, 15, 16, 26, 19, 8, 19, 
    26, 20, 13, 15, 31, 39, 39, 28, 26, 13, 11, 14, 29, 24, 20, 
    
    -- channel=258
    23, 23, 31, 26, 22, 32, 29, 28, 27, 24, 21, 26, 21, 21, 19, 
    20, 23, 25, 24, 21, 27, 21, 22, 30, 27, 25, 25, 22, 30, 25, 
    16, 25, 19, 18, 21, 30, 35, 30, 26, 12, 30, 23, 19, 21, 24, 
    22, 28, 17, 20, 22, 41, 31, 17, 21, 26, 30, 27, 21, 20, 12, 
    22, 29, 21, 16, 35, 31, 13, 29, 37, 33, 31, 27, 19, 15, 11, 
    16, 25, 23, 21, 28, 16, 21, 37, 26, 20, 19, 28, 19, 20, 18, 
    22, 22, 18, 21, 18, 15, 16, 6, 7, 14, 13, 7, 16, 21, 20, 
    17, 21, 14, 16, 22, 0, 8, 11, 17, 7, 0, 12, 6, 16, 8, 
    23, 21, 16, 18, 6, 16, 8, 8, 1, 0, 7, 5, 2, 17, 24, 
    18, 15, 15, 22, 20, 8, 10, 4, 2, 3, 2, 5, 7, 10, 21, 
    12, 28, 24, 27, 15, 17, 10, 3, 1, 0, 3, 5, 11, 18, 28, 
    22, 31, 28, 23, 25, 12, 13, 4, 0, 3, 5, 6, 15, 22, 26, 
    11, 21, 32, 30, 24, 31, 15, 2, 8, 7, 5, 2, 10, 15, 28, 
    19, 9, 25, 32, 29, 30, 24, 23, 11, 5, 7, 2, 7, 26, 28, 
    27, 33, 21, 29, 32, 28, 29, 22, 15, 12, 11, 10, 15, 20, 30, 
    
    -- channel=259
    4, 1, 11, 15, 0, 17, 3, 11, 9, 10, 2, 23, 0, 14, 10, 
    8, 8, 9, 16, 0, 14, 8, 17, 3, 13, 0, 28, 0, 16, 6, 
    10, 3, 13, 13, 0, 12, 11, 9, 12, 9, 7, 28, 0, 14, 8, 
    3, 19, 11, 0, 7, 16, 7, 0, 27, 0, 18, 24, 0, 12, 0, 
    5, 28, 0, 7, 8, 8, 0, 17, 4, 11, 6, 14, 7, 14, 0, 
    0, 30, 11, 0, 22, 2, 0, 2, 5, 6, 1, 21, 2, 16, 0, 
    0, 24, 24, 6, 0, 0, 0, 2, 0, 0, 0, 6, 3, 21, 0, 
    5, 20, 21, 12, 0, 2, 0, 0, 0, 0, 2, 0, 0, 16, 0, 
    10, 18, 15, 13, 12, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    16, 8, 9, 16, 4, 14, 0, 0, 0, 0, 0, 0, 0, 12, 19, 
    1, 11, 3, 14, 21, 0, 14, 0, 0, 0, 0, 0, 0, 9, 19, 
    6, 5, 0, 22, 5, 19, 2, 0, 0, 0, 0, 0, 0, 12, 15, 
    20, 11, 0, 3, 3, 15, 0, 0, 2, 0, 0, 0, 0, 17, 18, 
    1, 28, 15, 0, 0, 6, 6, 0, 17, 0, 0, 0, 0, 22, 9, 
    0, 0, 32, 15, 0, 2, 7, 10, 4, 0, 0, 0, 0, 13, 31, 
    
    -- channel=260
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=261
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 
    0, 9, 0, 0, 0, 7, 0, 0, 7, 0, 10, 15, 1, 0, 0, 
    0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 4, 0, 
    0, 39, 4, 0, 8, 0, 0, 9, 0, 0, 0, 6, 0, 9, 0, 
    0, 18, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 
    0, 11, 3, 5, 0, 0, 0, 0, 0, 0, 0, 9, 0, 3, 0, 
    0, 2, 0, 2, 19, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 2, 23, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 7, 0, 0, 28, 3, 0, 0, 0, 0, 0, 0, 11, 
    0, 3, 0, 2, 0, 6, 17, 6, 0, 0, 0, 0, 0, 2, 0, 
    18, 34, 0, 0, 0, 14, 11, 0, 13, 0, 5, 0, 0, 0, 1, 
    0, 12, 39, 1, 0, 0, 0, 0, 3, 8, 0, 0, 0, 0, 0, 
    0, 0, 23, 40, 4, 0, 0, 0, 0, 6, 7, 0, 0, 0, 36, 
    
    -- channel=262
    0, 20, 0, 0, 35, 0, 0, 0, 0, 0, 14, 0, 51, 0, 0, 
    0, 14, 1, 0, 45, 0, 0, 0, 0, 0, 13, 0, 44, 0, 3, 
    1, 0, 0, 3, 43, 0, 0, 1, 0, 24, 0, 0, 14, 0, 0, 
    18, 0, 6, 15, 9, 0, 0, 33, 0, 30, 0, 0, 0, 0, 25, 
    23, 0, 31, 12, 0, 0, 42, 0, 0, 0, 0, 0, 0, 0, 61, 
    41, 0, 0, 49, 0, 0, 17, 0, 1, 0, 3, 0, 7, 0, 71, 
    35, 0, 0, 0, 11, 0, 6, 0, 0, 0, 0, 0, 6, 0, 60, 
    17, 0, 0, 0, 0, 24, 0, 0, 5, 0, 0, 0, 23, 0, 63, 
    0, 0, 0, 0, 0, 26, 0, 0, 0, 0, 2, 0, 6, 10, 40, 
    0, 6, 14, 0, 0, 0, 0, 0, 0, 0, 2, 2, 26, 0, 0, 
    32, 0, 18, 0, 0, 9, 0, 0, 1, 2, 0, 0, 11, 0, 0, 
    0, 0, 30, 0, 6, 0, 0, 0, 0, 16, 0, 2, 15, 0, 0, 
    0, 0, 8, 12, 8, 0, 0, 14, 0, 0, 0, 17, 18, 0, 0, 
    15, 0, 0, 0, 15, 0, 0, 10, 0, 0, 0, 17, 49, 0, 0, 
    25, 7, 0, 0, 0, 8, 4, 0, 2, 0, 0, 11, 25, 0, 0, 
    
    -- channel=263
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=264
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=265
    11, 10, 15, 22, 12, 6, 8, 10, 7, 6, 8, 10, 2, 2, 7, 
    17, 15, 17, 22, 9, 6, 5, 8, 10, 15, 6, 11, 2, 15, 20, 
    7, 4, 14, 17, 7, 6, 16, 15, 14, 13, 0, 15, 10, 21, 10, 
    13, 13, 15, 10, 7, 17, 8, 2, 5, 9, 13, 16, 7, 18, 14, 
    16, 18, 23, 5, 6, 14, 7, 5, 15, 10, 7, 6, 10, 20, 11, 
    12, 14, 19, 23, 18, 0, 0, 13, 13, 2, 0, 10, 9, 23, 7, 
    16, 18, 22, 15, 0, 0, 0, 0, 0, 0, 0, 1, 7, 22, 7, 
    13, 16, 22, 11, 0, 0, 0, 0, 0, 0, 0, 0, 3, 17, 12, 
    16, 22, 19, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 11, 
    20, 13, 14, 8, 12, 0, 0, 0, 0, 0, 0, 0, 0, 12, 10, 
    17, 6, 12, 16, 15, 13, 0, 0, 0, 0, 0, 0, 0, 13, 32, 
    11, 19, 15, 20, 18, 6, 0, 0, 0, 0, 0, 0, 0, 11, 25, 
    6, 0, 5, 12, 12, 12, 0, 0, 0, 0, 0, 0, 0, 11, 19, 
    8, 0, 0, 1, 10, 12, 1, 2, 5, 0, 0, 0, 0, 7, 14, 
    3, 1, 0, 0, 1, 16, 14, 9, 0, 0, 0, 0, 7, 18, 13, 
    
    -- channel=266
    0, 0, 0, 0, 0, 12, 0, 3, 14, 19, 0, 23, 0, 22, 0, 
    0, 0, 0, 0, 0, 17, 4, 3, 0, 0, 0, 31, 0, 0, 0, 
    7, 14, 0, 0, 0, 0, 0, 0, 15, 0, 23, 25, 0, 0, 0, 
    0, 12, 0, 0, 0, 16, 4, 0, 20, 0, 16, 21, 15, 0, 0, 
    0, 45, 0, 0, 13, 4, 0, 0, 0, 1, 13, 30, 11, 4, 0, 
    0, 56, 10, 0, 10, 2, 0, 10, 0, 7, 4, 16, 5, 12, 0, 
    0, 22, 28, 0, 0, 10, 0, 3, 10, 13, 1, 4, 9, 11, 0, 
    0, 18, 2, 11, 0, 0, 23, 12, 0, 0, 0, 27, 0, 18, 0, 
    0, 0, 8, 14, 32, 0, 12, 8, 4, 15, 10, 9, 16, 15, 0, 
    0, 7, 0, 24, 11, 48, 1, 4, 10, 5, 4, 5, 0, 0, 10, 
    0, 20, 0, 13, 0, 0, 44, 8, 3, 10, 10, 7, 0, 0, 5, 
    0, 0, 0, 2, 0, 12, 22, 24, 12, 0, 9, 8, 6, 21, 8, 
    38, 79, 7, 0, 0, 26, 19, 24, 48, 6, 17, 0, 0, 23, 11, 
    0, 50, 94, 24, 0, 0, 13, 0, 0, 24, 13, 0, 0, 27, 5, 
    0, 0, 59, 84, 28, 0, 0, 4, 6, 35, 38, 10, 0, 0, 42, 
    
    -- channel=267
    12, 15, 12, 21, 20, 10, 13, 13, 8, 12, 18, 12, 11, 3, 19, 
    13, 21, 15, 21, 22, 4, 11, 15, 14, 14, 13, 8, 12, 11, 14, 
    20, 17, 22, 19, 22, 6, 13, 17, 13, 19, 10, 7, 13, 17, 21, 
    16, 7, 18, 17, 18, 5, 16, 12, 13, 19, 0, 14, 12, 19, 16, 
    22, 7, 24, 14, 11, 10, 11, 18, 3, 11, 9, 9, 12, 21, 20, 
    22, 6, 21, 24, 8, 5, 14, 3, 14, 7, 8, 16, 12, 20, 21, 
    24, 7, 17, 24, 4, 0, 0, 0, 4, 1, 1, 1, 14, 20, 24, 
    22, 13, 23, 19, 0, 2, 0, 1, 0, 0, 1, 1, 11, 18, 22, 
    19, 16, 19, 16, 4, 17, 0, 0, 0, 0, 2, 0, 5, 9, 25, 
    23, 14, 25, 18, 10, 0, 3, 3, 2, 0, 4, 1, 2, 18, 16, 
    18, 16, 19, 7, 18, 18, 0, 0, 6, 3, 0, 0, 4, 14, 19, 
    20, 3, 13, 15, 20, 11, 0, 0, 4, 8, 0, 0, 0, 13, 22, 
    12, 3, 11, 15, 14, 16, 0, 0, 1, 2, 0, 0, 1, 10, 26, 
    13, 6, 0, 11, 11, 11, 7, 11, 6, 0, 4, 2, 2, 24, 9, 
    15, 8, 0, 0, 9, 12, 14, 7, 13, 0, 0, 2, 17, 1, 5, 
    
    -- channel=268
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=269
    0, 3, 0, 12, 8, 8, 3, 11, 5, 15, 6, 15, 0, 9, 6, 
    5, 2, 7, 10, 9, 4, 12, 8, 5, 4, 5, 10, 0, 0, 0, 
    10, 16, 12, 12, 10, 2, 0, 4, 19, 6, 11, 9, 0, 5, 6, 
    7, 0, 0, 3, 10, 0, 7, 19, 4, 7, 0, 1, 6, 6, 0, 
    8, 10, 0, 4, 4, 4, 1, 3, 0, 0, 0, 23, 2, 9, 2, 
    9, 13, 17, 0, 0, 2, 0, 0, 0, 3, 3, 2, 2, 15, 0, 
    0, 3, 17, 11, 0, 0, 0, 0, 0, 0, 0, 0, 2, 10, 6, 
    10, 9, 7, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 9, 
    8, 2, 16, 17, 11, 0, 0, 0, 0, 0, 0, 0, 5, 7, 6, 
    6, 15, 10, 12, 3, 12, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    7, 6, 5, 10, 7, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 
    8, 0, 0, 4, 11, 13, 0, 0, 0, 0, 0, 0, 0, 0, 20, 
    14, 26, 0, 0, 0, 8, 2, 0, 10, 0, 0, 0, 0, 13, 17, 
    0, 17, 25, 6, 0, 0, 1, 0, 0, 0, 0, 0, 0, 7, 21, 
    5, 0, 12, 19, 6, 0, 0, 0, 2, 1, 0, 1, 0, 0, 0, 
    
    -- channel=270
    0, 0, 0, 0, 0, 5, 0, 0, 3, 0, 0, 0, 0, 19, 0, 
    0, 0, 0, 0, 0, 27, 0, 8, 0, 0, 0, 7, 0, 0, 0, 
    14, 0, 0, 4, 0, 0, 0, 1, 0, 24, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 34, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 14, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 
    0, 95, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 10, 0, 
    0, 0, 87, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 14, 
    
    -- channel=271
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 1, 0, 0, 
    0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 19, 1, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    0, 15, 8, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 8, 0, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 2, 1, 15, 0, 1, 0, 0, 0, 0, 8, 1, 1, 0, 
    0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 2, 0, 12, 12, 0, 6, 0, 0, 0, 0, 0, 
    0, 3, 0, 3, 0, 4, 8, 8, 10, 0, 1, 0, 0, 0, 8, 
    1, 11, 0, 0, 0, 0, 10, 3, 4, 0, 9, 0, 0, 0, 0, 
    0, 5, 0, 0, 0, 2, 0, 0, 4, 7, 0, 0, 0, 0, 0, 
    0, 0, 4, 1, 0, 0, 0, 0, 0, 5, 6, 0, 0, 2, 0, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=272
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    
    -- channel=273
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 19, 0, 0, 4, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 10, 0, 
    0, 8, 9, 3, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 26, 0, 0, 0, 0, 0, 20, 25, 0, 0, 0, 0, 5, 0, 
    0, 33, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 
    0, 0, 0, 16, 0, 0, 0, 0, 5, 11, 19, 10, 0, 0, 0, 
    
    -- channel=274
    4, 20, 14, 14, 25, 29, 9, 9, 0, 0, 0, 0, 0, 21, 11, 
    0, 0, 3, 8, 24, 29, 19, 15, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 6, 7, 26, 28, 7, 0, 4, 8, 3, 0, 0, 0, 0, 
    13, 10, 0, 9, 26, 0, 0, 23, 16, 5, 0, 0, 0, 0, 0, 
    7, 0, 0, 7, 0, 0, 2, 17, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 18, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 
    
    -- channel=275
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 14, 3, 0, 0, 0, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 2, 4, 4, 0, 3, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 1, 4, 0, 8, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 6, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 12, 7, 0, 0, 8, 4, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 6, 18, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 8, 0, 0, 0, 
    
    -- channel=276
    0, 7, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 
    0, 3, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 15, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 
    5, 0, 0, 2, 4, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 1, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 14, 
    5, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 
    
    -- channel=277
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=278
    0, 13, 6, 5, 16, 8, 9, 9, 11, 3, 4, 0, 9, 5, 1, 
    0, 13, 6, 1, 21, 15, 2, 10, 0, 7, 3, 0, 0, 2, 0, 
    11, 0, 0, 11, 19, 1, 8, 20, 0, 22, 0, 0, 0, 0, 0, 
    5, 0, 11, 4, 15, 4, 17, 16, 8, 0, 0, 7, 0, 0, 0, 
    14, 0, 0, 21, 0, 0, 10, 2, 0, 4, 4, 5, 0, 0, 4, 
    17, 0, 0, 0, 5, 5, 1, 0, 1, 2, 0, 4, 0, 0, 8, 
    6, 0, 0, 0, 5, 0, 0, 3, 0, 0, 0, 0, 0, 0, 1, 
    5, 0, 0, 0, 0, 21, 0, 0, 0, 0, 3, 0, 0, 0, 17, 
    0, 1, 5, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 10, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 6, 9, 0, 0, 3, 0, 0, 0, 0, 0, 8, 6, 
    3, 31, 0, 0, 1, 9, 7, 0, 8, 0, 0, 2, 7, 1, 0, 
    10, 5, 27, 0, 0, 0, 0, 2, 17, 0, 0, 0, 0, 0, 0, 
    
    -- channel=279
    33, 17, 16, 23, 53, 0, 27, 0, 30, 19, 56, 0, 105, 0, 13, 
    31, 19, 36, 28, 43, 0, 18, 0, 39, 16, 58, 0, 103, 0, 49, 
    38, 20, 26, 27, 28, 0, 16, 35, 14, 44, 23, 0, 95, 37, 56, 
    48, 0, 43, 33, 0, 18, 56, 30, 0, 33, 21, 6, 83, 46, 100, 
    38, 4, 85, 31, 0, 37, 72, 0, 41, 23, 51, 6, 63, 51, 115, 
    41, 0, 55, 65, 25, 24, 25, 22, 45, 36, 49, 0, 71, 48, 111, 
    41, 11, 22, 60, 41, 21, 23, 28, 29, 21, 18, 23, 55, 38, 89, 
    40, 16, 26, 56, 46, 17, 16, 28, 32, 27, 26, 20, 63, 44, 74, 
    24, 31, 38, 42, 17, 52, 15, 32, 36, 35, 38, 26, 53, 36, 57, 
    39, 42, 41, 27, 44, 11, 28, 36, 36, 53, 31, 45, 63, 32, 6, 
    73, 14, 47, 23, 24, 39, 7, 51, 53, 49, 34, 42, 46, 21, 49, 
    22, 50, 77, 22, 59, 19, 30, 46, 42, 52, 37, 40, 44, 18, 53, 
    34, 23, 76, 67, 56, 27, 37, 54, 4, 41, 41, 46, 53, 0, 52, 
    63, 0, 12, 57, 79, 52, 47, 49, 0, 36, 37, 48, 61, 0, 26, 
    68, 28, 0, 13, 61, 72, 69, 55, 39, 27, 33, 35, 38, 32, 7, 
    
    -- channel=280
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    5, 0, 0, 7, 0, 0, 0, 0, 0, 4, 0, 2, 0, 0, 0, 
    0, 0, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 1, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 2, 8, 3, 7, 0, 0, 0, 0, 0, 0, 0, 1, 3, 0, 
    4, 3, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 1, 0, 
    0, 12, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=281
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 5, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 18, 9, 0, 
    0, 1, 0, 3, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 27, 0, 0, 0, 0, 5, 32, 26, 0, 0, 0, 0, 0, 0, 
    0, 42, 29, 0, 0, 0, 0, 0, 0, 5, 0, 2, 8, 0, 0, 
    0, 0, 22, 19, 0, 0, 0, 0, 5, 23, 35, 0, 0, 0, 0, 
    
    -- channel=282
    24, 14, 24, 28, 7, 19, 19, 27, 30, 30, 20, 41, 11, 18, 19, 
    36, 28, 29, 31, 5, 15, 15, 24, 29, 33, 20, 45, 19, 37, 33, 
    23, 17, 25, 28, 2, 18, 31, 28, 31, 17, 22, 54, 41, 41, 38, 
    17, 33, 31, 13, 14, 40, 26, 5, 26, 15, 44, 48, 48, 48, 27, 
    22, 55, 32, 23, 30, 42, 12, 23, 42, 40, 41, 47, 49, 50, 13, 
    17, 52, 55, 26, 43, 28, 27, 48, 41, 35, 32, 46, 42, 54, 7, 
    20, 45, 58, 50, 32, 26, 22, 30, 26, 29, 32, 38, 40, 54, 18, 
    24, 43, 46, 49, 33, 28, 27, 33, 33, 32, 32, 46, 32, 45, 13, 
    40, 48, 47, 47, 51, 21, 44, 39, 36, 35, 36, 38, 36, 37, 11, 
    47, 38, 24, 33, 32, 55, 34, 43, 46, 40, 36, 34, 20, 22, 41, 
    28, 32, 27, 45, 44, 24, 54, 50, 43, 40, 33, 31, 28, 39, 56, 
    44, 60, 37, 46, 39, 48, 46, 43, 46, 37, 37, 33, 24, 41, 51, 
    45, 59, 52, 46, 35, 51, 49, 29, 38, 38, 49, 29, 19, 36, 43, 
    19, 25, 47, 54, 48, 41, 38, 27, 42, 40, 37, 30, 8, 24, 39, 
    20, 2, 36, 54, 59, 54, 48, 41, 29, 32, 34, 24, 19, 36, 61, 
    
    -- channel=283
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=284
    11, 4, 5, 15, 18, 4, 5, 4, 4, 9, 14, 3, 8, 10, 8, 
    9, 0, 12, 16, 11, 4, 17, 2, 11, 2, 14, 0, 15, 0, 7, 
    8, 12, 15, 11, 9, 4, 2, 3, 17, 9, 22, 0, 12, 8, 14, 
    20, 12, 5, 7, 2, 1, 7, 15, 3, 12, 5, 0, 20, 10, 20, 
    8, 15, 18, 4, 0, 5, 11, 0, 5, 0, 0, 4, 8, 14, 25, 
    4, 15, 21, 5, 2, 0, 0, 0, 0, 2, 8, 0, 3, 21, 18, 
    5, 9, 13, 13, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 17, 
    10, 13, 6, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 14, 
    9, 2, 9, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    6, 9, 11, 12, 14, 7, 0, 0, 0, 0, 0, 0, 0, 11, 12, 
    15, 12, 5, 16, 0, 2, 2, 0, 0, 0, 0, 0, 0, 6, 9, 
    10, 0, 0, 0, 20, 5, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    4, 15, 4, 0, 0, 10, 0, 0, 2, 0, 0, 0, 0, 0, 16, 
    14, 0, 17, 9, 0, 0, 3, 7, 0, 0, 0, 0, 0, 6, 19, 
    12, 4, 0, 6, 7, 0, 2, 5, 0, 0, 0, 3, 1, 11, 0, 
    
    -- channel=285
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=286
    1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 11, 0, 
    
    -- channel=287
    11, 11, 0, 3, 27, 0, 7, 0, 7, 4, 33, 0, 74, 0, 5, 
    20, 23, 13, 7, 31, 0, 0, 0, 16, 3, 32, 0, 77, 0, 29, 
    24, 12, 13, 13, 25, 0, 0, 16, 0, 25, 0, 0, 70, 25, 36, 
    20, 0, 27, 25, 0, 0, 27, 15, 0, 35, 0, 4, 54, 36, 62, 
    29, 0, 69, 15, 0, 18, 48, 0, 12, 11, 29, 2, 45, 39, 81, 
    41, 0, 41, 69, 0, 22, 38, 17, 39, 25, 30, 3, 59, 31, 85, 
    42, 0, 10, 55, 42, 24, 33, 22, 30, 26, 31, 27, 44, 27, 77, 
    35, 0, 25, 43, 44, 32, 14, 34, 42, 35, 37, 25, 71, 31, 61, 
    18, 22, 30, 29, 15, 78, 20, 40, 42, 38, 44, 39, 55, 35, 56, 
    33, 34, 34, 9, 26, 0, 53, 46, 47, 58, 44, 48, 53, 17, 0, 
    56, 0, 39, 0, 19, 45, 0, 61, 61, 52, 43, 43, 46, 21, 28, 
    29, 36, 69, 11, 39, 9, 28, 48, 52, 64, 38, 44, 46, 16, 36, 
    20, 10, 70, 60, 48, 12, 35, 50, 11, 52, 40, 56, 44, 0, 30, 
    34, 0, 0, 47, 69, 39, 28, 40, 5, 35, 47, 57, 52, 0, 12, 
    42, 11, 0, 0, 53, 67, 51, 31, 33, 22, 29, 36, 39, 1, 0, 
    
    -- channel=288
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=289
    0, 9, 0, 0, 31, 0, 0, 0, 0, 0, 15, 0, 50, 0, 0, 
    0, 0, 0, 0, 32, 0, 0, 0, 0, 0, 15, 0, 53, 0, 0, 
    0, 0, 0, 0, 29, 0, 0, 0, 0, 15, 0, 0, 19, 0, 0, 
    20, 0, 1, 13, 0, 0, 0, 33, 0, 23, 0, 0, 7, 0, 27, 
    10, 0, 30, 0, 0, 0, 45, 0, 0, 0, 0, 0, 0, 0, 60, 
    20, 0, 0, 38, 0, 0, 0, 0, 0, 0, 5, 0, 4, 0, 68, 
    19, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 5, 0, 51, 
    9, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 12, 0, 52, 
    0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 31, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 1, 0, 
    24, 0, 9, 0, 0, 4, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    0, 0, 23, 0, 5, 0, 0, 0, 0, 2, 0, 0, 2, 0, 0, 
    0, 0, 0, 2, 8, 0, 0, 0, 0, 0, 0, 7, 10, 0, 0, 
    15, 0, 0, 0, 6, 0, 0, 18, 0, 0, 0, 2, 35, 0, 0, 
    18, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 23, 0, 0, 
    
    -- channel=290
    0, 0, 0, 0, 4, 0, 0, 0, 0, 14, 0, 0, 0, 5, 0, 
    0, 0, 0, 0, 8, 0, 12, 0, 0, 0, 1, 0, 0, 0, 0, 
    6, 22, 0, 2, 14, 0, 0, 0, 17, 6, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 40, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 22, 0, 0, 10, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 2, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 6, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 
    0, 0, 10, 12, 0, 0, 0, 0, 0, 0, 0, 0, 11, 18, 3, 
    0, 20, 5, 0, 10, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    13, 37, 0, 0, 0, 0, 0, 14, 28, 0, 0, 0, 0, 16, 0, 
    0, 22, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 13, 
    0, 0, 0, 23, 0, 0, 0, 0, 0, 6, 18, 22, 0, 0, 0, 
    
    -- channel=291
    0, 0, 0, 0, 5, 0, 0, 0, 0, 8, 0, 0, 0, 5, 0, 
    0, 0, 0, 0, 8, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 7, 0, 8, 10, 0, 0, 0, 1, 24, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 34, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 8, 0, 0, 8, 0, 0, 0, 0, 13, 0, 0, 15, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 5, 0, 0, 0, 0, 0, 5, 0, 0, 0, 3, 0, 0, 
    3, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 36, 
    0, 0, 16, 9, 16, 0, 0, 0, 0, 5, 0, 0, 17, 15, 0, 
    0, 21, 13, 0, 2, 32, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    19, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    31, 24, 0, 0, 0, 0, 0, 32, 24, 0, 0, 0, 0, 23, 0, 
    0, 51, 23, 0, 0, 0, 1, 0, 0, 0, 0, 9, 33, 0, 0, 
    0, 0, 23, 12, 0, 0, 0, 0, 19, 7, 24, 10, 0, 0, 0, 
    
    -- channel=292
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=293
    14, 24, 23, 6, 1, 8, 6, 2, 0, 0, 0, 5, 2, 0, 9, 
    15, 32, 5, 5, 5, 0, 0, 10, 5, 11, 0, 10, 17, 43, 18, 
    0, 0, 0, 0, 3, 26, 42, 6, 0, 0, 0, 19, 9, 16, 6, 
    1, 27, 19, 6, 23, 29, 0, 0, 3, 19, 27, 18, 0, 9, 0, 
    13, 0, 27, 3, 16, 13, 5, 35, 24, 29, 1, 0, 0, 0, 0, 
    0, 0, 0, 58, 32, 2, 6, 28, 20, 2, 0, 26, 0, 0, 4, 
    29, 5, 0, 6, 0, 0, 21, 12, 0, 0, 12, 20, 0, 5, 5, 
    0, 0, 11, 0, 25, 11, 0, 1, 19, 38, 18, 0, 27, 0, 0, 
    18, 21, 0, 0, 0, 28, 9, 1, 14, 0, 0, 5, 0, 0, 13, 
    4, 0, 0, 0, 0, 0, 6, 18, 0, 3, 2, 0, 0, 9, 3, 
    0, 0, 11, 3, 12, 17, 0, 2, 4, 0, 0, 0, 3, 9, 21, 
    42, 79, 54, 19, 0, 0, 0, 0, 0, 2, 9, 0, 0, 0, 0, 
    0, 0, 11, 35, 17, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 33, 22, 0, 15, 31, 0, 0, 0, 0, 0, 1, 
    0, 16, 0, 0, 0, 41, 30, 11, 0, 0, 0, 0, 42, 38, 27, 
    
    -- channel=294
    20, 25, 27, 28, 27, 31, 28, 28, 32, 31, 29, 30, 24, 29, 28, 
    19, 31, 24, 26, 29, 31, 26, 34, 25, 30, 25, 31, 14, 25, 23, 
    34, 31, 26, 25, 29, 28, 30, 33, 24, 34, 25, 28, 15, 27, 25, 
    25, 24, 26, 26, 29, 33, 41, 30, 36, 21, 25, 39, 16, 22, 20, 
    29, 21, 20, 27, 30, 27, 26, 33, 23, 34, 32, 34, 21, 21, 17, 
    27, 23, 16, 23, 31, 28, 15, 17, 28, 29, 23, 38, 24, 19, 20, 
    25, 23, 22, 24, 23, 19, 16, 21, 20, 17, 14, 22, 18, 27, 17, 
    29, 24, 29, 22, 10, 21, 18, 15, 9, 13, 19, 7, 17, 22, 27, 
    22, 25, 24, 22, 22, 13, 12, 8, 15, 15, 12, 17, 11, 16, 28, 
    26, 25, 33, 32, 23, 13, 11, 10, 8, 9, 14, 14, 12, 25, 22, 
    24, 28, 27, 18, 31, 29, 12, 7, 9, 10, 13, 12, 15, 16, 25, 
    17, 17, 27, 33, 23, 23, 17, 10, 7, 11, 10, 14, 19, 24, 28, 
    35, 21, 23, 34, 33, 23, 18, 17, 12, 8, 5, 11, 20, 26, 39, 
    29, 45, 31, 24, 31, 37, 34, 18, 27, 12, 12, 16, 18, 39, 24, 
    27, 31, 42, 32, 21, 29, 37, 34, 34, 17, 16, 13, 22, 20, 36, 
    
    -- channel=295
    4, 0, 3, 2, 0, 4, 5, 6, 15, 14, 7, 11, 10, 10, 3, 
    7, 5, 7, 2, 0, 7, 4, 7, 8, 10, 7, 13, 10, 6, 7, 
    6, 7, 2, 3, 0, 5, 7, 9, 7, 6, 9, 14, 16, 11, 9, 
    3, 7, 6, 0, 0, 16, 16, 6, 7, 0, 18, 16, 18, 10, 7, 
    3, 13, 3, 8, 8, 18, 10, 4, 16, 14, 24, 23, 17, 10, 2, 
    1, 14, 10, 1, 17, 14, 6, 12, 16, 19, 17, 15, 19, 10, 0, 
    0, 12, 14, 9, 17, 17, 13, 17, 15, 13, 13, 20, 15, 12, 3, 
    6, 9, 10, 12, 12, 17, 21, 18, 17, 17, 16, 13, 14, 11, 4, 
    7, 12, 11, 13, 20, 4, 17, 16, 20, 21, 19, 16, 18, 14, 0, 
    9, 13, 5, 10, 8, 20, 13, 14, 18, 18, 18, 17, 10, 5, 12, 
    7, 8, 7, 11, 15, 4, 19, 18, 13, 17, 15, 16, 14, 7, 10, 
    7, 18, 14, 14, 8, 15, 18, 20, 15, 13, 18, 18, 19, 11, 16, 
    20, 28, 27, 22, 13, 12, 20, 21, 16, 13, 18, 17, 15, 18, 14, 
    9, 22, 30, 28, 27, 19, 20, 13, 15, 19, 14, 18, 12, 10, 15, 
    9, 3, 30, 31, 29, 28, 26, 23, 13, 17, 18, 15, 8, 14, 22, 
    
    -- channel=296
    34, 22, 25, 35, 39, 4, 30, 18, 34, 32, 49, 12, 65, 11, 27, 
    35, 29, 39, 37, 33, 6, 24, 15, 41, 30, 48, 7, 71, 19, 45, 
    36, 33, 37, 31, 27, 11, 30, 37, 31, 35, 36, 9, 72, 45, 55, 
    42, 24, 38, 33, 11, 33, 53, 31, 15, 38, 27, 32, 69, 50, 67, 
    39, 29, 70, 26, 17, 43, 50, 13, 42, 37, 53, 31, 58, 54, 72, 
    35, 24, 61, 58, 35, 26, 25, 30, 46, 39, 42, 24, 62, 54, 69, 
    40, 26, 39, 59, 30, 14, 21, 20, 25, 17, 19, 24, 49, 49, 65, 
    42, 33, 42, 55, 38, 11, 18, 23, 23, 21, 21, 23, 46, 48, 51, 
    37, 40, 42, 47, 22, 47, 11, 24, 25, 28, 29, 22, 36, 34, 51, 
    45, 43, 43, 39, 44, 15, 29, 30, 29, 36, 27, 31, 40, 36, 31, 
    55, 32, 45, 34, 36, 44, 19, 38, 39, 33, 26, 30, 33, 32, 53, 
    42, 47, 63, 38, 55, 30, 29, 33, 34, 37, 27, 26, 31, 31, 63, 
    37, 42, 72, 63, 55, 40, 30, 30, 16, 33, 26, 30, 32, 19, 60, 
    49, 8, 38, 65, 69, 54, 48, 51, 14, 26, 32, 29, 35, 29, 47, 
    51, 30, 0, 37, 67, 70, 68, 55, 35, 22, 22, 34, 40, 36, 28, 
    
    -- channel=297
    2, 15, 0, 1, 19, 0, 6, 3, 4, 6, 16, 0, 27, 0, 9, 
    4, 14, 7, 0, 26, 0, 6, 3, 6, 3, 13, 0, 24, 0, 2, 
    9, 7, 6, 5, 25, 0, 2, 8, 0, 17, 0, 0, 8, 2, 5, 
    13, 0, 10, 11, 15, 0, 16, 28, 0, 18, 0, 0, 5, 1, 10, 
    15, 0, 9, 18, 0, 5, 24, 1, 0, 2, 9, 10, 7, 0, 27, 
    23, 0, 0, 22, 0, 10, 18, 0, 5, 8, 13, 0, 14, 0, 32, 
    18, 0, 0, 6, 16, 9, 12, 6, 13, 6, 5, 4, 10, 0, 33, 
    14, 0, 0, 1, 0, 25, 1, 11, 7, 8, 12, 0, 11, 0, 34, 
    2, 0, 6, 3, 5, 7, 1, 5, 3, 8, 14, 4, 18, 9, 19, 
    1, 10, 15, 0, 0, 4, 4, 0, 8, 1, 10, 9, 11, 5, 1, 
    16, 0, 16, 0, 9, 5, 0, 2, 0, 12, 6, 10, 13, 4, 0, 
    7, 0, 20, 4, 5, 2, 0, 2, 4, 12, 0, 9, 20, 0, 7, 
    1, 0, 12, 18, 18, 0, 3, 16, 2, 4, 1, 16, 13, 10, 7, 
    11, 8, 0, 9, 19, 14, 13, 17, 1, 0, 2, 18, 25, 0, 3, 
    19, 10, 0, 0, 9, 13, 15, 12, 20, 6, 4, 15, 22, 0, 0, 
    
    -- channel=298
    18, 0, 2, 1, 0, 0, 9, 0, 23, 23, 26, 9, 45, 5, 10, 
    19, 1, 12, 9, 0, 0, 7, 0, 21, 10, 25, 14, 54, 4, 24, 
    30, 22, 17, 8, 0, 0, 0, 10, 14, 10, 28, 17, 73, 28, 44, 
    6, 12, 20, 12, 0, 12, 26, 0, 11, 8, 25, 30, 80, 46, 56, 
    4, 38, 41, 9, 10, 30, 23, 0, 21, 23, 43, 30, 67, 54, 41, 
    8, 39, 56, 13, 22, 47, 42, 40, 41, 46, 47, 29, 64, 51, 34, 
    7, 25, 42, 57, 54, 59, 54, 57, 62, 62, 57, 57, 61, 44, 32, 
    20, 29, 36, 63, 70, 36, 67, 75, 68, 62, 64, 79, 70, 57, 17, 
    24, 31, 38, 44, 64, 73, 62, 77, 78, 86, 80, 72, 85, 46, 18, 
    39, 37, 25, 39, 45, 63, 75, 82, 86, 92, 73, 79, 63, 26, 20, 
    37, 32, 22, 25, 24, 35, 76, 95, 93, 86, 79, 78, 62, 30, 38, 
    32, 55, 39, 24, 40, 40, 75, 102, 92, 77, 83, 80, 62, 46, 35, 
    56, 87, 79, 50, 38, 47, 69, 83, 74, 86, 87, 75, 64, 18, 34, 
    30, 18, 77, 80, 57, 38, 48, 43, 30, 86, 86, 76, 45, 18, 25, 
    28, 0, 9, 75, 87, 60, 48, 48, 51, 73, 74, 58, 18, 12, 42, 
    
    -- channel=299
    0, 0, 2, 0, 0, 30, 0, 9, 0, 2, 0, 39, 0, 21, 0, 
    0, 0, 0, 0, 0, 22, 0, 14, 0, 0, 0, 50, 0, 12, 0, 
    0, 0, 0, 0, 0, 17, 0, 0, 7, 0, 2, 45, 0, 0, 0, 
    0, 22, 0, 0, 0, 11, 0, 0, 25, 0, 9, 21, 0, 0, 0, 
    0, 36, 0, 0, 25, 0, 0, 19, 0, 0, 0, 14, 0, 0, 0, 
    0, 41, 0, 0, 6, 0, 0, 9, 0, 0, 0, 27, 0, 0, 0, 
    0, 19, 12, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 12, 1, 0, 0, 0, 13, 0, 0, 0, 0, 15, 0, 0, 0, 
    0, 0, 0, 0, 11, 0, 8, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 4, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 13, 0, 3, 0, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 13, 0, 
    5, 28, 0, 0, 0, 6, 0, 0, 30, 0, 0, 0, 0, 22, 0, 
    0, 30, 40, 0, 0, 0, 0, 0, 15, 3, 0, 0, 0, 25, 0, 
    0, 0, 46, 35, 0, 0, 0, 0, 0, 4, 5, 0, 0, 0, 34, 
    
    -- channel=300
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    
    -- channel=301
    7, 14, 0, 0, 38, 0, 1, 0, 0, 0, 24, 0, 65, 0, 0, 
    1, 2, 3, 0, 40, 0, 1, 0, 8, 0, 25, 0, 72, 0, 8, 
    0, 4, 1, 0, 36, 0, 0, 0, 0, 12, 0, 0, 36, 0, 8, 
    26, 0, 3, 21, 0, 0, 4, 32, 0, 41, 0, 0, 20, 0, 40, 
    18, 0, 50, 2, 0, 0, 50, 0, 0, 0, 0, 0, 1, 0, 77, 
    29, 0, 1, 58, 0, 0, 14, 0, 4, 0, 12, 0, 11, 0, 85, 
    32, 0, 0, 12, 12, 0, 13, 0, 1, 0, 5, 0, 10, 0, 72, 
    17, 0, 0, 0, 23, 0, 0, 0, 15, 4, 0, 0, 30, 0, 56, 
    0, 0, 0, 0, 0, 51, 0, 4, 0, 0, 5, 0, 10, 2, 51, 
    0, 2, 9, 0, 4, 0, 9, 0, 0, 9, 4, 6, 36, 5, 0, 
    35, 0, 19, 0, 0, 19, 0, 0, 10, 4, 3, 9, 14, 0, 0, 
    7, 0, 34, 0, 17, 0, 0, 0, 0, 20, 0, 3, 17, 0, 0, 
    0, 0, 30, 14, 11, 0, 0, 4, 0, 10, 0, 22, 22, 0, 0, 
    26, 0, 0, 10, 23, 0, 0, 27, 0, 0, 4, 11, 43, 0, 6, 
    32, 21, 0, 0, 10, 21, 12, 0, 0, 0, 0, 21, 31, 0, 0, 
    
    -- channel=302
    20, 15, 26, 8, 4, 5, 15, 0, 0, 0, 4, 0, 23, 0, 9, 
    15, 19, 10, 10, 2, 0, 0, 1, 15, 8, 8, 0, 41, 36, 22, 
    0, 0, 4, 0, 0, 21, 35, 9, 0, 0, 3, 4, 34, 16, 21, 
    4, 27, 13, 8, 10, 29, 1, 0, 0, 20, 29, 7, 9, 16, 4, 
    10, 10, 37, 0, 17, 19, 12, 27, 30, 28, 10, 0, 11, 8, 2, 
    0, 0, 11, 48, 27, 2, 21, 41, 27, 7, 7, 20, 7, 0, 21, 
    23, 8, 0, 13, 8, 8, 23, 9, 0, 6, 18, 14, 7, 10, 21, 
    0, 1, 6, 0, 41, 0, 0, 13, 30, 34, 11, 7, 29, 5, 0, 
    20, 20, 0, 0, 0, 45, 9, 11, 14, 0, 4, 7, 0, 0, 21, 
    7, 0, 0, 0, 0, 0, 18, 24, 6, 17, 3, 8, 12, 6, 8, 
    0, 7, 16, 12, 4, 17, 0, 13, 15, 0, 0, 6, 13, 15, 25, 
    39, 80, 52, 12, 8, 0, 8, 2, 1, 9, 20, 7, 1, 7, 0, 
    0, 0, 29, 39, 17, 7, 0, 0, 0, 14, 5, 8, 9, 0, 0, 
    3, 0, 0, 20, 42, 21, 0, 25, 11, 0, 9, 0, 0, 0, 10, 
    7, 21, 0, 0, 17, 48, 33, 13, 0, 0, 0, 0, 33, 29, 19, 
    
    -- channel=303
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 2, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 15, 13, 
    0, 1, 17, 0, 0, 1, 0, 0, 0, 0, 4, 0, 22, 18, 5, 
    0, 0, 21, 6, 0, 10, 8, 11, 13, 11, 10, 5, 18, 16, 3, 
    0, 0, 8, 24, 16, 14, 15, 13, 16, 17, 20, 21, 18, 12, 5, 
    0, 0, 9, 21, 33, 2, 19, 26, 26, 24, 21, 30, 33, 16, 0, 
    2, 5, 5, 9, 14, 40, 20, 30, 32, 33, 29, 25, 28, 4, 0, 
    8, 4, 0, 1, 9, 7, 33, 39, 36, 41, 29, 29, 19, 0, 0, 
    6, 0, 0, 0, 0, 11, 24, 45, 45, 33, 30, 28, 17, 2, 10, 
    14, 31, 13, 0, 9, 5, 30, 44, 39, 34, 35, 29, 14, 7, 5, 
    9, 24, 38, 18, 4, 8, 22, 21, 17, 38, 35, 29, 16, 0, 0, 
    0, 0, 13, 34, 24, 4, 4, 6, 1, 32, 37, 25, 0, 0, 2, 
    0, 0, 0, 14, 38, 30, 17, 10, 5, 15, 16, 13, 0, 0, 5, 
    
    -- channel=304
    18, 2, 11, 21, 8, 7, 18, 22, 40, 45, 34, 36, 31, 26, 20, 
    29, 17, 27, 25, 5, 13, 23, 20, 29, 30, 30, 40, 31, 11, 29, 
    45, 41, 29, 27, 4, 1, 13, 29, 38, 30, 34, 43, 52, 41, 42, 
    20, 21, 27, 19, 1, 30, 48, 25, 27, 15, 27, 56, 71, 50, 46, 
    20, 48, 34, 21, 23, 46, 26, 7, 31, 35, 54, 66, 64, 56, 33, 
    22, 54, 59, 15, 37, 47, 25, 34, 45, 52, 48, 43, 64, 60, 22, 
    15, 38, 63, 60, 47, 43, 34, 44, 49, 44, 38, 49, 57, 55, 27, 
    34, 43, 51, 63, 43, 35, 52, 49, 40, 36, 44, 57, 47, 55, 34, 
    32, 42, 56, 60, 71, 36, 46, 52, 53, 65, 56, 55, 63, 53, 20, 
    48, 55, 43, 50, 50, 71, 50, 53, 62, 58, 55, 54, 39, 28, 35, 
    46, 39, 29, 36, 43, 39, 64, 67, 61, 64, 56, 54, 41, 32, 45, 
    33, 33, 34, 44, 50, 50, 63, 72, 66, 53, 51, 52, 51, 44, 62, 
    75, 101, 75, 53, 47, 54, 65, 67, 73, 56, 60, 50, 39, 45, 60, 
    34, 60, 98, 80, 56, 53, 60, 38, 39, 64, 60, 53, 38, 37, 46, 
    31, 6, 50, 94, 84, 62, 57, 63, 56, 60, 66, 51, 16, 22, 59, 
    
    -- channel=305
    38, 32, 35, 27, 12, 14, 27, 22, 23, 17, 26, 31, 42, 2, 31, 
    48, 47, 35, 29, 14, 0, 4, 25, 41, 35, 29, 34, 72, 58, 46, 
    2, 1, 25, 18, 8, 35, 57, 28, 16, 6, 25, 47, 75, 52, 55, 
    24, 49, 43, 20, 28, 53, 29, 0, 21, 38, 58, 49, 57, 58, 29, 
    31, 43, 65, 27, 38, 55, 34, 47, 62, 63, 51, 34, 59, 52, 26, 
    19, 23, 61, 79, 56, 37, 50, 64, 60, 42, 44, 53, 55, 45, 38, 
    45, 38, 39, 61, 47, 41, 54, 45, 33, 38, 53, 57, 49, 55, 51, 
    28, 36, 48, 48, 70, 40, 38, 56, 66, 75, 55, 50, 67, 41, 14, 
    55, 58, 31, 35, 34, 66, 54, 57, 57, 46, 55, 47, 35, 22, 36, 
    45, 22, 17, 20, 25, 24, 57, 65, 64, 60, 51, 50, 38, 30, 52, 
    24, 32, 44, 48, 52, 39, 53, 67, 59, 48, 42, 48, 48, 52, 59, 
    88, 119, 92, 51, 42, 50, 50, 52, 54, 57, 60, 50, 42, 35, 49, 
    4, 19, 87, 87, 57, 44, 48, 13, 9, 58, 57, 53, 36, 18, 35, 
    23, 0, 1, 79, 95, 64, 47, 62, 57, 41, 50, 42, 5, 13, 52, 
    30, 23, 0, 20, 80, 104, 84, 61, 27, 21, 7, 30, 66, 66, 67, 
    
    -- channel=306
    6, 0, 9, 2, 4, 1, 12, 6, 11, 0, 2, 0, 10, 0, 0, 
    0, 6, 7, 4, 5, 6, 0, 0, 12, 12, 3, 0, 0, 15, 13, 
    8, 0, 0, 3, 0, 0, 7, 19, 0, 2, 0, 3, 9, 3, 10, 
    0, 0, 6, 0, 0, 16, 11, 0, 0, 0, 3, 2, 6, 9, 12, 
    8, 6, 9, 9, 13, 14, 0, 0, 17, 10, 17, 3, 0, 5, 2, 
    5, 4, 4, 1, 3, 0, 9, 34, 12, 1, 0, 6, 5, 4, 7, 
    6, 3, 0, 13, 14, 8, 0, 0, 0, 9, 11, 0, 0, 5, 7, 
    0, 0, 1, 5, 18, 0, 0, 7, 14, 0, 0, 10, 9, 0, 0, 
    2, 8, 4, 0, 8, 13, 13, 10, 1, 0, 0, 7, 1, 13, 0, 
    15, 0, 0, 2, 3, 8, 9, 9, 4, 9, 0, 3, 0, 0, 0, 
    0, 0, 1, 4, 1, 3, 0, 7, 7, 2, 0, 0, 0, 0, 25, 
    0, 27, 4, 0, 9, 0, 13, 1, 0, 5, 3, 9, 6, 8, 0, 
    8, 0, 14, 8, 0, 17, 21, 16, 0, 2, 12, 0, 11, 0, 10, 
    4, 0, 0, 7, 6, 1, 0, 0, 5, 8, 3, 5, 0, 3, 0, 
    14, 2, 3, 1, 15, 9, 7, 0, 1, 12, 22, 0, 0, 0, 10, 
    
    -- channel=307
    15, 21, 16, 10, 28, 1, 15, 5, 9, 2, 18, 0, 40, 2, 9, 
    11, 18, 15, 8, 27, 6, 9, 2, 14, 8, 21, 0, 37, 9, 19, 
    4, 2, 6, 7, 24, 12, 21, 16, 0, 20, 2, 0, 20, 10, 6, 
    24, 6, 16, 16, 14, 16, 19, 20, 0, 21, 13, 2, 6, 3, 21, 
    19, 0, 28, 14, 0, 9, 34, 5, 21, 13, 13, 0, 6, 0, 34, 
    17, 0, 0, 36, 17, 3, 0, 1, 12, 6, 11, 0, 12, 0, 41, 
    24, 0, 0, 1, 3, 2, 11, 7, 0, 0, 0, 0, 7, 0, 29, 
    13, 0, 0, 0, 11, 11, 0, 0, 7, 11, 3, 0, 13, 0, 30, 
    4, 4, 0, 0, 0, 7, 0, 0, 3, 0, 0, 0, 0, 0, 26, 
    0, 2, 12, 0, 9, 0, 0, 0, 0, 0, 0, 2, 19, 12, 0, 
    18, 0, 17, 1, 1, 14, 0, 0, 0, 0, 0, 3, 11, 0, 10, 
    1, 19, 40, 8, 12, 0, 0, 0, 0, 1, 0, 1, 9, 0, 6, 
    0, 0, 12, 26, 22, 0, 0, 0, 0, 0, 0, 5, 14, 0, 6, 
    22, 0, 0, 2, 28, 25, 15, 21, 0, 0, 0, 3, 22, 0, 4, 
    23, 28, 0, 0, 0, 21, 27, 20, 5, 0, 0, 3, 27, 22, 0, 
    
    -- channel=308
    4, 1, 1, 0, 16, 0, 3, 0, 0, 0, 9, 0, 33, 0, 0, 
    0, 0, 4, 0, 12, 0, 0, 0, 1, 0, 11, 0, 32, 0, 6, 
    0, 0, 0, 0, 6, 0, 1, 3, 0, 0, 0, 0, 16, 0, 6, 
    8, 0, 3, 7, 0, 0, 5, 1, 0, 8, 0, 0, 7, 0, 22, 
    5, 0, 20, 0, 0, 0, 18, 0, 1, 0, 0, 0, 3, 0, 34, 
    5, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 39, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 12, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    8, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 17, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 7, 0, 0, 8, 0, 0, 0, 0, 4, 0, 0, 
    14, 8, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 6, 4, 0, 
    
    -- channel=309
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 12, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 9, 0, 3, 10, 2, 0, 0, 
    0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 2, 5, 0, 
    0, 22, 7, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 
    0, 10, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 
    0, 10, 9, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 
    0, 1, 7, 11, 12, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 6, 0, 6, 1, 16, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 1, 0, 3, 4, 0, 17, 1, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 6, 0, 10, 3, 3, 4, 0, 0, 0, 0, 0, 11, 
    19, 30, 0, 0, 0, 1, 0, 0, 13, 0, 0, 0, 0, 10, 3, 
    0, 18, 35, 0, 0, 0, 6, 0, 0, 1, 0, 0, 0, 1, 9, 
    0, 0, 17, 26, 0, 0, 0, 4, 0, 0, 0, 0, 0, 1, 17, 
    
    -- channel=310
    9, 17, 0, 0, 51, 0, 6, 0, 0, 0, 31, 0, 93, 0, 0, 
    5, 9, 15, 0, 50, 0, 0, 0, 11, 0, 35, 0, 86, 0, 19, 
    3, 0, 0, 7, 35, 0, 0, 11, 0, 33, 0, 0, 51, 0, 13, 
    36, 0, 21, 15, 0, 0, 22, 30, 0, 21, 0, 0, 24, 0, 66, 
    25, 0, 53, 21, 0, 0, 69, 0, 9, 0, 6, 0, 13, 0, 103, 
    38, 0, 0, 56, 0, 0, 9, 0, 11, 0, 21, 0, 26, 0, 108, 
    32, 0, 0, 8, 11, 0, 0, 0, 0, 0, 0, 0, 19, 0, 80, 
    17, 0, 0, 0, 0, 15, 0, 0, 1, 0, 0, 0, 28, 0, 73, 
    0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 15, 5, 41, 
    0, 6, 11, 0, 0, 0, 0, 0, 0, 6, 0, 5, 39, 6, 0, 
    47, 0, 27, 0, 0, 0, 0, 0, 1, 7, 0, 3, 18, 0, 0, 
    0, 1, 54, 0, 18, 0, 0, 0, 0, 14, 0, 2, 18, 0, 6, 
    0, 0, 19, 30, 20, 0, 0, 17, 0, 0, 0, 17, 27, 0, 1, 
    37, 0, 0, 0, 43, 12, 0, 18, 0, 0, 0, 17, 55, 0, 0, 
    49, 16, 0, 0, 0, 28, 29, 8, 2, 0, 0, 5, 29, 12, 0, 
    
    -- channel=311
    19, 21, 16, 23, 33, 9, 24, 17, 25, 25, 38, 6, 49, 9, 23, 
    16, 25, 25, 21, 34, 8, 21, 16, 27, 21, 35, 0, 45, 7, 25, 
    29, 30, 26, 20, 32, 11, 23, 30, 18, 28, 25, 0, 36, 24, 31, 
    30, 6, 23, 26, 20, 18, 45, 35, 14, 31, 6, 21, 37, 22, 36, 
    30, 1, 37, 22, 16, 22, 35, 17, 21, 28, 39, 21, 32, 24, 48, 
    32, 2, 28, 37, 13, 17, 22, 4, 24, 19, 23, 16, 39, 24, 51, 
    31, 5, 13, 28, 17, 9, 14, 5, 16, 9, 6, 4, 25, 23, 49, 
    32, 14, 19, 26, 10, 8, 4, 12, 6, 4, 10, 1, 19, 23, 42, 
    19, 16, 23, 24, 9, 25, 0, 4, 4, 8, 15, 6, 24, 22, 43, 
    23, 28, 34, 24, 21, 1, 11, 1, 5, 8, 10, 13, 22, 21, 17, 
    34, 19, 35, 12, 23, 26, 0, 7, 8, 11, 9, 12, 21, 19, 20, 
    19, 6, 41, 26, 30, 12, 2, 8, 8, 14, 3, 10, 24, 20, 38, 
    24, 24, 39, 44, 43, 21, 11, 21, 6, 9, 0, 14, 19, 20, 41, 
    33, 17, 25, 37, 44, 42, 39, 39, 2, 4, 10, 19, 33, 29, 27, 
    42, 31, 5, 25, 38, 37, 43, 36, 30, 16, 12, 25, 31, 12, 3, 
    
    -- channel=312
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 7, 0, 
    0, 0, 0, 0, 0, 4, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 21, 0, 0, 0, 0, 0, 0, 10, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 8, 9, 11, 0, 0, 0, 0, 0, 0, 0, 18, 17, 0, 
    0, 14, 3, 6, 3, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 49, 0, 0, 0, 0, 0, 26, 36, 0, 0, 0, 0, 14, 1, 
    0, 47, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 
    0, 0, 23, 37, 0, 0, 0, 0, 4, 18, 33, 11, 0, 0, 0, 
    
    -- channel=313
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=314
    0, 0, 0, 0, 0, 24, 0, 14, 0, 9, 0, 37, 0, 14, 3, 
    0, 0, 0, 0, 0, 11, 0, 17, 0, 0, 0, 39, 0, 2, 0, 
    0, 15, 0, 0, 0, 14, 0, 0, 9, 0, 3, 32, 0, 0, 0, 
    0, 6, 0, 0, 17, 0, 0, 0, 11, 0, 0, 13, 0, 0, 0, 
    0, 11, 0, 0, 32, 0, 0, 25, 0, 0, 0, 23, 0, 0, 0, 
    0, 15, 0, 0, 0, 0, 4, 0, 0, 0, 0, 27, 0, 0, 0, 
    0, 0, 6, 0, 0, 11, 8, 0, 2, 12, 14, 3, 0, 0, 0, 
    0, 3, 0, 0, 0, 0, 17, 7, 5, 0, 0, 19, 0, 0, 0, 
    0, 0, 0, 0, 8, 1, 7, 7, 0, 4, 5, 4, 0, 0, 0, 
    0, 0, 0, 3, 0, 12, 13, 1, 2, 0, 8, 0, 0, 0, 10, 
    0, 12, 0, 0, 0, 0, 17, 0, 0, 0, 6, 0, 0, 2, 0, 
    4, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 13, 0, 
    0, 32, 0, 0, 0, 4, 0, 0, 36, 4, 0, 0, 0, 28, 0, 
    0, 20, 40, 0, 0, 0, 0, 0, 6, 3, 8, 0, 0, 19, 5, 
    0, 0, 25, 32, 0, 0, 0, 0, 0, 10, 10, 13, 0, 0, 6, 
    
    -- channel=315
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 
    3, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 17, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 2, 10, 4, 4, 14, 9, 2, 0, 0, 0, 4, 
    0, 0, 0, 0, 4, 0, 13, 10, 4, 1, 7, 1, 4, 0, 7, 
    0, 0, 0, 0, 1, 13, 0, 7, 8, 17, 10, 3, 22, 0, 0, 
    0, 0, 0, 0, 0, 0, 9, 2, 7, 10, 8, 11, 14, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 6, 9, 14, 15, 15, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 16, 8, 10, 11, 12, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 22, 14, 12, 6, 15, 14, 0, 0, 
    3, 0, 5, 0, 0, 0, 0, 0, 0, 13, 11, 16, 21, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 17, 15, 13, 0, 0, 0, 
    
    -- channel=316
    6, 0, 1, 3, 0, 0, 1, 0, 9, 6, 5, 1, 10, 0, 0, 
    9, 0, 7, 8, 0, 0, 0, 0, 8, 4, 6, 4, 10, 4, 10, 
    10, 1, 3, 8, 0, 0, 0, 6, 6, 7, 2, 8, 24, 10, 15, 
    3, 3, 9, 0, 0, 6, 5, 0, 0, 0, 13, 6, 28, 19, 26, 
    2, 20, 16, 7, 0, 12, 4, 0, 11, 3, 11, 9, 21, 23, 16, 
    2, 20, 23, 0, 9, 6, 5, 15, 11, 11, 11, 4, 18, 23, 10, 
    0, 15, 22, 22, 14, 7, 1, 11, 10, 12, 11, 12, 19, 20, 7, 
    3, 13, 14, 25, 15, 8, 11, 14, 11, 7, 9, 25, 14, 21, 6, 
    9, 15, 19, 19, 23, 6, 20, 19, 17, 18, 17, 15, 24, 15, 0, 
    18, 14, 6, 12, 16, 30, 11, 23, 23, 25, 15, 18, 14, 7, 5, 
    15, 7, 4, 14, 8, 3, 25, 27, 27, 24, 16, 15, 10, 8, 24, 
    4, 21, 5, 7, 19, 15, 22, 26, 25, 20, 18, 19, 8, 12, 17, 
    22, 28, 20, 8, 4, 21, 23, 24, 17, 20, 30, 13, 14, 2, 15, 
    10, 6, 19, 19, 12, 4, 9, 1, 7, 24, 19, 16, 8, 0, 0, 
    8, 0, 7, 20, 24, 15, 13, 8, 12, 18, 25, 7, 0, 5, 18, 
    
    -- channel=317
    4, 19, 0, 0, 13, 0, 0, 5, 0, 0, 6, 0, 19, 0, 6, 
    7, 15, 4, 0, 20, 0, 4, 0, 3, 0, 7, 0, 25, 0, 0, 
    0, 1, 2, 3, 20, 1, 2, 0, 0, 8, 0, 0, 9, 0, 0, 
    13, 0, 7, 7, 21, 0, 0, 21, 0, 22, 0, 0, 4, 0, 1, 
    9, 0, 8, 14, 0, 1, 21, 3, 2, 0, 0, 5, 5, 0, 19, 
    19, 0, 0, 20, 0, 6, 32, 0, 6, 5, 18, 0, 5, 0, 26, 
    19, 0, 0, 0, 18, 18, 28, 14, 20, 15, 19, 10, 19, 0, 28, 
    8, 0, 0, 0, 9, 35, 8, 22, 25, 24, 20, 14, 14, 1, 25, 
    6, 0, 4, 1, 0, 13, 17, 22, 13, 17, 30, 10, 23, 13, 14, 
    0, 4, 3, 0, 0, 11, 9, 9, 21, 14, 20, 18, 23, 7, 1, 
    11, 0, 12, 0, 0, 0, 0, 12, 14, 20, 15, 23, 24, 15, 0, 
    14, 1, 24, 0, 4, 0, 0, 14, 17, 23, 9, 21, 26, 6, 0, 
    0, 0, 14, 15, 7, 0, 0, 17, 10, 18, 18, 26, 22, 16, 0, 
    5, 0, 0, 9, 17, 6, 5, 19, 0, 8, 16, 25, 31, 0, 0, 
    12, 5, 0, 0, 9, 9, 8, 1, 14, 4, 8, 23, 24, 8, 0, 
    
    -- channel=318
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 5, 12, 1, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 2, 17, 26, 20, 18, 23, 29, 26, 19, 7, 0, 0, 
    0, 0, 0, 3, 31, 17, 30, 35, 32, 25, 25, 36, 30, 0, 0, 
    0, 0, 0, 0, 16, 36, 31, 38, 38, 40, 36, 31, 37, 5, 0, 
    0, 0, 0, 0, 0, 19, 34, 40, 40, 46, 35, 36, 27, 0, 0, 
    0, 0, 0, 0, 0, 0, 24, 41, 46, 41, 38, 36, 20, 0, 0, 
    0, 1, 0, 0, 0, 0, 29, 48, 40, 37, 40, 41, 25, 0, 0, 
    5, 12, 7, 0, 0, 0, 22, 44, 30, 40, 44, 37, 31, 0, 0, 
    0, 0, 3, 4, 0, 0, 0, 0, 0, 42, 41, 37, 18, 0, 0, 
    0, 0, 0, 0, 8, 0, 0, 0, 4, 31, 38, 17, 0, 0, 0, 
    
    -- channel=319
    0, 0, 24, 5, 0, 46, 0, 14, 11, 4, 0, 52, 0, 30, 1, 
    0, 0, 0, 7, 0, 34, 0, 29, 0, 16, 0, 74, 0, 43, 0, 
    0, 0, 0, 0, 0, 35, 23, 0, 9, 0, 17, 68, 0, 6, 0, 
    0, 54, 0, 0, 0, 48, 0, 0, 57, 0, 49, 51, 0, 1, 0, 
    0, 73, 0, 0, 37, 7, 0, 39, 12, 26, 5, 17, 0, 0, 0, 
    0, 72, 0, 0, 48, 9, 0, 32, 0, 3, 0, 50, 0, 2, 0, 
    0, 49, 25, 0, 0, 3, 0, 13, 0, 4, 0, 17, 0, 18, 0, 
    0, 30, 19, 0, 0, 0, 20, 4, 0, 6, 8, 14, 0, 4, 0, 
    4, 22, 0, 0, 26, 0, 21, 0, 7, 2, 0, 14, 0, 0, 0, 
    7, 0, 0, 22, 0, 27, 0, 12, 0, 0, 0, 0, 0, 0, 23, 
    0, 27, 0, 22, 17, 0, 55, 0, 0, 0, 0, 0, 0, 0, 22, 
    3, 34, 0, 25, 0, 25, 31, 3, 0, 0, 12, 0, 0, 15, 0, 
    18, 25, 0, 0, 0, 24, 9, 0, 16, 0, 5, 0, 0, 6, 0, 
    0, 36, 46, 0, 0, 0, 4, 0, 43, 12, 0, 0, 0, 39, 1, 
    0, 0, 72, 51, 0, 0, 0, 3, 0, 6, 0, 0, 0, 12, 89, 
    
    -- channel=320
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=321
    51, 43, 43, 39, 44, 43, 44, 38, 36, 24, 22, 23, 25, 24, 26, 
    36, 41, 44, 43, 45, 48, 49, 43, 45, 29, 19, 26, 26, 27, 28, 
    36, 35, 41, 43, 43, 48, 48, 47, 50, 47, 39, 36, 26, 27, 27, 
    36, 36, 41, 42, 45, 46, 46, 43, 39, 44, 41, 38, 25, 25, 26, 
    27, 33, 41, 41, 47, 42, 32, 33, 36, 31, 36, 36, 24, 26, 24, 
    10, 35, 36, 41, 38, 38, 32, 26, 25, 25, 25, 28, 19, 25, 24, 
    16, 24, 36, 32, 35, 31, 33, 31, 31, 28, 28, 22, 18, 25, 23, 
    30, 19, 32, 33, 26, 39, 41, 31, 28, 28, 32, 23, 17, 27, 31, 
    37, 21, 31, 30, 12, 22, 33, 23, 19, 15, 18, 16, 13, 20, 28, 
    31, 21, 23, 26, 14, 17, 34, 35, 39, 21, 22, 24, 17, 20, 32, 
    33, 22, 20, 36, 6, 4, 9, 10, 22, 16, 11, 17, 20, 15, 31, 
    34, 25, 25, 41, 46, 38, 38, 25, 15, 14, 12, 6, 12, 15, 22, 
    30, 31, 25, 28, 41, 28, 27, 39, 32, 25, 22, 21, 17, 17, 14, 
    26, 23, 34, 22, 27, 29, 28, 33, 33, 34, 37, 37, 38, 33, 30, 
    33, 29, 33, 35, 35, 35, 33, 31, 31, 30, 32, 34, 35, 34, 31, 
    
    -- channel=322
    14, 23, 12, 13, 12, 11, 14, 12, 11, 13, 11, 9, 8, 10, 12, 
    12, 14, 11, 11, 12, 13, 13, 14, 12, 7, 12, 12, 14, 9, 10, 
    5, 13, 10, 10, 9, 11, 9, 9, 18, 18, 20, 12, 7, 10, 10, 
    5, 13, 10, 12, 10, 10, 7, 10, 9, 11, 5, 6, 8, 6, 7, 
    11, 10, 11, 7, 10, 8, 3, 4, 1, 6, 7, 10, 14, 11, 9, 
    12, 0, 4, 7, 6, 13, 6, 6, 14, 7, 1, 1, 14, 12, 9, 
    11, 10, 5, 6, 7, 6, 9, 9, 11, 5, 3, 6, 12, 13, 8, 
    5, 10, 5, 6, 10, 9, 9, 7, 7, 8, 6, 12, 17, 18, 5, 
    7, 10, 3, 2, 8, 0, 0, 3, 6, 1, 2, 9, 14, 11, 4, 
    0, 3, 2, 0, 18, 9, 3, 23, 0, 3, 11, 18, 17, 15, 5, 
    1, 3, 0, 6, 0, 0, 0, 0, 4, 10, 10, 19, 13, 11, 10, 
    2, 0, 7, 14, 18, 23, 17, 5, 3, 12, 15, 10, 12, 3, 15, 
    4, 1, 0, 11, 14, 12, 5, 11, 17, 17, 16, 20, 15, 6, 0, 
    0, 0, 4, 1, 8, 5, 4, 4, 10, 16, 19, 22, 19, 17, 16, 
    3, 4, 2, 7, 9, 5, 3, 7, 6, 3, 9, 8, 6, 7, 10, 
    
    -- channel=323
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 8, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=324
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=325
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 19, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    0, 13, 0, 0, 34, 5, 0, 0, 0, 0, 0, 0, 0, 19, 0, 
    0, 1, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 29, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=326
    41, 0, 8, 1, 8, 5, 13, 1, 24, 5, 1, 8, 0, 0, 23, 
    6, 12, 10, 2, 1, 6, 17, 6, 27, 17, 0, 0, 0, 10, 5, 
    21, 0, 4, 2, 2, 8, 15, 1, 13, 34, 0, 19, 0, 3, 5, 
    25, 0, 3, 0, 4, 8, 11, 14, 0, 6, 14, 29, 7, 0, 0, 
    8, 0, 2, 1, 0, 7, 9, 0, 20, 0, 6, 44, 0, 2, 0, 
    0, 9, 0, 2, 11, 0, 23, 0, 24, 0, 13, 39, 0, 3, 0, 
    0, 0, 3, 8, 0, 0, 18, 22, 0, 0, 38, 32, 0, 0, 0, 
    14, 0, 9, 0, 0, 9, 14, 0, 0, 2, 43, 33, 0, 0, 30, 
    13, 0, 1, 28, 0, 0, 29, 0, 0, 6, 44, 18, 0, 0, 62, 
    21, 0, 0, 76, 0, 0, 44, 0, 38, 24, 12, 10, 0, 0, 69, 
    18, 0, 0, 77, 0, 0, 1, 0, 40, 22, 0, 0, 0, 0, 46, 
    18, 0, 0, 27, 30, 9, 1, 24, 22, 4, 7, 0, 0, 0, 0, 
    3, 0, 2, 0, 37, 18, 0, 29, 26, 15, 13, 0, 0, 6, 0, 
    8, 0, 21, 3, 21, 0, 0, 26, 8, 16, 12, 0, 14, 0, 9, 
    0, 0, 14, 1, 14, 0, 4, 9, 9, 9, 0, 0, 11, 17, 0, 
    
    -- channel=327
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=328
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=329
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=330
    0, 0, 11, 15, 12, 13, 10, 10, 0, 0, 2, 0, 0, 5, 0, 
    13, 14, 9, 13, 18, 11, 6, 11, 0, 0, 11, 7, 7, 0, 0, 
    4, 27, 13, 21, 19, 18, 9, 20, 13, 0, 0, 0, 8, 11, 0, 
    0, 22, 19, 24, 20, 23, 19, 15, 26, 17, 1, 0, 3, 6, 7, 
    16, 20, 17, 20, 22, 23, 9, 4, 0, 34, 19, 0, 12, 10, 8, 
    50, 2, 21, 19, 21, 31, 0, 31, 9, 20, 7, 0, 14, 6, 11, 
    34, 42, 17, 12, 10, 25, 10, 0, 0, 0, 0, 0, 0, 4, 7, 
    0, 53, 13, 22, 24, 4, 1, 25, 12, 6, 0, 0, 4, 4, 0, 
    0, 35, 8, 0, 50, 31, 4, 48, 43, 40, 13, 0, 12, 31, 0, 
    0, 47, 13, 0, 89, 32, 0, 22, 0, 0, 0, 0, 12, 48, 0, 
    0, 38, 23, 0, 0, 37, 24, 54, 13, 0, 6, 9, 0, 63, 0, 
    9, 13, 23, 0, 0, 0, 0, 0, 0, 0, 0, 5, 20, 28, 35, 
    8, 15, 7, 41, 0, 2, 6, 0, 0, 0, 0, 0, 4, 0, 31, 
    10, 30, 6, 10, 6, 3, 19, 0, 0, 0, 0, 0, 0, 0, 3, 
    8, 6, 1, 5, 0, 5, 14, 15, 7, 1, 8, 11, 0, 0, 0, 
    
    -- channel=331
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 7, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 6, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=332
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=333
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=334
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 15, 0, 0, 
    0, 2, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 59, 77, 2, 52, 0, 0, 18, 0, 0, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 22, 17, 7, 40, 2, 38, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 50, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=335
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 3, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=336
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=337
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 9, 12, 0, 0, 16, 0, 0, 0, 
    0, 4, 0, 0, 0, 0, 8, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 4, 11, 2, 28, 27, 38, 52, 20, 0, 0, 0, 
    0, 0, 0, 11, 20, 0, 15, 0, 0, 14, 0, 0, 0, 0, 0, 
    0, 0, 6, 15, 0, 44, 38, 25, 41, 11, 16, 3, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 11, 7, 1, 7, 6, 9, 8, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 
    0, 3, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=338
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 1, 4, 8, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 13, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 11, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 20, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 20, 16, 12, 0, 0, 
    0, 0, 0, 0, 31, 11, 0, 0, 0, 16, 21, 12, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 32, 38, 38, 36, 17, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 27, 37, 38, 19, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=339
    16, 3, 22, 24, 23, 25, 26, 25, 22, 24, 25, 26, 23, 22, 25, 
    12, 12, 22, 20, 21, 21, 27, 28, 30, 28, 23, 25, 24, 27, 26, 
    14, 7, 18, 20, 21, 22, 25, 27, 25, 16, 12, 27, 31, 30, 26, 
    16, 7, 17, 18, 17, 26, 28, 30, 26, 24, 29, 30, 31, 30, 28, 
    16, 11, 14, 21, 16, 28, 25, 22, 26, 31, 29, 24, 23, 27, 26, 
    18, 19, 12, 17, 22, 8, 2, 13, 21, 23, 29, 32, 19, 26, 26, 
    9, 16, 9, 13, 13, 3, 9, 10, 0, 6, 21, 27, 18, 21, 26, 
    28, 13, 11, 14, 2, 0, 14, 6, 1, 1, 11, 23, 17, 10, 26, 
    30, 17, 9, 21, 2, 17, 19, 25, 20, 27, 32, 29, 17, 11, 23, 
    39, 20, 4, 26, 6, 15, 24, 8, 30, 34, 21, 21, 18, 7, 8, 
    33, 28, 11, 24, 28, 32, 34, 41, 42, 35, 26, 22, 23, 14, 3, 
    36, 31, 16, 5, 19, 16, 19, 35, 31, 22, 21, 23, 24, 29, 12, 
    33, 33, 27, 13, 17, 30, 31, 27, 20, 18, 16, 11, 16, 30, 24, 
    36, 33, 29, 33, 22, 23, 26, 35, 25, 20, 17, 12, 16, 18, 21, 
    30, 27, 33, 28, 24, 24, 34, 34, 33, 35, 30, 28, 29, 28, 26, 
    
    -- channel=340
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 16, 
    0, 0, 0, 18, 0, 0, 0, 0, 3, 0, 3, 3, 0, 0, 15, 
    0, 0, 0, 3, 18, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 18, 8, 7, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 12, 17, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=341
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=342
    0, 13, 8, 0, 3, 9, 7, 11, 13, 13, 2, 6, 6, 7, 5, 
    0, 0, 5, 4, 1, 4, 10, 5, 9, 22, 5, 7, 0, 4, 6, 
    2, 0, 5, 1, 0, 4, 4, 11, 0, 6, 9, 15, 7, 1, 2, 
    1, 1, 1, 0, 3, 4, 3, 6, 1, 0, 9, 13, 4, 5, 3, 
    0, 0, 0, 3, 0, 1, 0, 0, 11, 0, 0, 7, 3, 5, 0, 
    0, 0, 0, 0, 4, 0, 0, 4, 0, 0, 1, 8, 5, 7, 3, 
    17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 8, 8, 7, 7, 
    11, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 13, 5, 0, 18, 
    0, 0, 0, 13, 0, 0, 2, 0, 0, 6, 4, 9, 10, 0, 7, 
    0, 0, 0, 12, 0, 0, 0, 0, 17, 8, 5, 9, 9, 0, 0, 
    0, 0, 0, 0, 20, 15, 0, 5, 1, 15, 14, 0, 11, 0, 0, 
    0, 0, 0, 0, 17, 4, 14, 10, 15, 14, 12, 18, 1, 18, 0, 
    0, 0, 7, 0, 7, 2, 0, 4, 11, 13, 17, 12, 17, 8, 9, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 5, 5, 5, 8, 13, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 4, 3, 0, 0, 1, 2, 2, 
    
    -- channel=343
    26, 0, 6, 3, 10, 3, 5, 0, 24, 0, 0, 3, 0, 0, 12, 
    15, 28, 0, 9, 8, 6, 5, 0, 21, 0, 0, 0, 0, 10, 0, 
    41, 17, 6, 7, 8, 11, 14, 0, 5, 21, 0, 1, 0, 0, 0, 
    22, 17, 13, 5, 13, 6, 10, 3, 0, 8, 2, 19, 1, 0, 0, 
    11, 11, 14, 8, 13, 11, 14, 15, 17, 0, 0, 45, 0, 0, 1, 
    0, 23, 14, 17, 16, 0, 54, 28, 29, 0, 19, 27, 0, 0, 0, 
    0, 0, 36, 34, 1, 31, 36, 41, 18, 19, 41, 17, 0, 0, 0, 
    14, 0, 39, 17, 13, 43, 20, 27, 39, 45, 62, 21, 0, 1, 18, 
    10, 0, 34, 26, 39, 5, 51, 20, 24, 28, 50, 7, 0, 0, 59, 
    19, 0, 40, 90, 0, 8, 48, 6, 39, 4, 0, 7, 0, 0, 100, 
    22, 0, 43, 78, 0, 0, 3, 0, 26, 0, 0, 0, 0, 0, 96, 
    7, 5, 18, 32, 15, 0, 0, 23, 2, 0, 0, 0, 0, 0, 28, 
    0, 8, 10, 8, 22, 14, 0, 18, 10, 2, 3, 0, 0, 0, 0, 
    16, 0, 26, 0, 32, 2, 0, 22, 1, 8, 2, 0, 4, 0, 18, 
    6, 1, 11, 0, 7, 13, 6, 6, 6, 0, 0, 0, 7, 15, 0, 
    
    -- channel=344
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=345
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 5, 5, 1, 
    7, 0, 0, 0, 0, 0, 0, 32, 9, 0, 2, 3, 7, 2, 3, 
    6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 2, 18, 2, 13, 36, 35, 49, 42, 7, 0, 0, 0, 
    0, 0, 0, 4, 50, 16, 10, 0, 0, 4, 0, 0, 3, 0, 0, 
    0, 9, 11, 0, 0, 42, 32, 40, 29, 6, 19, 6, 0, 16, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 13, 8, 26, 6, 
    0, 0, 0, 14, 0, 2, 0, 0, 0, 0, 0, 0, 1, 0, 17, 
    7, 12, 6, 4, 6, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 8, 1, 0, 0, 0, 0, 0, 0, 
    
    -- channel=346
    6, 14, 4, 3, 0, 0, 0, 1, 0, 0, 1, 0, 0, 8, 0, 
    15, 9, 4, 7, 4, 1, 0, 0, 0, 0, 1, 3, 5, 2, 2, 
    16, 13, 7, 7, 8, 4, 0, 1, 0, 0, 8, 0, 2, 2, 3, 
    14, 21, 9, 11, 10, 1, 2, 0, 5, 4, 3, 0, 0, 0, 4, 
    18, 15, 12, 9, 9, 7, 9, 11, 4, 3, 7, 0, 1, 4, 3, 
    12, 16, 17, 15, 10, 26, 32, 27, 3, 13, 8, 0, 5, 0, 3, 
    25, 22, 28, 18, 21, 35, 21, 14, 30, 29, 9, 0, 4, 0, 2, 
    3, 31, 25, 28, 37, 35, 23, 38, 41, 36, 12, 1, 8, 12, 4, 
    3, 31, 31, 19, 28, 26, 15, 16, 16, 17, 0, 0, 7, 23, 0, 
    0, 31, 39, 0, 36, 30, 6, 20, 6, 0, 0, 0, 9, 35, 7, 
    6, 24, 31, 0, 0, 2, 0, 6, 0, 0, 0, 0, 4, 36, 17, 
    7, 12, 25, 9, 7, 2, 6, 0, 0, 0, 0, 0, 0, 12, 18, 
    5, 12, 13, 27, 8, 3, 3, 0, 0, 0, 0, 0, 5, 0, 11, 
    4, 13, 9, 7, 4, 4, 13, 0, 4, 5, 2, 8, 3, 6, 8, 
    5, 11, 5, 11, 9, 11, 5, 4, 2, 0, 3, 8, 6, 1, 5, 
    
    -- channel=347
    0, 0, 0, 0, 0, 2, 4, 8, 1, 8, 10, 9, 12, 11, 1, 
    0, 0, 0, 0, 0, 0, 0, 5, 8, 11, 13, 9, 8, 5, 9, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 9, 5, 11, 9, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 12, 15, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 8, 7, 7, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 10, 8, 10, 
    15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 8, 9, 10, 
    4, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 5, 0, 
    5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 16, 7, 0, 
    7, 14, 0, 0, 14, 0, 0, 1, 0, 10, 7, 12, 15, 12, 0, 
    0, 8, 0, 0, 24, 19, 10, 25, 0, 9, 13, 14, 13, 16, 0, 
    1, 6, 0, 0, 0, 9, 8, 10, 13, 17, 15, 16, 18, 10, 0, 
    3, 8, 0, 0, 0, 0, 11, 3, 6, 11, 14, 17, 17, 12, 16, 
    6, 8, 0, 2, 0, 8, 11, 2, 8, 2, 4, 8, 2, 7, 7, 
    12, 8, 1, 5, 0, 3, 6, 4, 6, 9, 8, 6, 2, 1, 9, 
    
    -- channel=348
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=349
    15, 13, 12, 14, 14, 13, 13, 8, 7, 4, 6, 6, 6, 6, 9, 
    4, 6, 11, 11, 12, 17, 21, 15, 14, 8, 2, 7, 9, 9, 8, 
    1, 0, 10, 10, 11, 12, 17, 17, 17, 17, 14, 17, 12, 9, 10, 
    2, 1, 6, 8, 9, 14, 16, 16, 12, 13, 13, 13, 7, 9, 8, 
    0, 2, 8, 6, 10, 12, 11, 14, 13, 10, 11, 10, 6, 7, 6, 
    0, 2, 5, 8, 6, 0, 0, 0, 3, 5, 7, 5, 2, 6, 6, 
    0, 0, 0, 0, 3, 0, 0, 5, 6, 4, 4, 4, 1, 6, 6, 
    11, 0, 0, 0, 0, 0, 10, 0, 0, 0, 8, 6, 0, 5, 13, 
    18, 0, 1, 2, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 12, 
    13, 0, 0, 6, 0, 0, 6, 10, 17, 0, 9, 13, 1, 0, 8, 
    15, 0, 0, 3, 0, 0, 0, 0, 3, 4, 0, 1, 8, 0, 0, 
    11, 10, 0, 16, 16, 20, 22, 10, 0, 0, 0, 0, 0, 0, 0, 
    15, 9, 4, 0, 20, 12, 14, 19, 15, 9, 5, 2, 0, 2, 0, 
    12, 5, 11, 3, 0, 11, 8, 16, 13, 15, 16, 16, 17, 14, 4, 
    10, 14, 15, 16, 15, 14, 13, 11, 11, 14, 16, 13, 16, 14, 13, 
    
    -- channel=350
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 7, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=351
    46, 10, 18, 15, 20, 13, 16, 6, 28, 0, 0, 5, 0, 0, 22, 
    34, 36, 20, 20, 17, 20, 22, 11, 26, 1, 0, 0, 4, 16, 5, 
    43, 17, 22, 20, 21, 25, 26, 7, 21, 41, 1, 18, 3, 5, 10, 
    47, 17, 25, 20, 29, 26, 25, 22, 9, 22, 21, 29, 2, 0, 6, 
    21, 20, 28, 24, 27, 25, 25, 24, 29, 1, 21, 48, 0, 4, 5, 
    0, 32, 17, 29, 27, 13, 63, 27, 41, 1, 24, 29, 0, 1, 0, 
    0, 13, 46, 43, 24, 35, 54, 50, 15, 29, 49, 21, 0, 0, 0, 
    22, 0, 51, 30, 28, 57, 47, 37, 52, 52, 70, 27, 0, 0, 24, 
    27, 0, 46, 49, 24, 27, 64, 24, 29, 29, 42, 2, 0, 0, 67, 
    30, 0, 51, 93, 0, 24, 62, 7, 47, 11, 1, 0, 0, 0, 94, 
    38, 1, 46, 74, 0, 0, 0, 0, 29, 2, 0, 0, 0, 0, 86, 
    29, 20, 22, 53, 25, 9, 7, 17, 0, 0, 0, 0, 0, 0, 18, 
    20, 21, 27, 11, 54, 27, 8, 33, 19, 2, 0, 0, 0, 0, 0, 
    25, 3, 41, 16, 31, 9, 4, 37, 15, 20, 15, 6, 17, 5, 11, 
    17, 17, 31, 20, 32, 21, 21, 18, 20, 15, 10, 11, 23, 24, 5, 
    
    -- channel=352
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=353
    28, 0, 0, 0, 2, 0, 6, 0, 17, 0, 0, 6, 1, 0, 10, 
    0, 1, 0, 0, 0, 0, 4, 0, 27, 9, 0, 0, 0, 3, 0, 
    9, 0, 0, 0, 0, 0, 9, 0, 5, 24, 0, 3, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 21, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 5, 0, 0, 29, 0, 0, 0, 
    0, 6, 0, 0, 0, 0, 4, 0, 7, 0, 2, 31, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 8, 26, 0, 0, 24, 22, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 14, 0, 0, 12, 
    4, 0, 0, 0, 0, 0, 10, 0, 0, 0, 35, 18, 0, 0, 44, 
    17, 0, 0, 57, 0, 0, 29, 0, 21, 16, 8, 3, 0, 0, 61, 
    7, 0, 0, 73, 0, 0, 4, 0, 27, 8, 0, 0, 0, 0, 44, 
    5, 0, 0, 19, 15, 0, 0, 18, 20, 6, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 0, 19, 16, 12, 14, 0, 0, 2, 0, 
    0, 0, 6, 0, 17, 0, 0, 17, 2, 3, 3, 0, 4, 0, 6, 
    4, 0, 5, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 8, 0, 
    
    -- channel=354
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 2, 16, 0, 0, 17, 0, 0, 0, 
    0, 7, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 12, 0, 18, 20, 29, 54, 17, 0, 0, 0, 
    0, 0, 0, 0, 28, 0, 20, 0, 0, 16, 0, 0, 0, 0, 0, 
    0, 0, 0, 26, 0, 27, 28, 4, 37, 5, 9, 6, 0, 0, 1, 
    5, 0, 2, 0, 0, 0, 0, 0, 4, 3, 2, 0, 3, 0, 16, 
    0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=355
    0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 2, 0, 0, 0, 
    2, 0, 0, 0, 9, 0, 0, 18, 1, 0, 6, 23, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 5, 7, 0, 0, 1, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 2, 
    0, 0, 0, 12, 0, 20, 8, 28, 21, 45, 53, 17, 0, 0, 0, 
    0, 0, 0, 15, 24, 0, 15, 0, 1, 21, 0, 0, 0, 0, 0, 
    0, 2, 10, 22, 4, 60, 35, 37, 38, 13, 19, 0, 0, 0, 0, 
    8, 0, 3, 0, 0, 0, 0, 4, 18, 10, 4, 15, 5, 22, 0, 
    0, 0, 3, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 12, 
    1, 6, 1, 5, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=356
    9, 13, 20, 22, 21, 24, 23, 16, 7, 5, 7, 7, 5, 9, 5, 
    13, 14, 19, 21, 24, 24, 27, 28, 18, 5, 7, 11, 12, 11, 9, 
    9, 10, 19, 22, 21, 25, 26, 26, 23, 10, 13, 15, 15, 14, 12, 
    2, 10, 18, 21, 22, 28, 28, 24, 24, 23, 19, 15, 14, 13, 13, 
    9, 12, 17, 19, 23, 21, 15, 13, 18, 25, 18, 8, 8, 11, 12, 
    6, 12, 15, 17, 17, 0, 0, 5, 6, 11, 14, 1, 5, 9, 11, 
    7, 8, 7, 9, 6, 4, 5, 0, 0, 0, 3, 0, 0, 7, 10, 
    10, 10, 8, 6, 2, 6, 14, 2, 0, 0, 0, 0, 0, 4, 5, 
    19, 9, 5, 6, 0, 4, 15, 10, 9, 8, 2, 0, 0, 2, 0, 
    20, 10, 0, 3, 1, 6, 11, 14, 12, 1, 0, 3, 5, 0, 0, 
    21, 13, 0, 0, 0, 0, 11, 18, 12, 2, 0, 3, 7, 5, 0, 
    21, 18, 4, 5, 12, 12, 12, 6, 0, 0, 0, 0, 3, 11, 1, 
    25, 20, 12, 8, 9, 14, 18, 14, 3, 0, 0, 0, 0, 3, 3, 
    19, 19, 18, 14, 12, 13, 20, 22, 13, 12, 9, 10, 8, 11, 8, 
    19, 22, 22, 19, 15, 21, 22, 22, 20, 20, 21, 20, 19, 17, 14, 
    
    -- channel=357
    25, 52, 3, 8, 5, 6, 2, 7, 0, 0, 0, 11, 9, 7, 3, 
    4, 0, 8, 9, 8, 13, 14, 13, 12, 7, 0, 0, 2, 5, 2, 
    1, 0, 10, 2, 6, 5, 10, 3, 9, 47, 37, 22, 0, 0, 8, 
    0, 0, 0, 3, 0, 0, 0, 1, 0, 0, 14, 10, 0, 4, 0, 
    0, 2, 5, 3, 2, 0, 3, 21, 10, 0, 0, 0, 0, 0, 0, 
    0, 14, 11, 4, 0, 5, 24, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 0, 0, 0, 15, 2, 0, 40, 51, 32, 4, 2, 3, 2, 0, 
    9, 0, 0, 0, 11, 12, 23, 0, 0, 5, 18, 0, 0, 23, 15, 
    8, 10, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 14, 
    3, 0, 0, 0, 0, 0, 0, 21, 16, 0, 13, 20, 3, 0, 25, 
    5, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 
    0, 6, 0, 45, 36, 47, 39, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 4, 0, 18, 0, 7, 30, 37, 37, 32, 27, 8, 0, 0, 
    0, 0, 0, 0, 0, 10, 2, 5, 18, 30, 34, 44, 43, 32, 0, 
    0, 22, 4, 16, 25, 14, 0, 0, 0, 0, 9, 8, 13, 10, 17, 
    
    -- channel=358
    9, 25, 17, 17, 16, 19, 17, 19, 18, 20, 15, 18, 18, 18, 14, 
    22, 19, 18, 16, 16, 18, 18, 17, 15, 23, 18, 15, 12, 14, 14, 
    18, 18, 21, 17, 17, 17, 18, 20, 12, 14, 16, 16, 14, 12, 15, 
    16, 17, 18, 18, 18, 18, 15, 19, 17, 12, 16, 19, 15, 17, 14, 
    17, 19, 18, 19, 19, 16, 13, 11, 20, 16, 16, 17, 18, 15, 14, 
    23, 14, 19, 16, 20, 9, 12, 15, 14, 13, 15, 15, 19, 18, 16, 
    30, 14, 12, 14, 16, 16, 14, 7, 11, 13, 13, 16, 21, 19, 17, 
    14, 15, 11, 12, 13, 9, 15, 5, 8, 6, 14, 18, 19, 12, 17, 
    8, 11, 9, 20, 16, 14, 17, 15, 16, 19, 13, 19, 25, 13, 17, 
    7, 12, 7, 20, 9, 16, 8, 2, 12, 16, 18, 16, 21, 8, 8, 
    8, 12, 11, 5, 31, 27, 19, 18, 13, 21, 23, 14, 21, 12, 2, 
    5, 12, 7, 14, 10, 12, 14, 12, 24, 24, 22, 28, 20, 24, 3, 
    13, 3, 18, 10, 18, 11, 7, 8, 15, 17, 21, 22, 25, 20, 21, 
    11, 10, 8, 20, 12, 13, 10, 9, 10, 12, 12, 13, 15, 19, 7, 
    4, 12, 7, 8, 10, 9, 13, 8, 12, 12, 12, 10, 11, 12, 14, 
    
    -- channel=359
    22, 20, 26, 28, 29, 28, 24, 21, 13, 9, 11, 9, 9, 10, 6, 
    27, 30, 28, 30, 31, 31, 30, 27, 20, 8, 11, 11, 12, 12, 11, 
    27, 30, 31, 33, 33, 35, 33, 33, 29, 10, 13, 11, 16, 15, 12, 
    23, 31, 31, 33, 34, 35, 33, 30, 31, 29, 26, 17, 14, 15, 15, 
    21, 27, 32, 34, 35, 34, 28, 26, 25, 30, 28, 17, 14, 15, 14, 
    18, 28, 32, 32, 36, 27, 19, 24, 19, 22, 22, 13, 12, 14, 14, 
    19, 27, 30, 28, 27, 28, 20, 9, 15, 18, 13, 4, 8, 13, 13, 
    14, 24, 25, 27, 26, 26, 26, 22, 21, 19, 10, 3, 7, 13, 10, 
    16, 22, 23, 22, 27, 27, 26, 28, 22, 21, 12, 3, 8, 18, 5, 
    19, 24, 20, 13, 23, 23, 18, 18, 20, 8, 2, 3, 8, 20, 6, 
    19, 23, 20, 8, 8, 16, 13, 27, 13, 5, 4, 5, 8, 22, 10, 
    20, 21, 18, 12, 9, 3, 8, 13, 4, 0, 0, 4, 10, 17, 16, 
    19, 21, 21, 23, 17, 18, 17, 10, 0, 0, 0, 0, 6, 9, 22, 
    20, 22, 20, 18, 13, 17, 19, 17, 11, 7, 6, 7, 7, 10, 10, 
    17, 18, 18, 18, 15, 21, 21, 21, 18, 15, 19, 20, 18, 17, 13, 
    
    -- channel=360
    10, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 1, 
    6, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 7, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    14, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 2, 0, 0, 0, 0, 1, 3, 0, 0, 0, 16, 0, 0, 0, 
    0, 4, 3, 1, 0, 8, 29, 11, 12, 0, 2, 11, 0, 0, 0, 
    0, 0, 16, 15, 4, 16, 20, 25, 12, 12, 17, 7, 0, 0, 0, 
    0, 0, 19, 7, 13, 24, 4, 17, 25, 28, 32, 9, 0, 0, 0, 
    0, 0, 19, 11, 25, 7, 20, 3, 10, 8, 22, 3, 0, 0, 29, 
    0, 0, 29, 41, 0, 3, 19, 0, 3, 0, 0, 0, 0, 0, 53, 
    0, 0, 25, 36, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 54, 
    0, 0, 10, 18, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 17, 
    0, 0, 0, 2, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=361
    38, 10, 24, 20, 26, 25, 27, 19, 24, 15, 12, 14, 15, 7, 18, 
    20, 25, 29, 23, 23, 27, 31, 23, 29, 23, 9, 14, 8, 14, 17, 
    24, 17, 24, 24, 24, 29, 30, 30, 28, 25, 7, 19, 13, 15, 12, 
    33, 15, 24, 21, 27, 28, 30, 27, 23, 25, 27, 30, 17, 13, 14, 
    16, 15, 22, 25, 27, 24, 23, 16, 28, 18, 22, 31, 13, 13, 12, 
    5, 20, 18, 23, 28, 12, 12, 13, 22, 9, 19, 34, 7, 15, 12, 
    0, 11, 17, 17, 19, 7, 24, 12, 0, 7, 25, 21, 8, 13, 12, 
    17, 0, 17, 17, 3, 18, 21, 3, 7, 6, 23, 20, 7, 1, 23, 
    20, 0, 14, 25, 0, 18, 27, 16, 12, 17, 33, 20, 1, 0, 31, 
    21, 0, 6, 34, 0, 4, 36, 0, 25, 21, 16, 8, 0, 0, 27, 
    19, 3, 7, 43, 0, 14, 18, 7, 35, 20, 12, 10, 6, 0, 20, 
    24, 7, 7, 26, 22, 10, 7, 14, 21, 13, 7, 7, 7, 8, 5, 
    15, 16, 14, 10, 31, 16, 13, 22, 15, 10, 11, 4, 0, 16, 5, 
    15, 12, 22, 13, 18, 13, 7, 21, 16, 12, 14, 5, 13, 9, 10, 
    17, 5, 20, 13, 16, 13, 17, 21, 17, 21, 14, 14, 18, 19, 14, 
    
    -- channel=362
    56, 47, 69, 72, 73, 68, 64, 52, 48, 26, 34, 30, 29, 38, 36, 
    80, 82, 67, 75, 80, 76, 69, 68, 57, 18, 31, 40, 48, 48, 38, 
    78, 81, 74, 82, 84, 82, 81, 70, 73, 44, 41, 40, 49, 50, 46, 
    67, 75, 81, 84, 88, 89, 88, 74, 76, 80, 63, 53, 43, 43, 50, 
    61, 78, 83, 83, 90, 87, 76, 76, 63, 77, 74, 61, 39, 46, 50, 
    40, 74, 87, 87, 80, 83, 76, 80, 68, 63, 65, 39, 29, 36, 46, 
    33, 84, 96, 90, 70, 93, 86, 67, 56, 62, 55, 23, 15, 33, 41, 
    50, 69, 96, 81, 89, 97, 83, 100, 92, 90, 68, 25, 13, 45, 31, 
    69, 71, 93, 67, 107, 89, 98, 93, 94, 84, 62, 15, 9, 62, 45, 
    73, 75, 99, 70, 66, 80, 83, 82, 61, 27, 11, 13, 15, 68, 64, 
    81, 75, 96, 57, 8, 40, 50, 74, 57, 11, 13, 21, 19, 65, 87, 
    76, 77, 77, 58, 35, 28, 34, 38, 1, 0, 0, 0, 19, 40, 83, 
    72, 82, 69, 81, 61, 60, 63, 47, 16, 0, 0, 0, 9, 17, 51, 
    78, 72, 81, 57, 68, 58, 72, 73, 49, 39, 32, 35, 31, 34, 48, 
    74, 74, 77, 69, 62, 76, 76, 73, 65, 59, 62, 68, 65, 60, 47, 
    
    -- channel=363
    0, 6, 2, 10, 0, 6, 2, 14, 0, 9, 9, 2, 6, 17, 0, 
    2, 0, 6, 3, 6, 2, 0, 11, 0, 0, 18, 11, 12, 1, 6, 
    0, 5, 5, 7, 7, 2, 0, 14, 5, 0, 10, 0, 11, 11, 8, 
    0, 4, 3, 12, 3, 7, 1, 5, 16, 4, 3, 0, 6, 16, 10, 
    8, 7, 2, 7, 2, 7, 0, 2, 0, 24, 12, 0, 15, 10, 10, 
    64, 0, 5, 2, 0, 23, 0, 1, 0, 20, 0, 0, 17, 9, 14, 
    53, 30, 0, 0, 11, 6, 0, 0, 0, 0, 0, 0, 12, 9, 9, 
    0, 57, 0, 4, 17, 0, 0, 7, 0, 0, 0, 0, 20, 12, 0, 
    0, 45, 0, 0, 12, 17, 0, 12, 9, 4, 0, 0, 37, 30, 0, 
    0, 52, 0, 0, 56, 20, 0, 19, 0, 0, 0, 0, 34, 49, 0, 
    0, 40, 0, 0, 23, 22, 12, 34, 0, 3, 8, 11, 20, 66, 0, 
    3, 16, 10, 0, 0, 2, 5, 0, 0, 5, 1, 18, 30, 36, 5, 
    15, 9, 7, 17, 0, 0, 14, 0, 0, 0, 0, 3, 21, 13, 25, 
    2, 32, 0, 20, 0, 6, 21, 0, 4, 0, 0, 5, 0, 9, 0, 
    7, 15, 0, 11, 1, 2, 8, 8, 7, 6, 13, 13, 1, 0, 16, 
    
    -- channel=364
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=365
    45, 0, 5, 4, 13, 5, 15, 0, 23, 0, 3, 9, 2, 0, 21, 
    5, 18, 7, 6, 6, 9, 15, 9, 30, 4, 0, 0, 0, 10, 4, 
    18, 1, 3, 3, 4, 8, 19, 0, 16, 40, 0, 11, 0, 3, 4, 
    24, 0, 5, 0, 5, 7, 11, 10, 0, 12, 9, 23, 8, 0, 0, 
    2, 0, 5, 1, 5, 2, 14, 10, 12, 0, 1, 43, 0, 0, 1, 
    0, 10, 0, 2, 5, 0, 20, 0, 32, 0, 8, 36, 0, 0, 0, 
    0, 0, 7, 15, 0, 0, 23, 42, 0, 0, 33, 26, 0, 0, 0, 
    12, 0, 14, 0, 0, 19, 7, 0, 1, 13, 45, 24, 0, 0, 15, 
    14, 0, 8, 8, 0, 0, 23, 0, 0, 0, 44, 20, 0, 0, 61, 
    23, 0, 5, 70, 0, 0, 49, 0, 26, 16, 15, 11, 0, 0, 85, 
    18, 0, 3, 85, 0, 0, 6, 0, 36, 10, 0, 4, 0, 0, 71, 
    16, 0, 0, 41, 22, 14, 0, 20, 14, 1, 4, 0, 0, 0, 12, 
    1, 4, 0, 0, 26, 15, 6, 29, 26, 14, 13, 0, 0, 3, 0, 
    6, 0, 21, 0, 28, 3, 0, 29, 11, 16, 18, 2, 16, 0, 15, 
    11, 0, 18, 0, 15, 4, 0, 9, 7, 8, 0, 0, 11, 18, 0, 
    
    -- channel=366
    28, 45, 11, 15, 15, 10, 12, 10, 9, 0, 3, 9, 7, 8, 10, 
    12, 10, 10, 14, 16, 19, 19, 18, 23, 1, 0, 0, 11, 11, 5, 
    7, 6, 13, 8, 13, 10, 18, 3, 23, 50, 38, 22, 1, 0, 12, 
    0, 6, 6, 10, 7, 10, 6, 9, 1, 11, 12, 12, 0, 3, 2, 
    0, 9, 12, 7, 9, 12, 8, 26, 5, 0, 3, 9, 0, 0, 2, 
    0, 11, 14, 11, 0, 22, 27, 0, 0, 6, 0, 0, 0, 0, 0, 
    2, 0, 9, 12, 14, 8, 0, 50, 49, 30, 8, 2, 0, 4, 0, 
    12, 0, 9, 0, 19, 23, 26, 18, 12, 20, 29, 3, 0, 31, 10, 
    20, 14, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 20, 
    10, 0, 11, 7, 0, 0, 0, 46, 19, 0, 9, 23, 0, 13, 41, 
    14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 23, 
    0, 12, 0, 47, 35, 49, 42, 8, 0, 0, 0, 0, 0, 0, 0, 
    12, 6, 1, 0, 25, 10, 13, 33, 37, 31, 23, 22, 2, 0, 0, 
    2, 0, 4, 0, 0, 14, 7, 16, 22, 33, 37, 47, 43, 30, 12, 
    9, 25, 12, 21, 27, 19, 5, 0, 5, 3, 14, 15, 18, 16, 17, 
    
    -- channel=367
    11, 7, 11, 13, 13, 8, 6, 1, 0, 0, 0, 0, 0, 0, 0, 
    23, 21, 11, 16, 17, 15, 9, 9, 3, 0, 0, 0, 2, 2, 0, 
    22, 19, 16, 19, 20, 19, 17, 8, 12, 7, 1, 0, 0, 0, 1, 
    17, 18, 19, 21, 23, 22, 20, 13, 12, 18, 10, 1, 0, 0, 1, 
    11, 21, 23, 20, 24, 18, 19, 21, 10, 12, 15, 6, 0, 0, 1, 
    0, 22, 26, 24, 17, 22, 32, 17, 14, 9, 11, 0, 0, 0, 0, 
    0, 23, 35, 30, 21, 31, 30, 27, 18, 20, 11, 0, 0, 0, 0, 
    5, 13, 36, 23, 35, 42, 31, 39, 39, 39, 23, 0, 0, 4, 0, 
    14, 20, 37, 17, 36, 30, 34, 19, 25, 15, 1, 0, 0, 11, 7, 
    16, 17, 43, 19, 0, 23, 25, 28, 12, 0, 0, 0, 0, 14, 24, 
    22, 17, 35, 8, 0, 0, 0, 2, 0, 0, 0, 0, 0, 7, 34, 
    17, 21, 21, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 
    18, 22, 17, 21, 14, 8, 11, 5, 0, 0, 0, 0, 0, 0, 0, 
    17, 14, 22, 9, 14, 9, 15, 18, 5, 3, 0, 1, 0, 0, 1, 
    17, 21, 21, 18, 17, 21, 15, 12, 10, 7, 9, 14, 14, 10, 2, 
    
    -- channel=368
    24, 15, 30, 31, 31, 30, 25, 24, 18, 12, 13, 10, 10, 15, 11, 
    46, 45, 34, 36, 36, 31, 26, 25, 14, 5, 17, 17, 17, 16, 14, 
    46, 48, 39, 43, 42, 42, 33, 33, 29, 2, 5, 7, 18, 21, 16, 
    46, 47, 45, 45, 48, 44, 41, 33, 40, 37, 27, 19, 16, 16, 21, 
    45, 44, 45, 47, 47, 42, 40, 32, 31, 41, 38, 25, 19, 21, 22, 
    43, 42, 47, 48, 51, 49, 42, 56, 39, 32, 35, 22, 16, 17, 21, 
    23, 59, 58, 51, 43, 63, 58, 19, 20, 32, 28, 8, 9, 14, 18, 
    17, 47, 56, 53, 57, 57, 44, 56, 60, 54, 27, 9, 12, 15, 9, 
    20, 39, 53, 45, 72, 69, 55, 67, 64, 66, 48, 9, 11, 36, 13, 
    27, 48, 61, 33, 62, 58, 47, 25, 20, 15, 0, 0, 9, 42, 18, 
    30, 47, 63, 26, 6, 46, 39, 50, 35, 7, 13, 10, 4, 53, 40, 
    35, 33, 48, 17, 3, 0, 0, 8, 3, 0, 0, 5, 17, 35, 49, 
    28, 37, 38, 56, 24, 24, 22, 5, 0, 0, 0, 0, 4, 11, 36, 
    32, 42, 37, 33, 36, 22, 31, 24, 13, 5, 0, 0, 0, 4, 17, 
    29, 25, 29, 24, 21, 28, 30, 33, 27, 21, 21, 26, 23, 19, 15, 
    
    -- channel=369
    65, 62, 38, 40, 41, 33, 29, 27, 22, 9, 15, 18, 21, 21, 21, 
    46, 45, 42, 46, 45, 49, 43, 35, 34, 11, 6, 13, 23, 23, 21, 
    44, 43, 46, 44, 48, 46, 45, 37, 48, 56, 48, 32, 17, 17, 26, 
    43, 45, 42, 46, 45, 42, 41, 35, 33, 42, 43, 30, 14, 20, 21, 
    25, 44, 49, 46, 50, 46, 47, 60, 37, 23, 35, 26, 12, 16, 19, 
    5, 52, 59, 53, 41, 67, 64, 18, 21, 35, 27, 9, 8, 12, 16, 
    20, 33, 57, 50, 60, 51, 39, 71, 82, 67, 35, 13, 10, 17, 13, 
    28, 31, 52, 45, 64, 76, 66, 61, 61, 63, 53, 11, 10, 46, 28, 
    39, 46, 65, 35, 25, 33, 38, 4, 4, 0, 0, 0, 5, 36, 33, 
    33, 37, 59, 21, 0, 32, 30, 62, 40, 0, 19, 19, 7, 47, 59, 
    38, 27, 32, 24, 0, 0, 0, 0, 0, 0, 0, 1, 16, 19, 51, 
    29, 36, 35, 75, 48, 48, 45, 14, 0, 0, 0, 0, 0, 0, 25, 
    35, 39, 31, 28, 52, 26, 36, 46, 36, 27, 17, 16, 5, 2, 5, 
    24, 20, 33, 17, 17, 35, 33, 34, 39, 40, 43, 51, 49, 37, 23, 
    37, 43, 39, 46, 50, 45, 28, 24, 24, 26, 34, 39, 41, 35, 34, 
    
    -- channel=370
    0, 17, 7, 11, 2, 2, 0, 0, 0, 3, 1, 0, 0, 4, 2, 
    10, 10, 1, 1, 4, 4, 7, 4, 0, 0, 0, 5, 9, 3, 0, 
    9, 0, 5, 4, 4, 3, 1, 2, 7, 0, 7, 8, 6, 2, 5, 
    0, 10, 3, 6, 6, 6, 7, 7, 11, 2, 0, 0, 0, 0, 0, 
    9, 3, 7, 0, 3, 10, 6, 3, 5, 5, 6, 11, 5, 7, 3, 
    0, 0, 0, 9, 4, 0, 22, 21, 14, 7, 7, 0, 8, 3, 1, 
    14, 2, 10, 5, 0, 12, 0, 0, 4, 6, 3, 0, 0, 0, 3, 
    0, 4, 8, 4, 8, 13, 17, 6, 9, 6, 11, 9, 2, 6, 7, 
    5, 8, 7, 12, 7, 0, 14, 1, 4, 10, 0, 0, 0, 0, 5, 
    0, 0, 7, 12, 12, 26, 4, 23, 8, 0, 0, 11, 7, 0, 8, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 4, 7, 6, 3, 
    0, 4, 0, 1, 11, 9, 14, 2, 0, 0, 0, 0, 0, 6, 0, 
    7, 0, 0, 5, 27, 21, 0, 4, 1, 0, 0, 0, 5, 0, 0, 
    4, 0, 9, 0, 0, 0, 4, 1, 0, 11, 3, 10, 6, 10, 8, 
    0, 8, 0, 7, 4, 7, 4, 8, 3, 0, 7, 5, 5, 4, 3, 
    
    -- channel=371
    23, 18, 11, 11, 14, 15, 15, 10, 16, 7, 8, 15, 9, 4, 11, 
    6, 12, 12, 12, 13, 14, 18, 16, 27, 16, 3, 2, 3, 11, 6, 
    17, 5, 11, 10, 10, 15, 19, 9, 14, 28, 12, 14, 5, 3, 8, 
    4, 6, 9, 7, 8, 10, 9, 11, 5, 8, 15, 22, 12, 6, 5, 
    5, 3, 9, 10, 10, 11, 9, 12, 17, 0, 3, 23, 3, 6, 6, 
    0, 16, 5, 8, 11, 0, 17, 0, 6, 2, 10, 15, 4, 8, 3, 
    0, 0, 3, 9, 2, 2, 0, 20, 11, 6, 19, 17, 8, 9, 6, 
    12, 0, 3, 0, 0, 3, 7, 0, 0, 2, 21, 14, 1, 9, 19, 
    6, 0, 0, 7, 0, 0, 9, 0, 0, 0, 6, 11, 0, 0, 29, 
    14, 0, 0, 35, 0, 0, 7, 0, 23, 11, 12, 18, 0, 0, 38, 
    9, 0, 0, 32, 14, 0, 0, 0, 6, 13, 4, 4, 5, 0, 20, 
    1, 1, 0, 18, 22, 12, 9, 22, 19, 12, 14, 7, 0, 0, 0, 
    3, 0, 3, 0, 12, 12, 3, 20, 20, 22, 24, 16, 9, 8, 0, 
    5, 0, 5, 1, 10, 6, 0, 13, 8, 13, 13, 12, 17, 11, 11, 
    3, 4, 4, 2, 8, 7, 4, 2, 8, 4, 5, 3, 8, 14, 4, 
    
    -- channel=372
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 16, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 32, 
    0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 
    0, 0, 0, 2, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 8, 5, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=373
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 13, 0, 5, 0, 0, 0, 0, 0, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=374
    31, 0, 0, 0, 0, 0, 1, 0, 24, 0, 0, 0, 0, 0, 10, 
    0, 7, 0, 0, 0, 0, 3, 0, 27, 6, 0, 0, 0, 3, 0, 
    23, 0, 0, 0, 0, 0, 6, 0, 0, 25, 0, 5, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 21, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 45, 0, 0, 0, 
    0, 6, 0, 0, 1, 0, 25, 0, 10, 0, 6, 35, 0, 0, 0, 
    0, 0, 2, 4, 0, 0, 6, 24, 0, 0, 35, 22, 0, 0, 0, 
    12, 0, 5, 0, 0, 7, 0, 0, 0, 4, 49, 22, 0, 0, 26, 
    2, 0, 0, 11, 0, 0, 24, 0, 0, 0, 40, 9, 0, 0, 65, 
    13, 0, 0, 88, 0, 0, 36, 0, 45, 9, 0, 10, 0, 0, 98, 
    9, 0, 0, 89, 0, 0, 0, 0, 24, 3, 0, 0, 0, 0, 74, 
    0, 0, 0, 20, 26, 0, 0, 31, 12, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 14, 3, 0, 23, 20, 12, 14, 0, 0, 0, 0, 
    1, 0, 12, 0, 15, 0, 0, 15, 0, 5, 3, 0, 7, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 
    
    -- channel=375
    18, 0, 5, 2, 7, 4, 8, 1, 18, 5, 1, 3, 2, 0, 10, 
    13, 15, 7, 4, 3, 6, 7, 1, 15, 11, 0, 0, 0, 2, 3, 
    15, 9, 6, 5, 6, 6, 9, 3, 8, 14, 0, 2, 0, 1, 0, 
    21, 2, 8, 5, 8, 5, 6, 7, 0, 3, 4, 15, 2, 0, 0, 
    4, 5, 7, 7, 8, 8, 5, 2, 7, 0, 6, 26, 3, 1, 0, 
    0, 2, 4, 6, 9, 7, 10, 11, 18, 0, 5, 22, 0, 4, 0, 
    0, 2, 8, 11, 6, 2, 18, 13, 0, 0, 16, 14, 1, 3, 0, 
    2, 0, 10, 6, 0, 9, 3, 3, 6, 6, 23, 18, 0, 0, 8, 
    1, 0, 6, 15, 7, 6, 17, 10, 12, 13, 30, 18, 0, 0, 30, 
    0, 0, 8, 37, 0, 0, 21, 0, 6, 13, 7, 2, 0, 0, 34, 
    1, 0, 10, 35, 0, 9, 9, 0, 26, 13, 10, 3, 0, 0, 33, 
    0, 0, 2, 16, 0, 0, 0, 5, 16, 11, 10, 3, 0, 0, 9, 
    0, 0, 0, 1, 20, 3, 0, 5, 7, 5, 8, 3, 0, 4, 0, 
    0, 0, 5, 0, 11, 0, 0, 3, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, 
    
    -- channel=376
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 0, 0, 0, 0, 0, 0, 21, 12, 0, 0, 10, 0, 0, 0, 
    0, 9, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 10, 0, 30, 29, 45, 54, 13, 0, 0, 0, 
    0, 0, 0, 0, 55, 4, 11, 0, 0, 10, 0, 0, 0, 0, 0, 
    0, 0, 5, 1, 0, 46, 36, 28, 40, 6, 18, 6, 0, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 5, 2, 10, 9, 12, 12, 
    0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=377
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=378
    7, 10, 20, 25, 19, 20, 22, 24, 0, 19, 18, 10, 15, 19, 9, 
    22, 12, 28, 18, 21, 22, 21, 26, 5, 9, 23, 21, 21, 10, 19, 
    0, 18, 24, 26, 24, 23, 18, 32, 26, 0, 12, 12, 18, 24, 19, 
    17, 12, 22, 29, 21, 32, 24, 29, 32, 25, 21, 4, 17, 23, 20, 
    24, 21, 20, 24, 24, 25, 21, 15, 8, 38, 33, 0, 26, 20, 19, 
    78, 7, 17, 19, 23, 34, 0, 7, 17, 27, 10, 1, 21, 20, 22, 
    30, 48, 5, 8, 30, 0, 13, 0, 0, 0, 0, 2, 16, 17, 16, 
    3, 48, 6, 20, 23, 2, 14, 9, 0, 0, 0, 0, 29, 16, 0, 
    15, 39, 6, 9, 5, 36, 0, 19, 22, 16, 0, 11, 37, 26, 0, 
    10, 42, 3, 0, 49, 28, 2, 23, 0, 16, 12, 0, 33, 39, 0, 
    8, 40, 0, 0, 9, 20, 29, 28, 20, 16, 13, 22, 24, 49, 0, 
    25, 18, 18, 0, 0, 14, 11, 0, 6, 10, 5, 15, 37, 33, 17, 
    30, 20, 12, 33, 12, 14, 26, 1, 0, 0, 0, 3, 12, 27, 12, 
    11, 43, 9, 30, 9, 15, 22, 11, 16, 6, 10, 8, 6, 12, 4, 
    20, 17, 20, 22, 17, 9, 20, 25, 18, 24, 25, 24, 17, 9, 28, 
    
    -- channel=379
    20, 7, 32, 32, 36, 35, 36, 26, 28, 20, 24, 23, 23, 19, 23, 
    24, 31, 31, 32, 34, 35, 36, 36, 34, 18, 25, 26, 26, 27, 24, 
    24, 31, 29, 33, 33, 36, 41, 35, 32, 19, 15, 23, 31, 30, 24, 
    26, 22, 32, 30, 34, 41, 41, 35, 34, 37, 29, 31, 32, 28, 28, 
    19, 27, 30, 32, 36, 31, 31, 26, 31, 40, 30, 32, 27, 26, 28, 
    24, 25, 28, 27, 30, 12, 10, 23, 36, 24, 29, 32, 21, 25, 28, 
    4, 27, 24, 27, 16, 13, 29, 16, 1, 7, 24, 20, 16, 25, 27, 
    28, 14, 26, 18, 10, 16, 17, 15, 12, 14, 22, 17, 12, 14, 17, 
    34, 10, 19, 16, 32, 30, 36, 40, 39, 35, 47, 29, 11, 16, 26, 
    39, 14, 16, 38, 19, 17, 44, 20, 28, 27, 19, 15, 11, 8, 24, 
    37, 21, 25, 40, 17, 38, 48, 47, 46, 20, 23, 24, 14, 8, 30, 
    39, 30, 20, 20, 13, 13, 15, 28, 22, 17, 12, 16, 24, 20, 31, 
    33, 35, 26, 24, 20, 31, 35, 22, 11, 6, 7, 7, 11, 26, 28, 
    40, 34, 36, 27, 34, 32, 31, 40, 24, 17, 17, 11, 13, 14, 23, 
    38, 29, 38, 27, 24, 33, 36, 39, 34, 37, 31, 30, 29, 31, 22, 
    
    -- channel=380
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 3, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 4, 3, 0, 2, 18, 20, 1, 2, 4, 0, 0, 0, 0, 
    5, 4, 14, 8, 0, 17, 7, 1, 9, 8, 4, 0, 0, 0, 0, 
    0, 9, 14, 11, 13, 17, 6, 17, 21, 19, 8, 0, 0, 0, 0, 
    0, 9, 15, 6, 21, 7, 15, 10, 13, 17, 6, 0, 0, 6, 0, 
    0, 10, 22, 8, 24, 14, 6, 10, 2, 0, 0, 0, 0, 9, 10, 
    3, 7, 21, 1, 0, 3, 0, 7, 0, 0, 0, 0, 0, 13, 18, 
    1, 4, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 11, 
    0, 4, 3, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    5, 2, 6, 0, 6, 0, 4, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 3, 0, 0, 0, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=381
    61, 30, 44, 40, 46, 44, 49, 39, 41, 27, 26, 27, 29, 23, 34, 
    35, 39, 47, 45, 46, 49, 52, 47, 53, 35, 20, 30, 27, 32, 34, 
    39, 30, 41, 45, 45, 51, 51, 51, 53, 49, 32, 40, 30, 35, 31, 
    42, 30, 42, 42, 45, 48, 52, 49, 41, 48, 50, 46, 34, 30, 31, 
    33, 30, 39, 42, 46, 44, 38, 35, 41, 35, 41, 42, 23, 30, 29, 
    13, 40, 34, 40, 44, 31, 26, 24, 30, 25, 32, 43, 18, 28, 26, 
    0, 25, 33, 33, 36, 18, 41, 36, 19, 20, 37, 34, 18, 24, 25, 
    35, 10, 33, 36, 18, 38, 39, 26, 24, 25, 34, 29, 19, 20, 37, 
    43, 15, 31, 35, 0, 30, 37, 25, 21, 23, 38, 27, 9, 10, 38, 
    45, 17, 22, 34, 7, 11, 50, 27, 42, 36, 27, 23, 15, 7, 36, 
    42, 23, 22, 57, 3, 14, 23, 15, 47, 26, 15, 22, 20, 5, 37, 
    50, 27, 32, 41, 50, 38, 31, 33, 26, 17, 13, 4, 14, 15, 27, 
    38, 43, 29, 34, 42, 32, 35, 47, 36, 26, 23, 17, 9, 26, 7, 
    34, 31, 44, 27, 40, 30, 30, 45, 40, 36, 38, 30, 37, 27, 36, 
    45, 30, 46, 39, 41, 38, 40, 42, 39, 42, 37, 38, 42, 41, 35, 
    
    -- channel=382
    33, 32, 51, 56, 53, 52, 49, 38, 30, 20, 27, 24, 21, 30, 28, 
    50, 52, 48, 53, 58, 56, 56, 55, 41, 14, 25, 34, 40, 39, 29, 
    49, 47, 52, 58, 58, 60, 61, 55, 52, 28, 31, 36, 43, 41, 37, 
    36, 46, 55, 58, 61, 68, 67, 58, 59, 59, 46, 40, 36, 35, 40, 
    40, 50, 55, 54, 61, 61, 55, 52, 50, 62, 55, 42, 30, 37, 39, 
    22, 47, 54, 57, 55, 39, 45, 51, 46, 45, 50, 26, 23, 29, 36, 
    25, 51, 57, 55, 39, 50, 46, 35, 28, 33, 37, 17, 12, 25, 34, 
    38, 44, 58, 46, 47, 55, 56, 53, 47, 47, 41, 18, 9, 28, 26, 
    55, 46, 55, 43, 57, 48, 69, 57, 58, 54, 40, 9, 6, 34, 31, 
    59, 46, 53, 50, 36, 52, 59, 58, 49, 21, 11, 16, 15, 33, 35, 
    65, 51, 52, 34, 6, 24, 41, 55, 45, 11, 10, 17, 20, 37, 43, 
    61, 59, 43, 34, 28, 27, 33, 33, 2, 0, 0, 0, 14, 34, 43, 
    62, 61, 48, 51, 45, 50, 51, 39, 13, 0, 0, 0, 9, 16, 32, 
    64, 58, 62, 45, 50, 43, 57, 61, 38, 34, 26, 27, 24, 28, 34, 
    55, 61, 63, 56, 48, 61, 61, 59, 53, 50, 53, 54, 53, 49, 38, 
    
    -- channel=383
    0, 30, 0, 6, 0, 2, 0, 8, 0, 0, 2, 0, 4, 20, 0, 
    0, 0, 0, 1, 3, 0, 0, 4, 0, 0, 15, 3, 10, 0, 0, 
    0, 10, 2, 2, 2, 0, 0, 7, 0, 0, 23, 0, 7, 0, 3, 
    0, 11, 0, 7, 0, 0, 0, 0, 7, 0, 0, 0, 0, 13, 4, 
    0, 11, 2, 3, 1, 0, 0, 4, 0, 16, 0, 0, 12, 2, 3, 
    56, 0, 16, 1, 0, 21, 0, 0, 0, 19, 0, 0, 19, 2, 11, 
    90, 19, 0, 0, 6, 20, 0, 0, 27, 16, 0, 0, 13, 9, 6, 
    0, 69, 0, 0, 26, 0, 0, 13, 0, 0, 0, 0, 14, 22, 0, 
    0, 55, 0, 0, 28, 3, 0, 0, 0, 0, 0, 0, 43, 43, 0, 
    0, 61, 0, 0, 54, 21, 0, 30, 0, 0, 0, 0, 37, 65, 0, 
    0, 35, 0, 0, 36, 7, 0, 33, 0, 0, 0, 0, 25, 73, 0, 
    0, 17, 0, 0, 0, 5, 17, 0, 0, 0, 0, 19, 26, 34, 0, 
    8, 0, 7, 4, 0, 0, 7, 0, 0, 0, 0, 12, 33, 0, 37, 
    0, 20, 0, 9, 0, 9, 25, 0, 0, 0, 0, 18, 0, 19, 0, 
    0, 23, 0, 8, 0, 6, 1, 0, 0, 0, 9, 9, 0, 0, 11, 
    
    -- channel=384
    0, 0, 4, 3, 4, 2, 2, 0, 0, 4, 0, 0, 0, 0, 0, 
    4, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=385
    85, 82, 80, 81, 78, 70, 66, 65, 54, 48, 47, 40, 15, 16, 38, 
    70, 71, 66, 61, 56, 53, 51, 52, 49, 46, 38, 32, 25, 23, 39, 
    48, 44, 46, 47, 48, 47, 47, 50, 49, 48, 24, 16, 30, 36, 45, 
    41, 45, 46, 46, 48, 48, 45, 49, 51, 42, 21, 9, 35, 42, 42, 
    43, 45, 45, 45, 44, 44, 39, 34, 30, 28, 21, 18, 26, 38, 40, 
    45, 44, 45, 44, 36, 29, 31, 26, 12, 7, 7, 23, 11, 21, 36, 
    45, 45, 42, 37, 26, 4, 0, 0, 0, 0, 0, 15, 13, 5, 18, 
    44, 43, 35, 22, 12, 10, 10, 6, 26, 9, 0, 15, 10, 10, 9, 
    42, 32, 11, 2, 6, 0, 5, 0, 0, 0, 0, 15, 9, 13, 10, 
    37, 16, 19, 0, 9, 4, 0, 0, 0, 0, 0, 8, 7, 0, 0, 
    24, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    19, 0, 0, 11, 6, 0, 0, 0, 13, 0, 10, 0, 0, 5, 10, 
    18, 1, 0, 5, 0, 1, 0, 0, 12, 1, 10, 0, 0, 7, 7, 
    20, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 5, 9, 
    19, 6, 2, 7, 5, 4, 6, 6, 8, 3, 0, 8, 11, 11, 11, 
    
    -- channel=386
    21, 11, 9, 4, 2, 1, 3, 3, 1, 0, 8, 9, 2, 12, 13, 
    0, 0, 0, 0, 0, 0, 1, 2, 4, 9, 3, 2, 15, 17, 9, 
    0, 0, 0, 0, 2, 2, 3, 7, 8, 8, 5, 12, 17, 19, 10, 
    2, 3, 3, 3, 5, 4, 4, 4, 8, 6, 0, 14, 16, 6, 7, 
    5, 3, 2, 3, 3, 6, 7, 0, 0, 0, 3, 15, 4, 6, 7, 
    3, 2, 2, 3, 0, 0, 13, 24, 18, 18, 25, 0, 11, 7, 5, 
    2, 1, 2, 2, 3, 0, 0, 0, 0, 0, 0, 0, 3, 9, 8, 
    1, 0, 2, 0, 0, 13, 10, 6, 6, 11, 0, 1, 18, 13, 12, 
    0, 0, 0, 1, 9, 6, 8, 18, 0, 0, 0, 0, 0, 9, 8, 
    0, 4, 0, 7, 10, 18, 14, 0, 0, 0, 13, 12, 4, 0, 0, 
    0, 0, 5, 9, 14, 15, 1, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 12, 8, 18, 12, 4, 0, 0, 11, 11, 3, 2, 0, 17, 
    4, 7, 8, 3, 10, 2, 0, 0, 0, 15, 6, 7, 9, 6, 16, 
    8, 13, 14, 16, 7, 0, 0, 0, 9, 11, 1, 10, 8, 15, 18, 
    10, 3, 3, 12, 16, 15, 15, 14, 16, 11, 16, 17, 21, 21, 21, 
    
    -- channel=387
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 13, 13, 6, 36, 43, 0, 13, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 9, 25, 44, 28, 0, 0, 7, 1, 
    0, 0, 4, 9, 1, 15, 29, 31, 22, 21, 14, 0, 2, 20, 15, 
    0, 2, 0, 18, 0, 15, 40, 34, 28, 22, 6, 0, 19, 19, 12, 
    0, 19, 0, 8, 0, 18, 57, 30, 17, 0, 38, 43, 16, 15, 0, 
    0, 17, 15, 0, 9, 33, 44, 27, 0, 10, 6, 41, 20, 0, 0, 
    0, 15, 23, 4, 31, 28, 49, 31, 0, 16, 3, 16, 28, 0, 0, 
    0, 8, 16, 6, 28, 25, 25, 23, 0, 20, 6, 2, 17, 0, 2, 
    0, 2, 15, 11, 12, 12, 10, 8, 5, 21, 1, 0, 3, 3, 5, 
    
    -- channel=388
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=389
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 23, 11, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 17, 66, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 32, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 66, 41, 31, 15, 0, 0, 0, 23, 
    0, 9, 0, 0, 0, 0, 41, 48, 27, 27, 39, 0, 11, 12, 3, 
    0, 40, 0, 0, 0, 0, 43, 33, 12, 0, 14, 73, 12, 5, 0, 
    0, 0, 10, 0, 0, 25, 48, 27, 0, 0, 0, 34, 20, 0, 0, 
    0, 0, 21, 0, 6, 3, 48, 21, 0, 2, 0, 0, 43, 0, 0, 
    0, 0, 13, 0, 29, 33, 32, 28, 0, 15, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    
    -- channel=390
    12, 22, 13, 21, 25, 22, 14, 27, 13, 10, 17, 9, 21, 0, 16, 
    18, 23, 26, 23, 20, 21, 15, 20, 16, 18, 1, 25, 25, 0, 14, 
    17, 22, 19, 21, 15, 16, 15, 14, 14, 10, 0, 35, 16, 0, 19, 
    12, 13, 14, 17, 13, 13, 9, 11, 11, 8, 34, 0, 5, 11, 17, 
    11, 14, 15, 16, 9, 5, 1, 3, 0, 12, 32, 3, 10, 17, 12, 
    12, 16, 16, 16, 2, 0, 0, 3, 0, 10, 0, 100, 0, 18, 14, 
    14, 17, 19, 6, 0, 0, 0, 19, 0, 0, 0, 118, 29, 0, 12, 
    15, 18, 0, 7, 10, 0, 14, 0, 0, 0, 0, 77, 58, 0, 0, 
    17, 2, 10, 0, 26, 0, 0, 0, 0, 0, 15, 101, 0, 0, 0, 
    3, 0, 94, 0, 44, 0, 0, 0, 0, 10, 0, 42, 0, 0, 9, 
    0, 0, 52, 12, 25, 0, 0, 0, 22, 56, 0, 0, 14, 10, 62, 
    0, 4, 0, 46, 0, 0, 0, 0, 100, 0, 11, 0, 0, 67, 14, 
    0, 0, 0, 47, 0, 0, 0, 0, 103, 0, 25, 4, 0, 76, 0, 
    0, 0, 0, 18, 0, 0, 0, 0, 48, 0, 15, 32, 0, 19, 0, 
    1, 9, 0, 9, 2, 0, 2, 4, 6, 0, 12, 32, 2, 1, 0, 
    
    -- channel=391
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=392
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=393
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 31, 21, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 16, 41, 30, 19, 0, 0, 
    0, 0, 0, 0, 0, 0, 15, 23, 30, 59, 49, 26, 1, 8, 0, 
    0, 0, 0, 0, 15, 8, 13, 39, 44, 39, 43, 0, 0, 25, 26, 
    0, 0, 34, 18, 9, 6, 33, 43, 44, 36, 15, 31, 46, 38, 22, 
    0, 17, 23, 18, 2, 18, 45, 47, 38, 9, 17, 15, 42, 25, 5, 
    0, 18, 25, 17, 11, 31, 39, 50, 29, 13, 8, 20, 26, 25, 0, 
    0, 16, 30, 28, 35, 48, 54, 47, 30, 18, 20, 16, 14, 8, 0, 
    0, 6, 19, 15, 21, 11, 12, 10, 0, 16, 15, 9, 4, 0, 0, 
    0, 7, 19, 22, 21, 20, 17, 12, 6, 4, 9, 1, 2, 2, 2, 
    
    -- channel=394
    31, 39, 57, 57, 53, 45, 49, 35, 37, 35, 22, 17, 2, 6, 1, 
    50, 37, 37, 39, 37, 29, 31, 24, 20, 15, 14, 0, 0, 0, 2, 
    40, 34, 27, 22, 22, 15, 16, 15, 13, 13, 26, 0, 0, 0, 4, 
    14, 13, 11, 10, 12, 12, 10, 9, 10, 15, 0, 0, 0, 12, 10, 
    8, 11, 11, 12, 15, 20, 20, 14, 0, 0, 0, 0, 0, 8, 9, 
    10, 10, 10, 13, 18, 12, 6, 9, 44, 41, 0, 0, 24, 0, 4, 
    11, 10, 11, 15, 25, 31, 22, 1, 14, 23, 39, 0, 0, 20, 0, 
    11, 10, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 16, 0, 16, 0, 9, 13, 33, 15, 13, 0, 0, 0, 0, 0, 
    16, 20, 0, 0, 0, 7, 33, 25, 2, 18, 59, 0, 0, 0, 0, 
    47, 67, 0, 0, 0, 0, 13, 6, 0, 0, 25, 104, 0, 0, 0, 
    33, 0, 0, 0, 0, 11, 30, 0, 0, 0, 0, 39, 17, 0, 0, 
    16, 0, 9, 0, 0, 0, 5, 0, 0, 0, 0, 0, 58, 0, 0, 
    0, 10, 20, 0, 45, 66, 70, 66, 3, 17, 0, 0, 16, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 
    
    -- channel=395
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 3, 12, 24, 22, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 13, 21, 11, 18, 18, 46, 18, 0, 0, 
    0, 0, 0, 0, 0, 7, 9, 15, 17, 28, 34, 38, 23, 6, 4, 
    0, 0, 0, 17, 14, 12, 23, 18, 28, 34, 30, 34, 0, 24, 9, 
    0, 0, 30, 19, 22, 15, 23, 25, 42, 39, 26, 34, 24, 28, 28, 
    0, 0, 43, 20, 20, 14, 28, 34, 38, 32, 19, 25, 39, 36, 16, 
    0, 30, 21, 21, 16, 18, 31, 39, 33, 18, 20, 10, 32, 27, 16, 
    0, 17, 18, 33, 23, 29, 26, 42, 46, 15, 23, 20, 12, 31, 1, 
    0, 11, 18, 31, 19, 23, 26, 28, 32, 12, 21, 22, 3, 22, 5, 
    0, 6, 21, 26, 20, 20, 18, 16, 13, 7, 20, 17, 10, 9, 9, 
    
    -- channel=396
    38, 51, 59, 61, 57, 50, 48, 43, 31, 23, 18, 5, 0, 0, 2, 
    54, 43, 45, 43, 38, 31, 30, 27, 21, 16, 8, 0, 0, 0, 4, 
    30, 30, 29, 25, 22, 16, 16, 16, 13, 11, 0, 0, 0, 0, 3, 
    14, 12, 11, 12, 13, 12, 10, 9, 8, 0, 0, 0, 0, 7, 11, 
    7, 10, 11, 10, 11, 6, 4, 1, 0, 0, 0, 0, 4, 10, 9, 
    9, 10, 11, 12, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    10, 9, 8, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    9, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=397
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 9, 22, 10, 22, 3, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 8, 2, 0, 0, 
    0, 0, 0, 12, 3, 11, 26, 0, 8, 18, 0, 10, 0, 0, 0, 
    0, 0, 0, 8, 8, 11, 21, 12, 20, 18, 45, 0, 0, 3, 4, 
    0, 14, 20, 1, 10, 3, 9, 15, 3, 37, 13, 46, 20, 20, 21, 
    0, 7, 9, 4, 4, 2, 23, 13, 5, 2, 4, 17, 24, 6, 6, 
    0, 5, 11, 7, 0, 0, 0, 17, 4, 8, 0, 0, 18, 20, 0, 
    0, 0, 16, 27, 29, 44, 47, 48, 39, 8, 11, 2, 10, 14, 0, 
    0, 0, 6, 0, 3, 2, 0, 1, 0, 11, 8, 10, 1, 1, 1, 
    
    -- channel=398
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 18, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 8, 0, 0, 
    0, 0, 0, 0, 0, 21, 45, 69, 35, 14, 0, 0, 41, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 38, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 16, 0, 22, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    5, 31, 0, 9, 0, 0, 35, 0, 5, 3, 118, 18, 0, 0, 2, 
    12, 3, 0, 0, 0, 19, 0, 0, 0, 0, 0, 83, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 37, 33, 0, 16, 
    0, 3, 21, 1, 69, 74, 70, 68, 0, 15, 0, 10, 65, 0, 13, 
    0, 0, 0, 0, 0, 0, 1, 5, 8, 53, 0, 0, 8, 8, 4, 
    
    -- channel=399
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 15, 17, 22, 61, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 17, 51, 15, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 21, 20, 45, 43, 0, 3, 0, 16, 
    0, 0, 0, 3, 0, 0, 3, 62, 42, 45, 37, 0, 6, 20, 26, 
    0, 38, 0, 5, 0, 0, 32, 47, 41, 16, 38, 42, 35, 29, 13, 
    0, 12, 23, 0, 0, 14, 28, 43, 25, 0, 0, 44, 32, 16, 0, 
    0, 5, 33, 0, 0, 23, 48, 40, 0, 5, 0, 2, 42, 0, 0, 
    0, 11, 31, 0, 25, 34, 41, 36, 0, 13, 1, 0, 28, 0, 0, 
    0, 4, 10, 0, 8, 8, 10, 8, 0, 21, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    
    -- channel=400
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 29, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 29, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 23, 50, 41, 21, 2, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 9, 33, 8, 9, 0, 0, 11, 24, 23, 
    0, 3, 0, 0, 0, 0, 8, 15, 14, 0, 3, 26, 26, 15, 0, 
    0, 0, 0, 0, 0, 8, 21, 18, 0, 0, 0, 0, 4, 0, 0, 
    0, 0, 15, 0, 2, 10, 21, 21, 0, 0, 0, 0, 7, 0, 0, 
    0, 0, 14, 7, 25, 36, 25, 14, 2, 11, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 10, 6, 7, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=401
    0, 0, 0, 5, 8, 8, 6, 7, 8, 21, 9, 0, 3, 15, 0, 
    2, 0, 2, 8, 8, 6, 2, 4, 1, 0, 0, 0, 5, 0, 0, 
    13, 21, 13, 5, 1, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 15, 0, 1, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 14, 0, 0, 
    0, 0, 0, 0, 0, 18, 51, 65, 44, 0, 0, 0, 0, 12, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 9, 0, 0, 
    0, 0, 0, 16, 8, 14, 0, 0, 0, 0, 0, 36, 0, 0, 0, 
    0, 0, 0, 0, 15, 4, 0, 0, 0, 25, 38, 0, 0, 0, 8, 
    0, 30, 29, 0, 13, 0, 0, 0, 22, 74, 43, 48, 12, 27, 58, 
    1, 9, 0, 0, 0, 0, 0, 0, 11, 0, 0, 6, 12, 16, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 20, 38, 3, 
    0, 0, 19, 39, 49, 87, 99, 104, 78, 2, 14, 6, 21, 24, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 19, 16, 0, 0, 0, 
    
    -- channel=402
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 20, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 25, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 17, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 32, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 17, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 18, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 21, 25, 24, 0, 0, 36, 16, 11, 
    0, 0, 0, 0, 1, 4, 5, 28, 8, 0, 0, 0, 10, 36, 13, 
    0, 0, 2, 4, 6, 26, 14, 0, 0, 0, 0, 0, 19, 1, 0, 
    0, 0, 0, 23, 28, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 22, 41, 43, 4, 0, 0, 8, 25, 0, 0, 0, 0, 
    1, 19, 0, 23, 42, 15, 0, 0, 0, 29, 31, 22, 0, 0, 34, 
    15, 15, 0, 22, 24, 0, 0, 0, 0, 20, 17, 32, 0, 14, 39, 
    20, 11, 1, 12, 7, 0, 0, 0, 0, 20, 13, 34, 43, 44, 45, 
    12, 24, 39, 38, 43, 42, 42, 44, 45, 36, 14, 38, 50, 49, 44, 
    
    -- channel=403
    61, 73, 73, 79, 79, 78, 74, 74, 73, 60, 57, 55, 49, 25, 46, 
    84, 76, 79, 86, 83, 78, 73, 71, 66, 61, 57, 51, 25, 19, 54, 
    72, 78, 77, 78, 71, 67, 67, 61, 59, 58, 46, 22, 22, 27, 51, 
    64, 66, 66, 66, 64, 66, 65, 60, 53, 57, 38, 13, 31, 53, 58, 
    61, 69, 69, 69, 67, 61, 49, 57, 50, 40, 17, 10, 46, 57, 56, 
    67, 70, 68, 68, 68, 49, 8, 1, 5, 3, 0, 18, 20, 34, 54, 
    70, 69, 71, 66, 48, 36, 27, 30, 27, 15, 0, 0, 19, 19, 40, 
    69, 72, 61, 47, 28, 16, 14, 0, 0, 0, 0, 0, 15, 22, 0, 
    71, 71, 49, 17, 10, 17, 4, 0, 0, 0, 0, 26, 26, 3, 0, 
    76, 22, 15, 12, 18, 16, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    68, 18, 1, 10, 21, 9, 0, 0, 0, 29, 24, 0, 0, 0, 22, 
    66, 23, 0, 11, 13, 0, 0, 0, 0, 12, 11, 16, 0, 7, 17, 
    55, 17, 0, 12, 0, 0, 0, 0, 0, 3, 6, 20, 0, 18, 21, 
    41, 21, 3, 13, 11, 16, 18, 20, 16, 10, 13, 17, 19, 19, 19, 
    35, 33, 12, 5, 9, 8, 8, 13, 15, 14, 15, 20, 15, 15, 12, 
    
    -- channel=404
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 4, 4, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 11, 7, 3, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 0, 4, 2, 
    0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 23, 29, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 7, 0, 0, 
    0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 0, 
    0, 0, 22, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 15, 0, 0, 0, 0, 7, 0, 5, 0, 0, 9, 6, 
    0, 0, 0, 15, 0, 0, 0, 0, 17, 0, 11, 8, 0, 13, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 10, 6, 
    0, 2, 6, 18, 7, 8, 10, 11, 13, 0, 0, 12, 10, 10, 4, 
    
    -- channel=405
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=406
    35, 32, 23, 24, 20, 19, 17, 19, 18, 16, 17, 15, 8, 4, 18, 
    12, 13, 19, 15, 12, 13, 13, 14, 16, 15, 5, 10, 12, 19, 16, 
    12, 11, 11, 12, 14, 14, 15, 15, 17, 15, 0, 0, 10, 18, 17, 
    13, 15, 15, 15, 15, 15, 6, 9, 11, 13, 6, 14, 21, 21, 15, 
    15, 16, 15, 14, 12, 6, 3, 0, 0, 0, 0, 16, 5, 11, 15, 
    16, 14, 15, 14, 6, 0, 0, 0, 0, 0, 0, 42, 3, 1, 13, 
    14, 15, 14, 6, 0, 0, 0, 14, 1, 0, 0, 0, 32, 0, 7, 
    14, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 
    14, 0, 7, 0, 3, 4, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    2, 0, 3, 0, 18, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 9, 15, 0, 0, 0, 0, 1, 21, 0, 0, 0, 9, 
    4, 0, 0, 14, 1, 0, 0, 0, 0, 0, 7, 16, 0, 5, 9, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 12, 15, 
    10, 1, 3, 11, 13, 4, 0, 0, 0, 0, 0, 17, 17, 13, 15, 
    3, 0, 0, 1, 5, 2, 8, 10, 13, 15, 2, 13, 16, 16, 12, 
    
    -- channel=407
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 33, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 22, 31, 52, 64, 74, 0, 5, 0, 
    0, 0, 0, 0, 0, 6, 50, 33, 19, 0, 47, 153, 5, 3, 0, 
    0, 0, 0, 0, 24, 0, 30, 7, 0, 14, 79, 151, 44, 0, 0, 
    0, 0, 1, 7, 50, 0, 0, 34, 76, 83, 123, 89, 0, 0, 36, 
    0, 0, 92, 1, 29, 0, 0, 68, 71, 92, 47, 76, 42, 61, 73, 
    0, 32, 98, 31, 4, 0, 0, 70, 131, 55, 1, 0, 87, 79, 74, 
    0, 0, 58, 46, 0, 0, 0, 73, 163, 7, 18, 0, 45, 102, 0, 
    0, 5, 42, 36, 0, 35, 28, 72, 143, 0, 42, 0, 14, 64, 0, 
    0, 0, 33, 20, 7, 30, 35, 41, 74, 0, 42, 25, 0, 5, 0, 
    0, 6, 10, 21, 1, 4, 7, 5, 4, 0, 24, 12, 0, 0, 0, 
    
    -- channel=408
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 16, 27, 8, 19, 25, 0, 13, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 30, 20, 0, 1, 0, 
    0, 0, 0, 7, 8, 9, 18, 7, 25, 28, 24, 19, 0, 4, 10, 
    0, 0, 8, 17, 10, 10, 21, 28, 32, 39, 20, 0, 9, 21, 24, 
    0, 22, 9, 13, 3, 0, 32, 28, 31, 28, 35, 30, 29, 31, 19, 
    0, 14, 9, 11, 0, 16, 29, 29, 14, 5, 7, 32, 20, 20, 1, 
    0, 8, 14, 11, 7, 14, 29, 32, 13, 7, 7, 16, 19, 13, 0, 
    0, 6, 21, 20, 34, 40, 41, 42, 14, 12, 12, 7, 14, 4, 0, 
    0, 0, 8, 3, 5, 5, 6, 6, 3, 16, 7, 2, 0, 0, 0, 
    
    -- channel=409
    0, 8, 18, 22, 22, 20, 20, 16, 19, 24, 11, 7, 9, 16, 4, 
    13, 9, 20, 23, 21, 17, 17, 13, 11, 5, 0, 0, 0, 1, 3, 
    30, 30, 22, 16, 12, 9, 8, 4, 3, 0, 2, 0, 0, 0, 5, 
    13, 10, 8, 6, 6, 6, 0, 0, 0, 0, 7, 11, 10, 12, 8, 
    9, 9, 10, 9, 8, 4, 3, 0, 0, 0, 0, 0, 0, 6, 8, 
    9, 8, 8, 9, 0, 0, 0, 2, 51, 44, 0, 0, 21, 0, 7, 
    7, 10, 11, 2, 2, 32, 37, 41, 26, 0, 0, 0, 0, 26, 10, 
    10, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 
    12, 0, 0, 12, 12, 9, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 4, 12, 0, 0, 0, 56, 51, 0, 0, 0, 20, 
    14, 64, 1, 1, 0, 0, 0, 0, 35, 29, 42, 60, 15, 33, 42, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 7, 10, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 41, 14, 8, 
    0, 11, 39, 40, 69, 97, 103, 105, 55, 10, 3, 0, 27, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 24, 0, 0, 0, 0, 
    
    -- channel=410
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 11, 10, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 41, 53, 56, 58, 60, 10, 8, 0, 0, 
    0, 0, 0, 0, 1, 21, 18, 2, 0, 38, 101, 19, 8, 6, 0, 
    0, 0, 0, 4, 12, 16, 21, 20, 54, 92, 96, 54, 0, 8, 17, 
    0, 0, 5, 21, 19, 13, 43, 97, 97, 92, 71, 1, 17, 40, 70, 
    0, 35, 23, 23, 1, 12, 57, 91, 85, 79, 79, 54, 73, 68, 49, 
    0, 65, 19, 13, 0, 16, 70, 85, 57, 6, 19, 70, 68, 50, 9, 
    0, 14, 41, 11, 7, 43, 75, 90, 32, 9, 8, 42, 52, 23, 0, 
    0, 23, 48, 15, 42, 60, 87, 80, 23, 31, 17, 10, 43, 0, 0, 
    0, 18, 34, 16, 34, 36, 36, 34, 6, 23, 17, 0, 8, 0, 0, 
    0, 5, 14, 10, 11, 11, 9, 4, 0, 20, 10, 0, 0, 0, 1, 
    
    -- channel=411
    31, 31, 29, 30, 31, 33, 32, 32, 38, 31, 32, 35, 21, 8, 26, 
    35, 30, 29, 40, 40, 38, 36, 36, 35, 33, 35, 24, 15, 16, 31, 
    28, 34, 37, 40, 40, 38, 38, 35, 35, 35, 31, 0, 8, 19, 28, 
    38, 40, 39, 38, 38, 40, 37, 33, 29, 30, 15, 9, 18, 31, 34, 
    38, 41, 40, 40, 39, 33, 20, 25, 23, 13, 0, 0, 13, 28, 33, 
    41, 41, 39, 39, 43, 31, 0, 0, 0, 0, 0, 0, 11, 0, 29, 
    41, 40, 40, 41, 30, 7, 5, 3, 20, 28, 0, 0, 0, 15, 11, 
    39, 40, 38, 15, 0, 2, 0, 1, 0, 0, 0, 0, 0, 20, 3, 
    40, 46, 21, 5, 0, 10, 6, 0, 0, 0, 0, 0, 30, 0, 0, 
    52, 24, 0, 7, 0, 19, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    54, 0, 0, 0, 5, 21, 8, 0, 0, 0, 18, 16, 0, 0, 0, 
    56, 6, 0, 0, 15, 11, 0, 0, 0, 8, 3, 24, 0, 0, 5, 
    44, 13, 0, 0, 9, 0, 0, 0, 0, 8, 0, 6, 16, 0, 17, 
    33, 22, 0, 0, 6, 0, 0, 0, 0, 16, 0, 1, 25, 9, 18, 
    22, 18, 7, 0, 6, 6, 7, 10, 11, 24, 0, 1, 17, 15, 15, 
    
    -- channel=412
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 21, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 24, 25, 22, 13, 27, 22, 0, 9, 0, 
    0, 0, 0, 0, 0, 0, 9, 16, 3, 0, 20, 29, 3, 0, 2, 
    0, 0, 0, 19, 16, 13, 11, 8, 11, 27, 26, 19, 1, 0, 3, 
    0, 0, 1, 13, 11, 5, 3, 29, 28, 17, 32, 5, 0, 15, 11, 
    0, 15, 40, 12, 9, 13, 4, 29, 27, 33, 13, 48, 27, 24, 23, 
    0, 8, 38, 12, 9, 15, 19, 22, 35, 13, 14, 0, 36, 25, 7, 
    0, 12, 35, 16, 16, 20, 16, 30, 30, 15, 10, 0, 29, 22, 0, 
    0, 3, 20, 17, 19, 33, 36, 37, 44, 13, 28, 12, 15, 17, 2, 
    0, 0, 21, 13, 12, 13, 11, 10, 9, 7, 14, 10, 6, 4, 4, 
    
    -- channel=413
    61, 59, 59, 60, 59, 55, 52, 51, 42, 28, 29, 31, 13, 4, 28, 
    59, 59, 58, 58, 54, 50, 47, 45, 42, 38, 33, 23, 3, 15, 35, 
    40, 40, 46, 47, 43, 43, 43, 40, 40, 38, 18, 4, 14, 24, 34, 
    37, 42, 42, 43, 44, 44, 44, 44, 39, 34, 0, 0, 20, 30, 34, 
    41, 44, 44, 44, 44, 42, 31, 31, 29, 29, 10, 13, 31, 35, 34, 
    43, 45, 44, 42, 36, 27, 24, 15, 0, 0, 0, 18, 0, 27, 32, 
    44, 44, 44, 37, 26, 0, 0, 0, 0, 0, 0, 6, 3, 0, 21, 
    44, 44, 35, 29, 3, 0, 0, 0, 10, 0, 0, 0, 3, 0, 7, 
    44, 34, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 12, 0, 
    38, 20, 9, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=414
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 13, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 21, 13, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 42, 56, 40, 16, 0, 0, 5, 19, 
    0, 0, 0, 0, 0, 0, 14, 14, 1, 5, 8, 0, 15, 28, 12, 
    0, 10, 10, 8, 0, 0, 12, 13, 10, 0, 0, 13, 29, 14, 0, 
    0, 0, 0, 4, 0, 23, 30, 14, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 13, 3, 11, 18, 20, 13, 0, 9, 5, 3, 6, 0, 0, 
    0, 6, 15, 15, 35, 41, 30, 15, 1, 15, 14, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 5, 0, 0, 0, 0, 
    0, 5, 19, 19, 14, 15, 14, 10, 6, 0, 0, 0, 3, 2, 3, 
    
    -- channel=415
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 30, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 11, 45, 49, 57, 67, 94, 0, 9, 0, 
    0, 0, 0, 0, 0, 8, 29, 20, 0, 0, 19, 166, 4, 0, 0, 
    0, 0, 0, 4, 19, 0, 20, 5, 0, 25, 91, 140, 63, 0, 0, 
    0, 0, 2, 0, 29, 0, 0, 24, 89, 97, 117, 109, 0, 3, 29, 
    0, 0, 105, 0, 27, 0, 0, 54, 84, 96, 58, 113, 52, 65, 74, 
    0, 10, 95, 17, 2, 0, 0, 68, 111, 64, 0, 0, 93, 77, 63, 
    0, 14, 20, 37, 0, 0, 0, 84, 142, 0, 5, 0, 39, 84, 0, 
    0, 0, 7, 43, 0, 28, 19, 80, 140, 0, 36, 0, 0, 67, 0, 
    0, 0, 11, 25, 0, 12, 21, 29, 61, 0, 24, 13, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 13, 9, 0, 0, 0, 
    
    -- channel=416
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=417
    0, 3, 0, 3, 10, 7, 1, 13, 4, 3, 15, 7, 5, 0, 7, 
    5, 8, 7, 8, 7, 6, 2, 8, 5, 6, 2, 15, 23, 0, 7, 
    0, 11, 7, 7, 4, 6, 4, 5, 4, 2, 0, 14, 8, 0, 8, 
    6, 2, 2, 4, 2, 2, 3, 3, 2, 0, 30, 0, 0, 3, 11, 
    0, 2, 2, 3, 0, 0, 0, 2, 8, 27, 28, 0, 1, 7, 5, 
    2, 3, 3, 4, 0, 0, 0, 0, 0, 0, 0, 54, 0, 8, 4, 
    2, 4, 6, 1, 0, 0, 15, 26, 14, 0, 0, 101, 8, 0, 0, 
    2, 5, 0, 0, 6, 0, 13, 15, 0, 0, 0, 44, 36, 0, 0, 
    3, 0, 2, 0, 15, 0, 0, 0, 0, 0, 18, 91, 0, 0, 0, 
    0, 0, 57, 0, 27, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 
    0, 0, 47, 5, 17, 0, 0, 0, 13, 51, 0, 0, 0, 0, 46, 
    0, 0, 0, 30, 0, 0, 0, 0, 85, 0, 11, 0, 0, 51, 8, 
    0, 0, 0, 34, 0, 0, 0, 0, 84, 0, 20, 0, 0, 54, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 22, 23, 0, 17, 0, 
    0, 10, 11, 12, 0, 1, 3, 6, 7, 0, 0, 21, 1, 0, 0, 
    
    -- channel=418
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 
    1, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 53, 0, 0, 16, 0, 0, 
    0, 0, 0, 0, 0, 18, 35, 48, 29, 0, 0, 0, 0, 11, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 11, 0, 0, 
    0, 0, 0, 15, 13, 15, 3, 0, 0, 6, 0, 34, 0, 0, 0, 
    0, 0, 0, 0, 16, 0, 0, 0, 0, 16, 62, 0, 0, 0, 0, 
    0, 41, 28, 0, 14, 0, 0, 0, 0, 76, 16, 48, 16, 15, 66, 
    0, 0, 0, 1, 0, 0, 0, 0, 20, 0, 0, 3, 11, 18, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 13, 43, 0, 
    0, 0, 15, 38, 40, 76, 85, 90, 83, 0, 18, 2, 16, 21, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 18, 0, 0, 0, 
    
    -- channel=419
    0, 0, 1, 9, 11, 11, 9, 9, 12, 32, 10, 2, 11, 11, 0, 
    8, 0, 10, 13, 11, 8, 6, 6, 4, 0, 0, 1, 3, 0, 0, 
    16, 26, 13, 8, 4, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 12, 0, 5, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 8, 17, 0, 1, 
    0, 0, 0, 0, 0, 35, 59, 78, 43, 0, 0, 0, 9, 17, 5, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 
    0, 0, 16, 17, 20, 22, 0, 0, 0, 3, 11, 50, 0, 0, 0, 
    0, 0, 0, 4, 21, 3, 0, 0, 0, 40, 23, 0, 0, 0, 13, 
    0, 58, 0, 3, 11, 0, 0, 0, 26, 75, 63, 40, 15, 25, 70, 
    10, 4, 0, 10, 0, 0, 0, 0, 26, 0, 0, 29, 0, 34, 0, 
    4, 0, 0, 0, 0, 0, 0, 2, 9, 0, 0, 9, 17, 38, 5, 
    0, 0, 21, 30, 54, 89, 96, 102, 59, 0, 24, 14, 35, 16, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 10, 10, 0, 0, 0, 
    
    -- channel=420
    86, 86, 90, 90, 85, 79, 75, 70, 63, 44, 47, 35, 5, 11, 34, 
    84, 77, 78, 77, 72, 64, 63, 57, 53, 50, 38, 19, 0, 16, 41, 
    59, 60, 62, 61, 56, 54, 54, 51, 50, 48, 9, 0, 6, 29, 38, 
    50, 53, 53, 53, 55, 56, 55, 50, 47, 36, 0, 0, 34, 40, 44, 
    51, 55, 56, 55, 55, 48, 38, 41, 29, 12, 0, 0, 30, 42, 41, 
    54, 55, 54, 53, 47, 21, 0, 0, 0, 0, 0, 0, 0, 21, 36, 
    55, 56, 53, 46, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 
    55, 54, 33, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    55, 39, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=421
    28, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 3, 0, 20, 8, 
    0, 0, 0, 0, 0, 0, 0, 2, 5, 8, 0, 0, 26, 23, 3, 
    0, 0, 2, 4, 6, 6, 14, 18, 16, 7, 0, 0, 7, 0, 0, 
    5, 3, 2, 1, 2, 3, 0, 9, 46, 63, 43, 37, 6, 0, 0, 
    4, 4, 3, 0, 3, 24, 42, 14, 0, 0, 51, 62, 0, 11, 0, 
    4, 3, 0, 0, 0, 0, 0, 0, 0, 0, 2, 60, 36, 0, 0, 
    2, 1, 7, 24, 0, 5, 8, 87, 144, 125, 10, 0, 6, 14, 56, 
    0, 5, 0, 0, 0, 0, 0, 33, 0, 0, 0, 0, 31, 89, 32, 
    7, 58, 44, 0, 0, 0, 3, 0, 0, 0, 0, 59, 69, 14, 0, 
    0, 0, 0, 2, 0, 30, 41, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 17, 10, 3, 6, 0, 7, 4, 0, 0, 0, 0, 
    0, 0, 0, 32, 57, 75, 38, 0, 6, 10, 36, 7, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 7, 20, 44, 26, 27, 24, 16, 10, 0, 0, 0, 6, 7, 8, 
    
    -- channel=422
    21, 21, 22, 23, 20, 20, 19, 18, 17, 12, 17, 16, 15, 20, 18, 
    17, 16, 16, 14, 12, 13, 14, 14, 14, 15, 14, 14, 15, 26, 15, 
    15, 13, 14, 11, 12, 12, 12, 13, 14, 13, 8, 10, 16, 21, 13, 
    14, 12, 11, 12, 12, 11, 10, 12, 12, 13, 7, 27, 23, 18, 14, 
    12, 11, 11, 10, 10, 10, 10, 8, 6, 7, 8, 24, 17, 14, 15, 
    11, 10, 11, 11, 9, 1, 0, 0, 2, 0, 0, 27, 19, 15, 14, 
    9, 10, 10, 8, 8, 7, 13, 25, 22, 13, 0, 1, 28, 16, 17, 
    10, 9, 3, 8, 6, 16, 5, 7, 0, 7, 0, 0, 16, 16, 13, 
    9, 3, 14, 9, 13, 22, 11, 0, 0, 0, 0, 13, 0, 8, 0, 
    2, 0, 4, 17, 22, 22, 15, 0, 0, 7, 0, 0, 0, 0, 12, 
    8, 0, 6, 20, 24, 14, 16, 0, 11, 15, 33, 1, 0, 11, 13, 
    5, 18, 1, 16, 18, 13, 7, 0, 0, 19, 18, 22, 1, 11, 24, 
    7, 10, 1, 15, 8, 0, 4, 0, 7, 9, 13, 27, 9, 18, 25, 
    12, 10, 13, 21, 22, 19, 19, 18, 10, 17, 10, 23, 22, 26, 23, 
    11, 11, 14, 20, 19, 19, 20, 21, 22, 19, 18, 23, 24, 24, 23, 
    
    -- channel=423
    52, 58, 68, 69, 65, 58, 57, 50, 42, 39, 32, 20, 11, 10, 18, 
    63, 57, 56, 52, 47, 42, 42, 37, 33, 30, 26, 16, 0, 5, 19, 
    44, 40, 36, 35, 33, 30, 31, 30, 29, 28, 14, 6, 5, 15, 22, 
    26, 26, 26, 26, 28, 28, 27, 31, 30, 26, 7, 0, 12, 22, 24, 
    23, 25, 25, 26, 27, 29, 28, 29, 25, 19, 0, 1, 20, 25, 21, 
    23, 25, 26, 26, 24, 22, 15, 16, 18, 10, 0, 0, 7, 17, 18, 
    25, 25, 26, 24, 17, 16, 4, 0, 0, 0, 7, 0, 0, 4, 15, 
    25, 25, 20, 15, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 22, 10, 2, 0, 0, 0, 3, 5, 3, 0, 0, 0, 0, 1, 
    23, 13, 0, 0, 0, 0, 0, 4, 0, 2, 0, 0, 0, 0, 0, 
    20, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=424
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 30, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 9, 20, 24, 44, 66, 36, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 35, 24, 15, 0, 52, 101, 3, 0, 0, 
    0, 0, 0, 0, 17, 2, 24, 26, 25, 34, 73, 90, 30, 0, 9, 
    0, 0, 0, 19, 32, 8, 0, 45, 67, 77, 87, 53, 0, 9, 31, 
    0, 0, 58, 11, 20, 0, 0, 64, 72, 67, 53, 68, 43, 54, 53, 
    0, 22, 77, 23, 9, 4, 1, 68, 86, 45, 9, 25, 71, 62, 42, 
    0, 16, 50, 29, 3, 14, 25, 70, 96, 14, 18, 0, 52, 60, 4, 
    0, 13, 41, 34, 15, 45, 41, 71, 92, 9, 32, 2, 23, 41, 0, 
    0, 3, 26, 23, 13, 28, 34, 37, 53, 8, 32, 17, 1, 10, 0, 
    0, 5, 20, 23, 11, 13, 12, 9, 6, 0, 19, 12, 0, 0, 0, 
    
    -- channel=425
    47, 58, 58, 64, 62, 57, 52, 54, 43, 37, 38, 28, 16, 19, 26, 
    59, 56, 55, 52, 48, 44, 40, 41, 37, 34, 25, 27, 19, 7, 28, 
    40, 44, 42, 40, 37, 34, 33, 34, 32, 30, 1, 20, 21, 12, 27, 
    33, 32, 31, 32, 32, 31, 31, 31, 32, 24, 18, 12, 18, 28, 33, 
    28, 31, 32, 31, 30, 26, 22, 23, 21, 20, 17, 4, 26, 32, 30, 
    30, 31, 31, 32, 22, 11, 0, 0, 0, 0, 0, 36, 8, 22, 28, 
    31, 31, 30, 23, 7, 0, 2, 21, 7, 0, 0, 26, 12, 1, 22, 
    31, 30, 18, 13, 14, 2, 2, 0, 0, 0, 0, 17, 15, 0, 0, 
    30, 17, 12, 2, 5, 0, 0, 0, 0, 0, 0, 52, 0, 0, 0, 
    19, 0, 25, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 9, 0, 15, 0, 0, 0, 0, 30, 0, 0, 0, 0, 26, 
    5, 1, 0, 16, 0, 0, 0, 0, 27, 0, 8, 0, 0, 18, 14, 
    10, 0, 0, 15, 0, 0, 0, 0, 31, 0, 5, 1, 0, 31, 4, 
    9, 0, 0, 4, 0, 0, 0, 0, 21, 0, 4, 14, 0, 16, 4, 
    8, 2, 2, 1, 0, 0, 1, 3, 6, 0, 0, 17, 6, 5, 2, 
    
    -- channel=426
    105, 110, 117, 116, 113, 100, 97, 88, 79, 78, 62, 51, 25, 14, 35, 
    110, 103, 97, 95, 88, 77, 75, 70, 62, 56, 51, 35, 7, 8, 43, 
    83, 82, 74, 70, 64, 63, 63, 61, 58, 54, 60, 16, 7, 36, 52, 
    55, 56, 58, 58, 59, 64, 66, 65, 62, 59, 34, 0, 41, 54, 51, 
    52, 58, 60, 62, 62, 69, 68, 69, 63, 62, 14, 0, 40, 45, 46, 
    59, 60, 61, 60, 59, 60, 68, 68, 87, 87, 75, 1, 12, 37, 39, 
    61, 62, 63, 54, 60, 54, 65, 27, 27, 8, 104, 66, 0, 23, 20, 
    62, 63, 54, 44, 36, 20, 21, 1, 12, 53, 109, 97, 16, 0, 20, 
    63, 56, 33, 33, 20, 4, 4, 96, 116, 126, 123, 44, 25, 12, 62, 
    53, 78, 25, 4, 0, 0, 11, 105, 102, 104, 108, 71, 54, 71, 76, 
    55, 82, 58, 4, 0, 0, 11, 94, 106, 32, 20, 87, 89, 77, 37, 
    47, 12, 49, 0, 0, 14, 51, 93, 71, 1, 0, 3, 74, 37, 0, 
    26, 19, 43, 0, 0, 29, 64, 94, 56, 5, 8, 0, 53, 10, 0, 
    20, 23, 33, 12, 28, 60, 69, 73, 48, 16, 24, 0, 0, 0, 0, 
    23, 8, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 
    
    -- channel=427
    29, 28, 34, 34, 28, 30, 33, 23, 36, 13, 19, 19, 4, 18, 11, 
    37, 26, 25, 32, 32, 29, 30, 25, 25, 21, 28, 7, 0, 17, 15, 
    31, 26, 28, 28, 29, 26, 25, 24, 23, 25, 29, 0, 0, 16, 11, 
    24, 27, 26, 24, 27, 25, 26, 19, 20, 26, 0, 19, 9, 16, 16, 
    25, 27, 27, 26, 30, 27, 23, 23, 18, 0, 0, 1, 7, 15, 20, 
    27, 27, 25, 25, 37, 33, 14, 7, 17, 0, 0, 0, 28, 0, 16, 
    28, 26, 21, 31, 36, 29, 0, 0, 3, 72, 22, 0, 0, 11, 10, 
    28, 24, 36, 13, 0, 13, 0, 0, 0, 27, 0, 0, 0, 18, 8, 
    26, 39, 15, 13, 0, 19, 51, 30, 0, 0, 0, 0, 10, 19, 0, 
    43, 53, 0, 12, 0, 28, 86, 1, 0, 0, 11, 0, 0, 0, 0, 
    79, 31, 0, 0, 0, 28, 71, 0, 0, 0, 29, 75, 0, 0, 0, 
    51, 9, 0, 0, 13, 32, 56, 0, 0, 4, 0, 71, 2, 0, 0, 
    39, 14, 0, 0, 28, 0, 24, 0, 0, 21, 0, 9, 36, 0, 13, 
    23, 21, 3, 0, 33, 22, 21, 14, 0, 33, 0, 0, 16, 0, 10, 
    13, 3, 0, 0, 0, 0, 0, 0, 0, 29, 0, 0, 2, 3, 10, 
    
    -- channel=428
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 15, 23, 0, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 19, 22, 3, 0, 3, 18, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 44, 5, 0, 0, 
    0, 0, 0, 4, 9, 0, 0, 0, 25, 28, 31, 23, 0, 0, 0, 
    0, 0, 14, 1, 6, 0, 0, 18, 28, 49, 29, 2, 0, 14, 23, 
    0, 22, 23, 3, 0, 0, 0, 21, 43, 31, 16, 20, 36, 32, 27, 
    0, 2, 0, 5, 0, 0, 1, 23, 33, 0, 0, 0, 14, 26, 0, 
    0, 0, 0, 4, 0, 0, 2, 26, 31, 0, 0, 0, 5, 21, 0, 
    0, 0, 13, 21, 24, 40, 46, 49, 33, 0, 9, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    
    -- channel=429
    5, 11, 8, 13, 19, 15, 9, 20, 1, 10, 15, 2, 5, 3, 12, 
    11, 17, 16, 14, 13, 13, 9, 14, 9, 14, 3, 8, 29, 0, 11, 
    7, 15, 12, 13, 8, 11, 9, 10, 9, 5, 0, 35, 13, 0, 15, 
    10, 8, 8, 11, 8, 9, 11, 10, 7, 0, 29, 0, 8, 6, 14, 
    7, 8, 8, 10, 4, 1, 2, 7, 7, 21, 39, 0, 9, 13, 8, 
    7, 9, 10, 10, 0, 0, 0, 0, 0, 12, 33, 62, 0, 27, 8, 
    7, 10, 12, 3, 0, 0, 5, 11, 2, 0, 0, 150, 0, 0, 10, 
    8, 11, 0, 0, 15, 0, 19, 22, 0, 0, 0, 74, 69, 0, 0, 
    9, 0, 0, 0, 23, 0, 0, 0, 0, 0, 33, 102, 0, 0, 0, 
    0, 0, 80, 0, 33, 0, 0, 0, 0, 0, 0, 65, 0, 0, 5, 
    0, 0, 81, 9, 20, 0, 0, 0, 25, 56, 0, 0, 17, 11, 56, 
    0, 0, 6, 39, 0, 0, 0, 0, 114, 0, 12, 0, 0, 64, 16, 
    0, 0, 0, 44, 0, 0, 0, 0, 113, 0, 31, 0, 0, 72, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 62, 0, 22, 22, 0, 20, 0, 
    0, 8, 8, 14, 1, 2, 2, 4, 5, 0, 10, 30, 0, 0, 0, 
    
    -- channel=430
    36, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 7, 
    0, 4, 0, 0, 0, 0, 0, 0, 0, 4, 10, 5, 1, 9, 9, 
    0, 0, 0, 0, 0, 2, 4, 6, 11, 12, 17, 0, 16, 21, 13, 
    0, 2, 5, 6, 8, 9, 14, 21, 19, 17, 0, 0, 8, 0, 0, 
    6, 5, 4, 5, 6, 14, 8, 9, 32, 51, 36, 16, 1, 0, 2, 
    7, 6, 5, 3, 7, 27, 59, 39, 0, 0, 84, 29, 0, 10, 0, 
    6, 5, 6, 5, 14, 0, 0, 0, 0, 0, 18, 75, 6, 0, 0, 
    3, 6, 16, 24, 0, 3, 12, 69, 115, 105, 20, 0, 20, 7, 51, 
    4, 13, 0, 0, 0, 0, 0, 58, 5, 0, 2, 0, 29, 69, 39, 
    13, 73, 34, 0, 0, 0, 0, 0, 0, 0, 0, 80, 64, 17, 0, 
    0, 0, 0, 0, 0, 25, 13, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 2, 14, 10, 4, 16, 4, 4, 3, 0, 0, 0, 0, 
    0, 0, 5, 17, 44, 63, 26, 0, 18, 11, 31, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 7, 9, 33, 16, 18, 14, 8, 3, 0, 0, 0, 3, 3, 5, 
    
    -- channel=431
    15, 11, 12, 10, 8, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 8, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 6, 10, 15, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 22, 26, 28, 32, 53, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 58, 56, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 15, 44, 73, 51, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 59, 72, 79, 78, 20, 0, 5, 33, 
    0, 27, 11, 0, 0, 0, 0, 60, 65, 53, 51, 57, 37, 42, 35, 
    0, 16, 27, 0, 0, 0, 1, 58, 55, 0, 0, 24, 53, 34, 0, 
    0, 0, 14, 0, 0, 0, 26, 62, 38, 0, 0, 0, 34, 10, 0, 
    0, 0, 10, 0, 0, 24, 39, 60, 34, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 8, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=432
    10, 20, 30, 31, 28, 23, 24, 17, 18, 26, 14, 1, 4, 15, 0, 
    27, 21, 20, 15, 14, 10, 11, 8, 5, 3, 0, 3, 0, 0, 0, 
    23, 22, 12, 6, 5, 2, 1, 3, 0, 0, 9, 11, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 1, 1, 4, 4, 15, 15, 4, 4, 2, 
    0, 0, 0, 0, 0, 4, 14, 14, 11, 5, 0, 0, 5, 2, 0, 
    0, 0, 0, 0, 1, 7, 14, 33, 64, 74, 29, 0, 19, 5, 0, 
    0, 0, 0, 0, 9, 47, 61, 48, 32, 28, 81, 15, 0, 16, 4, 
    0, 0, 0, 2, 21, 13, 13, 0, 0, 24, 84, 69, 0, 0, 0, 
    0, 0, 16, 33, 22, 21, 26, 60, 96, 104, 93, 33, 0, 0, 36, 
    0, 12, 7, 14, 2, 3, 34, 88, 87, 96, 99, 25, 27, 55, 62, 
    9, 81, 38, 7, 0, 0, 30, 79, 83, 51, 49, 98, 76, 70, 47, 
    8, 13, 30, 0, 0, 18, 56, 77, 45, 3, 0, 35, 60, 33, 0, 
    2, 13, 34, 0, 0, 14, 57, 82, 31, 8, 0, 2, 55, 16, 0, 
    0, 11, 37, 28, 54, 86, 96, 98, 50, 22, 24, 0, 16, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 14, 0, 0, 0, 0, 
    
    -- channel=433
    41, 28, 21, 16, 13, 9, 9, 9, 1, 0, 0, 10, 0, 0, 4, 
    21, 25, 13, 3, 3, 3, 3, 4, 4, 6, 20, 12, 0, 6, 10, 
    0, 0, 0, 0, 1, 5, 7, 10, 12, 16, 20, 14, 24, 20, 9, 
    0, 3, 6, 8, 9, 12, 23, 28, 28, 23, 0, 0, 2, 2, 3, 
    6, 6, 5, 6, 10, 21, 22, 34, 70, 85, 55, 27, 20, 6, 4, 
    6, 7, 7, 6, 12, 57, 93, 73, 23, 18, 110, 50, 0, 22, 3, 
    8, 7, 5, 9, 26, 0, 0, 0, 0, 21, 87, 99, 12, 0, 0, 
    6, 8, 32, 43, 23, 21, 29, 88, 157, 140, 94, 40, 9, 8, 64, 
    4, 20, 9, 1, 0, 0, 33, 102, 78, 77, 63, 25, 51, 93, 82, 
    18, 101, 60, 3, 0, 0, 20, 66, 70, 21, 21, 118, 105, 69, 28, 
    9, 0, 19, 2, 0, 29, 53, 70, 21, 0, 0, 0, 39, 14, 0, 
    0, 4, 35, 14, 13, 22, 52, 82, 45, 5, 10, 0, 26, 11, 0, 
    0, 9, 30, 37, 65, 99, 79, 69, 52, 26, 42, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 11, 26, 35, 18, 20, 15, 7, 1, 0, 0, 0, 0, 0, 1, 
    
    -- channel=434
    10, 7, 10, 6, 4, 3, 5, 2, 1, 0, 0, 0, 12, 1, 2, 
    3, 6, 10, 4, 4, 3, 5, 1, 1, 1, 0, 4, 0, 3, 3, 
    12, 0, 0, 2, 0, 0, 0, 0, 1, 1, 14, 18, 3, 10, 6, 
    0, 0, 0, 0, 2, 1, 2, 0, 3, 6, 0, 0, 0, 0, 0, 
    3, 1, 1, 1, 3, 11, 13, 0, 0, 0, 0, 24, 17, 6, 2, 
    1, 1, 1, 1, 0, 0, 45, 89, 80, 46, 27, 15, 0, 21, 3, 
    1, 2, 2, 0, 18, 8, 0, 0, 0, 0, 11, 15, 4, 5, 14, 
    2, 0, 1, 22, 0, 10, 0, 0, 0, 43, 9, 36, 10, 0, 1, 
    2, 0, 0, 0, 11, 0, 0, 50, 34, 2, 0, 0, 0, 10, 29, 
    0, 13, 21, 0, 0, 2, 7, 5, 2, 40, 25, 36, 38, 15, 16, 
    4, 25, 0, 7, 0, 0, 0, 4, 18, 0, 0, 0, 15, 10, 0, 
    0, 0, 2, 5, 0, 10, 0, 16, 9, 0, 0, 0, 0, 6, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 4, 1, 3, 3, 0, 0, 2, 
    0, 3, 15, 9, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    8, 0, 0, 2, 4, 2, 0, 0, 0, 0, 17, 0, 0, 0, 0, 
    
    -- channel=435
    24, 25, 23, 23, 24, 22, 20, 24, 18, 8, 18, 12, 18, 5, 18, 
    20, 23, 23, 19, 18, 18, 17, 19, 18, 19, 13, 23, 15, 6, 17, 
    14, 13, 14, 17, 16, 16, 17, 19, 18, 17, 1, 14, 20, 13, 20, 
    14, 14, 14, 16, 15, 15, 14, 19, 19, 15, 19, 0, 9, 13, 16, 
    13, 13, 13, 13, 11, 10, 10, 11, 16, 29, 21, 13, 17, 18, 15, 
    12, 13, 15, 14, 10, 2, 0, 0, 0, 0, 0, 46, 0, 18, 15, 
    13, 13, 14, 11, 0, 0, 0, 0, 0, 0, 0, 45, 25, 0, 12, 
    11, 14, 4, 12, 6, 0, 12, 19, 15, 0, 0, 9, 15, 8, 7, 
    12, 9, 12, 0, 13, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 
    9, 0, 37, 0, 16, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 4, 11, 12, 1, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    1, 0, 0, 22, 6, 0, 0, 0, 31, 6, 10, 0, 0, 22, 7, 
    2, 0, 0, 19, 0, 1, 0, 0, 31, 0, 18, 6, 0, 16, 7, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 20, 0, 9, 11, 
    7, 11, 10, 21, 13, 13, 15, 14, 16, 0, 1, 14, 15, 15, 11, 
    
    -- channel=436
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 20, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 6, 3, 0, 0, 29, 17, 0, 0, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 8, 19, 0, 0, 0, 
    0, 0, 27, 0, 4, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 
    0, 0, 25, 2, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 6, 
    0, 0, 11, 12, 0, 0, 0, 0, 46, 0, 3, 0, 0, 22, 0, 
    0, 0, 0, 8, 0, 5, 0, 0, 42, 0, 14, 0, 0, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 3, 4, 0, 0, 0, 
    0, 0, 0, 8, 0, 1, 2, 2, 1, 0, 0, 2, 0, 0, 0, 
    
    -- channel=437
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 26, 22, 13, 34, 43, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 6, 16, 14, 26, 38, 28, 0, 0, 0, 1, 
    0, 0, 0, 2, 0, 0, 23, 42, 34, 21, 26, 0, 0, 13, 8, 
    0, 26, 0, 0, 0, 0, 32, 34, 19, 17, 37, 64, 20, 16, 0, 
    0, 0, 6, 0, 0, 10, 38, 25, 0, 0, 0, 29, 26, 0, 0, 
    0, 0, 16, 0, 4, 7, 38, 37, 0, 0, 0, 0, 30, 0, 0, 
    0, 0, 7, 0, 27, 44, 47, 47, 1, 11, 2, 0, 8, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    
    -- channel=438
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 16, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 2, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 39, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 104, 0, 8, 0, 
    0, 0, 0, 0, 0, 0, 10, 15, 0, 0, 0, 146, 21, 0, 0, 
    0, 0, 0, 0, 15, 0, 19, 0, 0, 0, 0, 111, 40, 0, 0, 
    0, 0, 3, 0, 37, 0, 0, 0, 0, 0, 41, 101, 0, 0, 0, 
    0, 0, 103, 0, 37, 0, 0, 0, 0, 14, 0, 35, 0, 1, 17, 
    0, 0, 63, 17, 12, 0, 0, 0, 56, 42, 0, 0, 18, 19, 64, 
    0, 0, 6, 55, 0, 0, 0, 0, 150, 0, 16, 0, 0, 92, 0, 
    0, 0, 0, 44, 0, 0, 0, 0, 135, 0, 38, 0, 0, 71, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 46, 0, 24, 31, 0, 7, 0, 
    0, 8, 7, 21, 3, 3, 6, 7, 9, 0, 4, 21, 0, 0, 0, 
    
    -- channel=439
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 16, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 5, 26, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 17, 24, 16, 0, 0, 48, 2, 3, 0, 
    0, 0, 0, 0, 11, 1, 7, 0, 0, 0, 0, 39, 28, 0, 0, 
    0, 0, 1, 9, 15, 5, 0, 0, 0, 4, 10, 38, 0, 0, 0, 
    0, 0, 26, 0, 21, 2, 0, 0, 5, 14, 9, 15, 0, 0, 15, 
    0, 0, 42, 10, 19, 0, 0, 0, 26, 39, 3, 0, 14, 22, 32, 
    0, 11, 6, 18, 3, 0, 0, 0, 46, 5, 13, 0, 9, 28, 15, 
    0, 0, 0, 17, 0, 0, 0, 5, 49, 0, 12, 2, 0, 39, 1, 
    0, 0, 7, 22, 3, 16, 20, 23, 44, 0, 13, 18, 3, 23, 5, 
    0, 2, 6, 9, 4, 4, 5, 7, 9, 0, 13, 22, 9, 8, 6, 
    
    -- channel=440
    0, 0, 0, 1, 2, 2, 2, 0, 0, 22, 0, 0, 5, 17, 0, 
    0, 0, 0, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 16, 6, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 10, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 33, 58, 0, 0, 31, 0, 0, 
    0, 0, 0, 0, 0, 27, 43, 54, 34, 0, 0, 0, 0, 27, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 
    0, 0, 0, 22, 13, 19, 0, 0, 0, 1, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 8, 9, 0, 0, 0, 40, 70, 0, 0, 0, 6, 
    0, 64, 14, 0, 8, 0, 0, 0, 12, 60, 36, 75, 14, 26, 57, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 13, 10, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 29, 5, 
    0, 2, 30, 43, 62, 103, 114, 117, 79, 3, 12, 0, 25, 18, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 21, 10, 0, 0, 0, 
    
    -- channel=441
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=442
    61, 67, 74, 78, 72, 69, 69, 61, 60, 34, 40, 42, 9, 31, 31, 
    79, 66, 64, 68, 65, 59, 57, 53, 49, 45, 47, 15, 2, 26, 34, 
    57, 56, 60, 54, 52, 48, 47, 44, 44, 48, 22, 9, 10, 24, 27, 
    46, 48, 47, 46, 48, 47, 47, 41, 40, 42, 0, 25, 29, 35, 39, 
    43, 48, 48, 47, 52, 47, 38, 43, 38, 0, 0, 12, 26, 37, 39, 
    47, 48, 46, 46, 54, 44, 16, 11, 12, 11, 0, 0, 37, 13, 34, 
    48, 47, 43, 52, 36, 16, 0, 0, 5, 65, 0, 0, 0, 11, 28, 
    49, 47, 53, 20, 0, 20, 0, 0, 0, 0, 0, 0, 0, 18, 5, 
    47, 56, 6, 15, 0, 15, 54, 0, 0, 0, 0, 0, 12, 12, 0, 
    67, 35, 0, 5, 0, 23, 68, 0, 0, 0, 24, 0, 0, 0, 0, 
    81, 0, 0, 0, 7, 19, 35, 0, 0, 0, 4, 50, 0, 0, 0, 
    43, 14, 0, 0, 14, 0, 35, 0, 0, 2, 0, 39, 0, 0, 16, 
    37, 5, 0, 0, 10, 0, 0, 0, 0, 12, 0, 4, 4, 0, 15, 
    22, 9, 0, 7, 9, 10, 13, 11, 0, 14, 0, 0, 0, 9, 10, 
    19, 2, 0, 0, 0, 0, 0, 0, 0, 11, 0, 3, 3, 5, 9, 
    
    -- channel=443
    81, 89, 97, 98, 98, 91, 88, 83, 75, 70, 62, 49, 24, 36, 49, 
    93, 86, 90, 92, 87, 79, 78, 73, 67, 61, 50, 31, 23, 30, 54, 
    76, 84, 81, 76, 71, 69, 69, 65, 61, 55, 21, 15, 18, 38, 54, 
    67, 66, 65, 64, 65, 66, 63, 58, 54, 45, 20, 21, 49, 58, 60, 
    63, 66, 67, 66, 65, 56, 49, 48, 34, 22, 0, 0, 45, 54, 56, 
    67, 67, 66, 65, 55, 29, 0, 0, 0, 4, 0, 0, 18, 44, 51, 
    66, 67, 67, 56, 29, 20, 34, 37, 35, 0, 0, 14, 0, 27, 40, 
    67, 66, 39, 19, 19, 4, 0, 0, 0, 0, 0, 13, 24, 0, 4, 
    68, 48, 15, 12, 7, 7, 0, 0, 0, 0, 5, 38, 10, 0, 0, 
    49, 0, 0, 0, 11, 0, 0, 0, 0, 0, 2, 0, 0, 0, 6, 
    30, 0, 22, 4, 12, 0, 0, 0, 14, 37, 15, 4, 0, 10, 34, 
    33, 2, 1, 3, 0, 0, 0, 0, 20, 3, 5, 0, 5, 15, 18, 
    27, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 7, 24, 14, 
    26, 4, 4, 9, 7, 28, 32, 36, 42, 3, 13, 9, 13, 19, 8, 
    22, 6, 0, 0, 0, 0, 0, 0, 3, 0, 11, 14, 3, 3, 0, 
    
    -- channel=444
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 21, 32, 42, 43, 30, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 21, 6, 1, 0, 66, 22, 0, 9, 0, 
    0, 0, 0, 0, 4, 2, 8, 0, 5, 41, 60, 56, 0, 0, 0, 
    0, 0, 0, 11, 16, 2, 2, 59, 65, 61, 60, 6, 3, 5, 41, 
    0, 9, 16, 8, 0, 0, 14, 61, 55, 66, 55, 29, 38, 43, 38, 
    0, 52, 21, 8, 0, 0, 20, 56, 58, 5, 12, 47, 51, 41, 16, 
    0, 0, 31, 5, 0, 20, 31, 57, 40, 0, 0, 11, 34, 27, 0, 
    0, 9, 33, 1, 7, 26, 48, 50, 29, 9, 6, 0, 31, 3, 0, 
    0, 8, 26, 9, 24, 34, 37, 36, 17, 9, 14, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 9, 0, 0, 0, 0, 
    
    -- channel=445
    97, 101, 97, 101, 98, 92, 85, 87, 71, 71, 63, 51, 29, 24, 48, 
    96, 92, 89, 87, 82, 77, 72, 72, 66, 65, 53, 46, 32, 19, 53, 
    68, 71, 71, 73, 69, 67, 67, 67, 64, 62, 28, 28, 34, 36, 55, 
    61, 65, 65, 67, 65, 67, 65, 65, 64, 52, 36, 14, 40, 56, 60, 
    59, 66, 67, 66, 64, 59, 49, 52, 48, 36, 32, 14, 36, 55, 55, 
    64, 67, 66, 65, 57, 42, 18, 8, 0, 11, 0, 31, 14, 25, 51, 
    67, 67, 64, 57, 31, 11, 4, 11, 5, 0, 0, 30, 16, 7, 29, 
    66, 66, 54, 28, 18, 10, 18, 7, 8, 0, 0, 26, 16, 17, 0, 
    64, 56, 26, 7, 10, 0, 5, 0, 0, 0, 0, 54, 18, 2, 0, 
    65, 2, 31, 0, 20, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 
    32, 0, 7, 0, 17, 0, 0, 0, 0, 22, 0, 0, 0, 0, 24, 
    34, 7, 0, 19, 3, 0, 0, 0, 28, 0, 11, 0, 0, 18, 18, 
    30, 2, 0, 19, 0, 0, 0, 0, 29, 0, 8, 0, 0, 29, 7, 
    26, 9, 0, 0, 0, 0, 0, 0, 19, 0, 12, 18, 0, 16, 7, 
    25, 16, 7, 2, 2, 0, 3, 5, 9, 0, 0, 17, 9, 8, 7, 
    
    -- channel=446
    115, 120, 129, 129, 126, 116, 112, 103, 93, 75, 67, 56, 29, 22, 51, 
    125, 117, 118, 117, 110, 99, 96, 87, 79, 71, 60, 40, 5, 23, 60, 
    99, 98, 97, 92, 85, 82, 83, 76, 73, 70, 47, 16, 13, 45, 64, 
    75, 78, 79, 79, 80, 83, 82, 78, 73, 65, 17, 0, 52, 65, 66, 
    75, 82, 83, 83, 84, 81, 71, 72, 56, 46, 0, 8, 54, 62, 62, 
    81, 83, 82, 80, 74, 51, 46, 51, 57, 43, 19, 5, 7, 49, 57, 
    83, 84, 83, 72, 58, 39, 27, 7, 7, 0, 31, 34, 0, 18, 37, 
    84, 84, 60, 47, 18, 11, 2, 0, 0, 11, 33, 48, 13, 0, 8, 
    85, 67, 28, 10, 6, 0, 0, 33, 46, 45, 53, 25, 14, 0, 24, 
    71, 46, 11, 0, 0, 0, 0, 32, 32, 49, 40, 31, 19, 23, 34, 
    60, 39, 17, 0, 0, 0, 0, 26, 46, 4, 0, 22, 33, 28, 16, 
    49, 0, 6, 0, 0, 0, 1, 28, 28, 0, 0, 0, 18, 15, 0, 
    32, 1, 3, 0, 0, 0, 10, 25, 21, 0, 0, 0, 10, 1, 0, 
    26, 9, 6, 0, 2, 19, 25, 27, 17, 0, 3, 0, 0, 0, 0, 
    28, 2, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    
    -- channel=447
    18, 0, 7, 0, 0, 0, 1, 0, 4, 0, 0, 0, 0, 5, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 7, 0, 0, 34, 0, 
    0, 0, 0, 0, 0, 0, 1, 1, 2, 5, 19, 0, 0, 26, 0, 
    1, 3, 3, 0, 6, 4, 6, 5, 5, 7, 0, 16, 9, 0, 0, 
    7, 4, 3, 0, 7, 9, 11, 5, 14, 0, 0, 18, 0, 0, 0, 
    5, 2, 1, 0, 12, 25, 36, 11, 11, 0, 6, 0, 16, 0, 0, 
    4, 1, 0, 6, 29, 6, 0, 0, 0, 71, 74, 0, 0, 6, 0, 
    3, 0, 10, 9, 0, 13, 0, 14, 60, 104, 8, 0, 0, 10, 40, 
    1, 8, 0, 0, 0, 11, 46, 91, 9, 0, 0, 0, 21, 51, 36, 
    10, 81, 0, 17, 0, 28, 94, 29, 0, 0, 0, 0, 29, 1, 0, 
    54, 12, 0, 0, 0, 39, 111, 10, 0, 0, 33, 71, 0, 0, 0, 
    22, 0, 6, 0, 14, 63, 83, 1, 0, 7, 0, 82, 4, 0, 0, 
    13, 11, 23, 0, 58, 30, 75, 0, 0, 31, 0, 12, 51, 0, 13, 
    12, 16, 7, 0, 27, 0, 0, 0, 0, 44, 0, 0, 17, 0, 9, 
    6, 0, 0, 0, 4, 5, 3, 0, 0, 40, 0, 0, 2, 4, 12, 
    
    -- channel=448
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=449
    10, 10, 9, 10, 16, 23, 22, 14, 13, 13, 13, 13, 13, 12, 14, 
    10, 11, 10, 15, 25, 32, 34, 33, 20, 15, 19, 20, 23, 21, 20, 
    10, 11, 14, 13, 30, 38, 42, 46, 39, 24, 22, 22, 19, 14, 15, 
    12, 12, 16, 24, 34, 39, 43, 49, 44, 34, 27, 26, 17, 19, 23, 
    19, 22, 24, 28, 37, 35, 41, 47, 51, 50, 44, 39, 27, 28, 29, 
    12, 10, 18, 26, 32, 34, 39, 41, 45, 50, 51, 43, 34, 26, 25, 
    5, 6, 15, 19, 24, 25, 39, 45, 41, 42, 50, 47, 35, 21, 17, 
    10, 12, 15, 28, 31, 29, 38, 44, 41, 41, 48, 47, 38, 27, 24, 
    13, 11, 19, 30, 25, 26, 28, 45, 39, 39, 45, 50, 43, 34, 24, 
    19, 14, 12, 16, 23, 31, 30, 42, 41, 39, 44, 50, 42, 32, 26, 
    1, 3, 6, 12, 22, 31, 28, 33, 40, 40, 38, 45, 44, 34, 32, 
    0, 0, 9, 20, 27, 34, 37, 25, 27, 36, 36, 42, 43, 32, 32, 
    7, 6, 10, 17, 30, 33, 29, 34, 35, 36, 34, 40, 41, 33, 31, 
    14, 19, 21, 20, 21, 26, 29, 35, 35, 29, 27, 35, 40, 35, 29, 
    19, 18, 24, 29, 27, 27, 29, 33, 34, 33, 31, 31, 35, 33, 29, 
    
    -- channel=450
    15, 14, 13, 14, 20, 24, 19, 19, 17, 18, 18, 18, 19, 18, 17, 
    15, 15, 15, 14, 29, 32, 37, 30, 20, 18, 17, 19, 21, 20, 19, 
    15, 16, 15, 25, 31, 38, 38, 39, 34, 25, 21, 19, 15, 13, 13, 
    17, 15, 11, 21, 38, 35, 36, 39, 33, 29, 29, 19, 12, 14, 18, 
    15, 18, 19, 25, 37, 41, 38, 37, 41, 40, 39, 34, 19, 16, 18, 
    9, 5, 9, 15, 32, 33, 29, 38, 37, 38, 39, 36, 22, 13, 10, 
    3, 2, 8, 7, 17, 33, 39, 40, 35, 34, 40, 40, 26, 13, 8, 
    8, 7, 8, 22, 20, 16, 26, 36, 38, 36, 40, 40, 33, 19, 15, 
    8, 1, 1, 0, 23, 13, 26, 31, 34, 35, 39, 42, 38, 26, 14, 
    4, 2, 0, 15, 15, 21, 23, 33, 36, 36, 38, 42, 37, 17, 13, 
    0, 0, 0, 1, 22, 29, 30, 28, 37, 36, 33, 36, 32, 23, 14, 
    0, 0, 7, 20, 15, 32, 32, 16, 25, 32, 32, 33, 26, 20, 15, 
    6, 9, 7, 14, 27, 30, 28, 29, 38, 38, 32, 34, 32, 17, 20, 
    12, 17, 19, 15, 11, 19, 20, 27, 30, 25, 28, 32, 27, 19, 15, 
    17, 13, 14, 15, 16, 18, 20, 18, 19, 22, 23, 21, 20, 16, 14, 
    
    -- channel=451
    9, 8, 9, 6, 2, 0, 2, 2, 4, 4, 3, 3, 2, 4, 2, 
    9, 7, 8, 5, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 
    9, 7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 7, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 10, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 9, 3, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 9, 5, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 12, 8, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 14, 11, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 11, 0, 8, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 9, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    8, 7, 5, 1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    4, 2, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=452
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=453
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 28, 26, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=454
    0, 0, 0, 0, 0, 0, 3, 0, 3, 0, 3, 6, 5, 0, 5, 
    0, 1, 0, 4, 0, 0, 3, 1, 3, 0, 1, 0, 0, 0, 4, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 8, 
    0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 6, 6, 
    0, 0, 16, 38, 0, 0, 0, 12, 0, 0, 0, 0, 0, 4, 3, 
    0, 0, 28, 37, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 59, 0, 0, 8, 0, 0, 4, 3, 0, 0, 0, 12, 
    0, 0, 0, 10, 48, 0, 5, 0, 0, 7, 6, 0, 0, 0, 3, 
    0, 0, 0, 20, 0, 21, 0, 12, 0, 0, 3, 3, 0, 0, 15, 
    0, 0, 0, 42, 0, 20, 0, 22, 0, 0, 0, 9, 0, 16, 8, 
    0, 0, 72, 0, 0, 2, 0, 0, 0, 0, 1, 5, 0, 2, 16, 
    8, 6, 23, 11, 23, 0, 0, 23, 0, 0, 0, 4, 12, 0, 26, 
    0, 0, 0, 0, 15, 13, 0, 9, 0, 0, 0, 3, 18, 0, 0, 
    0, 0, 0, 9, 2, 0, 4, 0, 0, 0, 0, 1, 4, 8, 0, 
    5, 8, 4, 8, 0, 0, 6, 13, 8, 1, 0, 0, 9, 3, 5, 
    
    -- channel=455
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=456
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=457
    13, 12, 9, 10, 0, 0, 2, 5, 8, 6, 5, 5, 4, 4, 4, 
    13, 12, 8, 3, 0, 0, 0, 0, 0, 3, 1, 1, 2, 3, 3, 
    11, 10, 3, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 
    9, 10, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 18, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 16, 11, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 13, 10, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 12, 10, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 17, 20, 16, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28, 31, 25, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 26, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 10, 4, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 9, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=458
    0, 0, 0, 0, 6, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 25, 10, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 10, 15, 23, 21, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 14, 11, 12, 22, 22, 28, 11, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 26, 8, 2, 23, 22, 30, 15, 0, 0, 0, 
    1, 6, 0, 0, 0, 22, 13, 10, 19, 17, 22, 28, 16, 7, 1, 
    11, 7, 0, 0, 16, 40, 16, 19, 20, 7, 17, 28, 15, 20, 2, 
    2, 0, 0, 0, 0, 0, 0, 22, 25, 5, 11, 19, 21, 6, 0, 
    2, 0, 0, 0, 0, 0, 13, 4, 27, 11, 9, 12, 23, 6, 5, 
    0, 0, 19, 0, 32, 5, 24, 3, 23, 16, 13, 9, 18, 0, 0, 
    13, 11, 0, 36, 33, 35, 28, 27, 26, 22, 19, 12, 8, 0, 0, 
    40, 32, 0, 0, 0, 21, 19, 0, 30, 23, 13, 4, 0, 20, 0, 
    11, 9, 3, 0, 0, 0, 25, 0, 13, 23, 8, 9, 0, 10, 14, 
    0, 1, 9, 12, 12, 5, 0, 11, 15, 29, 39, 14, 10, 8, 18, 
    6, 11, 8, 0, 9, 16, 2, 1, 4, 6, 16, 19, 7, 7, 9, 
    
    -- channel=459
    17, 17, 14, 15, 7, 5, 10, 12, 14, 13, 13, 13, 12, 10, 11, 
    17, 17, 12, 13, 2, 0, 0, 0, 8, 8, 8, 9, 9, 7, 8, 
    16, 15, 13, 7, 0, 0, 0, 0, 0, 5, 6, 4, 6, 6, 5, 
    14, 12, 11, 3, 0, 0, 0, 0, 0, 0, 0, 0, 5, 6, 1, 
    15, 15, 12, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 16, 15, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 17, 16, 19, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    16, 15, 14, 12, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    13, 12, 17, 22, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 20, 21, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 27, 24, 8, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 21, 32, 8, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 14, 12, 11, 8, 2, 0, 1, 0, 0, 1, 0, 0, 0, 0, 
    11, 8, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=460
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 13, 12, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 8, 8, 10, 14, 10, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 9, 18, 16, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 8, 15, 18, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 6, 0, 3, 15, 12, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 12, 14, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 12, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 4, 0, 0, 
    0, 0, 0, 0, 0, 6, 0, 2, 0, 0, 1, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 0, 0, 3, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=461
    6, 6, 5, 4, 3, 0, 0, 4, 3, 2, 4, 4, 3, 1, 0, 
    6, 4, 2, 9, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    7, 6, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 5, 5, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 1, 7, 13, 6, 7, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    21, 28, 13, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 9, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=462
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 24, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 26, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 7, 0, 6, 19, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 23, 0, 0, 0, 0, 4, 
    0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 12, 6, 0, 0, 0, 
    
    -- channel=463
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 10, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 12, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 10, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 10, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 19, 22, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 36, 17, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    37, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 8, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=464
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 15, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=465
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 37, 35, 22, 24, 8, 8, 0, 0, 0, 0, 0, 0, 0, 
    48, 57, 18, 0, 0, 1, 0, 0, 3, 0, 0, 0, 0, 0, 0, 
    21, 11, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 18, 16, 0, 0, 0, 0, 6, 14, 0, 0, 0, 0, 
    6, 19, 11, 0, 0, 0, 0, 0, 0, 0, 0, 8, 7, 0, 0, 
    
    -- channel=466
    0, 0, 0, 0, 0, 0, 0, 2, 7, 9, 15, 20, 26, 29, 31, 
    0, 0, 0, 3, 0, 0, 0, 0, 10, 11, 16, 15, 14, 11, 10, 
    1, 1, 4, 4, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    4, 4, 13, 16, 8, 9, 3, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 3, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 6, 
    0, 0, 0, 0, 0, 6, 0, 5, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 7, 5, 0, 0, 1, 5, 7, 8, 1, 3, 6, 4, 
    
    -- channel=467
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 5, 6, 9, 9, 
    0, 0, 0, 1, 0, 0, 0, 0, 2, 1, 2, 1, 0, 2, 4, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 8, 11, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 6, 7, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 14, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 25, 
    0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 21, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 12, 
    0, 0, 0, 9, 16, 7, 5, 0, 0, 0, 0, 0, 0, 15, 20, 
    5, 15, 16, 19, 22, 13, 7, 14, 19, 11, 6, 3, 9, 21, 28, 
    
    -- channel=468
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 11, 6, 10, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 2, 0, 0, 10, 2, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 3, 0, 0, 3, 0, 5, 5, 0, 0, 0, 0, 
    0, 0, 0, 27, 0, 0, 0, 0, 0, 4, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 11, 2, 3, 0, 0, 0, 5, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 3, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 6, 0, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 1, 0, 4, 
    0, 0, 0, 0, 15, 3, 0, 17, 0, 0, 0, 1, 3, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=469
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=470
    0, 0, 0, 0, 5, 2, 10, 4, 3, 4, 8, 10, 11, 9, 9, 
    0, 0, 0, 10, 10, 18, 11, 18, 13, 3, 6, 4, 4, 3, 4, 
    1, 0, 11, 7, 18, 23, 27, 25, 11, 2, 0, 1, 4, 1, 5, 
    1, 0, 0, 25, 22, 21, 22, 24, 26, 13, 8, 11, 0, 4, 7, 
    0, 0, 0, 21, 26, 4, 9, 25, 24, 28, 26, 13, 4, 4, 5, 
    0, 0, 0, 23, 6, 12, 20, 19, 15, 23, 26, 19, 12, 0, 0, 
    0, 0, 0, 4, 17, 7, 12, 19, 12, 18, 22, 27, 15, 0, 1, 
    0, 0, 0, 0, 0, 12, 11, 17, 9, 14, 23, 27, 13, 10, 4, 
    0, 0, 0, 4, 0, 0, 0, 22, 13, 12, 18, 24, 19, 20, 14, 
    0, 0, 0, 0, 0, 0, 8, 17, 14, 14, 15, 25, 25, 19, 9, 
    0, 0, 6, 0, 13, 14, 20, 10, 12, 17, 15, 19, 24, 4, 18, 
    0, 0, 0, 0, 17, 20, 3, 22, 12, 14, 8, 12, 24, 8, 9, 
    0, 0, 0, 0, 0, 13, 12, 9, 19, 11, 3, 17, 16, 18, 1, 
    0, 2, 9, 13, 10, 1, 14, 16, 21, 22, 6, 15, 20, 15, 14, 
    11, 12, 11, 15, 13, 5, 13, 16, 16, 15, 20, 17, 15, 17, 13, 
    
    -- channel=471
    28, 27, 18, 29, 26, 27, 29, 24, 23, 21, 17, 16, 11, 3, 7, 
    28, 30, 24, 11, 29, 14, 30, 23, 16, 17, 13, 11, 9, 9, 13, 
    25, 27, 28, 8, 22, 13, 13, 10, 3, 20, 22, 23, 18, 21, 20, 
    22, 21, 35, 3, 12, 11, 6, 7, 10, 15, 24, 29, 17, 21, 14, 
    19, 27, 77, 20, 6, 6, 24, 23, 14, 13, 12, 21, 13, 16, 12, 
    41, 49, 97, 16, 17, 2, 31, 30, 17, 15, 16, 9, 5, 15, 19, 
    46, 48, 56, 61, 8, 5, 37, 21, 20, 25, 24, 0, 16, 13, 25, 
    40, 40, 54, 40, 63, 0, 31, 11, 22, 39, 26, 14, 20, 10, 15, 
    39, 39, 59, 51, 68, 66, 33, 27, 21, 37, 29, 26, 10, 11, 18, 
    52, 66, 80, 124, 49, 92, 18, 38, 23, 30, 31, 32, 12, 17, 0, 
    86, 105, 97, 63, 36, 44, 20, 14, 23, 25, 30, 28, 10, 11, 3, 
    92, 78, 56, 49, 43, 8, 8, 25, 11, 12, 20, 32, 13, 0, 21, 
    43, 36, 32, 27, 36, 19, 11, 30, 11, 3, 40, 35, 25, 0, 6, 
    23, 21, 28, 23, 6, 14, 4, 18, 7, 5, 25, 29, 23, 0, 0, 
    22, 15, 6, 0, 0, 5, 12, 5, 0, 1, 0, 5, 9, 0, 0, 
    
    -- channel=472
    4, 4, 4, 5, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 
    4, 3, 1, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 2, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 8, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 4, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 1, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 6, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 17, 19, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 22, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 7, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=473
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 10, 0, 0, 0, 0, 0, 0, 0, 6, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 14, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 5, 16, 16, 11, 2, 2, 0, 0, 0, 0, 0, 0, 0, 
    54, 40, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 20, 9, 0, 0, 0, 0, 10, 9, 0, 0, 2, 5, 
    14, 18, 7, 0, 0, 0, 0, 1, 0, 0, 2, 11, 4, 3, 3, 
    
    -- channel=474
    30, 27, 29, 31, 27, 21, 22, 21, 20, 18, 14, 11, 8, 7, 5, 
    29, 26, 26, 23, 20, 19, 15, 13, 14, 16, 13, 13, 15, 17, 16, 
    26, 25, 19, 14, 11, 6, 6, 3, 14, 26, 26, 22, 20, 18, 12, 
    23, 24, 11, 13, 5, 3, 3, 6, 5, 18, 23, 16, 16, 16, 10, 
    39, 49, 36, 8, 7, 19, 20, 9, 4, 5, 11, 12, 17, 14, 13, 
    56, 57, 37, 13, 9, 26, 23, 9, 8, 5, 2, 9, 14, 14, 14, 
    52, 49, 47, 8, 17, 23, 14, 12, 17, 12, 6, 9, 9, 15, 13, 
    48, 51, 49, 44, 19, 23, 15, 15, 24, 19, 8, 4, 8, 12, 11, 
    55, 61, 65, 54, 44, 25, 25, 18, 23, 21, 13, 7, 13, 11, 1, 
    85, 93, 92, 53, 55, 32, 34, 12, 22, 23, 19, 10, 8, 0, 0, 
    96, 87, 38, 31, 24, 19, 11, 14, 20, 19, 15, 6, 3, 2, 0, 
    69, 50, 31, 34, 12, 6, 15, 8, 11, 14, 20, 13, 0, 9, 0, 
    33, 33, 30, 29, 24, 15, 19, 9, 17, 25, 31, 21, 0, 0, 5, 
    24, 26, 22, 10, 3, 8, 10, 9, 6, 13, 22, 13, 3, 0, 1, 
    16, 5, 0, 0, 0, 8, 3, 0, 0, 0, 2, 2, 0, 0, 0, 
    
    -- channel=475
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 3, 5, 11, 3, 0, 0, 6, 3, 0, 0, 0, 9, 13, 
    
    -- channel=476
    10, 9, 7, 8, 1, 1, 1, 6, 7, 7, 6, 7, 7, 5, 5, 
    10, 10, 7, 2, 0, 0, 0, 0, 1, 5, 1, 0, 0, 0, 0, 
    10, 11, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 8, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 9, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 4, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 3, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 12, 3, 21, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 28, 16, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 10, 9, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=477
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 
    0, 0, 0, 4, 4, 0, 0, 3, 5, 0, 0, 0, 0, 7, 7, 
    
    -- channel=478
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 4, 4, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 9, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=479
    19, 20, 12, 21, 17, 17, 21, 15, 13, 9, 7, 5, 0, 0, 0, 
    19, 20, 11, 12, 13, 0, 17, 11, 7, 5, 3, 4, 4, 6, 10, 
    15, 15, 15, 2, 2, 0, 0, 0, 1, 16, 19, 18, 16, 17, 14, 
    11, 11, 25, 0, 0, 0, 0, 0, 0, 0, 17, 23, 13, 18, 11, 
    17, 28, 62, 25, 0, 0, 6, 8, 0, 0, 0, 9, 9, 19, 15, 
    44, 52, 77, 24, 0, 0, 12, 13, 0, 0, 0, 0, 0, 18, 21, 
    47, 49, 53, 73, 0, 0, 19, 0, 0, 8, 0, 0, 6, 5, 21, 
    40, 43, 55, 49, 64, 0, 16, 0, 1, 20, 5, 0, 0, 0, 13, 
    42, 45, 65, 77, 64, 63, 19, 19, 0, 16, 8, 1, 0, 5, 13, 
    70, 87, 99, 127, 38, 68, 8, 33, 1, 10, 11, 10, 0, 9, 0, 
    103, 114, 118, 33, 23, 22, 5, 1, 2, 7, 9, 6, 0, 3, 5, 
    95, 74, 67, 37, 26, 0, 0, 17, 0, 0, 2, 13, 4, 0, 25, 
    39, 31, 28, 26, 33, 17, 0, 17, 0, 0, 20, 18, 18, 0, 0, 
    17, 18, 23, 18, 5, 5, 0, 0, 0, 0, 1, 11, 6, 0, 0, 
    17, 9, 1, 0, 0, 0, 10, 4, 0, 0, 0, 0, 1, 0, 0, 
    
    -- channel=480
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=481
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 2, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 2, 3, 0, 3, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 4, 1, 0, 0, 
    0, 0, 6, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 30, 9, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 1, 0, 0, 7, 
    0, 0, 0, 20, 0, 22, 0, 8, 0, 0, 0, 3, 0, 17, 7, 
    0, 0, 44, 6, 0, 0, 0, 0, 0, 0, 0, 6, 1, 5, 7, 
    0, 7, 10, 0, 12, 0, 0, 10, 0, 0, 0, 2, 8, 0, 18, 
    0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 13, 0, 0, 
    0, 0, 0, 1, 3, 0, 0, 0, 0, 0, 0, 0, 3, 4, 0, 
    0, 2, 5, 4, 0, 0, 0, 7, 2, 0, 0, 0, 7, 0, 0, 
    
    -- channel=482
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 8, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 14, 6, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 9, 6, 2, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 37, 28, 18, 28, 8, 19, 0, 0, 2, 0, 0, 0, 0, 
    50, 56, 16, 0, 0, 8, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    18, 14, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 18, 17, 0, 0, 0, 5, 9, 22, 7, 0, 1, 0, 
    6, 19, 11, 0, 0, 0, 0, 2, 0, 0, 1, 10, 10, 0, 0, 
    
    -- channel=483
    0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 11, 0, 4, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    1, 0, 8, 3, 4, 0, 4, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 3, 0, 0, 0, 0, 3, 8, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 4, 0, 0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 4, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 8, 0, 15, 0, 1, 0, 0, 0, 0, 0, 0, 8, 0, 
    0, 2, 62, 47, 26, 31, 10, 11, 0, 0, 1, 0, 0, 0, 0, 
    57, 65, 6, 0, 5, 8, 0, 1, 11, 0, 0, 0, 2, 0, 0, 
    22, 16, 11, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 
    2, 0, 5, 22, 20, 0, 0, 0, 0, 12, 16, 0, 3, 3, 4, 
    9, 22, 12, 2, 0, 0, 0, 3, 0, 0, 4, 9, 6, 2, 2, 
    
    -- channel=484
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 
    0, 0, 1, 5, 8, 1, 0, 5, 7, 2, 0, 0, 1, 11, 11, 
    
    -- channel=485
    0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 5, 12, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 5, 17, 27, 33, 32, 26, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 26, 19, 13, 3, 0, 0, 
    0, 5, 25, 14, 0, 7, 11, 4, 0, 0, 0, 0, 0, 5, 9, 
    47, 56, 37, 14, 1, 0, 20, 16, 0, 0, 0, 0, 8, 17, 19, 
    14, 0, 0, 21, 18, 17, 0, 0, 4, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 49, 0, 0, 0, 0, 4, 10, 1, 0, 0, 0, 0, 
    1, 9, 4, 1, 62, 44, 20, 5, 1, 7, 4, 1, 0, 0, 8, 
    14, 27, 59, 65, 23, 32, 4, 15, 0, 0, 9, 6, 0, 0, 0, 
    66, 42, 0, 0, 0, 0, 0, 4, 0, 0, 6, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 11, 15, 
    0, 0, 0, 0, 2, 0, 0, 16, 0, 0, 7, 11, 4, 0, 13, 
    0, 0, 0, 0, 6, 23, 0, 0, 7, 6, 11, 0, 11, 0, 0, 
    0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=486
    19, 20, 18, 18, 26, 26, 24, 20, 21, 22, 22, 22, 23, 22, 21, 
    19, 20, 20, 24, 31, 36, 32, 30, 23, 21, 22, 21, 19, 18, 18, 
    21, 20, 23, 30, 38, 43, 46, 44, 28, 20, 20, 19, 19, 18, 19, 
    21, 20, 19, 35, 44, 46, 47, 45, 42, 30, 27, 24, 17, 18, 20, 
    14, 11, 15, 33, 44, 36, 37, 46, 46, 46, 43, 32, 19, 18, 19, 
    10, 10, 6, 32, 34, 37, 40, 46, 44, 47, 48, 42, 28, 17, 17, 
    11, 11, 7, 25, 34, 35, 40, 43, 38, 43, 45, 47, 35, 19, 17, 
    13, 11, 14, 7, 14, 31, 35, 41, 37, 41, 46, 49, 37, 26, 20, 
    11, 6, 1, 22, 12, 23, 23, 39, 40, 41, 45, 47, 40, 33, 23, 
    0, 0, 2, 8, 18, 12, 27, 39, 41, 42, 43, 47, 44, 32, 21, 
    0, 0, 20, 26, 40, 35, 43, 37, 40, 42, 41, 46, 41, 23, 20, 
    8, 10, 18, 17, 37, 46, 32, 36, 42, 42, 38, 39, 36, 22, 21, 
    20, 18, 17, 19, 17, 30, 31, 32, 39, 39, 33, 40, 35, 28, 18, 
    20, 21, 24, 25, 23, 21, 28, 32, 38, 41, 34, 42, 38, 26, 24, 
    23, 24, 24, 25, 23, 20, 28, 27, 26, 29, 33, 33, 30, 27, 22, 
    
    -- channel=487
    1, 1, 1, 2, 12, 12, 5, 1, 1, 1, 0, 0, 0, 0, 0, 
    1, 1, 3, 6, 16, 22, 18, 12, 3, 3, 2, 1, 0, 0, 0, 
    2, 1, 4, 8, 21, 26, 31, 29, 11, 7, 7, 7, 5, 4, 4, 
    2, 2, 0, 13, 24, 29, 31, 35, 31, 19, 15, 13, 5, 4, 6, 
    2, 3, 6, 13, 23, 25, 28, 34, 38, 34, 31, 20, 11, 10, 11, 
    8, 10, 7, 10, 18, 26, 30, 31, 35, 39, 39, 30, 19, 16, 14, 
    8, 8, 7, 1, 19, 26, 28, 31, 29, 32, 37, 34, 23, 17, 11, 
    7, 8, 10, 8, 6, 16, 27, 33, 30, 29, 35, 34, 25, 15, 7, 
    10, 10, 9, 14, 15, 14, 21, 32, 31, 29, 33, 34, 28, 16, 13, 
    8, 11, 16, 13, 26, 19, 28, 31, 30, 29, 33, 34, 27, 15, 10, 
    12, 13, 12, 24, 22, 30, 26, 29, 31, 29, 32, 32, 24, 13, 11, 
    13, 12, 3, 13, 23, 27, 20, 19, 29, 28, 27, 29, 22, 19, 12, 
    5, 5, 6, 7, 9, 16, 23, 16, 24, 26, 25, 28, 21, 20, 17, 
    6, 7, 11, 12, 12, 11, 17, 22, 23, 24, 25, 27, 24, 20, 19, 
    9, 12, 13, 12, 14, 17, 16, 17, 18, 17, 20, 20, 18, 17, 16, 
    
    -- channel=488
    31, 29, 23, 28, 27, 29, 27, 25, 23, 22, 19, 17, 13, 9, 10, 
    30, 31, 25, 18, 27, 19, 28, 21, 17, 19, 15, 14, 12, 11, 13, 
    28, 29, 23, 16, 23, 18, 17, 16, 14, 21, 21, 20, 16, 17, 14, 
    25, 25, 29, 8, 21, 20, 16, 11, 11, 19, 25, 22, 16, 16, 10, 
    29, 33, 51, 20, 16, 21, 28, 23, 17, 16, 17, 22, 12, 10, 6, 
    40, 46, 68, 19, 23, 16, 33, 33, 23, 18, 19, 17, 7, 8, 11, 
    44, 44, 49, 43, 12, 17, 36, 25, 25, 27, 24, 12, 15, 11, 17, 
    41, 41, 45, 37, 41, 8, 27, 18, 30, 38, 27, 19, 22, 12, 13, 
    41, 43, 58, 46, 55, 45, 30, 24, 30, 39, 32, 28, 19, 12, 3, 
    56, 61, 63, 89, 42, 61, 20, 34, 32, 36, 35, 32, 19, 10, 0, 
    75, 81, 67, 52, 37, 37, 26, 22, 29, 30, 29, 31, 15, 6, 0, 
    69, 64, 54, 40, 35, 21, 21, 20, 21, 24, 29, 31, 8, 0, 7, 
    41, 34, 31, 26, 31, 17, 11, 30, 20, 21, 42, 33, 17, 0, 1, 
    25, 21, 20, 13, 3, 10, 7, 15, 12, 13, 31, 33, 18, 0, 0, 
    14, 7, 1, 0, 0, 1, 7, 0, 0, 0, 0, 3, 2, 0, 0, 
    
    -- channel=489
    0, 3, 0, 1, 7, 10, 11, 5, 4, 4, 6, 7, 7, 4, 7, 
    1, 2, 0, 13, 11, 16, 19, 18, 12, 5, 8, 6, 5, 1, 4, 
    2, 2, 8, 5, 22, 25, 27, 29, 16, 2, 5, 6, 6, 6, 10, 
    3, 1, 12, 14, 23, 25, 28, 29, 27, 17, 11, 17, 8, 8, 10, 
    0, 0, 1, 27, 21, 11, 17, 33, 32, 31, 26, 22, 11, 12, 11, 
    0, 0, 9, 27, 15, 7, 25, 30, 27, 33, 32, 25, 18, 12, 13, 
    0, 0, 2, 23, 10, 9, 24, 26, 19, 28, 33, 27, 23, 11, 14, 
    0, 0, 0, 10, 15, 9, 21, 22, 17, 25, 32, 30, 21, 17, 13, 
    0, 0, 0, 14, 0, 12, 7, 28, 19, 24, 29, 32, 23, 21, 18, 
    0, 0, 0, 7, 8, 15, 13, 32, 20, 22, 25, 33, 27, 28, 19, 
    0, 0, 33, 19, 18, 28, 23, 25, 20, 24, 25, 32, 29, 17, 21, 
    0, 9, 14, 5, 25, 25, 14, 22, 17, 23, 18, 25, 32, 13, 24, 
    7, 1, 6, 5, 12, 12, 8, 23, 16, 14, 12, 26, 31, 20, 15, 
    7, 4, 9, 16, 17, 11, 17, 18, 19, 14, 14, 24, 29, 26, 15, 
    10, 16, 19, 20, 16, 9, 18, 25, 21, 19, 17, 19, 24, 22, 19, 
    
    -- channel=490
    26, 23, 28, 31, 30, 33, 27, 23, 16, 14, 10, 4, 0, 0, 0, 
    25, 23, 27, 13, 26, 27, 30, 21, 16, 13, 9, 8, 6, 10, 11, 
    23, 23, 22, 12, 15, 12, 16, 22, 24, 27, 28, 33, 30, 31, 25, 
    19, 20, 15, 0, 3, 8, 10, 20, 28, 41, 38, 37, 34, 27, 22, 
    28, 39, 54, 0, 2, 20, 25, 16, 24, 24, 31, 37, 38, 38, 36, 
    68, 76, 74, 0, 9, 18, 29, 23, 24, 20, 24, 27, 42, 54, 49, 
    72, 72, 69, 23, 19, 29, 33, 24, 30, 22, 22, 18, 38, 50, 41, 
    62, 67, 74, 59, 29, 9, 29, 26, 35, 29, 19, 17, 30, 27, 30, 
    69, 78, 85, 57, 83, 62, 54, 27, 33, 30, 22, 17, 20, 26, 38, 
    96, 116, 124, 118, 77, 87, 44, 35, 30, 29, 29, 20, 16, 24, 24, 
    139, 141, 79, 75, 51, 49, 35, 32, 33, 33, 32, 22, 18, 32, 21, 
    122, 103, 66, 45, 18, 7, 26, 10, 19, 22, 28, 27, 23, 38, 34, 
    57, 49, 47, 43, 37, 14, 27, 27, 10, 19, 39, 30, 29, 32, 43, 
    35, 37, 42, 41, 35, 37, 16, 26, 19, 25, 40, 26, 30, 31, 36, 
    35, 34, 31, 24, 23, 39, 32, 29, 24, 22, 19, 29, 29, 26, 30, 
    
    -- channel=491
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 4, 6, 0, 0, 
    0, 0, 0, 0, 2, 15, 0, 0, 0, 0, 0, 6, 0, 7, 0, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 5, 0, 0, 0, 0, 15, 0, 
    0, 0, 0, 0, 0, 0, 7, 0, 0, 9, 0, 0, 0, 8, 5, 
    0, 0, 0, 0, 4, 0, 1, 0, 0, 10, 0, 0, 0, 2, 15, 
    0, 0, 0, 0, 18, 9, 0, 0, 5, 2, 9, 2, 0, 8, 10, 
    
    -- channel=492
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 24, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 25, 28, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    39, 31, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=493
    0, 1, 0, 0, 0, 2, 1, 2, 4, 1, 3, 5, 4, 0, 7, 
    0, 4, 0, 0, 0, 0, 8, 1, 1, 4, 4, 5, 3, 1, 6, 
    0, 1, 1, 0, 2, 0, 0, 0, 0, 0, 2, 2, 0, 4, 7, 
    0, 0, 29, 0, 0, 0, 0, 0, 0, 0, 0, 6, 4, 7, 8, 
    0, 0, 29, 26, 0, 0, 0, 8, 0, 0, 0, 0, 0, 8, 5, 
    0, 0, 53, 17, 9, 0, 0, 12, 0, 2, 0, 0, 0, 3, 6, 
    0, 0, 14, 62, 0, 0, 14, 0, 0, 6, 7, 0, 0, 0, 9, 
    0, 0, 0, 16, 58, 0, 11, 0, 0, 12, 8, 0, 0, 0, 7, 
    0, 0, 13, 5, 25, 30, 8, 4, 0, 7, 8, 6, 0, 0, 12, 
    0, 0, 0, 64, 0, 42, 0, 21, 0, 0, 4, 11, 0, 17, 9, 
    0, 8, 53, 1, 0, 5, 0, 0, 0, 0, 5, 11, 0, 12, 9, 
    2, 12, 31, 19, 23, 0, 0, 15, 0, 0, 0, 12, 8, 0, 29, 
    2, 0, 1, 0, 23, 12, 0, 17, 0, 0, 2, 4, 22, 0, 3, 
    0, 0, 0, 5, 3, 5, 0, 1, 0, 0, 0, 7, 6, 7, 0, 
    1, 6, 7, 7, 0, 0, 6, 13, 5, 3, 0, 0, 14, 0, 2, 
    
    -- channel=494
    3, 1, 0, 0, 0, 5, 4, 1, 4, 2, 0, 0, 0, 4, 9, 
    2, 4, 0, 0, 1, 0, 4, 7, 2, 5, 14, 23, 30, 31, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 21, 31, 21, 18, 9, 0, 0, 
    2, 6, 21, 0, 0, 5, 8, 5, 0, 0, 3, 0, 5, 7, 11, 
    43, 55, 49, 4, 2, 11, 26, 11, 5, 2, 0, 7, 13, 19, 22, 
    21, 8, 17, 3, 19, 14, 0, 3, 10, 7, 6, 0, 1, 9, 7, 
    0, 0, 10, 37, 0, 0, 1, 6, 13, 9, 6, 0, 1, 0, 0, 
    7, 15, 13, 16, 60, 25, 19, 9, 13, 12, 7, 4, 2, 0, 10, 
    19, 28, 59, 44, 43, 38, 18, 12, 1, 5, 12, 10, 4, 2, 0, 
    68, 53, 0, 15, 0, 12, 0, 8, 6, 6, 12, 10, 1, 0, 1, 
    10, 2, 0, 0, 0, 0, 0, 0, 3, 1, 0, 4, 6, 21, 11, 
    0, 0, 0, 11, 0, 0, 12, 5, 0, 0, 12, 13, 4, 1, 17, 
    0, 0, 0, 3, 21, 27, 0, 6, 7, 10, 20, 2, 15, 1, 5, 
    0, 5, 0, 0, 0, 7, 6, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 4, 0, 2, 3, 0, 0, 0, 0, 0, 
    
    -- channel=495
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 18, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    32, 36, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 5, 
    30, 31, 30, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 31, 33, 23, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    33, 44, 56, 34, 40, 25, 12, 0, 0, 0, 0, 0, 0, 0, 0, 
    67, 77, 72, 66, 24, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    88, 85, 38, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    57, 42, 28, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 9, 9, 8, 5, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=496
    29, 28, 30, 32, 37, 36, 29, 25, 19, 18, 15, 10, 5, 2, 0, 
    29, 26, 29, 28, 32, 42, 36, 28, 20, 16, 10, 4, 1, 1, 3, 
    29, 27, 26, 24, 32, 31, 37, 36, 22, 18, 22, 24, 23, 23, 21, 
    24, 23, 9, 12, 29, 27, 27, 33, 39, 44, 39, 35, 24, 19, 14, 
    19, 22, 25, 13, 24, 32, 31, 32, 37, 38, 43, 38, 27, 20, 17, 
    53, 63, 50, 14, 18, 33, 46, 41, 36, 35, 36, 42, 37, 32, 28, 
    65, 64, 54, 11, 28, 47, 45, 39, 38, 35, 36, 38, 38, 38, 32, 
    55, 54, 56, 44, 7, 14, 29, 37, 44, 41, 36, 35, 37, 31, 20, 
    56, 60, 52, 41, 53, 35, 39, 36, 49, 46, 37, 34, 36, 31, 26, 
    59, 77, 102, 83, 81, 59, 51, 43, 46, 47, 43, 38, 37, 23, 6, 
    108, 108, 85, 84, 67, 66, 52, 47, 46, 48, 46, 39, 30, 14, 4, 
    118, 107, 57, 40, 30, 36, 31, 20, 42, 43, 37, 37, 26, 26, 11, 
    58, 51, 46, 37, 24, 13, 35, 28, 28, 39, 42, 44, 27, 21, 23, 
    35, 32, 39, 40, 31, 21, 19, 30, 28, 42, 56, 44, 35, 21, 22, 
    32, 33, 24, 11, 13, 23, 23, 19, 12, 15, 23, 30, 21, 12, 12, 
    
    -- channel=497
    28, 25, 24, 22, 23, 30, 26, 20, 20, 16, 10, 7, 5, 7, 13, 
    26, 26, 20, 18, 24, 17, 26, 25, 16, 22, 28, 35, 40, 40, 34, 
    20, 21, 9, 3, 17, 21, 18, 24, 36, 49, 44, 39, 28, 19, 11, 
    22, 27, 38, 18, 17, 28, 33, 32, 23, 17, 30, 27, 23, 24, 24, 
    73, 89, 72, 26, 20, 35, 53, 42, 33, 27, 23, 31, 34, 40, 40, 
    66, 58, 58, 30, 37, 44, 37, 34, 38, 38, 31, 26, 28, 34, 32, 
    42, 43, 57, 54, 14, 11, 28, 34, 42, 42, 35, 28, 25, 17, 12, 
    52, 62, 57, 63, 78, 55, 49, 39, 45, 45, 38, 28, 25, 21, 28, 
    68, 86, 123, 104, 83, 64, 50, 48, 37, 42, 43, 37, 31, 21, 0, 
    135, 123, 75, 66, 47, 51, 39, 43, 38, 42, 45, 40, 24, 11, 7, 
    98, 83, 26, 8, 6, 8, 12, 16, 35, 33, 31, 34, 26, 31, 22, 
    9, 0, 31, 42, 29, 13, 35, 24, 12, 28, 44, 44, 24, 20, 28, 
    13, 14, 23, 33, 43, 39, 19, 29, 32, 42, 54, 41, 33, 15, 23, 
    24, 29, 16, 0, 0, 24, 26, 20, 14, 3, 8, 26, 22, 11, 8, 
    6, 0, 0, 9, 10, 18, 19, 12, 10, 12, 6, 2, 6, 6, 4, 
    
    -- channel=498
    4, 4, 1, 6, 2, 0, 0, 0, 4, 3, 0, 0, 0, 0, 0, 
    3, 3, 4, 0, 10, 5, 4, 0, 0, 0, 0, 0, 3, 8, 8, 
    1, 2, 7, 6, 0, 0, 0, 0, 0, 11, 13, 9, 8, 8, 2, 
    0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 2, 0, 0, 0, 1, 
    0, 13, 30, 8, 7, 10, 13, 10, 3, 0, 0, 0, 0, 0, 7, 
    13, 9, 5, 6, 0, 0, 0, 4, 4, 6, 2, 0, 0, 3, 6, 
    5, 1, 0, 0, 3, 15, 10, 0, 1, 7, 5, 0, 4, 3, 3, 
    0, 0, 11, 16, 13, 0, 6, 5, 7, 9, 5, 2, 0, 0, 0, 
    4, 0, 0, 11, 20, 15, 9, 9, 0, 3, 5, 4, 0, 10, 6, 
    20, 34, 36, 28, 6, 13, 3, 4, 0, 1, 5, 6, 1, 0, 0, 
    9, 16, 0, 0, 0, 0, 1, 6, 6, 6, 4, 0, 0, 2, 5, 
    14, 0, 1, 19, 0, 0, 0, 0, 0, 0, 5, 6, 1, 3, 1, 
    0, 0, 0, 2, 19, 24, 10, 0, 6, 5, 10, 9, 8, 0, 1, 
    0, 5, 9, 0, 0, 0, 0, 3, 2, 0, 0, 0, 4, 2, 0, 
    10, 0, 0, 0, 1, 2, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=499
    2, 3, 0, 1, 5, 12, 12, 5, 7, 8, 8, 10, 11, 10, 14, 
    3, 6, 3, 3, 16, 10, 19, 21, 10, 11, 14, 14, 14, 12, 12, 
    3, 4, 6, 8, 21, 26, 27, 25, 14, 10, 10, 9, 5, 5, 7, 
    5, 6, 21, 21, 27, 30, 29, 28, 26, 9, 10, 13, 5, 9, 12, 
    6, 4, 21, 25, 23, 14, 26, 35, 31, 31, 21, 18, 9, 10, 12, 
    0, 0, 15, 22, 26, 16, 22, 30, 27, 32, 33, 23, 8, 5, 7, 
    0, 0, 0, 35, 6, 2, 24, 26, 22, 30, 34, 22, 17, 3, 7, 
    0, 0, 0, 0, 40, 14, 26, 22, 19, 28, 34, 32, 22, 14, 10, 
    0, 0, 0, 12, 9, 22, 10, 29, 18, 25, 32, 36, 22, 13, 11, 
    0, 0, 0, 5, 0, 18, 6, 30, 21, 21, 27, 35, 25, 20, 12, 
    0, 0, 11, 0, 6, 13, 13, 12, 19, 18, 23, 31, 24, 17, 20, 
    0, 0, 0, 9, 26, 23, 12, 29, 18, 19, 19, 29, 24, 5, 22, 
    0, 0, 0, 0, 9, 17, 12, 22, 22, 13, 20, 24, 30, 15, 9, 
    2, 2, 4, 5, 4, 9, 17, 17, 16, 9, 6, 21, 23, 15, 8, 
    4, 5, 9, 14, 8, 7, 14, 15, 17, 16, 11, 9, 15, 14, 13, 
    
    -- channel=500
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=501
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 11, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 13, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 7, 16, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 24, 13, 27, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=502
    0, 1, 0, 0, 0, 0, 5, 0, 4, 2, 2, 6, 3, 0, 5, 
    0, 4, 0, 0, 5, 0, 4, 3, 1, 1, 2, 1, 0, 0, 4, 
    0, 0, 9, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 
    0, 0, 26, 1, 1, 0, 0, 0, 0, 0, 0, 7, 0, 5, 3, 
    0, 0, 45, 26, 0, 0, 2, 15, 1, 0, 0, 0, 0, 1, 0, 
    0, 0, 61, 24, 4, 0, 9, 13, 0, 6, 5, 0, 0, 0, 2, 
    0, 0, 9, 60, 0, 0, 13, 1, 0, 11, 13, 0, 0, 0, 7, 
    0, 0, 3, 5, 61, 0, 17, 0, 0, 17, 15, 0, 0, 0, 0, 
    0, 0, 3, 22, 12, 36, 0, 17, 0, 11, 12, 14, 0, 0, 8, 
    0, 0, 0, 56, 0, 48, 0, 23, 0, 1, 8, 20, 0, 12, 0, 
    0, 13, 68, 14, 0, 11, 0, 0, 0, 0, 8, 15, 0, 0, 10, 
    6, 9, 13, 20, 38, 0, 0, 23, 0, 0, 0, 14, 8, 0, 21, 
    0, 0, 0, 0, 17, 10, 0, 14, 0, 0, 7, 11, 14, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 3, 0, 0, 0, 7, 10, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 5, 0, 0, 
    
    -- channel=503
    14, 15, 10, 13, 21, 25, 23, 19, 15, 15, 16, 16, 14, 9, 11, 
    14, 16, 11, 18, 26, 30, 37, 30, 21, 13, 12, 11, 8, 4, 7, 
    16, 16, 17, 19, 35, 37, 38, 40, 27, 14, 11, 12, 10, 10, 13, 
    15, 12, 18, 17, 37, 37, 36, 33, 34, 31, 27, 24, 13, 12, 11, 
    3, 1, 20, 30, 31, 27, 32, 39, 42, 42, 40, 34, 13, 9, 8, 
    4, 9, 29, 24, 26, 19, 39, 47, 38, 38, 43, 35, 18, 9, 10, 
    11, 12, 15, 29, 15, 22, 43, 40, 34, 39, 43, 36, 30, 14, 16, 
    11, 8, 13, 17, 21, 6, 27, 31, 35, 43, 44, 42, 35, 19, 14, 
    4, 0, 3, 16, 21, 26, 20, 33, 38, 43, 44, 46, 35, 24, 14, 
    0, 0, 7, 43, 20, 37, 19, 44, 39, 41, 42, 48, 37, 25, 9, 
    4, 15, 40, 39, 38, 48, 40, 33, 36, 39, 38, 45, 32, 16, 8, 
    25, 30, 32, 18, 35, 35, 26, 27, 30, 36, 34, 35, 26, 7, 18, 
    24, 15, 16, 14, 22, 17, 16, 38, 30, 28, 34, 39, 34, 12, 12, 
    15, 13, 17, 18, 14, 15, 15, 22, 26, 25, 34, 40, 32, 16, 7, 
    14, 15, 14, 12, 3, 8, 18, 15, 11, 15, 13, 16, 18, 9, 8, 
    
    -- channel=504
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 8, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 1, 21, 2, 0, 0, 0, 0, 0, 0, 3, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 2, 1, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 23, 36, 25, 31, 14, 19, 0, 0, 0, 0, 0, 0, 0, 
    60, 60, 14, 0, 0, 8, 0, 0, 7, 0, 0, 0, 0, 0, 0, 
    21, 13, 2, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 19, 13, 0, 0, 0, 2, 13, 26, 3, 0, 0, 0, 
    9, 19, 8, 0, 0, 0, 0, 0, 0, 0, 1, 10, 5, 0, 0, 
    
    -- channel=505
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=506
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 8, 0, 9, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 15, 2, 8, 8, 11, 12, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 3, 8, 5, 11, 13, 11, 9, 3, 0, 3, 0, 2, 
    0, 0, 0, 4, 8, 16, 1, 2, 10, 9, 12, 5, 4, 3, 5, 
    0, 0, 0, 1, 2, 9, 0, 3, 8, 10, 8, 13, 14, 11, 6, 
    0, 0, 0, 0, 4, 24, 1, 6, 4, 2, 3, 19, 8, 12, 2, 
    0, 0, 0, 2, 0, 7, 0, 13, 5, 0, 2, 8, 4, 6, 2, 
    0, 0, 0, 0, 0, 0, 4, 0, 5, 0, 0, 0, 9, 6, 6, 
    0, 0, 0, 0, 0, 0, 7, 0, 3, 0, 0, 0, 7, 1, 17, 
    0, 0, 0, 0, 4, 1, 10, 20, 7, 4, 3, 1, 6, 8, 5, 
    0, 0, 0, 0, 0, 12, 10, 0, 12, 12, 5, 0, 6, 22, 2, 
    0, 0, 0, 0, 0, 0, 10, 0, 7, 17, 0, 0, 3, 16, 17, 
    1, 0, 0, 4, 17, 8, 10, 2, 12, 13, 9, 3, 0, 20, 21, 
    1, 9, 15, 14, 27, 14, 8, 14, 18, 13, 16, 15, 12, 22, 20, 
    
    -- channel=507
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 2, 3, 2, 2, 
    0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 
    0, 0, 5, 1, 2, 0, 0, 4, 0, 0, 0, 0, 3, 7, 12, 
    0, 0, 6, 0, 0, 0, 0, 0, 4, 5, 0, 8, 10, 7, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 4, 7, 10, 9, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 1, 0, 10, 17, 15, 
    0, 0, 0, 5, 1, 0, 0, 0, 0, 0, 0, 0, 10, 17, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 11, 
    0, 0, 0, 0, 0, 4, 5, 0, 0, 0, 0, 0, 0, 5, 26, 
    0, 0, 0, 9, 0, 14, 0, 0, 0, 0, 0, 0, 0, 21, 28, 
    0, 0, 15, 22, 8, 11, 6, 5, 0, 0, 0, 0, 3, 16, 18, 
    12, 25, 11, 0, 2, 0, 0, 1, 2, 0, 0, 0, 11, 16, 24, 
    9, 4, 8, 3, 1, 0, 0, 6, 0, 0, 0, 0, 12, 19, 21, 
    5, 1, 8, 22, 24, 17, 3, 8, 4, 3, 4, 0, 12, 26, 22, 
    13, 25, 28, 24, 19, 17, 16, 26, 21, 17, 12, 19, 26, 28, 28, 
    
    -- channel=508
    11, 10, 10, 13, 6, 0, 2, 4, 5, 3, 0, 0, 0, 0, 0, 
    11, 9, 10, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 9, 8, 0, 0, 0, 0, 0, 0, 3, 5, 5, 5, 7, 2, 
    6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 0, 
    9, 16, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28, 31, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 
    30, 28, 25, 0, 3, 1, 0, 0, 0, 0, 0, 0, 0, 4, 6, 
    22, 24, 27, 18, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 27, 30, 18, 22, 12, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    43, 54, 61, 42, 27, 24, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    62, 62, 25, 18, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    55, 39, 20, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 17, 12, 11, 8, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    6, 7, 7, 2, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=509
    2, 3, 1, 7, 7, 11, 13, 9, 6, 6, 8, 9, 9, 9, 12, 
    2, 4, 1, 15, 11, 12, 19, 18, 15, 10, 14, 14, 14, 12, 13, 
    3, 4, 7, 7, 18, 19, 21, 23, 22, 10, 12, 12, 13, 12, 15, 
    5, 4, 15, 18, 16, 16, 21, 25, 23, 20, 14, 18, 15, 17, 20, 
    6, 4, 6, 28, 13, 8, 14, 26, 26, 26, 23, 21, 19, 25, 25, 
    0, 1, 16, 28, 14, 7, 17, 20, 19, 26, 25, 20, 21, 24, 24, 
    0, 3, 11, 23, 9, 5, 19, 20, 16, 21, 26, 20, 17, 16, 19, 
    2, 4, 4, 26, 28, 15, 19, 20, 14, 18, 25, 20, 17, 19, 22, 
    2, 3, 11, 16, 8, 13, 15, 27, 13, 16, 21, 23, 17, 18, 24, 
    0, 0, 2, 12, 10, 22, 17, 29, 14, 14, 18, 24, 17, 24, 30, 
    0, 0, 27, 12, 8, 23, 11, 21, 15, 15, 19, 23, 21, 25, 34, 
    0, 4, 14, 11, 17, 15, 10, 17, 11, 15, 14, 19, 30, 24, 33, 
    7, 3, 9, 11, 22, 13, 11, 22, 14, 9, 9, 18, 28, 27, 29, 
    11, 10, 12, 19, 24, 23, 23, 21, 20, 7, 12, 15, 21, 32, 26, 
    13, 21, 26, 30, 27, 23, 23, 31, 33, 27, 21, 21, 29, 31, 31, 
    
    -- channel=510
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 3, 7, 9, 11, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 10, 8, 7, 
    0, 1, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 17, 18, 
    20, 23, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 29, 28, 
    22, 23, 18, 6, 0, 0, 0, 0, 0, 0, 0, 0, 2, 21, 20, 
    13, 17, 24, 17, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    18, 22, 23, 14, 25, 23, 15, 0, 0, 0, 0, 0, 0, 0, 25, 
    32, 47, 54, 47, 16, 28, 2, 0, 0, 0, 0, 0, 0, 5, 21, 
    54, 59, 28, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 19, 
    49, 34, 23, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 22, 
    13, 10, 8, 11, 10, 0, 0, 0, 0, 0, 0, 0, 2, 18, 23, 
    4, 8, 13, 18, 15, 14, 0, 2, 0, 0, 0, 0, 0, 19, 23, 
    15, 17, 16, 17, 18, 20, 14, 18, 16, 9, 3, 10, 14, 22, 25, 
    
    -- channel=511
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 7, 0, 0, 10, 0, 0, 0, 0, 0, 2, 6, 8, 1, 
    0, 0, 0, 2, 0, 3, 6, 6, 8, 7, 2, 1, 0, 0, 0, 
    0, 3, 0, 8, 2, 7, 9, 11, 9, 7, 1, 0, 0, 0, 0, 
    18, 21, 0, 0, 10, 23, 7, 0, 3, 6, 10, 0, 4, 0, 1, 
    13, 3, 0, 0, 2, 39, 0, 0, 5, 1, 2, 12, 13, 0, 0, 
    0, 0, 0, 0, 17, 19, 0, 1, 10, 0, 0, 18, 2, 4, 0, 
    4, 6, 0, 0, 0, 30, 0, 12, 12, 0, 0, 5, 4, 3, 0, 
    13, 17, 3, 0, 0, 0, 3, 0, 11, 0, 0, 0, 12, 2, 0, 
    29, 25, 0, 0, 0, 0, 13, 0, 10, 0, 0, 0, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 2, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 4, 18, 0, 13, 9, 6, 0, 0, 17, 0, 
    0, 0, 0, 0, 0, 0, 17, 0, 11, 25, 2, 0, 0, 9, 0, 
    0, 5, 0, 0, 0, 0, 1, 0, 2, 17, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 13, 10, 0, 0, 0, 1, 11, 2, 0, 2, 0, 
    
    -- channel=512
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=513
    9, 2, 22, 27, 18, 26, 30, 29, 29, 23, 8, 27, 33, 34, 35, 
    9, 0, 12, 22, 10, 18, 18, 22, 23, 28, 8, 21, 26, 28, 29, 
    10, 4, 7, 21, 2, 12, 7, 6, 8, 14, 9, 11, 16, 18, 23, 
    32, 26, 22, 25, 0, 13, 19, 17, 13, 6, 8, 13, 16, 15, 13, 
    35, 21, 21, 27, 2, 3, 12, 14, 7, 3, 11, 12, 14, 26, 18, 
    23, 20, 20, 25, 11, 6, 7, 12, 8, 4, 4, 9, 14, 27, 28, 
    24, 21, 25, 13, 7, 4, 11, 10, 14, 5, 7, 10, 16, 23, 30, 
    25, 19, 23, 11, 17, 4, 11, 6, 8, 19, 8, 13, 7, 16, 18, 
    25, 17, 20, 12, 11, 12, 10, 14, 14, 15, 18, 17, 7, 11, 13, 
    28, 24, 13, 11, 8, 3, 4, 15, 15, 16, 20, 19, 20, 22, 9, 
    21, 20, 9, 13, 15, 15, 5, 5, 15, 19, 16, 20, 14, 18, 19, 
    19, 23, 9, 9, 10, 19, 14, 14, 14, 23, 17, 17, 13, 20, 20, 
    20, 28, 15, 6, 9, 9, 10, 15, 17, 19, 14, 16, 13, 14, 17, 
    22, 28, 18, 7, 21, 17, 19, 15, 18, 19, 16, 16, 18, 13, 18, 
    19, 25, 22, 1, 12, 16, 19, 16, 19, 14, 17, 17, 20, 18, 15, 
    
    -- channel=514
    16, 13, 15, 3, 0, 7, 6, 7, 6, 0, 12, 8, 6, 7, 6, 
    16, 11, 16, 2, 1, 0, 9, 10, 3, 7, 14, 3, 0, 1, 2, 
    17, 13, 17, 0, 0, 0, 0, 0, 0, 8, 2, 0, 0, 0, 1, 
    9, 18, 21, 4, 0, 0, 3, 1, 3, 3, 3, 5, 0, 1, 5, 
    18, 18, 6, 3, 0, 0, 0, 0, 4, 1, 5, 4, 0, 2, 7, 
    8, 6, 8, 5, 4, 0, 0, 0, 4, 0, 0, 2, 0, 5, 11, 
    6, 4, 0, 5, 0, 0, 0, 8, 3, 4, 0, 4, 0, 5, 7, 
    6, 5, 0, 5, 0, 0, 0, 0, 10, 3, 3, 7, 8, 0, 8, 
    6, 1, 0, 0, 3, 1, 0, 0, 2, 1, 9, 1, 0, 0, 10, 
    9, 8, 0, 1, 0, 0, 0, 0, 0, 5, 1, 6, 5, 6, 0, 
    6, 2, 2, 0, 1, 0, 0, 0, 3, 1, 6, 5, 2, 0, 5, 
    4, 8, 2, 0, 0, 2, 3, 0, 0, 1, 9, 3, 5, 4, 5, 
    6, 11, 8, 0, 0, 0, 0, 0, 0, 4, 7, 3, 0, 5, 4, 
    7, 12, 9, 0, 0, 4, 0, 0, 1, 5, 6, 4, 4, 6, 7, 
    7, 15, 9, 0, 0, 0, 4, 7, 4, 9, 6, 7, 7, 8, 5, 
    
    -- channel=515
    3, 22, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 
    4, 17, 0, 0, 5, 3, 0, 0, 0, 0, 23, 0, 0, 0, 0, 
    2, 9, 5, 3, 15, 0, 5, 7, 0, 0, 21, 8, 3, 0, 0, 
    0, 12, 17, 0, 17, 0, 0, 0, 5, 20, 6, 12, 4, 2, 5, 
    0, 6, 3, 0, 24, 10, 0, 0, 6, 15, 10, 13, 5, 0, 10, 
    0, 5, 0, 0, 12, 8, 0, 0, 7, 16, 15, 19, 7, 0, 3, 
    0, 2, 0, 0, 11, 16, 3, 6, 3, 11, 15, 16, 9, 0, 1, 
    0, 0, 0, 11, 3, 7, 3, 7, 0, 10, 2, 12, 3, 5, 4, 
    0, 6, 0, 16, 2, 6, 10, 0, 14, 0, 0, 0, 26, 2, 12, 
    0, 4, 4, 2, 14, 13, 4, 0, 0, 4, 0, 0, 0, 0, 9, 
    4, 2, 10, 7, 6, 0, 15, 11, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 18, 7, 3, 0, 5, 2, 0, 0, 5, 0, 0, 0, 0, 
    4, 0, 12, 9, 0, 3, 5, 0, 0, 0, 2, 0, 1, 0, 0, 
    1, 0, 13, 12, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 
    0, 0, 12, 15, 3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    
    -- channel=516
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=517
    0, 22, 7, 0, 0, 0, 0, 0, 0, 0, 16, 5, 0, 0, 0, 
    0, 1, 28, 0, 0, 0, 4, 4, 1, 0, 38, 4, 0, 0, 0, 
    0, 0, 35, 0, 27, 0, 0, 12, 0, 0, 30, 17, 8, 7, 1, 
    0, 0, 31, 0, 39, 0, 0, 0, 0, 24, 18, 30, 14, 11, 20, 
    0, 13, 7, 0, 35, 15, 0, 0, 0, 16, 22, 37, 15, 0, 19, 
    3, 10, 7, 0, 25, 13, 0, 0, 1, 11, 19, 44, 18, 0, 3, 
    3, 4, 0, 8, 2, 5, 0, 5, 1, 15, 13, 41, 22, 5, 0, 
    0, 8, 0, 39, 1, 11, 0, 0, 12, 6, 8, 37, 36, 18, 10, 
    0, 5, 0, 24, 8, 11, 0, 0, 16, 0, 6, 0, 34, 12, 34, 
    0, 2, 16, 8, 20, 23, 15, 0, 0, 5, 0, 0, 0, 0, 15, 
    9, 0, 23, 8, 10, 0, 25, 16, 0, 0, 0, 3, 4, 0, 0, 
    12, 0, 33, 17, 12, 0, 13, 7, 3, 0, 8, 0, 9, 0, 0, 
    7, 0, 26, 17, 0, 0, 19, 5, 0, 0, 7, 0, 4, 0, 0, 
    2, 0, 20, 24, 0, 0, 1, 0, 0, 0, 2, 0, 0, 2, 0, 
    0, 0, 9, 33, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=518
    3, 0, 0, 2, 0, 0, 0, 0, 15, 44, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 5, 0, 0, 0, 59, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 43, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    36, 0, 0, 18, 0, 13, 24, 15, 0, 0, 0, 0, 0, 6, 0, 
    15, 0, 0, 42, 0, 0, 9, 34, 0, 0, 0, 0, 0, 25, 0, 
    0, 0, 0, 22, 0, 0, 17, 15, 0, 0, 0, 0, 0, 24, 0, 
    0, 0, 17, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 14, 
    4, 0, 42, 0, 5, 0, 2, 4, 0, 0, 0, 0, 0, 0, 0, 
    18, 0, 0, 0, 0, 0, 6, 26, 0, 14, 0, 24, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 11, 24, 0, 10, 0, 0, 0, 0, 
    0, 13, 0, 0, 0, 19, 0, 0, 9, 13, 0, 0, 0, 11, 0, 
    0, 16, 0, 0, 0, 17, 0, 0, 1, 36, 0, 0, 0, 10, 11, 
    0, 5, 0, 0, 18, 4, 0, 0, 9, 19, 0, 0, 0, 0, 1, 
    2, 8, 0, 0, 18, 3, 1, 0, 9, 10, 0, 0, 11, 0, 0, 
    4, 0, 0, 0, 3, 5, 22, 0, 18, 0, 0, 0, 7, 0, 0, 
    
    -- channel=519
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=520
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=521
    4, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 13, 1, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    2, 2, 0, 0, 15, 17, 0, 0, 0, 0, 16, 3, 3, 1, 0, 
    15, 6, 10, 0, 11, 15, 14, 7, 0, 7, 12, 8, 18, 16, 6, 
    0, 14, 5, 0, 11, 15, 10, 8, 3, 9, 8, 12, 14, 5, 1, 
    3, 6, 2, 0, 12, 15, 8, 5, 11, 14, 14, 9, 16, 7, 1, 
    1, 0, 0, 0, 13, 12, 11, 12, 16, 18, 13, 10, 14, 12, 13, 
    1, 0, 0, 0, 14, 19, 13, 14, 3, 8, 7, 0, 0, 11, 9, 
    5, 0, 0, 11, 15, 25, 26, 10, 0, 0, 0, 0, 0, 0, 0, 
    6, 8, 6, 13, 13, 12, 15, 18, 13, 0, 0, 0, 0, 0, 0, 
    9, 11, 7, 12, 12, 11, 7, 11, 4, 0, 0, 0, 0, 0, 0, 
    9, 6, 10, 14, 11, 1, 6, 7, 4, 0, 0, 0, 0, 0, 0, 
    8, 0, 7, 16, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 3, 14, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 12, 12, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=522
    0, 39, 39, 11, 8, 24, 12, 17, 0, 0, 34, 12, 12, 14, 12, 
    0, 12, 66, 21, 0, 0, 24, 19, 9, 0, 35, 8, 8, 14, 14, 
    0, 0, 65, 9, 23, 0, 7, 42, 30, 6, 20, 26, 12, 11, 4, 
    0, 0, 14, 0, 43, 0, 0, 0, 1, 28, 20, 29, 3, 7, 31, 
    0, 0, 8, 0, 34, 11, 0, 0, 6, 19, 29, 33, 11, 0, 34, 
    10, 15, 16, 0, 21, 9, 0, 0, 0, 5, 19, 51, 17, 0, 16, 
    13, 14, 7, 24, 0, 4, 0, 4, 0, 7, 12, 44, 23, 4, 0, 
    11, 19, 0, 58, 0, 2, 0, 0, 26, 7, 13, 71, 59, 23, 19, 
    0, 15, 0, 23, 3, 0, 0, 0, 28, 0, 14, 0, 65, 48, 59, 
    3, 0, 11, 8, 18, 27, 14, 0, 0, 14, 5, 17, 0, 6, 34, 
    15, 0, 27, 3, 6, 0, 30, 18, 0, 0, 12, 11, 10, 0, 10, 
    19, 0, 33, 12, 9, 1, 12, 7, 4, 0, 20, 9, 18, 0, 0, 
    14, 12, 32, 11, 0, 9, 35, 16, 10, 0, 24, 8, 20, 16, 1, 
    12, 10, 36, 20, 0, 0, 12, 16, 9, 3, 17, 6, 0, 18, 10, 
    20, 15, 25, 35, 0, 2, 5, 20, 0, 12, 10, 9, 0, 9, 16, 
    
    -- channel=523
    11, 0, 0, 0, 0, 0, 0, 0, 0, 12, 1, 0, 0, 0, 0, 
    11, 6, 0, 0, 12, 8, 1, 0, 1, 13, 0, 0, 0, 0, 0, 
    10, 9, 0, 1, 15, 22, 5, 2, 2, 11, 3, 9, 10, 8, 4, 
    7, 8, 0, 7, 7, 22, 17, 6, 6, 8, 10, 12, 16, 13, 10, 
    13, 6, 7, 10, 6, 18, 17, 14, 11, 10, 8, 6, 16, 13, 5, 
    9, 8, 7, 14, 8, 17, 14, 18, 12, 15, 11, 7, 15, 16, 6, 
    7, 8, 4, 4, 10, 20, 18, 18, 12, 13, 16, 5, 15, 16, 13, 
    10, 7, 6, 0, 19, 15, 22, 18, 8, 14, 10, 3, 5, 13, 18, 
    11, 7, 5, 0, 21, 16, 24, 14, 1, 12, 4, 4, 0, 8, 5, 
    12, 13, 8, 12, 12, 18, 22, 18, 15, 9, 0, 0, 5, 1, 0, 
    13, 17, 10, 13, 17, 13, 10, 17, 15, 1, 4, 0, 3, 5, 4, 
    12, 14, 8, 17, 15, 13, 6, 11, 10, 7, 0, 4, 4, 8, 3, 
    12, 9, 7, 17, 12, 8, 3, 6, 5, 7, 0, 6, 2, 3, 3, 
    11, 7, 7, 16, 14, 10, 0, 2, 4, 3, 0, 5, 5, 0, 4, 
    9, 4, 10, 12, 18, 10, 6, 0, 1, 4, 0, 2, 3, 2, 0, 
    
    -- channel=524
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=525
    1, 5, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    1, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 1, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 3, 0, 0, 12, 10, 0, 4, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 11, 7, 
    0, 0, 0, 0, 0, 5, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 1, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=526
    3, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 21, 0, 0, 0, 0, 7, 14, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 66, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=527
    0, 0, 6, 0, 0, 0, 0, 0, 2, 0, 10, 2, 0, 0, 0, 
    0, 0, 10, 0, 22, 0, 5, 8, 3, 0, 24, 8, 0, 0, 0, 
    0, 0, 11, 0, 36, 7, 0, 0, 1, 12, 21, 12, 12, 13, 9, 
    0, 0, 16, 0, 36, 22, 8, 0, 2, 14, 24, 26, 24, 15, 16, 
    1, 14, 8, 0, 25, 23, 15, 0, 9, 13, 19, 28, 19, 0, 2, 
    6, 7, 6, 0, 22, 19, 11, 0, 17, 17, 17, 28, 19, 0, 0, 
    0, 2, 0, 20, 10, 13, 10, 15, 15, 21, 15, 28, 19, 17, 0, 
    0, 4, 0, 31, 12, 22, 16, 12, 23, 0, 14, 0, 30, 14, 13, 
    0, 0, 13, 17, 28, 30, 17, 9, 0, 0, 14, 0, 0, 2, 12, 
    3, 0, 18, 21, 13, 19, 31, 19, 3, 12, 0, 1, 3, 0, 0, 
    9, 0, 22, 16, 18, 5, 17, 18, 14, 0, 0, 5, 11, 0, 0, 
    7, 2, 20, 24, 20, 5, 18, 15, 10, 0, 6, 2, 15, 0, 0, 
    4, 0, 11, 24, 10, 0, 20, 5, 0, 0, 5, 0, 0, 2, 0, 
    0, 0, 0, 26, 7, 12, 2, 0, 0, 0, 1, 0, 0, 1, 4, 
    0, 0, 0, 31, 14, 5, 0, 0, 0, 0, 0, 1, 0, 0, 1, 
    
    -- channel=528
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 21, 15, 0, 0, 8, 5, 0, 0, 0, 0, 1, 4, 0, 0, 
    1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 12, 6, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=529
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 19, 24, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 34, 1, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 19, 0, 0, 4, 2, 0, 0, 3, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 8, 4, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 10, 3, 5, 0, 0, 0, 0, 0, 0, 
    
    -- channel=530
    39, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    36, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=531
    16, 13, 0, 10, 5, 4, 4, 2, 0, 17, 2, 0, 0, 0, 1, 
    16, 18, 0, 13, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 
    17, 18, 0, 11, 0, 0, 12, 9, 11, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 5, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 7, 4, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 8, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 2, 5, 0, 7, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 5, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 1, 0, 1, 5, 
    0, 0, 0, 0, 0, 25, 0, 0, 1, 7, 1, 4, 4, 5, 3, 
    0, 0, 0, 0, 0, 4, 2, 4, 7, 11, 2, 5, 7, 6, 0, 
    0, 0, 0, 0, 0, 0, 5, 8, 12, 8, 5, 2, 5, 2, 5, 
    
    -- channel=532
    5, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=533
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=534
    10, 12, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 
    11, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=535
    0, 0, 25, 33, 34, 23, 32, 26, 51, 47, 0, 40, 38, 37, 39, 
    0, 0, 12, 11, 49, 41, 32, 36, 53, 72, 0, 57, 53, 46, 45, 
    0, 0, 0, 12, 38, 90, 33, 25, 44, 21, 35, 51, 62, 59, 60, 
    42, 0, 9, 53, 26, 78, 54, 50, 25, 0, 67, 35, 72, 88, 53, 
    68, 26, 62, 67, 14, 58, 72, 67, 26, 5, 44, 50, 82, 94, 41, 
    64, 51, 70, 51, 35, 57, 75, 40, 39, 15, 39, 46, 85, 100, 57, 
    65, 50, 64, 47, 54, 37, 74, 17, 64, 39, 35, 47, 77, 91, 70, 
    70, 45, 72, 16, 68, 59, 60, 49, 43, 30, 59, 27, 51, 94, 61, 
    89, 38, 54, 25, 65, 69, 64, 90, 1, 38, 60, 43, 6, 62, 28, 
    83, 45, 55, 62, 55, 65, 65, 69, 58, 31, 61, 33, 19, 48, 26, 
    73, 74, 45, 60, 62, 82, 40, 51, 76, 69, 25, 29, 41, 50, 36, 
    68, 89, 31, 66, 75, 60, 46, 53, 66, 65, 12, 40, 44, 48, 42, 
    72, 76, 33, 68, 97, 6, 49, 52, 63, 46, 23, 35, 41, 35, 39, 
    72, 71, 23, 63, 83, 27, 57, 44, 46, 23, 26, 30, 39, 11, 34, 
    60, 65, 20, 51, 71, 70, 53, 32, 45, 6, 24, 30, 32, 23, 30, 
    
    -- channel=536
    3, 11, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    3, 11, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 6, 0, 0, 10, 5, 7, 4, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 3, 0, 0, 0, 10, 4, 1, 6, 5, 0, 
    0, 0, 0, 0, 10, 13, 5, 1, 3, 10, 6, 0, 3, 0, 0, 
    0, 0, 0, 0, 3, 12, 8, 5, 2, 10, 10, 1, 2, 0, 0, 
    0, 0, 1, 0, 7, 13, 6, 5, 6, 6, 12, 3, 3, 0, 0, 
    0, 0, 0, 0, 5, 8, 7, 14, 0, 11, 6, 11, 0, 2, 0, 
    0, 0, 0, 9, 3, 2, 11, 2, 10, 0, 0, 0, 13, 3, 0, 
    0, 0, 2, 0, 11, 17, 9, 5, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 2, 5, 2, 5, 9, 12, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 7, 8, 1, 1, 3, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 5, 15, 0, 2, 0, 0, 0, 0, 4, 0, 0, 
    0, 0, 0, 6, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 5, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=537
    0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 17, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 0, 0, 0, 0, 8, 28, 26, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 49, 11, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 29, 28, 8, 
    0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 3, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 1, 1, 0, 3, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 11, 1, 3, 5, 0, 0, 0, 14, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 12, 8, 2, 0, 0, 0, 0, 0, 1, 
    
    -- channel=538
    2, 29, 31, 32, 34, 32, 31, 36, 31, 14, 40, 50, 40, 40, 36, 
    2, 15, 32, 37, 55, 46, 44, 49, 47, 19, 60, 59, 51, 46, 43, 
    2, 6, 36, 36, 68, 43, 33, 36, 32, 38, 69, 64, 64, 65, 62, 
    13, 28, 65, 39, 67, 58, 43, 33, 33, 56, 66, 75, 82, 72, 70, 
    50, 61, 62, 32, 62, 65, 55, 34, 36, 51, 70, 80, 79, 59, 61, 
    59, 63, 59, 38, 65, 64, 46, 34, 43, 52, 65, 82, 82, 59, 55, 
    59, 57, 44, 43, 50, 54, 48, 53, 57, 56, 64, 82, 83, 77, 65, 
    57, 55, 25, 64, 64, 60, 56, 46, 51, 58, 53, 68, 74, 76, 70, 
    51, 49, 46, 70, 68, 73, 64, 45, 53, 38, 48, 22, 53, 49, 70, 
    62, 59, 64, 62, 68, 69, 68, 64, 40, 46, 43, 33, 38, 43, 45, 
    69, 56, 67, 67, 68, 54, 62, 64, 58, 43, 32, 45, 46, 37, 36, 
    69, 53, 71, 73, 68, 54, 61, 60, 55, 30, 42, 44, 48, 39, 31, 
    65, 55, 66, 70, 49, 35, 56, 52, 43, 29, 39, 37, 41, 35, 34, 
    61, 48, 57, 73, 56, 46, 50, 37, 30, 26, 36, 32, 27, 34, 39, 
    51, 45, 49, 72, 63, 52, 33, 30, 20, 23, 32, 33, 29, 35, 36, 
    
    -- channel=539
    12, 16, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    13, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 12, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=540
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 9, 2, 0, 0, 1, 4, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 9, 11, 0, 0, 1, 0, 7, 0, 0, 0, 1, 
    0, 0, 0, 0, 2, 9, 4, 0, 3, 0, 6, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 3, 5, 5, 3, 0, 1, 5, 3, 0, 0, 
    0, 0, 0, 0, 1, 10, 6, 2, 2, 4, 2, 0, 2, 4, 0, 
    0, 0, 0, 0, 0, 1, 14, 0, 10, 0, 0, 0, 3, 2, 1, 
    0, 0, 0, 0, 9, 3, 0, 10, 0, 0, 2, 0, 0, 10, 0, 
    2, 0, 0, 0, 2, 8, 12, 5, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 7, 0, 0, 0, 5, 2, 7, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 6, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 12, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=541
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=542
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 2, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    23, 25, 6, 0, 0, 1, 6, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 4, 0, 1, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 9, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=543
    0, 0, 23, 42, 40, 28, 41, 35, 57, 57, 0, 43, 52, 52, 54, 
    0, 0, 0, 29, 55, 53, 40, 47, 61, 85, 0, 68, 65, 59, 59, 
    0, 0, 0, 29, 44, 102, 34, 19, 43, 34, 29, 57, 73, 71, 74, 
    45, 0, 0, 67, 27, 91, 75, 49, 21, 6, 64, 51, 94, 98, 65, 
    77, 41, 65, 80, 12, 68, 81, 74, 26, 18, 44, 57, 95, 104, 48, 
    72, 61, 72, 75, 38, 69, 81, 53, 37, 29, 45, 46, 95, 106, 58, 
    71, 61, 72, 50, 57, 47, 74, 36, 66, 43, 48, 50, 90, 100, 85, 
    78, 58, 90, 6, 81, 69, 68, 68, 45, 48, 68, 30, 63, 98, 81, 
    91, 45, 63, 37, 81, 79, 82, 86, 10, 63, 52, 60, 0, 58, 36, 
    86, 62, 64, 74, 62, 73, 82, 87, 79, 39, 60, 36, 39, 48, 29, 
    79, 85, 49, 75, 76, 90, 42, 67, 85, 69, 38, 35, 48, 58, 40, 
    75, 91, 36, 80, 87, 80, 58, 68, 76, 75, 17, 48, 46, 62, 50, 
    77, 76, 41, 78, 96, 39, 48, 64, 69, 56, 23, 44, 40, 41, 43, 
    78, 71, 31, 66, 93, 62, 60, 51, 52, 34, 22, 38, 44, 16, 38, 
    64, 58, 32, 51, 84, 77, 63, 35, 45, 14, 27, 33, 40, 26, 33, 
    
    -- channel=544
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=545
    0, 0, 0, 0, 0, 0, 0, 0, 14, 26, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    36, 0, 0, 0, 0, 6, 7, 9, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 29, 0, 0, 0, 19, 0, 0, 0, 0, 0, 11, 0, 
    0, 0, 0, 9, 0, 0, 9, 10, 0, 0, 0, 0, 0, 13, 0, 
    0, 0, 3, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 2, 0, 0, 0, 0, 23, 0, 0, 0, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 10, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 16, 0, 0, 0, 1, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 0, 0, 0, 1, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 10, 0, 0, 0, 0, 0, 0, 
    
    -- channel=546
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 9, 22, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 26, 19, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 6, 32, 7, 
    0, 0, 0, 0, 0, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 0, 0, 0, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 18, 0, 0, 6, 3, 0, 0, 0, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 4, 10, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 12, 4, 3, 0, 0, 0, 0, 0, 0, 
    
    -- channel=547
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 24, 25, 25, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 0, 5, 0, 0, 0, 0, 0, 4, 4, 
    0, 0, 0, 0, 0, 0, 8, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 20, 0, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 40, 0, 2, 0, 
    0, 7, 0, 0, 0, 0, 0, 0, 10, 3, 0, 0, 43, 34, 3, 
    0, 0, 0, 0, 8, 15, 0, 0, 0, 0, 11, 0, 0, 0, 19, 
    0, 0, 0, 0, 0, 3, 4, 6, 0, 6, 1, 0, 0, 5, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 12, 37, 0, 7, 12, 6, 0, 4, 14, 6, 0, 
    0, 1, 4, 0, 0, 0, 5, 11, 13, 13, 0, 0, 4, 0, 0, 
    15, 0, 13, 0, 0, 0, 17, 5, 11, 0, 2, 0, 0, 0, 4, 
    
    -- channel=548
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=549
    2, 0, 0, 0, 1, 0, 5, 5, 27, 29, 0, 21, 14, 12, 9, 
    2, 0, 0, 0, 19, 13, 0, 2, 0, 11, 34, 14, 12, 8, 5, 
    3, 0, 0, 11, 0, 15, 0, 0, 0, 0, 24, 0, 1, 9, 16, 
    103, 78, 64, 0, 0, 11, 51, 23, 3, 0, 0, 2, 13, 0, 0, 
    28, 50, 9, 7, 0, 0, 0, 0, 0, 0, 0, 4, 2, 0, 0, 
    1, 0, 0, 11, 1, 0, 0, 0, 18, 12, 0, 0, 0, 11, 2, 
    0, 0, 0, 0, 4, 0, 2, 5, 10, 5, 1, 0, 0, 10, 27, 
    0, 0, 3, 0, 8, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 10, 10, 2, 33, 32, 9, 0, 0, 0, 22, 0, 0, 0, 
    5, 17, 1, 3, 0, 0, 0, 21, 52, 4, 0, 0, 21, 5, 0, 
    0, 3, 0, 10, 9, 1, 0, 0, 0, 0, 0, 8, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 8, 1, 0, 0, 6, 0, 0, 2, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 5, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 4, 0, 
    
    -- channel=550
    19, 28, 14, 9, 16, 14, 14, 12, 4, 20, 14, 9, 10, 12, 12, 
    20, 31, 15, 5, 2, 14, 10, 9, 8, 6, 15, 8, 9, 11, 10, 
    20, 26, 15, 12, 0, 7, 15, 17, 11, 4, 11, 10, 7, 5, 6, 
    18, 14, 16, 14, 0, 0, 7, 9, 10, 11, 4, 4, 0, 6, 8, 
    7, 14, 11, 12, 5, 1, 3, 8, 11, 10, 5, 6, 5, 14, 20, 
    11, 12, 12, 14, 2, 3, 5, 8, 8, 10, 10, 6, 7, 16, 22, 
    15, 14, 16, 8, 8, 7, 6, 3, 2, 6, 10, 6, 7, 5, 15, 
    17, 13, 11, 0, 3, 5, 0, 14, 3, 11, 12, 15, 5, 9, 13, 
    17, 16, 0, 1, 0, 0, 3, 2, 14, 13, 7, 22, 21, 15, 15, 
    12, 14, 4, 3, 7, 5, 0, 0, 17, 10, 9, 10, 12, 11, 20, 
    11, 16, 4, 5, 4, 7, 7, 6, 1, 11, 11, 9, 8, 9, 14, 
    13, 13, 8, 1, 3, 2, 5, 4, 8, 9, 14, 10, 6, 11, 11, 
    16, 17, 12, 3, 6, 12, 5, 9, 9, 14, 13, 12, 11, 9, 12, 
    17, 22, 18, 3, 0, 9, 5, 13, 14, 14, 13, 14, 13, 14, 10, 
    19, 21, 23, 3, 5, 10, 13, 12, 15, 20, 14, 13, 12, 15, 11, 
    
    -- channel=551
    0, 9, 28, 20, 23, 27, 27, 26, 17, 7, 11, 25, 28, 28, 29, 
    0, 2, 29, 14, 9, 17, 19, 21, 17, 3, 14, 24, 27, 28, 27, 
    0, 0, 25, 13, 7, 4, 12, 19, 17, 8, 19, 21, 20, 22, 23, 
    0, 0, 19, 16, 10, 3, 3, 7, 7, 10, 16, 15, 15, 18, 20, 
    13, 14, 20, 12, 10, 8, 8, 4, 5, 7, 18, 20, 20, 22, 25, 
    20, 20, 21, 12, 10, 8, 9, 3, 4, 5, 16, 23, 24, 24, 26, 
    24, 21, 21, 14, 12, 7, 7, 2, 7, 6, 12, 24, 22, 23, 24, 
    24, 19, 14, 19, 10, 8, 3, 5, 9, 10, 14, 26, 25, 24, 21, 
    22, 18, 11, 19, 8, 7, 4, 6, 17, 10, 14, 13, 27, 24, 26, 
    23, 16, 15, 13, 15, 13, 6, 7, 9, 12, 18, 17, 12, 17, 23, 
    23, 16, 15, 16, 13, 12, 12, 11, 11, 17, 13, 16, 15, 14, 14, 
    23, 17, 16, 13, 15, 11, 14, 13, 14, 13, 15, 14, 14, 12, 12, 
    24, 24, 17, 13, 11, 12, 17, 17, 15, 12, 16, 12, 15, 13, 13, 
    24, 26, 20, 14, 11, 8, 20, 16, 15, 12, 15, 12, 11, 13, 13, 
    23, 25, 17, 14, 12, 16, 15, 15, 13, 11, 13, 13, 11, 13, 15, 
    
    -- channel=552
    4, 0, 18, 23, 26, 18, 22, 23, 37, 28, 0, 26, 24, 25, 24, 
    3, 0, 9, 15, 44, 32, 29, 31, 36, 45, 1, 45, 39, 33, 30, 
    1, 0, 0, 14, 42, 61, 23, 22, 33, 30, 36, 50, 55, 52, 50, 
    26, 0, 16, 36, 33, 62, 42, 33, 22, 11, 56, 44, 60, 65, 52, 
    56, 31, 52, 46, 24, 50, 54, 44, 26, 18, 44, 51, 69, 70, 43, 
    54, 46, 56, 43, 34, 47, 53, 35, 35, 25, 40, 52, 74, 79, 52, 
    55, 46, 43, 42, 44, 41, 53, 27, 47, 38, 41, 50, 70, 78, 62, 
    58, 42, 43, 23, 54, 49, 52, 37, 41, 30, 47, 27, 55, 74, 64, 
    69, 37, 40, 24, 60, 58, 53, 59, 9, 34, 45, 31, 13, 52, 41, 
    69, 44, 46, 52, 48, 55, 59, 58, 43, 32, 36, 26, 22, 33, 23, 
    65, 60, 47, 52, 54, 57, 39, 47, 58, 41, 26, 25, 32, 35, 27, 
    61, 69, 38, 57, 58, 45, 40, 44, 48, 42, 17, 31, 36, 36, 30, 
    62, 62, 39, 59, 62, 10, 40, 40, 43, 33, 22, 28, 28, 29, 29, 
    61, 58, 34, 59, 60, 25, 37, 32, 31, 19, 21, 25, 27, 14, 29, 
    52, 55, 29, 52, 58, 51, 35, 23, 28, 13, 20, 25, 25, 19, 24, 
    
    -- channel=553
    3, 0, 0, 11, 9, 11, 14, 10, 11, 22, 0, 0, 11, 12, 15, 
    3, 0, 0, 6, 0, 8, 1, 0, 4, 26, 0, 2, 9, 10, 12, 
    4, 0, 0, 7, 0, 9, 6, 1, 8, 1, 0, 0, 0, 0, 3, 
    15, 0, 0, 15, 0, 0, 5, 4, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 24, 0, 0, 0, 10, 0, 0, 0, 0, 0, 18, 1, 
    4, 0, 3, 18, 0, 0, 5, 10, 0, 0, 0, 0, 0, 16, 10, 
    8, 6, 18, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 11, 
    12, 5, 22, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 2, 
    14, 6, 4, 0, 0, 0, 0, 6, 0, 11, 0, 13, 0, 8, 0, 
    9, 4, 0, 0, 0, 0, 0, 0, 7, 0, 8, 5, 4, 2, 0, 
    2, 10, 0, 0, 0, 7, 0, 0, 3, 7, 9, 0, 0, 11, 5, 
    2, 11, 0, 0, 0, 6, 0, 0, 1, 21, 0, 3, 0, 8, 10, 
    5, 14, 0, 0, 6, 15, 0, 4, 9, 14, 0, 6, 2, 6, 5, 
    8, 16, 0, 0, 8, 1, 4, 8, 13, 15, 0, 6, 12, 0, 1, 
    13, 11, 8, 0, 0, 5, 16, 5, 15, 4, 5, 3, 9, 0, 2, 
    
    -- channel=554
    0, 3, 93, 86, 76, 83, 85, 85, 78, 37, 43, 94, 101, 100, 101, 
    0, 0, 87, 80, 82, 70, 86, 91, 99, 63, 57, 105, 107, 107, 107, 
    0, 0, 56, 74, 102, 82, 61, 82, 89, 66, 85, 107, 113, 111, 107, 
    2, 0, 58, 80, 102, 98, 61, 55, 54, 64, 107, 109, 120, 118, 112, 
    84, 69, 97, 72, 85, 103, 98, 70, 58, 62, 97, 119, 128, 107, 97, 
    102, 96, 105, 79, 91, 97, 93, 60, 64, 63, 87, 124, 129, 110, 89, 
    102, 97, 94, 105, 85, 82, 87, 64, 81, 75, 84, 120, 131, 125, 89, 
    101, 98, 92, 107, 97, 92, 88, 73, 90, 74, 95, 104, 133, 134, 111, 
    100, 84, 100, 93, 108, 101, 87, 86, 63, 76, 97, 61, 86, 115, 109, 
    105, 83, 105, 104, 104, 117, 115, 92, 67, 85, 86, 83, 68, 82, 84, 
    110, 94, 105, 105, 107, 97, 100, 106, 106, 90, 72, 77, 87, 80, 74, 
    109, 102, 99, 117, 117, 100, 99, 101, 102, 77, 69, 81, 93, 80, 67, 
    104, 98, 94, 114, 113, 73, 112, 101, 97, 72, 74, 74, 82, 78, 71, 
    101, 90, 83, 114, 103, 78, 94, 89, 80, 56, 68, 68, 63, 61, 77, 
    91, 87, 68, 111, 105, 101, 81, 77, 64, 50, 61, 68, 59, 62, 72, 
    
    -- channel=555
    0, 75, 11, 0, 0, 5, 0, 1, 0, 0, 53, 0, 0, 0, 0, 
    2, 47, 32, 16, 0, 0, 2, 2, 0, 0, 60, 0, 0, 0, 0, 
    2, 17, 56, 14, 12, 0, 0, 13, 0, 5, 14, 0, 0, 0, 0, 
    0, 19, 27, 0, 29, 0, 0, 0, 0, 39, 0, 13, 0, 0, 0, 
    0, 8, 0, 0, 31, 0, 0, 0, 3, 26, 5, 10, 0, 0, 5, 
    0, 0, 0, 0, 12, 0, 0, 0, 0, 15, 6, 17, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 11, 0, 4, 3, 15, 0, 0, 0, 
    0, 0, 0, 39, 0, 0, 0, 0, 4, 0, 0, 25, 14, 0, 0, 
    0, 0, 0, 20, 0, 0, 0, 0, 27, 0, 0, 0, 39, 0, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 2, 0, 15, 
    0, 0, 3, 0, 0, 0, 11, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 
    0, 0, 14, 0, 0, 12, 5, 0, 0, 0, 11, 0, 0, 0, 0, 
    0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 15, 0, 
    0, 0, 11, 6, 0, 0, 0, 0, 0, 13, 1, 0, 0, 4, 2, 
    
    -- channel=556
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 12, 3, 1, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 1, 6, 0, 0, 0, 0, 1, 0, 6, 11, 1, 
    0, 0, 0, 1, 0, 9, 8, 7, 0, 0, 0, 0, 5, 3, 0, 
    0, 0, 0, 0, 0, 11, 10, 2, 0, 0, 1, 0, 5, 0, 0, 
    0, 0, 4, 0, 1, 3, 8, 1, 0, 0, 0, 0, 4, 1, 0, 
    0, 0, 2, 0, 6, 7, 8, 7, 0, 1, 4, 11, 1, 9, 1, 
    0, 0, 0, 0, 5, 0, 6, 4, 0, 0, 0, 0, 0, 9, 0, 
    0, 0, 0, 2, 7, 17, 13, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 0, 1, 1, 8, 0, 10, 6, 2, 0, 0, 0, 0, 0, 
    1, 1, 0, 9, 10, 9, 0, 2, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 13, 7, 0, 3, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 4, 7, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=557
    3, 0, 0, 5, 2, 0, 4, 0, 32, 29, 0, 0, 3, 1, 6, 
    0, 0, 0, 0, 7, 0, 0, 0, 3, 66, 0, 1, 5, 3, 6, 
    0, 0, 0, 0, 0, 48, 0, 0, 4, 7, 0, 0, 1, 0, 5, 
    39, 0, 0, 8, 0, 33, 28, 18, 0, 0, 0, 0, 0, 9, 0, 
    32, 0, 0, 39, 0, 0, 18, 34, 0, 0, 0, 0, 2, 30, 0, 
    5, 0, 5, 24, 0, 0, 26, 18, 0, 0, 0, 0, 2, 38, 0, 
    2, 0, 12, 2, 0, 0, 19, 0, 7, 0, 0, 0, 0, 21, 16, 
    6, 0, 49, 0, 8, 0, 14, 0, 0, 0, 0, 0, 0, 4, 0, 
    28, 0, 21, 0, 10, 6, 8, 43, 0, 12, 5, 24, 0, 0, 0, 
    21, 0, 0, 4, 0, 0, 6, 25, 23, 0, 12, 2, 0, 1, 0, 
    4, 13, 0, 0, 0, 23, 0, 0, 25, 12, 5, 0, 0, 14, 0, 
    0, 29, 0, 0, 5, 19, 0, 0, 7, 40, 0, 0, 0, 12, 17, 
    2, 13, 0, 0, 31, 0, 0, 0, 14, 20, 0, 0, 0, 5, 6, 
    8, 15, 0, 0, 32, 0, 1, 3, 10, 6, 0, 0, 12, 0, 0, 
    6, 14, 0, 0, 12, 10, 18, 0, 20, 0, 0, 0, 11, 0, 0, 
    
    -- channel=558
    1, 0, 7, 13, 3, 3, 13, 15, 39, 18, 0, 27, 24, 21, 19, 
    1, 0, 0, 2, 29, 9, 2, 15, 13, 24, 28, 22, 17, 15, 14, 
    2, 0, 0, 10, 13, 20, 0, 0, 0, 11, 24, 0, 14, 21, 25, 
    76, 56, 58, 6, 0, 28, 48, 23, 6, 0, 7, 17, 27, 10, 0, 
    46, 50, 18, 12, 2, 0, 12, 8, 2, 0, 2, 20, 14, 7, 0, 
    16, 9, 7, 18, 16, 1, 0, 2, 25, 11, 0, 3, 11, 22, 7, 
    9, 6, 0, 17, 4, 0, 12, 12, 23, 12, 2, 8, 10, 30, 29, 
    5, 0, 14, 11, 21, 10, 9, 15, 0, 1, 0, 0, 0, 1, 8, 
    15, 0, 26, 12, 22, 44, 31, 20, 0, 2, 17, 16, 0, 0, 0, 
    21, 22, 14, 15, 0, 0, 3, 31, 38, 15, 0, 4, 22, 15, 0, 
    12, 10, 5, 16, 23, 10, 0, 0, 11, 2, 0, 16, 11, 0, 1, 
    4, 15, 4, 10, 8, 5, 20, 12, 8, 2, 11, 2, 9, 11, 9, 
    5, 4, 1, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    4, 3, 0, 7, 20, 40, 0, 0, 0, 0, 1, 0, 0, 0, 10, 
    0, 6, 0, 0, 10, 4, 0, 0, 0, 0, 0, 5, 11, 9, 0, 
    
    -- channel=559
    0, 0, 33, 31, 28, 28, 31, 30, 34, 7, 8, 43, 45, 43, 43, 
    0, 0, 21, 26, 45, 30, 35, 41, 45, 27, 21, 55, 52, 50, 49, 
    0, 0, 4, 24, 54, 48, 18, 23, 29, 27, 43, 54, 62, 60, 57, 
    0, 0, 25, 30, 48, 59, 37, 22, 15, 24, 57, 58, 73, 67, 57, 
    45, 37, 50, 30, 37, 56, 53, 31, 19, 23, 50, 64, 75, 57, 41, 
    51, 48, 51, 37, 43, 51, 47, 24, 28, 28, 46, 63, 76, 63, 38, 
    50, 47, 41, 49, 41, 41, 44, 30, 41, 36, 44, 63, 75, 76, 51, 
    48, 46, 45, 46, 54, 49, 46, 38, 41, 33, 46, 37, 67, 74, 62, 
    50, 34, 51, 44, 63, 64, 54, 47, 19, 34, 45, 26, 22, 47, 50, 
    55, 41, 55, 56, 53, 59, 64, 57, 40, 38, 35, 30, 29, 35, 30, 
    59, 48, 54, 59, 61, 52, 46, 55, 58, 38, 25, 31, 39, 33, 26, 
    57, 51, 48, 67, 65, 53, 51, 53, 52, 33, 23, 33, 42, 35, 25, 
    54, 44, 42, 64, 58, 29, 51, 47, 43, 26, 24, 27, 28, 28, 26, 
    51, 39, 30, 63, 57, 43, 40, 35, 28, 13, 20, 23, 19, 16, 30, 
    38, 37, 18, 58, 59, 50, 30, 24, 17, 9, 16, 22, 19, 18, 24, 
    
    -- channel=560
    0, 25, 61, 52, 54, 59, 55, 55, 41, 19, 42, 60, 62, 64, 63, 
    0, 12, 65, 55, 51, 53, 63, 65, 66, 30, 43, 75, 74, 72, 70, 
    0, 0, 50, 51, 70, 53, 55, 71, 71, 47, 65, 91, 83, 79, 75, 
    0, 0, 35, 61, 78, 62, 31, 33, 38, 56, 80, 85, 85, 90, 95, 
    52, 48, 74, 54, 66, 79, 67, 46, 43, 55, 79, 93, 99, 87, 90, 
    79, 79, 84, 57, 65, 75, 68, 45, 39, 50, 74, 103, 105, 86, 81, 
    84, 81, 78, 67, 66, 68, 58, 49, 52, 59, 71, 99, 107, 94, 76, 
    85, 81, 55, 71, 68, 69, 63, 50, 69, 63, 74, 104, 112, 108, 96, 
    80, 74, 57, 67, 77, 65, 60, 53, 61, 59, 63, 44, 89, 103, 101, 
    83, 67, 76, 76, 86, 96, 86, 61, 42, 58, 64, 56, 44, 55, 77, 
    91, 78, 83, 79, 78, 72, 82, 84, 74, 63, 55, 52, 60, 58, 53, 
    94, 80, 82, 87, 87, 72, 68, 73, 73, 54, 50, 60, 63, 54, 46, 
    90, 84, 84, 87, 82, 64, 78, 78, 72, 52, 56, 56, 64, 59, 49, 
    88, 79, 82, 88, 69, 42, 69, 68, 59, 46, 50, 50, 45, 48, 52, 
    85, 74, 74, 89, 79, 73, 63, 55, 45, 39, 47, 48, 40, 43, 56, 
    
    -- channel=561
    0, 0, 50, 55, 54, 54, 62, 66, 81, 42, 37, 83, 79, 75, 72, 
    0, 0, 24, 45, 79, 63, 51, 67, 63, 57, 70, 89, 84, 78, 75, 
    0, 0, 29, 54, 68, 67, 22, 12, 15, 55, 79, 70, 84, 92, 95, 
    90, 81, 97, 53, 46, 86, 89, 57, 42, 47, 67, 86, 101, 77, 70, 
    99, 92, 82, 59, 52, 64, 67, 44, 36, 41, 69, 89, 95, 82, 60, 
    79, 73, 70, 69, 66, 60, 50, 46, 60, 55, 60, 80, 97, 95, 72, 
    77, 71, 48, 59, 58, 58, 62, 55, 71, 57, 66, 83, 94, 109, 102, 
    73, 61, 56, 64, 82, 61, 65, 53, 47, 58, 49, 18, 59, 80, 83, 
    77, 55, 81, 74, 85, 104, 89, 70, 41, 49, 62, 48, 11, 25, 54, 
    92, 81, 76, 73, 63, 51, 66, 94, 82, 61, 47, 48, 65, 60, 29, 
    85, 72, 69, 86, 86, 67, 51, 57, 73, 49, 41, 62, 57, 50, 42, 
    78, 75, 67, 80, 74, 62, 75, 71, 64, 51, 51, 49, 56, 56, 49, 
    77, 70, 64, 74, 54, 23, 55, 53, 45, 38, 40, 42, 31, 36, 48, 
    72, 64, 54, 75, 86, 84, 55, 38, 33, 30, 40, 40, 36, 36, 52, 
    50, 62, 45, 61, 74, 62, 33, 30, 27, 29, 36, 42, 48, 43, 36, 
    
    -- channel=562
    0, 5, 10, 6, 10, 10, 10, 7, 6, 2, 0, 15, 11, 9, 8, 
    0, 4, 6, 0, 7, 14, 18, 14, 9, 1, 10, 11, 7, 7, 10, 
    2, 2, 0, 0, 2, 10, 0, 0, 0, 0, 11, 0, 6, 12, 14, 
    0, 0, 33, 15, 2, 6, 12, 5, 0, 4, 9, 5, 20, 20, 2, 
    17, 29, 9, 2, 0, 0, 12, 9, 1, 2, 7, 8, 5, 2, 0, 
    7, 7, 8, 1, 13, 13, 0, 0, 4, 2, 6, 1, 7, 6, 3, 
    5, 3, 4, 0, 0, 0, 4, 14, 13, 6, 0, 5, 4, 11, 11, 
    7, 8, 6, 3, 18, 11, 1, 17, 0, 8, 10, 19, 5, 9, 2, 
    4, 0, 4, 10, 6, 14, 5, 3, 4, 0, 10, 0, 0, 0, 4, 
    6, 12, 11, 8, 0, 1, 6, 4, 8, 3, 9, 0, 3, 13, 0, 
    6, 7, 0, 4, 10, 4, 0, 0, 10, 16, 0, 9, 8, 0, 9, 
    5, 4, 2, 11, 14, 13, 9, 6, 8, 0, 6, 6, 7, 9, 0, 
    6, 4, 3, 2, 1, 0, 1, 5, 1, 3, 3, 2, 5, 0, 2, 
    7, 4, 0, 5, 7, 23, 10, 0, 0, 0, 2, 0, 0, 0, 5, 
    2, 2, 0, 3, 4, 8, 11, 5, 1, 0, 1, 3, 0, 10, 1, 
    
    -- channel=563
    10, 0, 0, 0, 0, 0, 4, 0, 14, 25, 0, 0, 1, 2, 3, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 
    10, 3, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    46, 7, 0, 3, 0, 0, 9, 12, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 15, 0, 0, 0, 7, 0, 0, 0, 0, 0, 5, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 15, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 3, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 1, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 5, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 2, 0, 0, 
    
    -- channel=564
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 0, 0, 0, 0, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 2, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=565
    0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 
    0, 0, 8, 0, 1, 0, 0, 0, 0, 0, 13, 2, 0, 0, 0, 
    0, 0, 17, 0, 19, 0, 6, 14, 5, 0, 17, 19, 8, 5, 0, 
    0, 0, 0, 0, 26, 0, 0, 0, 0, 15, 15, 18, 9, 9, 20, 
    0, 0, 6, 0, 25, 19, 2, 0, 1, 14, 19, 23, 20, 4, 18, 
    4, 9, 7, 0, 10, 12, 6, 0, 0, 10, 20, 32, 21, 0, 6, 
    6, 7, 0, 4, 16, 23, 1, 0, 1, 11, 19, 30, 23, 7, 0, 
    4, 4, 0, 19, 0, 10, 6, 0, 12, 6, 8, 24, 27, 20, 15, 
    0, 10, 0, 16, 9, 6, 6, 0, 13, 0, 0, 0, 37, 23, 25, 
    2, 0, 9, 9, 25, 27, 16, 3, 0, 1, 0, 0, 0, 0, 16, 
    11, 2, 19, 12, 8, 4, 25, 20, 2, 0, 0, 0, 1, 0, 0, 
    15, 0, 22, 15, 11, 0, 7, 8, 5, 0, 0, 0, 3, 0, 0, 
    12, 4, 18, 20, 8, 13, 15, 7, 2, 0, 3, 0, 5, 1, 0, 
    8, 0, 15, 20, 0, 0, 3, 2, 0, 0, 0, 0, 0, 2, 0, 
    8, 0, 8, 26, 10, 3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    
    -- channel=566
    1, 0, 0, 0, 0, 0, 0, 0, 21, 45, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 61, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    55, 0, 0, 14, 0, 22, 24, 24, 0, 0, 0, 0, 0, 14, 0, 
    26, 0, 0, 41, 0, 0, 15, 37, 0, 0, 0, 0, 0, 38, 0, 
    0, 0, 4, 12, 0, 0, 24, 10, 0, 0, 0, 0, 0, 40, 0, 
    2, 0, 20, 0, 2, 0, 26, 0, 15, 0, 0, 0, 0, 15, 19, 
    10, 0, 40, 0, 10, 0, 6, 0, 0, 0, 0, 0, 0, 9, 0, 
    33, 0, 3, 0, 0, 1, 9, 49, 0, 0, 0, 16, 0, 0, 0, 
    21, 0, 0, 0, 0, 0, 0, 17, 23, 0, 19, 0, 0, 4, 0, 
    0, 16, 0, 0, 0, 29, 0, 0, 15, 25, 0, 0, 0, 11, 0, 
    0, 29, 0, 0, 2, 8, 0, 0, 6, 38, 0, 0, 0, 7, 10, 
    2, 17, 0, 0, 37, 0, 0, 0, 13, 13, 0, 0, 0, 0, 1, 
    8, 18, 0, 0, 30, 0, 8, 0, 7, 0, 0, 0, 10, 0, 0, 
    3, 9, 0, 0, 5, 14, 15, 0, 19, 0, 0, 0, 2, 0, 0, 
    
    -- channel=567
    7, 0, 3, 10, 7, 7, 9, 9, 12, 18, 0, 0, 6, 8, 10, 
    6, 0, 0, 4, 1, 6, 6, 4, 8, 28, 0, 7, 9, 8, 8, 
    6, 1, 0, 1, 0, 19, 4, 6, 15, 7, 0, 9, 10, 9, 10, 
    11, 0, 0, 17, 0, 12, 8, 6, 1, 0, 8, 0, 4, 16, 12, 
    24, 0, 13, 24, 0, 3, 12, 17, 3, 0, 2, 0, 15, 33, 15, 
    18, 12, 18, 22, 0, 3, 15, 13, 1, 0, 0, 0, 17, 35, 24, 
    20, 15, 18, 11, 6, 4, 13, 0, 5, 0, 3, 0, 16, 23, 21, 
    26, 13, 20, 0, 10, 4, 10, 5, 6, 4, 13, 4, 12, 23, 23, 
    32, 11, 6, 0, 10, 0, 4, 16, 0, 14, 9, 15, 0, 25, 8, 
    28, 13, 5, 8, 5, 10, 10, 9, 10, 4, 10, 8, 3, 6, 2, 
    20, 24, 4, 5, 8, 16, 0, 6, 15, 12, 13, 0, 3, 12, 9, 
    20, 31, 0, 6, 8, 10, 0, 6, 11, 22, 0, 7, 4, 13, 12, 
    23, 31, 7, 9, 16, 0, 2, 10, 16, 18, 3, 9, 7, 10, 8, 
    25, 33, 11, 8, 15, 0, 6, 12, 17, 12, 3, 9, 14, 0, 7, 
    27, 30, 13, 3, 13, 15, 18, 9, 17, 7, 6, 8, 10, 3, 6, 
    
    -- channel=568
    0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 26, 28, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 48, 19, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 39, 14, 
    0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 0, 0, 3, 0, 0, 0, 7, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 4, 4, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 11, 5, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=569
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=570
    1, 62, 18, 6, 4, 19, 8, 12, 0, 0, 53, 0, 6, 6, 5, 
    3, 41, 22, 23, 0, 0, 12, 7, 0, 0, 38, 0, 0, 2, 4, 
    4, 15, 39, 14, 2, 0, 0, 12, 5, 21, 0, 1, 0, 0, 0, 
    0, 18, 0, 0, 13, 0, 0, 0, 0, 27, 0, 11, 0, 0, 6, 
    0, 1, 0, 0, 9, 0, 0, 0, 3, 21, 2, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 2, 5, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 17, 0, 0, 2, 1, 0, 0, 0, 
    0, 4, 0, 19, 0, 0, 0, 0, 8, 1, 0, 21, 19, 0, 3, 
    0, 3, 0, 1, 0, 0, 0, 0, 20, 7, 0, 0, 19, 2, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 7, 11, 0, 10, 
    0, 0, 3, 0, 0, 0, 1, 0, 0, 0, 17, 1, 0, 0, 0, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 
    0, 0, 8, 0, 0, 30, 0, 0, 0, 0, 9, 4, 0, 9, 0, 
    0, 0, 17, 0, 0, 8, 0, 1, 0, 12, 3, 4, 0, 15, 3, 
    0, 0, 13, 0, 0, 0, 0, 8, 0, 20, 6, 2, 1, 3, 5, 
    
    -- channel=571
    5, 0, 22, 12, 12, 14, 13, 9, 8, 8, 0, 4, 12, 11, 16, 
    5, 0, 26, 8, 0, 0, 7, 2, 9, 15, 0, 0, 7, 10, 13, 
    5, 4, 10, 3, 0, 7, 12, 20, 26, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 1, 0, 2, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 1, 5, 9, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 14, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 12, 13, 3, 2, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 27, 0, 0, 0, 1, 1, 6, 0, 6, 2, 3, 0, 0, 
    0, 1, 13, 0, 0, 0, 0, 10, 0, 7, 9, 11, 8, 22, 0, 
    0, 0, 0, 0, 0, 5, 2, 0, 0, 4, 12, 16, 1, 4, 8, 
    0, 0, 0, 0, 0, 4, 2, 2, 7, 11, 14, 2, 5, 12, 9, 
    0, 1, 0, 0, 2, 6, 0, 0, 6, 17, 0, 6, 7, 8, 11, 
    0, 0, 0, 0, 20, 19, 10, 9, 16, 15, 8, 9, 13, 15, 9, 
    0, 1, 0, 0, 5, 0, 7, 17, 19, 12, 8, 10, 14, 7, 8, 
    3, 2, 0, 0, 0, 9, 17, 17, 20, 9, 9, 10, 9, 4, 11, 
    
    -- channel=572
    0, 0, 16, 16, 18, 15, 14, 15, 14, 5, 7, 26, 18, 17, 16, 
    0, 0, 20, 14, 32, 24, 25, 24, 28, 11, 18, 32, 27, 25, 23, 
    0, 0, 14, 12, 41, 31, 21, 25, 24, 15, 36, 36, 38, 37, 33, 
    0, 0, 28, 21, 40, 37, 19, 18, 17, 24, 42, 38, 48, 47, 38, 
    23, 24, 33, 17, 33, 41, 38, 24, 19, 23, 39, 43, 46, 33, 28, 
    31, 32, 34, 15, 36, 41, 33, 17, 23, 24, 36, 46, 48, 33, 24, 
    30, 28, 27, 25, 28, 28, 34, 26, 34, 31, 32, 44, 48, 44, 30, 
    31, 28, 19, 37, 39, 37, 35, 27, 29, 28, 32, 43, 41, 49, 34, 
    29, 24, 28, 37, 39, 43, 36, 33, 24, 17, 31, 7, 29, 33, 35, 
    33, 26, 37, 36, 40, 47, 43, 35, 19, 24, 28, 18, 13, 26, 24, 
    38, 30, 37, 38, 39, 34, 36, 39, 38, 30, 13, 22, 26, 21, 20, 
    37, 31, 36, 46, 45, 35, 33, 34, 35, 18, 17, 24, 29, 21, 14, 
    35, 29, 30, 43, 40, 15, 36, 31, 29, 16, 19, 20, 27, 19, 18, 
    33, 23, 23, 44, 37, 19, 32, 22, 18, 9, 18, 15, 14, 14, 20, 
    26, 22, 18, 43, 38, 33, 22, 17, 13, 5, 14, 16, 11, 16, 19, 
    
    -- channel=573
    9, 0, 10, 26, 15, 23, 26, 24, 27, 26, 2, 15, 28, 29, 31, 
    9, 0, 0, 24, 7, 12, 12, 12, 16, 42, 0, 13, 21, 23, 26, 
    10, 3, 0, 17, 0, 16, 12, 4, 11, 19, 0, 4, 9, 10, 15, 
    26, 19, 0, 18, 0, 16, 17, 17, 11, 0, 0, 0, 6, 7, 6, 
    25, 0, 8, 32, 0, 2, 11, 20, 5, 0, 3, 0, 7, 23, 3, 
    13, 8, 10, 23, 0, 3, 11, 21, 0, 0, 0, 0, 4, 18, 12, 
    13, 13, 23, 5, 6, 7, 10, 10, 7, 0, 2, 0, 4, 10, 18, 
    14, 10, 28, 0, 10, 0, 15, 0, 7, 12, 1, 4, 0, 4, 9, 
    15, 11, 22, 2, 7, 3, 7, 18, 9, 19, 9, 18, 0, 9, 0, 
    15, 11, 3, 9, 1, 0, 3, 16, 11, 8, 19, 17, 17, 14, 2, 
    8, 11, 0, 7, 7, 14, 0, 4, 16, 14, 21, 11, 9, 22, 15, 
    6, 15, 0, 3, 4, 24, 4, 10, 10, 32, 7, 14, 7, 18, 21, 
    9, 16, 0, 1, 11, 27, 4, 13, 19, 23, 7, 17, 10, 17, 16, 
    12, 16, 3, 0, 20, 14, 17, 16, 21, 25, 10, 15, 21, 10, 14, 
    14, 13, 8, 0, 10, 11, 23, 16, 23, 11, 15, 13, 21, 11, 13, 
    
    -- channel=574
    0, 0, 50, 44, 41, 45, 46, 41, 37, 21, 14, 47, 55, 52, 54, 
    0, 0, 45, 37, 35, 34, 43, 42, 47, 30, 17, 45, 51, 53, 57, 
    0, 0, 22, 33, 41, 40, 31, 41, 45, 25, 29, 39, 47, 47, 45, 
    0, 0, 18, 36, 41, 41, 27, 26, 23, 25, 42, 38, 50, 49, 39, 
    27, 22, 33, 29, 31, 43, 45, 34, 25, 24, 35, 40, 47, 34, 27, 
    35, 32, 38, 30, 36, 43, 42, 24, 24, 23, 34, 41, 44, 34, 20, 
    33, 34, 43, 44, 31, 28, 38, 28, 31, 27, 29, 40, 44, 42, 24, 
    32, 38, 55, 47, 40, 38, 34, 37, 35, 26, 39, 44, 47, 49, 32, 
    31, 28, 51, 42, 41, 39, 34, 39, 26, 34, 42, 29, 32, 44, 35, 
    29, 25, 43, 43, 37, 48, 47, 35, 32, 37, 42, 39, 31, 39, 36, 
    33, 31, 37, 42, 42, 40, 38, 44, 46, 45, 30, 35, 41, 38, 36, 
    33, 31, 32, 49, 53, 50, 41, 43, 46, 37, 29, 37, 42, 38, 30, 
    31, 26, 25, 44, 55, 43, 51, 46, 45, 35, 32, 34, 39, 35, 33, 
    32, 24, 18, 42, 43, 45, 45, 43, 39, 24, 30, 30, 29, 26, 34, 
    27, 23, 13, 40, 42, 45, 41, 39, 33, 21, 26, 30, 25, 29, 32, 
    
    -- channel=575
    0, 88, 25, 0, 0, 6, 0, 5, 0, 0, 61, 18, 2, 2, 0, 
    1, 53, 53, 4, 0, 0, 6, 10, 0, 0, 99, 1, 0, 0, 0, 
    0, 19, 82, 19, 27, 0, 0, 15, 0, 0, 54, 8, 0, 0, 0, 
    0, 43, 86, 0, 39, 0, 0, 0, 7, 54, 4, 33, 0, 0, 5, 
    0, 38, 2, 0, 55, 0, 0, 0, 8, 33, 20, 39, 0, 0, 20, 
    0, 5, 0, 0, 30, 0, 0, 0, 12, 30, 20, 43, 0, 0, 0, 
    0, 0, 0, 7, 0, 4, 0, 10, 0, 16, 17, 44, 0, 0, 0, 
    0, 0, 0, 58, 0, 0, 0, 2, 2, 8, 0, 25, 15, 0, 0, 
    0, 3, 0, 41, 0, 1, 0, 0, 37, 0, 1, 0, 50, 0, 34, 
    0, 1, 8, 0, 9, 0, 0, 0, 0, 18, 0, 0, 8, 0, 22, 
    0, 0, 17, 0, 0, 0, 24, 2, 0, 0, 0, 15, 7, 0, 0, 
    0, 0, 37, 0, 0, 0, 16, 0, 0, 0, 32, 0, 8, 0, 0, 
    0, 0, 26, 0, 0, 0, 18, 0, 0, 0, 20, 0, 0, 0, 0, 
    0, 0, 26, 8, 0, 7, 0, 0, 0, 0, 14, 0, 0, 20, 3, 
    0, 0, 16, 22, 0, 0, 0, 0, 0, 15, 2, 3, 0, 15, 2, 
    
    -- channel=576
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=577
    9, 8, 6, 11, 8, 9, 16, 15, 9, 10, 10, 9, 16, 20, 19, 
    4, 4, 8, 4, 0, 0, 0, 0, 0, 0, 8, 3, 7, 16, 16, 
    0, 0, 5, 1, 0, 0, 0, 0, 0, 0, 0, 7, 8, 13, 13, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 8, 23, 13, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 17, 
    0, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 14, 0, 5, 0, 0, 0, 1, 13, 15, 15, 17, 5, 0, 0, 
    3, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 3, 0, 0, 0, 9, 7, 4, 0, 0, 
    0, 0, 0, 0, 0, 3, 6, 4, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 6, 0, 0, 
    
    -- channel=578
    0, 0, 0, 0, 2, 4, 13, 15, 5, 0, 0, 0, 1, 5, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 3, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 9, 5, 9, 13, 17, 11, 1, 0, 0, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 1, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 10, 1, 2, 4, 0, 3, 7, 7, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 13, 11, 5, 28, 14, 7, 4, 8, 0, 
    0, 0, 0, 0, 0, 5, 13, 12, 14, 0, 0, 0, 6, 6, 0, 
    0, 0, 0, 0, 0, 6, 7, 5, 2, 0, 0, 0, 5, 5, 0, 
    
    -- channel=579
    11, 14, 11, 6, 6, 7, 6, 12, 16, 10, 10, 10, 4, 12, 3, 
    15, 16, 10, 3, 21, 27, 31, 28, 22, 15, 10, 16, 11, 2, 9, 
    17, 18, 8, 0, 34, 36, 34, 32, 40, 44, 26, 13, 10, 0, 18, 
    17, 15, 16, 0, 42, 20, 24, 37, 31, 32, 34, 24, 4, 0, 7, 
    17, 13, 15, 9, 38, 43, 28, 38, 37, 39, 28, 30, 15, 1, 10, 
    20, 8, 2, 11, 36, 34, 35, 33, 32, 38, 33, 31, 33, 17, 17, 
    19, 3, 11, 2, 31, 34, 23, 26, 29, 23, 17, 32, 33, 24, 16, 
    2, 1, 10, 1, 31, 23, 34, 22, 17, 17, 19, 17, 28, 40, 36, 
    2, 0, 18, 0, 24, 15, 6, 0, 13, 15, 0, 8, 30, 21, 35, 
    5, 0, 10, 2, 26, 16, 31, 35, 18, 38, 28, 30, 28, 18, 49, 
    12, 0, 13, 7, 14, 16, 19, 18, 26, 24, 24, 27, 23, 17, 43, 
    19, 0, 10, 12, 0, 16, 30, 0, 35, 0, 11, 25, 0, 25, 45, 
    22, 0, 25, 15, 2, 5, 6, 9, 17, 24, 3, 0, 2, 13, 50, 
    27, 17, 11, 8, 14, 0, 6, 11, 13, 35, 30, 0, 0, 24, 44, 
    25, 23, 14, 11, 14, 3, 9, 12, 16, 20, 26, 0, 3, 21, 49, 
    
    -- channel=580
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=581
    15, 17, 14, 0, 11, 10, 12, 19, 32, 23, 18, 24, 0, 13, 0, 
    25, 26, 18, 0, 22, 32, 26, 32, 44, 33, 20, 31, 23, 2, 24, 
    28, 29, 13, 0, 20, 14, 8, 2, 11, 20, 39, 31, 13, 0, 30, 
    28, 26, 11, 0, 52, 38, 15, 27, 22, 22, 26, 45, 8, 0, 9, 
    30, 22, 7, 0, 45, 32, 11, 28, 31, 28, 19, 46, 33, 1, 0, 
    37, 18, 0, 0, 28, 19, 13, 20, 20, 25, 30, 34, 51, 28, 29, 
    30, 0, 6, 0, 10, 19, 11, 5, 20, 24, 2, 33, 54, 44, 39, 
    17, 0, 17, 0, 6, 0, 0, 0, 7, 5, 0, 12, 31, 30, 67, 
    0, 0, 32, 0, 13, 13, 2, 0, 0, 0, 0, 0, 13, 14, 68, 
    3, 0, 24, 0, 19, 0, 12, 25, 13, 21, 12, 16, 28, 0, 59, 
    15, 0, 0, 0, 0, 2, 3, 0, 23, 0, 0, 12, 0, 8, 43, 
    18, 0, 13, 0, 0, 0, 22, 0, 39, 0, 10, 32, 0, 21, 43, 
    20, 0, 0, 13, 0, 0, 0, 0, 0, 48, 12, 0, 0, 0, 52, 
    24, 14, 0, 7, 0, 0, 0, 0, 1, 44, 24, 0, 0, 11, 45, 
    19, 11, 0, 0, 0, 0, 0, 0, 0, 3, 19, 0, 0, 6, 52, 
    
    -- channel=582
    0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 10, 
    0, 0, 0, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 
    0, 0, 8, 86, 0, 0, 0, 4, 0, 0, 0, 0, 0, 14, 0, 
    0, 0, 2, 82, 0, 0, 19, 0, 0, 0, 0, 0, 0, 11, 0, 
    0, 0, 31, 56, 0, 0, 8, 0, 0, 0, 0, 0, 0, 12, 0, 
    0, 4, 33, 63, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 23, 2, 34, 0, 0, 8, 2, 0, 0, 9, 0, 0, 0, 0, 
    0, 49, 0, 28, 3, 5, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    10, 69, 0, 58, 0, 0, 5, 29, 0, 0, 28, 2, 0, 0, 0, 
    10, 84, 0, 50, 0, 11, 0, 0, 3, 0, 0, 0, 0, 27, 0, 
    0, 97, 0, 15, 9, 0, 0, 32, 0, 7, 0, 0, 25, 0, 0, 
    0, 104, 0, 0, 47, 0, 0, 41, 0, 5, 0, 0, 73, 0, 0, 
    0, 59, 0, 0, 33, 27, 1, 0, 0, 0, 3, 46, 38, 0, 0, 
    0, 5, 28, 0, 0, 42, 1, 0, 0, 0, 0, 42, 33, 0, 0, 
    0, 0, 17, 24, 0, 19, 3, 0, 0, 0, 0, 14, 33, 0, 0, 
    
    -- channel=583
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=584
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=585
    25, 27, 24, 18, 13, 20, 26, 32, 32, 25, 22, 19, 24, 21, 19, 
    32, 32, 26, 29, 28, 30, 30, 25, 20, 18, 12, 17, 19, 14, 10, 
    32, 31, 29, 37, 48, 62, 66, 68, 61, 46, 20, 21, 19, 7, 5, 
    32, 32, 29, 41, 47, 52, 68, 68, 67, 64, 53, 11, 17, 12, 11, 
    29, 29, 37, 39, 54, 60, 56, 66, 63, 66, 59, 33, 30, 27, 25, 
    22, 24, 31, 50, 41, 55, 58, 57, 55, 55, 50, 44, 27, 32, 32, 
    20, 17, 15, 27, 61, 60, 59, 53, 51, 52, 39, 32, 23, 19, 27, 
    12, 11, 2, 31, 49, 43, 38, 32, 25, 27, 23, 21, 29, 40, 26, 
    17, 23, 12, 14, 30, 28, 38, 42, 35, 41, 46, 39, 47, 46, 34, 
    23, 26, 6, 19, 27, 28, 31, 25, 38, 36, 36, 35, 33, 33, 34, 
    24, 27, 17, 20, 20, 18, 37, 38, 24, 37, 33, 37, 35, 30, 43, 
    36, 29, 9, 29, 27, 18, 14, 8, 14, 18, 31, 25, 19, 19, 27, 
    43, 40, 42, 29, 27, 18, 9, 12, 16, 22, 42, 34, 20, 16, 43, 
    43, 41, 37, 26, 28, 19, 11, 13, 20, 27, 25, 23, 12, 20, 43, 
    47, 47, 39, 28, 25, 18, 17, 18, 21, 24, 27, 18, 18, 20, 42, 
    
    -- channel=586
    0, 0, 0, 0, 7, 0, 0, 0, 7, 10, 8, 18, 0, 1, 0, 
    5, 5, 1, 0, 18, 28, 28, 42, 56, 48, 27, 25, 18, 6, 27, 
    10, 11, 0, 0, 0, 0, 0, 0, 0, 0, 44, 17, 5, 8, 48, 
    9, 7, 0, 0, 18, 0, 0, 0, 0, 0, 0, 55, 3, 0, 11, 
    14, 4, 0, 0, 9, 0, 0, 0, 0, 0, 0, 28, 16, 0, 0, 
    33, 6, 0, 0, 11, 0, 0, 0, 0, 0, 4, 14, 44, 9, 10, 
    21, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 22, 57, 54, 28, 
    11, 0, 25, 0, 0, 0, 0, 0, 1, 0, 0, 13, 31, 13, 67, 
    0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 55, 
    0, 0, 35, 0, 10, 0, 2, 24, 0, 10, 2, 7, 19, 0, 46, 
    1, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 16, 
    0, 0, 22, 0, 0, 0, 32, 0, 42, 1, 0, 21, 0, 22, 40, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 0, 0, 0, 0, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 26, 0, 0, 4, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 24, 
    
    -- channel=587
    24, 22, 23, 23, 21, 20, 21, 24, 19, 22, 21, 20, 25, 16, 21, 
    27, 26, 26, 36, 28, 32, 34, 31, 28, 21, 19, 18, 19, 17, 15, 
    28, 28, 28, 47, 40, 43, 51, 49, 42, 35, 24, 14, 20, 16, 9, 
    28, 27, 31, 50, 40, 42, 51, 58, 56, 53, 30, 20, 20, 19, 9, 
    26, 28, 36, 56, 36, 49, 57, 53, 52, 55, 48, 23, 21, 23, 24, 
    23, 27, 42, 47, 31, 47, 53, 49, 45, 47, 44, 28, 25, 28, 27, 
    17, 23, 22, 41, 46, 48, 51, 46, 47, 41, 37, 31, 21, 30, 24, 
    13, 24, 18, 25, 46, 37, 40, 41, 30, 28, 34, 26, 23, 36, 19, 
    22, 34, 5, 29, 33, 33, 33, 27, 29, 30, 26, 24, 28, 37, 13, 
    25, 40, 7, 39, 18, 32, 26, 41, 25, 39, 37, 34, 34, 39, 26, 
    26, 43, 15, 26, 25, 23, 29, 33, 19, 34, 32, 27, 35, 36, 24, 
    33, 44, 16, 27, 27, 20, 20, 31, 16, 26, 24, 23, 40, 12, 33, 
    36, 48, 28, 22, 34, 23, 16, 16, 19, 21, 25, 29, 25, 19, 26, 
    39, 36, 40, 23, 30, 27, 16, 17, 21, 7, 34, 31, 28, 18, 30, 
    41, 42, 38, 28, 26, 24, 19, 20, 21, 23, 25, 25, 23, 18, 31, 
    
    -- channel=588
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=589
    0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 4, 0, 0, 1, 
    2, 2, 0, 10, 17, 21, 25, 30, 28, 20, 10, 1, 1, 0, 1, 
    4, 4, 5, 0, 19, 8, 12, 7, 12, 17, 14, 0, 0, 1, 7, 
    4, 1, 9, 7, 19, 20, 11, 30, 22, 25, 8, 12, 4, 0, 0, 
    5, 2, 10, 25, 17, 25, 31, 28, 27, 28, 21, 10, 0, 0, 0, 
    8, 3, 6, 6, 26, 23, 20, 26, 28, 25, 30, 25, 12, 4, 4, 
    1, 6, 5, 13, 8, 19, 24, 20, 22, 20, 19, 19, 22, 27, 10, 
    0, 7, 10, 0, 19, 15, 14, 13, 22, 25, 19, 24, 32, 22, 17, 
    0, 0, 0, 21, 17, 11, 15, 2, 0, 0, 0, 0, 0, 5, 21, 
    0, 0, 8, 8, 12, 14, 14, 26, 17, 22, 24, 22, 17, 22, 23, 
    2, 2, 0, 4, 4, 17, 6, 0, 21, 3, 9, 3, 7, 11, 15, 
    8, 4, 14, 0, 0, 2, 20, 25, 13, 20, 5, 5, 21, 13, 30, 
    15, 0, 0, 1, 7, 0, 4, 5, 10, 3, 0, 0, 6, 12, 10, 
    8, 12, 9, 3, 10, 3, 0, 3, 3, 13, 28, 7, 8, 6, 20, 
    17, 15, 7, 11, 9, 7, 1, 2, 4, 7, 12, 14, 1, 6, 16, 
    
    -- channel=590
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 17, 15, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 31, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 22, 0, 0, 
    0, 0, 0, 0, 0, 7, 37, 22, 24, 17, 27, 27, 22, 24, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 27, 0, 49, 13, 0, 35, 18, 20, 0, 1, 17, 
    0, 0, 3, 0, 19, 0, 0, 30, 1, 16, 8, 0, 38, 0, 13, 
    0, 0, 0, 0, 0, 28, 75, 0, 50, 0, 0, 16, 0, 55, 14, 
    0, 0, 0, 0, 0, 0, 1, 4, 9, 0, 0, 0, 0, 0, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 7, 0, 0, 11, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 10, 20, 0, 0, 7, 1, 
    
    -- channel=591
    27, 26, 30, 4, 23, 27, 29, 35, 34, 27, 21, 28, 23, 13, 12, 
    37, 36, 31, 3, 32, 41, 27, 27, 37, 29, 15, 30, 25, 6, 20, 
    37, 37, 29, 8, 54, 56, 54, 52, 45, 36, 32, 33, 18, 5, 7, 
    37, 37, 26, 14, 65, 59, 51, 63, 63, 58, 37, 34, 25, 10, 3, 
    37, 35, 16, 27, 64, 51, 52, 60, 59, 58, 60, 42, 42, 30, 25, 
    39, 30, 29, 18, 35, 52, 45, 49, 48, 53, 45, 44, 49, 37, 38, 
    33, 14, 15, 25, 47, 48, 58, 44, 50, 53, 29, 30, 34, 31, 48, 
    25, 0, 30, 24, 38, 30, 20, 18, 18, 21, 15, 20, 39, 41, 60, 
    23, 0, 31, 0, 43, 24, 42, 28, 31, 31, 36, 26, 39, 36, 49, 
    29, 0, 23, 0, 22, 20, 18, 28, 39, 32, 31, 32, 40, 15, 47, 
    32, 0, 13, 14, 0, 13, 37, 2, 37, 17, 28, 43, 0, 50, 32, 
    41, 0, 23, 34, 0, 1, 8, 5, 17, 30, 36, 28, 2, 14, 38, 
    47, 35, 19, 38, 16, 0, 0, 3, 5, 60, 41, 30, 0, 16, 44, 
    46, 39, 29, 30, 24, 1, 0, 4, 17, 27, 33, 21, 0, 18, 46, 
    45, 45, 34, 6, 21, 7, 4, 8, 11, 18, 26, 23, 0, 17, 56, 
    
    -- channel=592
    6, 2, 5, 0, 1, 12, 18, 20, 10, 3, 0, 0, 6, 2, 0, 
    9, 8, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 6, 5, 0, 30, 41, 42, 39, 29, 9, 2, 7, 0, 0, 0, 
    6, 3, 2, 5, 39, 40, 26, 34, 42, 49, 12, 0, 1, 1, 0, 
    5, 5, 0, 3, 32, 20, 20, 36, 34, 29, 32, 22, 7, 10, 18, 
    0, 0, 9, 13, 15, 26, 28, 24, 22, 22, 23, 12, 12, 6, 6, 
    0, 0, 0, 15, 36, 32, 34, 30, 33, 30, 10, 1, 0, 0, 2, 
    0, 0, 6, 1, 11, 14, 15, 9, 3, 4, 4, 0, 2, 5, 14, 
    7, 0, 0, 0, 21, 19, 26, 35, 45, 46, 46, 43, 40, 32, 16, 
    4, 0, 0, 0, 6, 1, 0, 6, 0, 0, 0, 0, 5, 0, 14, 
    4, 1, 5, 1, 0, 8, 28, 6, 8, 13, 13, 24, 11, 24, 19, 
    8, 0, 9, 23, 7, 0, 0, 0, 4, 1, 18, 5, 0, 0, 8, 
    19, 31, 22, 13, 11, 3, 0, 0, 5, 40, 32, 19, 0, 8, 19, 
    21, 15, 13, 12, 11, 4, 2, 5, 8, 0, 0, 0, 0, 7, 21, 
    18, 21, 18, 6, 8, 7, 4, 5, 5, 6, 4, 12, 0, 5, 25, 
    
    -- channel=593
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 23, 27, 37, 49, 43, 25, 4, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    0, 0, 0, 7, 0, 0, 0, 3, 0, 0, 0, 10, 0, 0, 0, 
    0, 0, 16, 32, 0, 8, 22, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 16, 5, 2, 13, 18, 13, 17, 10, 0, 0, 0, 
    0, 17, 17, 0, 0, 0, 0, 0, 0, 0, 9, 13, 30, 32, 0, 
    0, 34, 0, 0, 18, 13, 9, 18, 35, 35, 27, 38, 35, 19, 0, 
    0, 0, 0, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 11, 14, 14, 4, 17, 21, 24, 22, 29, 37, 32, 22, 31, 0, 
    0, 0, 0, 0, 5, 7, 0, 0, 15, 0, 3, 0, 0, 0, 0, 
    0, 31, 3, 0, 0, 5, 40, 44, 0, 17, 0, 0, 45, 24, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 12, 36, 18, 10, 0, 0, 
    1, 0, 0, 5, 1, 0, 0, 0, 0, 0, 11, 11, 0, 0, 0, 
    
    -- channel=594
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 18, 9, 11, 15, 14, 8, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 10, 7, 12, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 10, 23, 19, 6, 4, 8, 0, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 27, 14, 9, 4, 0, 0, 0, 0, 9, 0, 
    0, 0, 0, 0, 2, 24, 34, 33, 28, 0, 0, 0, 15, 23, 0, 
    0, 0, 0, 0, 0, 12, 33, 29, 11, 0, 0, 0, 24, 22, 0, 
    0, 0, 0, 0, 4, 11, 24, 23, 20, 11, 0, 0, 23, 24, 0, 
    
    -- channel=595
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 11, 13, 17, 12, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 18, 12, 6, 10, 10, 14, 12, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 0, 0, 9, 7, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 21, 7, 14, 14, 10, 6, 9, 0, 0, 0, 0, 0, 
    0, 0, 1, 20, 22, 18, 16, 17, 17, 14, 6, 4, 0, 0, 0, 
    0, 5, 14, 12, 12, 15, 13, 17, 11, 5, 15, 11, 5, 0, 0, 
    2, 29, 5, 12, 24, 27, 26, 21, 24, 27, 21, 22, 27, 19, 0, 
    0, 15, 7, 33, 10, 6, 6, 6, 0, 0, 0, 0, 0, 3, 0, 
    0, 21, 11, 26, 19, 24, 27, 16, 22, 22, 22, 22, 10, 26, 5, 
    0, 13, 14, 19, 24, 20, 11, 20, 18, 19, 18, 8, 21, 7, 7, 
    4, 27, 10, 5, 17, 23, 25, 25, 12, 11, 2, 4, 31, 21, 16, 
    6, 4, 6, 6, 15, 16, 18, 19, 19, 0, 0, 0, 22, 18, 11, 
    3, 7, 12, 7, 14, 16, 16, 14, 11, 18, 16, 9, 22, 17, 13, 
    9, 8, 7, 18, 14, 16, 16, 16, 17, 18, 19, 11, 21, 17, 8, 
    
    -- channel=596
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 16, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 
    
    -- channel=597
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=598
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 8, 0, 0, 13, 0, 0, 0, 0, 11, 0, 0, 
    0, 3, 0, 0, 5, 10, 9, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 6, 3, 1, 0, 0, 0, 14, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 2, 0, 0, 0, 0, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 
    
    -- channel=599
    76, 70, 84, 73, 55, 49, 53, 54, 66, 81, 78, 70, 82, 66, 69, 
    83, 82, 100, 82, 56, 47, 38, 53, 59, 60, 64, 65, 77, 89, 54, 
    85, 84, 98, 108, 27, 49, 43, 57, 49, 37, 25, 70, 85, 83, 34, 
    85, 95, 74, 122, 14, 50, 81, 64, 65, 49, 55, 45, 76, 86, 47, 
    81, 97, 83, 86, 34, 39, 68, 52, 54, 47, 77, 32, 64, 98, 59, 
    60, 103, 70, 89, 10, 39, 52, 46, 48, 43, 50, 34, 43, 85, 84, 
    54, 88, 49, 59, 22, 40, 61, 40, 28, 52, 41, 15, 36, 46, 76, 
    71, 63, 2, 84, 41, 45, 31, 44, 25, 19, 28, 17, 0, 18, 34, 
    69, 61, 19, 56, 15, 23, 32, 47, 22, 6, 66, 30, 13, 44, 0, 
    80, 84, 29, 26, 8, 33, 13, 0, 63, 36, 55, 45, 56, 47, 0, 
    68, 94, 24, 31, 12, 0, 4, 52, 0, 49, 38, 24, 42, 26, 0, 
    72, 100, 5, 35, 43, 1, 0, 45, 0, 36, 42, 43, 49, 24, 0, 
    61, 87, 20, 64, 47, 28, 2, 0, 0, 0, 64, 113, 28, 0, 0, 
    56, 76, 71, 66, 33, 46, 1, 0, 0, 10, 31, 116, 18, 0, 0, 
    63, 61, 77, 46, 30, 30, 8, 8, 6, 11, 16, 70, 20, 0, 0, 
    
    -- channel=600
    8, 8, 10, 13, 3, 10, 5, 3, 9, 9, 9, 8, 3, 5, 0, 
    16, 16, 15, 20, 27, 31, 40, 39, 30, 19, 7, 11, 10, 4, 0, 
    20, 20, 16, 20, 37, 43, 42, 41, 46, 46, 16, 8, 13, 1, 4, 
    20, 18, 24, 23, 42, 39, 46, 55, 50, 48, 44, 16, 8, 0, 4, 
    19, 18, 29, 35, 43, 57, 49, 56, 55, 56, 42, 28, 12, 2, 0, 
    20, 18, 18, 40, 48, 45, 55, 53, 53, 54, 52, 42, 25, 20, 19, 
    23, 21, 24, 21, 36, 53, 45, 45, 43, 40, 35, 35, 36, 30, 18, 
    12, 24, 10, 8, 48, 44, 46, 42, 38, 36, 38, 36, 37, 45, 28, 
    10, 14, 15, 29, 32, 28, 24, 16, 4, 10, 0, 1, 20, 35, 38, 
    15, 22, 12, 16, 30, 27, 37, 38, 36, 45, 44, 41, 33, 41, 41, 
    20, 14, 19, 14, 23, 22, 21, 34, 30, 35, 34, 26, 41, 21, 44, 
    30, 27, 8, 15, 17, 18, 36, 14, 29, 17, 18, 30, 22, 32, 38, 
    36, 11, 23, 21, 16, 13, 9, 11, 19, 5, 10, 7, 21, 13, 37, 
    36, 37, 30, 18, 24, 13, 6, 10, 11, 35, 37, 23, 11, 18, 40, 
    41, 37, 30, 29, 23, 14, 10, 13, 18, 25, 34, 20, 15, 16, 36, 
    
    -- channel=601
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 16, 35, 39, 45, 58, 58, 26, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 8, 0, 0, 8, 0, 0, 0, 16, 0, 0, 0, 
    0, 0, 23, 13, 10, 22, 18, 9, 12, 8, 0, 0, 0, 0, 0, 
    3, 5, 0, 0, 23, 4, 8, 22, 22, 15, 29, 14, 0, 0, 0, 
    4, 15, 17, 0, 0, 9, 13, 5, 13, 23, 13, 27, 45, 40, 0, 
    11, 21, 0, 0, 14, 0, 0, 16, 40, 31, 31, 50, 39, 25, 10, 
    0, 0, 8, 29, 1, 15, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 30, 0, 23, 9, 22, 34, 22, 27, 32, 27, 32, 16, 10, 
    0, 0, 0, 0, 2, 8, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    4, 6, 10, 0, 0, 9, 52, 20, 38, 18, 0, 35, 16, 35, 12, 
    1, 0, 0, 4, 0, 0, 2, 1, 0, 0, 0, 0, 3, 0, 0, 
    0, 6, 0, 8, 2, 0, 0, 0, 1, 38, 32, 11, 0, 2, 2, 
    7, 0, 0, 7, 5, 0, 0, 0, 0, 4, 20, 8, 0, 0, 0, 
    
    -- channel=602
    82, 79, 77, 61, 59, 70, 77, 84, 90, 87, 80, 81, 74, 78, 64, 
    93, 93, 86, 54, 54, 59, 62, 66, 70, 74, 70, 80, 81, 68, 73, 
    93, 93, 84, 31, 59, 69, 67, 65, 64, 64, 76, 85, 74, 54, 70, 
    93, 88, 79, 45, 80, 93, 79, 79, 79, 87, 78, 76, 75, 65, 56, 
    92, 87, 69, 41, 72, 74, 66, 77, 80, 81, 78, 91, 90, 77, 73, 
    86, 80, 57, 44, 53, 58, 62, 61, 60, 63, 72, 73, 91, 93, 93, 
    75, 60, 51, 41, 62, 68, 61, 55, 62, 69, 48, 58, 74, 83, 90, 
    62, 34, 50, 44, 50, 35, 37, 31, 29, 28, 26, 30, 43, 60, 95, 
    65, 36, 51, 27, 45, 56, 55, 47, 47, 60, 53, 47, 64, 68, 98, 
    68, 27, 40, 9, 42, 25, 34, 51, 51, 53, 50, 50, 57, 38, 81, 
    73, 31, 30, 20, 16, 28, 43, 30, 41, 39, 35, 48, 43, 43, 83, 
    74, 20, 34, 41, 19, 13, 29, 6, 47, 42, 53, 61, 10, 36, 61, 
    74, 39, 51, 49, 24, 12, 8, 12, 22, 71, 78, 45, 16, 22, 71, 
    75, 70, 47, 44, 36, 13, 10, 17, 28, 55, 54, 33, 5, 29, 69, 
    72, 67, 52, 38, 32, 20, 17, 19, 24, 32, 43, 35, 12, 26, 70, 
    
    -- channel=603
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 2, 14, 2, 13, 16, 8, 11, 19, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 19, 0, 12, 3, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 6, 18, 6, 0, 25, 1, 7, 10, 0, 0, 0, 
    0, 0, 15, 0, 0, 12, 20, 0, 19, 0, 0, 0, 0, 18, 12, 
    0, 0, 0, 0, 0, 0, 13, 15, 15, 1, 0, 0, 0, 16, 15, 
    0, 0, 0, 0, 0, 0, 11, 11, 6, 12, 0, 0, 0, 23, 11, 
    0, 0, 0, 0, 1, 0, 5, 7, 9, 10, 9, 0, 0, 21, 17, 
    
    -- channel=604
    7, 3, 10, 1, 8, 4, 4, 0, 0, 7, 2, 8, 6, 0, 3, 
    10, 9, 11, 6, 26, 32, 25, 31, 31, 21, 10, 7, 7, 2, 4, 
    12, 12, 16, 12, 43, 36, 34, 34, 37, 30, 24, 7, 2, 4, 2, 
    12, 14, 12, 30, 30, 27, 23, 47, 43, 37, 11, 22, 10, 0, 0, 
    12, 14, 13, 42, 39, 31, 48, 43, 39, 36, 42, 16, 7, 13, 0, 
    13, 14, 12, 22, 32, 41, 39, 39, 41, 41, 40, 24, 22, 12, 12, 
    6, 15, 8, 25, 20, 29, 42, 31, 31, 32, 19, 19, 23, 25, 16, 
    3, 4, 11, 3, 37, 34, 35, 29, 26, 29, 25, 21, 29, 29, 31, 
    0, 0, 0, 18, 28, 10, 15, 18, 5, 0, 6, 2, 0, 11, 11, 
    11, 4, 20, 8, 21, 25, 23, 23, 28, 35, 37, 37, 40, 26, 15, 
    12, 13, 3, 18, 9, 21, 20, 6, 34, 23, 30, 30, 15, 26, 0, 
    20, 14, 27, 14, 6, 6, 15, 31, 2, 18, 18, 10, 13, 26, 14, 
    28, 25, 0, 26, 22, 7, 9, 11, 9, 15, 0, 16, 5, 15, 5, 
    22, 28, 23, 28, 21, 15, 7, 7, 6, 16, 36, 38, 12, 9, 14, 
    30, 31, 29, 19, 21, 17, 9, 12, 13, 16, 19, 37, 4, 13, 16, 
    
    -- channel=605
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 13, 14, 12, 15, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    
    -- channel=606
    2, 4, 3, 0, 0, 3, 3, 4, 1, 0, 0, 0, 0, 0, 0, 
    2, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 1, 0, 9, 37, 46, 43, 44, 39, 19, 1, 0, 0, 0, 0, 
    1, 0, 2, 10, 27, 19, 24, 32, 36, 33, 14, 0, 0, 0, 0, 
    0, 0, 0, 13, 30, 22, 24, 32, 27, 28, 25, 10, 2, 7, 14, 
    0, 0, 9, 19, 21, 32, 30, 25, 25, 27, 17, 11, 7, 1, 1, 
    1, 0, 0, 15, 34, 30, 26, 27, 23, 17, 9, 5, 0, 0, 0, 
    0, 0, 4, 5, 27, 31, 31, 16, 4, 9, 6, 0, 9, 17, 7, 
    2, 2, 2, 0, 19, 4, 16, 29, 39, 36, 36, 40, 42, 17, 5, 
    4, 0, 0, 4, 13, 13, 14, 5, 11, 14, 10, 12, 10, 10, 16, 
    4, 3, 10, 12, 11, 12, 32, 15, 23, 26, 25, 37, 15, 21, 17, 
    9, 0, 8, 23, 11, 7, 0, 0, 0, 0, 15, 0, 0, 7, 13, 
    18, 28, 28, 15, 14, 9, 5, 8, 12, 19, 15, 10, 3, 13, 27, 
    19, 14, 14, 10, 13, 7, 10, 10, 8, 7, 6, 4, 3, 15, 25, 
    18, 21, 19, 9, 12, 8, 12, 14, 14, 14, 12, 7, 7, 16, 31, 
    
    -- channel=607
    92, 87, 94, 90, 65, 65, 68, 73, 80, 95, 93, 85, 101, 78, 86, 
    102, 101, 111, 109, 50, 42, 46, 52, 54, 63, 73, 73, 89, 99, 64, 
    104, 103, 112, 137, 25, 53, 59, 68, 47, 33, 27, 76, 96, 90, 37, 
    104, 108, 100, 133, 16, 70, 105, 76, 79, 69, 64, 45, 93, 95, 60, 
    101, 111, 102, 105, 25, 57, 83, 63, 66, 70, 83, 38, 83, 110, 81, 
    77, 114, 111, 103, 8, 45, 60, 55, 54, 51, 57, 49, 49, 105, 103, 
    68, 99, 64, 87, 38, 55, 70, 51, 41, 54, 53, 18, 29, 58, 92, 
    80, 85, 19, 87, 49, 48, 25, 42, 23, 18, 28, 17, 1, 29, 28, 
    90, 97, 18, 73, 17, 39, 59, 60, 34, 35, 74, 37, 26, 61, 14, 
    99, 112, 7, 55, 0, 35, 6, 9, 62, 36, 54, 42, 41, 64, 0, 
    85, 125, 23, 31, 14, 0, 14, 56, 0, 51, 36, 22, 51, 36, 2, 
    87, 124, 0, 38, 52, 0, 0, 49, 0, 52, 43, 36, 86, 0, 0, 
    78, 114, 29, 47, 54, 25, 0, 0, 0, 0, 83, 107, 38, 0, 0, 
    69, 86, 86, 47, 35, 47, 0, 0, 0, 0, 33, 95, 25, 0, 0, 
    76, 74, 78, 49, 25, 30, 5, 3, 3, 8, 16, 54, 27, 0, 0, 
    
    -- channel=608
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=609
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 68, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 67, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 44, 0, 0, 2, 0, 0, 0, 0, 0, 0, 7, 0, 
    0, 0, 15, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 26, 0, 17, 2, 20, 9, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 28, 0, 40, 0, 0, 0, 14, 0, 0, 11, 0, 0, 0, 0, 
    1, 48, 0, 26, 0, 8, 0, 0, 3, 0, 0, 0, 0, 15, 0, 
    0, 61, 0, 12, 2, 0, 0, 12, 0, 16, 7, 0, 13, 0, 0, 
    0, 65, 0, 0, 22, 0, 0, 34, 0, 0, 0, 0, 40, 0, 0, 
    0, 46, 0, 0, 22, 13, 0, 0, 0, 0, 0, 29, 14, 0, 0, 
    0, 0, 14, 0, 0, 26, 0, 0, 0, 0, 0, 44, 19, 0, 0, 
    0, 0, 11, 9, 0, 9, 0, 0, 0, 0, 0, 19, 13, 0, 0, 
    
    -- channel=610
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 20, 21, 23, 33, 46, 40, 31, 12, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 8, 3, 
    0, 0, 0, 12, 0, 0, 0, 3, 0, 0, 0, 8, 0, 0, 0, 
    0, 0, 19, 34, 0, 1, 23, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 15, 4, 0, 9, 15, 2, 14, 10, 0, 0, 0, 
    0, 19, 12, 6, 0, 0, 3, 0, 0, 0, 12, 11, 27, 38, 0, 
    0, 31, 0, 0, 14, 7, 0, 2, 27, 33, 12, 27, 35, 9, 0, 
    0, 0, 0, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 5, 14, 8, 6, 10, 11, 13, 25, 15, 28, 24, 13, 28, 0, 
    0, 10, 0, 0, 0, 12, 0, 0, 17, 0, 0, 0, 0, 0, 0, 
    0, 25, 12, 0, 0, 0, 23, 47, 0, 27, 0, 0, 47, 18, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 10, 30, 11, 10, 0, 0, 
    3, 0, 0, 10, 0, 1, 0, 0, 0, 0, 3, 16, 0, 0, 0, 
    
    -- channel=611
    0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 29, 23, 24, 45, 56, 38, 23, 12, 0, 0, 5, 0, 
    0, 0, 0, 11, 0, 0, 0, 0, 0, 15, 0, 0, 0, 9, 10, 
    0, 0, 8, 17, 0, 0, 0, 3, 0, 0, 0, 10, 0, 0, 3, 
    0, 0, 38, 28, 0, 18, 19, 3, 1, 5, 0, 0, 0, 0, 0, 
    1, 4, 0, 11, 31, 8, 9, 17, 24, 14, 26, 21, 0, 0, 0, 
    5, 31, 28, 0, 0, 0, 0, 0, 0, 0, 9, 17, 39, 36, 0, 
    6, 52, 0, 0, 24, 26, 29, 23, 39, 40, 27, 35, 35, 26, 0, 
    0, 1, 0, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 26, 16, 6, 20, 16, 36, 21, 30, 40, 45, 41, 25, 40, 2, 
    0, 8, 0, 0, 15, 13, 0, 15, 17, 17, 10, 0, 39, 0, 1, 
    3, 43, 1, 0, 0, 12, 49, 30, 6, 0, 0, 6, 33, 44, 9, 
    3, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 16, 0, 0, 
    0, 10, 0, 0, 0, 0, 0, 0, 0, 34, 36, 16, 9, 0, 0, 
    9, 0, 0, 22, 2, 0, 0, 0, 0, 5, 19, 10, 2, 0, 0, 
    
    -- channel=612
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=613
    15, 21, 10, 0, 0, 13, 29, 49, 24, 1, 0, 0, 25, 24, 18, 
    5, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 17, 0, 30, 37, 41, 14, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 8, 0, 4, 15, 11, 0, 0, 20, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 24, 62, 
    0, 0, 10, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 21, 0, 0, 0, 0, 7, 52, 103, 106, 105, 114, 87, 20, 0, 
    1, 5, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 16, 10, 0, 0, 0, 32, 21, 0, 9, 0, 23, 3, 7, 10, 
    0, 0, 0, 35, 29, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    0, 58, 63, 0, 13, 20, 0, 0, 1, 26, 49, 28, 0, 0, 14, 
    0, 0, 0, 0, 0, 10, 14, 11, 8, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 14, 11, 5, 0, 0, 0, 17, 0, 9, 
    
    -- channel=614
    0, 3, 0, 8, 1, 0, 0, 1, 2, 1, 6, 1, 1, 9, 8, 
    0, 0, 0, 4, 0, 0, 2, 1, 0, 6, 8, 4, 2, 12, 8, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 5, 4, 0, 5, 14, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 3, 0, 6, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 7, 3, 0, 0, 
    0, 8, 0, 0, 0, 0, 0, 6, 5, 3, 9, 9, 0, 1, 0, 
    0, 2, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 2, 15, 0, 6, 8, 7, 0, 0, 0, 0, 0, 1, 4, 
    0, 0, 8, 6, 14, 4, 0, 13, 0, 2, 2, 0, 4, 0, 2, 
    0, 10, 0, 0, 10, 19, 17, 7, 14, 0, 0, 5, 11, 4, 9, 
    0, 0, 5, 0, 3, 15, 16, 14, 11, 0, 0, 0, 13, 6, 3, 
    0, 0, 0, 0, 1, 9, 15, 13, 11, 3, 0, 0, 16, 8, 0, 
    0, 0, 0, 0, 4, 8, 12, 10, 9, 6, 3, 0, 15, 8, 0, 
    
    -- channel=615
    11, 11, 9, 10, 4, 5, 4, 6, 12, 13, 15, 14, 11, 17, 13, 
    10, 11, 11, 0, 0, 0, 0, 4, 6, 15, 15, 16, 15, 20, 16, 
    10, 10, 7, 0, 0, 0, 0, 0, 0, 0, 9, 14, 17, 19, 24, 
    10, 9, 5, 0, 0, 0, 0, 0, 0, 0, 2, 12, 12, 14, 17, 
    10, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 10, 9, 8, 
    10, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 10, 10, 
    10, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 7, 10, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    4, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=616
    70, 64, 70, 57, 51, 47, 52, 55, 61, 71, 67, 66, 72, 59, 64, 
    74, 73, 79, 61, 47, 47, 42, 50, 56, 59, 62, 61, 67, 71, 57, 
    75, 74, 77, 73, 40, 48, 47, 54, 48, 43, 44, 62, 66, 66, 43, 
    75, 78, 65, 81, 30, 51, 65, 63, 61, 54, 49, 53, 67, 66, 42, 
    72, 79, 63, 68, 38, 45, 63, 52, 53, 53, 70, 41, 63, 79, 58, 
    59, 78, 62, 58, 19, 43, 48, 44, 44, 46, 48, 40, 54, 75, 74, 
    47, 61, 38, 53, 29, 38, 53, 37, 35, 44, 36, 28, 40, 54, 72, 
    47, 41, 20, 50, 41, 37, 29, 34, 19, 18, 24, 16, 15, 32, 47, 
    53, 44, 18, 36, 25, 26, 35, 38, 29, 22, 50, 31, 23, 36, 23, 
    62, 54, 23, 28, 13, 30, 17, 16, 48, 39, 48, 43, 48, 40, 8, 
    58, 64, 19, 27, 11, 9, 20, 29, 17, 37, 35, 32, 27, 36, 3, 
    60, 62, 15, 34, 28, 4, 4, 36, 0, 37, 38, 32, 40, 17, 0, 
    55, 71, 20, 46, 39, 19, 5, 4, 0, 20, 52, 71, 18, 6, 0, 
    51, 59, 55, 44, 31, 32, 6, 4, 7, 14, 39, 73, 18, 0, 5, 
    56, 55, 58, 33, 27, 25, 12, 13, 12, 15, 19, 49, 15, 4, 8, 
    
    -- channel=617
    0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 
    0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 
    0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 18, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 25, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 30, 0, 0, 7, 0, 0, 13, 0, 0, 0, 0, 21, 0, 0, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 9, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 2, 12, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 
    
    -- channel=618
    115, 110, 121, 93, 95, 87, 86, 91, 110, 122, 118, 122, 108, 98, 91, 
    130, 130, 133, 82, 83, 87, 81, 98, 116, 112, 113, 124, 127, 112, 112, 
    136, 136, 129, 70, 50, 52, 46, 45, 48, 57, 90, 124, 120, 106, 100, 
    135, 137, 116, 84, 66, 86, 80, 75, 70, 63, 67, 122, 118, 103, 83, 
    136, 137, 103, 70, 65, 66, 77, 64, 71, 69, 82, 90, 122, 119, 94, 
    134, 137, 89, 50, 39, 54, 53, 54, 55, 62, 72, 74, 122, 136, 136, 
    118, 114, 89, 61, 31, 48, 56, 36, 44, 57, 42, 58, 102, 122, 140, 
    116, 75, 75, 81, 50, 37, 33, 35, 31, 27, 28, 31, 46, 64, 123, 
    102, 49, 73, 49, 43, 49, 46, 25, 20, 18, 32, 14, 33, 57, 90, 
    112, 52, 64, 15, 30, 30, 30, 49, 76, 69, 72, 69, 83, 46, 62, 
    113, 53, 30, 24, 4, 16, 23, 21, 44, 43, 42, 49, 31, 52, 42, 
    107, 46, 39, 40, 4, 1, 30, 28, 26, 59, 57, 74, 29, 42, 42, 
    94, 55, 23, 71, 25, 0, 0, 0, 0, 61, 75, 73, 3, 9, 34, 
    89, 92, 64, 64, 36, 10, 0, 0, 11, 55, 80, 80, 0, 10, 40, 
    86, 76, 67, 33, 31, 14, 1, 6, 11, 26, 45, 58, 0, 11, 48, 
    
    -- channel=619
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 9, 5, 8, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 0, 0, 0, 0, 1, 29, 0, 0, 0, 17, 
    0, 0, 0, 0, 35, 2, 0, 0, 0, 0, 0, 19, 0, 0, 0, 
    0, 0, 0, 0, 22, 8, 0, 0, 0, 1, 0, 23, 0, 0, 0, 
    5, 0, 0, 0, 27, 2, 0, 0, 0, 5, 3, 18, 25, 0, 0, 
    4, 0, 0, 0, 4, 0, 0, 0, 5, 0, 0, 25, 27, 17, 0, 
    0, 0, 30, 0, 0, 0, 0, 0, 6, 9, 0, 16, 39, 26, 42, 
    0, 0, 25, 0, 14, 4, 0, 0, 0, 0, 0, 0, 9, 0, 59, 
    0, 0, 16, 0, 20, 0, 17, 39, 0, 8, 0, 0, 1, 0, 78, 
    0, 0, 0, 0, 0, 19, 15, 0, 36, 0, 0, 12, 0, 4, 60, 
    0, 0, 24, 0, 0, 13, 37, 0, 60, 0, 0, 6, 0, 15, 84, 
    0, 0, 0, 0, 0, 0, 3, 10, 21, 51, 0, 0, 0, 20, 78, 
    0, 0, 0, 0, 0, 0, 0, 8, 20, 37, 15, 0, 0, 36, 65, 
    0, 0, 0, 0, 0, 0, 0, 1, 7, 11, 19, 0, 0, 28, 71, 
    
    -- channel=620
    7, 6, 10, 15, 6, 3, 0, 0, 2, 9, 11, 9, 5, 0, 1, 
    16, 15, 19, 39, 31, 34, 39, 42, 36, 20, 11, 8, 12, 9, 0, 
    20, 20, 23, 34, 18, 23, 26, 27, 31, 29, 7, 5, 14, 10, 0, 
    20, 22, 24, 44, 17, 24, 40, 45, 38, 31, 25, 13, 9, 2, 2, 
    19, 21, 43, 48, 24, 44, 50, 42, 41, 43, 36, 12, 10, 8, 0, 
    17, 26, 24, 37, 24, 33, 39, 42, 41, 38, 42, 29, 14, 20, 20, 
    15, 27, 22, 19, 21, 37, 41, 32, 31, 34, 26, 20, 26, 31, 17, 
    14, 27, 1, 19, 36, 23, 20, 24, 25, 22, 23, 25, 24, 34, 12, 
    11, 19, 0, 33, 11, 16, 15, 3, 0, 0, 0, 0, 0, 21, 11, 
    17, 32, 8, 16, 13, 22, 20, 26, 32, 35, 40, 35, 34, 34, 11, 
    19, 28, 0, 8, 8, 5, 0, 22, 7, 19, 15, 2, 25, 8, 11, 
    30, 41, 1, 0, 8, 4, 19, 20, 4, 17, 10, 21, 31, 15, 11, 
    31, 15, 2, 14, 12, 1, 0, 0, 0, 0, 4, 15, 11, 0, 5, 
    26, 31, 28, 16, 14, 7, 0, 0, 0, 15, 31, 29, 6, 0, 11, 
    34, 31, 25, 21, 11, 6, 0, 0, 1, 7, 17, 17, 3, 0, 3, 
    
    -- channel=621
    3, 0, 8, 14, 1, 0, 0, 0, 0, 0, 0, 0, 24, 0, 21, 
    0, 0, 11, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 
    0, 0, 20, 80, 0, 0, 0, 12, 0, 0, 0, 0, 4, 22, 0, 
    0, 2, 5, 83, 0, 0, 12, 0, 2, 0, 0, 0, 14, 21, 0, 
    0, 8, 12, 62, 0, 0, 16, 0, 0, 0, 14, 0, 0, 35, 8, 
    0, 14, 39, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 26, 0, 46, 0, 0, 17, 1, 0, 0, 4, 0, 0, 0, 0, 
    3, 29, 0, 27, 5, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 54, 0, 34, 0, 0, 10, 40, 8, 0, 48, 17, 0, 0, 0, 
    21, 62, 0, 38, 0, 13, 0, 0, 11, 0, 0, 0, 0, 19, 0, 
    2, 88, 0, 21, 0, 0, 0, 9, 0, 5, 1, 0, 0, 0, 0, 
    4, 84, 0, 9, 36, 0, 0, 51, 0, 14, 1, 0, 62, 0, 0, 
    0, 85, 0, 4, 41, 19, 0, 0, 0, 0, 9, 63, 20, 0, 0, 
    0, 11, 33, 9, 4, 43, 0, 0, 0, 0, 0, 67, 26, 0, 0, 
    0, 7, 29, 14, 0, 21, 2, 0, 0, 0, 0, 37, 20, 0, 0, 
    
    -- channel=622
    25, 27, 23, 1, 14, 25, 46, 63, 38, 16, 13, 10, 37, 28, 28, 
    20, 20, 17, 0, 0, 0, 0, 0, 0, 0, 0, 6, 5, 1, 12, 
    9, 9, 9, 21, 6, 28, 32, 31, 5, 0, 0, 18, 5, 0, 0, 
    9, 9, 0, 14, 11, 18, 18, 0, 14, 23, 0, 0, 11, 33, 0, 
    7, 11, 0, 0, 0, 0, 0, 0, 0, 0, 8, 1, 19, 38, 61, 
    0, 2, 23, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 9, 
    0, 0, 0, 16, 43, 1, 4, 2, 5, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 17, 2, 0, 3, 2, 23, 49, 94, 94, 106, 101, 76, 23, 0, 
    15, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 19, 10, 4, 0, 0, 29, 1, 0, 0, 0, 17, 0, 23, 0, 
    0, 0, 0, 43, 19, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 
    0, 65, 44, 6, 16, 11, 0, 0, 0, 52, 65, 53, 0, 1, 0, 
    7, 0, 5, 3, 0, 10, 10, 10, 12, 0, 0, 0, 0, 0, 0, 
    0, 2, 13, 0, 0, 3, 11, 9, 2, 0, 0, 0, 6, 0, 6, 
    
    -- channel=623
    74, 69, 75, 52, 50, 51, 55, 63, 71, 76, 69, 72, 70, 58, 54, 
    85, 84, 83, 46, 37, 42, 38, 45, 55, 58, 57, 71, 74, 62, 59, 
    87, 86, 81, 44, 30, 40, 39, 41, 35, 35, 47, 73, 70, 55, 44, 
    86, 86, 73, 51, 38, 61, 59, 54, 54, 51, 48, 63, 72, 60, 39, 
    86, 85, 59, 43, 35, 44, 49, 45, 49, 51, 62, 55, 78, 80, 65, 
    78, 82, 60, 34, 9, 33, 34, 32, 31, 37, 39, 43, 71, 87, 87, 
    66, 62, 42, 38, 25, 31, 40, 23, 26, 35, 22, 25, 47, 64, 86, 
    63, 31, 33, 41, 28, 19, 11, 9, 0, 0, 0, 0, 8, 34, 70, 
    61, 29, 30, 7, 20, 20, 29, 23, 21, 21, 35, 18, 25, 36, 51, 
    69, 28, 15, 0, 1, 6, 1, 17, 38, 32, 35, 32, 40, 21, 34, 
    68, 35, 5, 2, 0, 0, 11, 4, 11, 20, 18, 28, 9, 28, 26, 
    67, 25, 3, 21, 0, 0, 0, 0, 0, 24, 29, 30, 9, 0, 17, 
    60, 50, 14, 33, 11, 0, 0, 0, 0, 31, 54, 45, 0, 0, 15, 
    57, 56, 40, 26, 12, 0, 0, 0, 0, 11, 36, 42, 0, 0, 19, 
    54, 51, 42, 9, 5, 0, 0, 0, 0, 0, 12, 24, 0, 0, 24, 
    
    -- channel=624
    86, 84, 86, 75, 68, 60, 57, 58, 83, 96, 95, 97, 77, 78, 72, 
    99, 98, 96, 67, 70, 75, 83, 98, 105, 107, 101, 98, 100, 95, 91, 
    105, 106, 96, 40, 30, 28, 24, 23, 34, 58, 87, 92, 95, 88, 98, 
    105, 104, 93, 46, 45, 59, 51, 57, 47, 40, 65, 106, 89, 71, 75, 
    105, 102, 87, 47, 45, 59, 59, 49, 55, 57, 56, 79, 93, 81, 56, 
    105, 101, 57, 23, 43, 40, 38, 43, 48, 51, 63, 76, 103, 105, 105, 
    91, 87, 72, 30, 8, 33, 31, 24, 26, 38, 39, 59, 101, 113, 109, 
    79, 62, 55, 41, 37, 32, 29, 26, 32, 32, 26, 36, 51, 62, 106, 
    63, 28, 51, 51, 26, 32, 25, 4, 0, 0, 0, 0, 1, 34, 89, 
    75, 34, 52, 10, 28, 26, 38, 51, 62, 65, 67, 64, 67, 46, 69, 
    81, 27, 17, 12, 9, 18, 8, 15, 42, 31, 30, 31, 31, 23, 53, 
    77, 36, 30, 9, 0, 8, 45, 24, 33, 44, 33, 58, 30, 45, 56, 
    68, 13, 6, 41, 10, 0, 0, 0, 5, 29, 35, 25, 6, 7, 38, 
    63, 65, 39, 39, 23, 2, 0, 0, 6, 59, 75, 47, 1, 10, 44, 
    64, 54, 40, 29, 22, 8, 0, 2, 8, 21, 40, 34, 0, 10, 42, 
    
    -- channel=625
    102, 99, 94, 67, 66, 85, 102, 118, 105, 95, 87, 87, 108, 99, 93, 
    102, 103, 95, 41, 13, 8, 2, 0, 7, 35, 61, 79, 82, 77, 80, 
    94, 93, 88, 57, 39, 66, 68, 69, 49, 30, 55, 93, 80, 58, 55, 
    94, 89, 78, 53, 46, 73, 59, 40, 57, 72, 54, 47, 89, 98, 55, 
    91, 92, 39, 22, 31, 20, 25, 35, 39, 40, 58, 74, 94, 114, 129, 
    70, 75, 71, 39, 0, 22, 27, 9, 7, 15, 13, 26, 72, 95, 94, 
    62, 45, 28, 52, 59, 34, 26, 27, 30, 28, 20, 10, 10, 29, 81, 
    52, 13, 41, 51, 3, 13, 11, 0, 0, 0, 0, 0, 0, 6, 59, 
    85, 55, 35, 0, 23, 31, 48, 76, 114, 120, 124, 121, 99, 57, 48, 
    78, 33, 1, 12, 0, 2, 0, 0, 13, 2, 0, 0, 9, 6, 28, 
    72, 56, 31, 14, 0, 0, 48, 19, 0, 28, 19, 47, 24, 40, 43, 
    60, 16, 9, 62, 32, 0, 0, 0, 0, 19, 46, 19, 0, 0, 10, 
    53, 97, 67, 34, 32, 18, 0, 0, 7, 76, 103, 72, 5, 10, 33, 
    61, 48, 41, 28, 20, 21, 11, 13, 15, 0, 4, 27, 1, 7, 28, 
    45, 50, 53, 18, 12, 16, 18, 17, 13, 9, 1, 20, 15, 7, 42, 
    
    -- channel=626
    8, 8, 5, 7, 11, 21, 31, 39, 30, 16, 13, 6, 9, 17, 5, 
    13, 12, 16, 21, 13, 10, 5, 6, 14, 11, 0, 5, 5, 6, 3, 
    6, 6, 10, 0, 0, 0, 0, 0, 0, 0, 4, 9, 10, 3, 0, 
    6, 6, 0, 6, 20, 40, 21, 2, 8, 17, 21, 0, 0, 19, 13, 
    5, 7, 15, 0, 8, 4, 0, 6, 9, 6, 9, 24, 19, 7, 10, 
    0, 13, 2, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 6, 
    0, 0, 0, 0, 29, 16, 17, 11, 24, 40, 18, 12, 5, 5, 5, 
    14, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    16, 18, 13, 0, 0, 29, 25, 13, 14, 31, 39, 21, 19, 31, 17, 
    4, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 10, 2, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 12, 
    10, 2, 0, 9, 13, 0, 0, 0, 21, 15, 17, 29, 0, 0, 0, 
    0, 2, 25, 5, 1, 7, 3, 0, 0, 31, 52, 38, 7, 0, 5, 
    9, 5, 0, 11, 4, 6, 1, 5, 21, 0, 0, 0, 0, 1, 0, 
    2, 3, 6, 2, 0, 2, 2, 1, 0, 0, 0, 0, 4, 0, 0, 
    
    -- channel=627
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 0, 0, 0, 0, 0, 3, 5, 0, 19, 15, 0, 0, 0, 
    0, 12, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 15, 0, 0, 1, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 18, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 0, 0, 2, 14, 4, 0, 0, 0, 0, 14, 7, 0, 0, 
    0, 0, 0, 0, 0, 13, 7, 0, 0, 0, 0, 2, 7, 0, 0, 
    0, 0, 0, 0, 0, 2, 3, 0, 0, 0, 0, 0, 12, 0, 0, 
    
    -- channel=628
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 27, 0, 3, 0, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 32, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 5, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 18, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 0, 0, 0, 0, 1, 13, 10, 1, 27, 14, 1, 0, 0, 
    0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 23, 0, 3, 0, 0, 0, 4, 0, 6, 1, 0, 0, 1, 0, 
    0, 14, 0, 8, 9, 0, 0, 6, 0, 0, 0, 0, 1, 0, 0, 
    0, 26, 0, 6, 8, 5, 0, 0, 0, 0, 9, 32, 2, 0, 0, 
    0, 0, 8, 4, 0, 10, 0, 0, 0, 0, 0, 20, 0, 0, 0, 
    0, 0, 6, 0, 0, 2, 0, 0, 0, 0, 0, 13, 1, 0, 0, 
    
    -- channel=629
    17, 17, 18, 9, 5, 3, 0, 0, 13, 20, 18, 22, 5, 10, 2, 
    24, 24, 18, 0, 20, 30, 35, 40, 37, 36, 24, 27, 25, 15, 18, 
    31, 32, 20, 0, 29, 26, 20, 18, 28, 38, 35, 23, 18, 9, 28, 
    31, 29, 27, 0, 30, 19, 16, 37, 29, 23, 30, 42, 19, 0, 7, 
    32, 26, 17, 5, 35, 40, 29, 35, 35, 36, 27, 33, 23, 9, 0, 
    37, 21, 1, 0, 40, 32, 28, 31, 36, 42, 42, 48, 50, 31, 32, 
    32, 18, 20, 0, 0, 20, 14, 13, 11, 9, 9, 27, 49, 43, 37, 
    12, 8, 16, 0, 26, 33, 33, 18, 20, 24, 15, 18, 39, 42, 59, 
    1, 0, 16, 7, 15, 1, 0, 0, 0, 0, 0, 0, 0, 5, 51, 
    13, 0, 17, 0, 18, 8, 29, 28, 29, 43, 38, 39, 32, 20, 53, 
    20, 0, 0, 0, 0, 10, 6, 0, 40, 23, 26, 31, 15, 8, 36, 
    23, 0, 9, 0, 0, 0, 30, 0, 16, 1, 2, 16, 0, 30, 45, 
    30, 0, 0, 13, 0, 0, 0, 0, 1, 6, 0, 0, 0, 0, 34, 
    25, 24, 7, 7, 3, 0, 0, 0, 0, 39, 41, 3, 0, 4, 37, 
    29, 23, 8, 4, 5, 0, 0, 0, 0, 10, 24, 6, 0, 5, 40, 
    
    -- channel=630
    0, 0, 5, 20, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 11, 
    0, 0, 14, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 
    0, 0, 19, 90, 0, 0, 0, 10, 0, 0, 0, 0, 8, 22, 0, 
    0, 1, 0, 94, 0, 0, 21, 0, 0, 0, 0, 0, 3, 27, 0, 
    0, 7, 23, 49, 0, 0, 1, 0, 0, 0, 5, 0, 0, 28, 0, 
    0, 18, 15, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 28, 0, 28, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 38, 0, 41, 0, 9, 0, 8, 0, 0, 0, 0, 0, 0, 0, 
    11, 50, 0, 46, 0, 0, 0, 30, 0, 0, 46, 16, 0, 0, 0, 
    14, 76, 0, 20, 0, 4, 0, 0, 8, 0, 0, 0, 0, 15, 0, 
    0, 90, 0, 11, 0, 0, 0, 36, 0, 15, 0, 0, 26, 0, 0, 
    0, 97, 0, 0, 46, 0, 0, 30, 0, 0, 0, 0, 38, 0, 0, 
    0, 64, 0, 9, 31, 30, 0, 0, 0, 0, 8, 76, 27, 0, 0, 
    0, 11, 29, 17, 0, 43, 0, 0, 0, 0, 0, 78, 18, 0, 0, 
    0, 0, 31, 25, 0, 17, 0, 0, 0, 0, 0, 35, 24, 0, 0, 
    
    -- channel=631
    9, 3, 8, 15, 8, 0, 0, 0, 0, 10, 12, 9, 15, 8, 20, 
    3, 2, 11, 21, 0, 0, 0, 0, 0, 7, 18, 4, 10, 24, 15, 
    4, 4, 10, 29, 0, 0, 0, 0, 0, 0, 0, 1, 11, 27, 8, 
    4, 6, 7, 26, 0, 0, 0, 0, 0, 0, 0, 0, 11, 18, 8, 
    3, 9, 9, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 
    0, 11, 14, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 3, 
    0, 11, 1, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 18, 0, 2, 0, 0, 0, 2, 1, 0, 5, 1, 0, 0, 0, 
    2, 16, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 28, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    0, 30, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 33, 0, 0, 6, 0, 0, 26, 0, 5, 0, 0, 28, 0, 0, 
    0, 14, 0, 0, 8, 6, 3, 0, 0, 0, 0, 14, 9, 0, 0, 
    0, 0, 7, 0, 0, 13, 1, 0, 0, 0, 0, 22, 13, 0, 0, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 11, 6, 0, 0, 
    
    -- channel=632
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 15, 31, 39, 51, 66, 61, 40, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 0, 0, 4, 8, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 19, 0, 0, 0, 
    0, 0, 20, 20, 0, 12, 19, 0, 2, 3, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 21, 2, 0, 12, 16, 5, 20, 13, 0, 0, 0, 
    0, 15, 11, 0, 0, 0, 2, 0, 0, 9, 14, 27, 49, 51, 0, 
    0, 26, 1, 0, 12, 0, 0, 5, 34, 34, 20, 40, 43, 21, 10, 
    0, 0, 0, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 0, 26, 0, 16, 7, 19, 32, 21, 26, 34, 30, 27, 22, 10, 
    0, 0, 0, 0, 0, 11, 0, 0, 12, 0, 0, 0, 0, 0, 0, 
    0, 10, 15, 0, 0, 0, 45, 37, 19, 21, 0, 12, 30, 30, 21, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 38, 7, 2, 0, 0, 
    1, 0, 0, 4, 0, 0, 0, 0, 0, 0, 11, 12, 0, 0, 0, 
    
    -- channel=633
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=634
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 1, 2, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 13, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 5, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 9, 17, 0, 
    0, 0, 33, 0, 0, 0, 0, 0, 0, 1, 0, 2, 22, 10, 18, 
    0, 0, 2, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 
    0, 0, 1, 0, 0, 0, 0, 33, 0, 0, 0, 0, 0, 0, 54, 
    0, 0, 0, 0, 0, 12, 5, 0, 18, 0, 0, 0, 0, 0, 38, 
    0, 0, 18, 0, 0, 2, 15, 0, 31, 7, 0, 0, 0, 0, 73, 
    0, 0, 0, 0, 0, 0, 1, 5, 16, 26, 0, 0, 0, 17, 43, 
    0, 0, 0, 0, 0, 0, 0, 4, 12, 0, 11, 0, 0, 17, 39, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 37, 
    
    -- channel=635
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 9, 10, 7, 13, 14, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 
    0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 16, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    2, 15, 13, 7, 0, 0, 0, 0, 0, 0, 0, 0, 5, 3, 0, 
    9, 22, 6, 0, 4, 10, 6, 12, 14, 14, 15, 15, 12, 4, 0, 
    0, 0, 3, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 10, 15, 8, 1, 12, 8, 0, 14, 12, 16, 15, 11, 13, 0, 
    0, 6, 3, 8, 4, 2, 0, 0, 10, 5, 10, 0, 0, 2, 0, 
    0, 19, 5, 0, 0, 3, 14, 29, 0, 7, 0, 0, 21, 14, 0, 
    0, 0, 0, 7, 4, 1, 5, 3, 0, 0, 0, 0, 3, 0, 0, 
    0, 1, 6, 7, 2, 8, 0, 0, 0, 3, 15, 29, 9, 0, 0, 
    0, 0, 2, 3, 5, 5, 0, 0, 0, 2, 4, 19, 0, 0, 0, 
    
    -- channel=636
    48, 46, 50, 38, 37, 39, 42, 44, 51, 52, 47, 49, 42, 41, 31, 
    59, 58, 59, 43, 49, 53, 50, 57, 61, 51, 41, 48, 50, 41, 38, 
    60, 60, 59, 27, 40, 47, 46, 47, 49, 49, 45, 53, 49, 36, 35, 
    60, 61, 49, 45, 52, 62, 59, 61, 57, 58, 53, 50, 44, 39, 30, 
    59, 60, 56, 38, 54, 56, 54, 58, 60, 56, 62, 58, 56, 51, 38, 
    56, 60, 33, 36, 36, 44, 48, 48, 47, 47, 54, 48, 57, 60, 60, 
    50, 49, 36, 23, 41, 49, 53, 41, 46, 55, 35, 41, 56, 59, 59, 
    48, 27, 24, 41, 35, 24, 25, 26, 23, 20, 21, 23, 30, 45, 64, 
    43, 21, 33, 21, 26, 35, 30, 26, 17, 19, 29, 17, 28, 46, 58, 
    47, 23, 33, 2, 29, 20, 25, 32, 45, 44, 46, 43, 53, 28, 40, 
    50, 24, 17, 13, 6, 13, 20, 23, 21, 26, 24, 25, 28, 27, 38, 
    57, 23, 22, 23, 11, 5, 19, 8, 25, 28, 36, 48, 7, 29, 23, 
    54, 27, 28, 41, 17, 5, 0, 2, 3, 35, 46, 41, 7, 7, 32, 
    53, 54, 36, 40, 25, 9, 0, 3, 14, 40, 42, 41, 0, 11, 33, 
    54, 50, 43, 28, 22, 12, 5, 8, 11, 19, 30, 33, 2, 10, 33, 
    
    -- channel=637
    2, 0, 1, 14, 2, 2, 2, 0, 0, 0, 0, 0, 10, 2, 11, 
    0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 2, 0, 1, 11, 1, 
    0, 0, 7, 20, 0, 0, 0, 0, 0, 0, 0, 0, 3, 10, 0, 
    0, 0, 5, 25, 0, 0, 0, 0, 0, 0, 0, 0, 10, 13, 3, 
    0, 0, 5, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 8, 
    0, 0, 15, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 15, 6, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 26, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 32, 0, 34, 0, 0, 0, 15, 2, 0, 9, 5, 0, 0, 0, 
    8, 29, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    2, 42, 0, 6, 3, 2, 0, 1, 0, 3, 0, 0, 19, 0, 0, 
    0, 31, 0, 0, 14, 0, 0, 18, 0, 0, 0, 0, 19, 0, 0, 
    0, 18, 0, 0, 10, 12, 4, 1, 2, 0, 0, 4, 15, 0, 0, 
    0, 0, 3, 0, 0, 14, 7, 1, 0, 0, 0, 5, 17, 0, 0, 
    0, 0, 0, 10, 0, 10, 4, 0, 0, 0, 0, 11, 15, 0, 0, 
    
    -- channel=638
    41, 39, 48, 38, 38, 36, 31, 32, 39, 43, 41, 43, 37, 30, 25, 
    51, 51, 55, 43, 43, 46, 44, 49, 55, 44, 35, 46, 48, 38, 32, 
    53, 54, 54, 34, 17, 20, 19, 20, 23, 29, 33, 46, 51, 40, 27, 
    53, 56, 46, 41, 28, 37, 35, 31, 29, 24, 32, 48, 45, 40, 30, 
    54, 55, 52, 36, 27, 32, 35, 27, 31, 29, 38, 40, 50, 48, 35, 
    56, 61, 39, 25, 11, 23, 25, 24, 24, 24, 28, 29, 47, 53, 54, 
    55, 56, 44, 24, 18, 26, 31, 21, 24, 33, 23, 27, 46, 53, 55, 
    63, 41, 34, 46, 21, 12, 8, 13, 11, 8, 10, 13, 18, 34, 51, 
    52, 30, 38, 22, 17, 22, 19, 11, 4, 2, 14, 0, 8, 29, 36, 
    52, 31, 32, 8, 13, 15, 14, 24, 37, 33, 36, 33, 44, 22, 23, 
    53, 29, 13, 11, 1, 0, 4, 14, 9, 14, 13, 12, 12, 20, 18, 
    55, 31, 15, 16, 5, 0, 10, 11, 12, 26, 25, 40, 17, 15, 12, 
    44, 28, 14, 33, 13, 0, 0, 0, 0, 18, 32, 37, 2, 0, 12, 
    44, 43, 31, 31, 16, 6, 0, 0, 6, 23, 36, 41, 0, 0, 13, 
    39, 37, 34, 16, 12, 6, 0, 0, 2, 9, 20, 26, 0, 0, 12, 
    
    -- channel=639
    0, 4, 0, 0, 0, 3, 6, 24, 25, 0, 0, 0, 0, 8, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 4, 4, 0, 17, 0, 0, 14, 
    0, 0, 0, 0, 16, 11, 3, 0, 0, 18, 46, 12, 0, 0, 29, 
    0, 0, 0, 0, 65, 14, 0, 0, 0, 1, 18, 34, 0, 0, 2, 
    0, 0, 0, 0, 42, 13, 0, 2, 5, 2, 0, 52, 15, 0, 3, 
    13, 0, 0, 0, 26, 0, 0, 0, 0, 9, 0, 18, 49, 0, 0, 
    16, 0, 0, 0, 16, 7, 0, 0, 11, 0, 0, 33, 37, 11, 8, 
    0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 4, 23, 25, 69, 
    0, 0, 53, 0, 22, 10, 0, 0, 21, 34, 0, 13, 57, 8, 76, 
    0, 0, 18, 0, 22, 0, 15, 34, 0, 6, 0, 0, 2, 0, 92, 
    0, 0, 9, 0, 0, 11, 22, 0, 30, 0, 0, 27, 0, 14, 73, 
    0, 0, 17, 6, 0, 13, 33, 0, 80, 0, 3, 28, 0, 17, 80, 
    0, 0, 30, 0, 0, 0, 0, 8, 20, 93, 0, 0, 0, 16, 101, 
    9, 0, 0, 0, 0, 0, 3, 14, 27, 50, 4, 0, 0, 45, 75, 
    0, 0, 0, 0, 0, 0, 0, 6, 12, 16, 23, 0, 0, 33, 96, 
    
    
    others => 0);
end gold_package;
