library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 35, 0, 0, 0, 0, 6, 12, 14, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 9, 2, 0, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 5, 24, 16, 
    79, 28, 0, 0, 39, 68, 63, 60, 37, 27, 28, 34, 31, 33, 31, 
    38, 69, 16, 0, 41, 23, 26, 28, 27, 25, 27, 22, 32, 38, 22, 
    42, 40, 63, 34, 20, 26, 20, 26, 28, 28, 40, 48, 43, 30, 64, 
    36, 41, 50, 70, 41, 47, 42, 25, 16, 19, 30, 36, 14, 19, 36, 
    
    -- channel=1
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 
    9, 0, 0, 0, 16, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 23, 0, 0, 35, 0, 23, 0, 0, 0, 11, 0, 0, 0, 0, 
    0, 42, 0, 0, 0, 0, 33, 3, 7, 0, 15, 0, 0, 0, 0, 
    0, 38, 0, 0, 0, 14, 26, 3, 2, 0, 14, 0, 0, 0, 0, 
    18, 23, 0, 7, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    35, 18, 31, 0, 0, 0, 0, 20, 0, 0, 9, 0, 0, 0, 0, 
    39, 12, 31, 0, 38, 0, 10, 43, 23, 0, 0, 0, 0, 0, 0, 
    20, 35, 13, 16, 68, 26, 11, 8, 10, 5, 10, 13, 16, 13, 16, 
    19, 4, 0, 58, 35, 11, 11, 8, 8, 7, 12, 12, 21, 22, 19, 
    28, 13, 0, 103, 19, 9, 11, 6, 10, 13, 18, 24, 22, 16, 42, 
    29, 22, 11, 32, 9, 10, 19, 15, 11, 15, 15, 11, 10, 34, 30, 
    
    -- channel=2
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 4, 0, 0, 
    17, 19, 0, 0, 0, 47, 1, 6, 0, 0, 0, 0, 0, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 5, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 6, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 22, 23, 0, 0, 0, 0, 0, 6, 0, 
    0, 0, 0, 0, 0, 42, 0, 0, 0, 0, 27, 35, 11, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 29, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 
    67, 6, 0, 0, 64, 51, 34, 32, 4, 0, 0, 0, 0, 0, 0, 
    0, 49, 0, 4, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 41, 46, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 35, 
    0, 0, 0, 55, 13, 18, 17, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=3
    9, 2, 4, 6, 6, 0, 7, 8, 6, 8, 9, 5, 2, 6, 8, 
    5, 1, 2, 7, 2, 0, 10, 5, 8, 0, 0, 0, 0, 5, 9, 
    12, 6, 10, 6, 8, 0, 3, 0, 0, 0, 0, 0, 0, 7, 0, 
    0, 0, 11, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 
    0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 18, 9, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 5, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 8, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 6, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=4
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 13, 20, 14, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 16, 42, 26, 18, 8, 5, 0, 
    4, 19, 0, 0, 0, 2, 22, 13, 15, 39, 8, 17, 7, 2, 8, 
    16, 45, 0, 7, 49, 29, 19, 11, 11, 32, 28, 9, 20, 7, 6, 
    22, 42, 0, 0, 50, 19, 23, 14, 8, 72, 18, 2, 25, 15, 10, 
    20, 37, 0, 0, 34, 38, 40, 16, 11, 71, 12, 13, 20, 29, 9, 
    33, 42, 10, 3, 21, 68, 7, 16, 7, 39, 10, 9, 28, 20, 0, 
    41, 59, 11, 37, 12, 14, 8, 23, 25, 1, 28, 0, 14, 2, 0, 
    41, 48, 16, 54, 28, 14, 29, 41, 20, 14, 0, 17, 30, 5, 0, 
    74, 48, 17, 88, 35, 50, 72, 51, 24, 21, 42, 53, 53, 50, 41, 
    84, 64, 37, 88, 32, 26, 49, 48, 46, 53, 58, 61, 64, 61, 60, 
    59, 72, 60, 65, 14, 55, 55, 52, 51, 57, 63, 69, 66, 67, 75, 
    61, 64, 89, 42, 40, 58, 52, 56, 58, 63, 64, 66, 61, 83, 66, 
    59, 68, 59, 51, 44, 56, 55, 54, 61, 63, 59, 59, 78, 75, 50, 
    
    -- channel=5
    36, 37, 42, 43, 42, 34, 44, 48, 42, 22, 15, 21, 32, 36, 36, 
    44, 43, 44, 43, 44, 41, 39, 25, 3, 0, 0, 0, 0, 20, 33, 
    0, 22, 43, 45, 40, 0, 6, 0, 0, 0, 0, 0, 0, 0, 21, 
    0, 8, 36, 43, 26, 21, 1, 0, 0, 0, 0, 0, 0, 0, 3, 
    7, 0, 40, 42, 31, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 9, 31, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 29, 
    0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 19, 27, 
    0, 0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=6
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 23, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 24, 23, 0, 0, 
    51, 0, 0, 0, 0, 0, 25, 13, 11, 0, 34, 0, 15, 7, 0, 
    62, 23, 5, 0, 75, 27, 29, 25, 7, 0, 24, 32, 14, 34, 0, 
    4, 15, 17, 0, 0, 0, 56, 27, 47, 0, 24, 21, 0, 23, 29, 
    18, 31, 0, 15, 0, 0, 14, 35, 38, 0, 31, 23, 2, 8, 22, 
    20, 50, 7, 28, 0, 0, 24, 0, 23, 0, 21, 17, 0, 0, 6, 
    34, 15, 38, 10, 0, 0, 3, 14, 1, 0, 0, 6, 0, 1, 0, 
    13, 4, 63, 0, 18, 0, 0, 53, 0, 0, 13, 0, 5, 0, 0, 
    0, 7, 48, 0, 129, 46, 0, 12, 43, 28, 19, 30, 11, 0, 0, 
    0, 0, 37, 0, 5, 0, 0, 0, 8, 8, 13, 11, 20, 13, 19, 
    25, 0, 0, 5, 24, 20, 18, 15, 15, 16, 20, 21, 16, 13, 30, 
    30, 17, 0, 42, 20, 14, 28, 15, 14, 17, 12, 7, 19, 14, 7, 
    36, 21, 3, 0, 1, 0, 1, 21, 23, 29, 21, 14, 22, 39, 45, 
    
    -- channel=7
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 9, 6, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 6, 4, 0, 0, 1, 4, 6, 0, 
    13, 0, 0, 0, 0, 0, 1, 7, 10, 0, 0, 7, 4, 9, 0, 
    27, 0, 0, 0, 0, 0, 0, 5, 14, 0, 9, 8, 4, 9, 6, 
    23, 10, 0, 0, 0, 0, 0, 0, 14, 0, 7, 11, 5, 3, 7, 
    15, 11, 5, 0, 0, 0, 13, 0, 0, 0, 0, 14, 5, 1, 0, 
    20, 14, 26, 0, 0, 0, 0, 3, 0, 0, 0, 7, 0, 0, 0, 
    6, 15, 24, 1, 16, 1, 0, 3, 18, 0, 3, 6, 0, 0, 0, 
    0, 8, 22, 0, 11, 30, 13, 16, 18, 15, 29, 31, 34, 18, 17, 
    50, 9, 12, 0, 34, 38, 41, 43, 48, 52, 57, 60, 63, 66, 66, 
    79, 47, 0, 19, 54, 55, 57, 55, 58, 61, 65, 70, 69, 66, 71, 
    84, 67, 39, 32, 49, 59, 59, 59, 58, 65, 72, 74, 72, 81, 81, 
    84, 75, 58, 55, 59, 60, 59, 57, 57, 64, 72, 68, 65, 88, 81, 
    
    -- channel=8
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 7, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 4, 1, 0, 
    20, 0, 0, 0, 0, 0, 0, 4, 4, 0, 0, 3, 0, 10, 0, 
    5, 0, 0, 0, 0, 0, 9, 0, 22, 0, 3, 5, 0, 2, 3, 
    1, 28, 0, 0, 0, 0, 0, 0, 12, 0, 10, 8, 0, 0, 0, 
    6, 21, 0, 0, 0, 0, 3, 0, 0, 0, 3, 8, 0, 0, 0, 
    20, 8, 30, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    4, 3, 41, 0, 2, 0, 0, 12, 0, 0, 4, 0, 0, 0, 0, 
    0, 0, 33, 0, 56, 15, 0, 11, 28, 19, 23, 30, 32, 19, 23, 
    13, 7, 5, 0, 41, 44, 33, 33, 47, 43, 50, 51, 58, 57, 60, 
    76, 14, 0, 19, 50, 50, 49, 48, 50, 53, 58, 60, 59, 58, 65, 
    82, 64, 0, 59, 46, 47, 56, 49, 49, 55, 62, 63, 69, 68, 73, 
    81, 70, 58, 38, 47, 44, 46, 48, 50, 59, 62, 57, 53, 80, 84, 
    
    -- channel=9
    34, 40, 35, 38, 38, 34, 38, 42, 40, 34, 29, 26, 29, 36, 38, 
    33, 39, 36, 41, 31, 32, 47, 41, 35, 10, 15, 22, 18, 17, 33, 
    46, 7, 36, 41, 34, 46, 47, 30, 4, 0, 21, 15, 26, 3, 18, 
    62, 0, 34, 35, 48, 12, 27, 15, 7, 0, 42, 14, 25, 15, 0, 
    34, 0, 45, 0, 27, 17, 49, 34, 26, 0, 23, 35, 12, 25, 0, 
    19, 6, 49, 29, 3, 20, 48, 33, 47, 0, 46, 41, 3, 17, 12, 
    13, 40, 19, 67, 0, 0, 34, 29, 49, 0, 47, 30, 4, 0, 19, 
    12, 37, 10, 37, 0, 0, 61, 24, 30, 0, 33, 39, 0, 9, 24, 
    26, 8, 43, 0, 19, 12, 28, 23, 0, 39, 13, 46, 0, 6, 20, 
    18, 6, 59, 0, 32, 7, 0, 28, 15, 23, 38, 4, 0, 6, 34, 
    0, 9, 58, 0, 40, 6, 0, 22, 31, 20, 0, 0, 0, 0, 0, 
    0, 0, 10, 0, 74, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 38, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=10
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 24, 0, 0, 0, 19, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 4, 0, 0, 0, 0, 0, 0, 0, 52, 0, 0, 0, 0, 32, 
    0, 0, 0, 14, 0, 0, 0, 0, 0, 31, 0, 0, 0, 0, 1, 
    0, 9, 0, 0, 67, 0, 0, 0, 0, 68, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 46, 0, 0, 0, 0, 76, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 11, 50, 0, 0, 0, 47, 0, 0, 0, 0, 0, 
    0, 2, 0, 7, 0, 26, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 4, 0, 22, 0, 0, 1, 0, 0, 0, 0, 0, 5, 0, 0, 
    38, 0, 0, 52, 0, 0, 31, 15, 0, 0, 0, 0, 0, 1, 0, 
    90, 44, 0, 57, 0, 0, 6, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 68, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 0, 
    0, 0, 107, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 12, 
    0, 0, 3, 19, 0, 9, 10, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=11
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 15, 14, 0, 7, 0, 5, 0, 
    0, 50, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 20, 9, 
    0, 13, 0, 0, 0, 0, 0, 0, 0, 51, 0, 0, 11, 14, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 58, 0, 0, 4, 7, 36, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 15, 13, 7, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 19, 13, 0, 
    0, 0, 0, 13, 0, 8, 13, 0, 0, 0, 0, 23, 43, 0, 0, 
    0, 0, 0, 44, 0, 0, 0, 0, 0, 11, 49, 56, 38, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 22, 31, 38, 38, 44, 39, 35, 
    47, 10, 23, 0, 0, 38, 34, 39, 41, 48, 53, 50, 32, 34, 56, 
    42, 52, 23, 0, 9, 41, 40, 39, 42, 43, 40, 33, 42, 56, 6, 
    35, 51, 41, 0, 24, 34, 28, 41, 46, 45, 36, 52, 65, 24, 39, 
    
    -- channel=12
    18, 14, 21, 20, 21, 16, 19, 20, 22, 15, 10, 13, 16, 15, 17, 
    23, 16, 19, 18, 21, 32, 18, 17, 0, 16, 12, 10, 10, 15, 19, 
    10, 12, 23, 19, 23, 0, 8, 0, 18, 9, 0, 0, 0, 8, 13, 
    0, 36, 18, 22, 23, 20, 9, 9, 5, 0, 0, 0, 0, 6, 6, 
    0, 8, 14, 26, 12, 13, 0, 6, 0, 24, 0, 1, 5, 0, 13, 
    2, 0, 15, 27, 0, 0, 0, 0, 0, 39, 0, 0, 0, 0, 10, 
    12, 0, 6, 7, 0, 29, 0, 6, 0, 11, 0, 3, 6, 9, 4, 
    15, 0, 9, 7, 7, 0, 0, 0, 0, 4, 0, 0, 1, 0, 5, 
    0, 0, 8, 2, 30, 0, 0, 7, 7, 0, 0, 0, 3, 5, 18, 
    0, 0, 0, 0, 0, 19, 13, 0, 10, 0, 0, 0, 6, 18, 14, 
    0, 0, 0, 33, 9, 13, 7, 0, 0, 0, 11, 15, 6, 3, 8, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    
    -- channel=13
    40, 38, 38, 40, 41, 35, 43, 46, 40, 31, 22, 23, 27, 37, 39, 
    41, 41, 41, 42, 38, 18, 41, 29, 21, 6, 7, 15, 17, 26, 35, 
    22, 20, 42, 43, 44, 27, 21, 19, 9, 0, 1, 0, 12, 21, 24, 
    21, 14, 46, 38, 32, 12, 11, 5, 3, 0, 0, 7, 5, 17, 18, 
    0, 3, 42, 11, 0, 0, 2, 3, 6, 0, 5, 11, 2, 10, 17, 
    0, 0, 35, 23, 0, 0, 0, 9, 13, 0, 0, 3, 1, 1, 10, 
    0, 0, 25, 34, 0, 0, 0, 0, 11, 0, 0, 6, 2, 0, 12, 
    0, 0, 10, 22, 9, 0, 0, 0, 7, 0, 0, 11, 0, 3, 21, 
    0, 0, 0, 0, 8, 0, 13, 5, 0, 21, 13, 2, 5, 19, 35, 
    0, 0, 0, 0, 8, 0, 0, 0, 6, 0, 0, 3, 2, 18, 27, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=14
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 22, 19, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 12, 27, 0, 0, 0, 22, 16, 0, 
    36, 41, 0, 0, 0, 35, 15, 10, 0, 0, 0, 0, 0, 24, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 4, 0, 4, 21, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 15, 
    0, 5, 0, 0, 63, 4, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 33, 0, 9, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 22, 24, 1, 0, 0, 0, 0, 9, 0, 
    0, 0, 0, 0, 0, 31, 0, 0, 0, 0, 31, 34, 14, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 43, 31, 5, 0, 0, 1, 
    10, 0, 0, 0, 0, 0, 0, 36, 14, 0, 0, 0, 0, 22, 16, 
    67, 29, 0, 0, 46, 54, 31, 29, 13, 0, 0, 0, 0, 0, 0, 
    0, 48, 2, 11, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 46, 59, 1, 0, 0, 0, 0, 0, 0, 6, 0, 0, 28, 
    0, 0, 3, 45, 9, 17, 17, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 6, 20, 0, 0, 0, 13, 0, 0, 4, 6, 0, 
    0, 25, 0, 0, 4, 10, 0, 0, 6, 49, 0, 0, 0, 6, 16, 
    0, 68, 0, 4, 0, 16, 0, 0, 0, 58, 0, 0, 0, 0, 51, 
    0, 26, 0, 53, 0, 0, 0, 0, 0, 86, 0, 0, 1, 0, 17, 
    0, 11, 0, 0, 68, 0, 0, 0, 0, 148, 0, 0, 11, 0, 0, 
    0, 0, 0, 0, 62, 46, 0, 0, 0, 118, 0, 0, 6, 14, 0, 
    0, 0, 0, 0, 32, 48, 0, 0, 0, 79, 0, 0, 20, 0, 0, 
    0, 0, 0, 26, 0, 7, 0, 0, 22, 0, 11, 0, 25, 29, 9, 
    0, 1, 0, 56, 0, 0, 35, 0, 0, 0, 0, 0, 28, 23, 0, 
    54, 0, 0, 138, 0, 0, 21, 0, 0, 0, 1, 4, 2, 0, 0, 
    46, 27, 0, 84, 0, 0, 2, 1, 0, 0, 0, 3, 4, 1, 0, 
    0, 45, 72, 0, 0, 0, 0, 0, 0, 2, 6, 4, 0, 0, 13, 
    0, 0, 93, 0, 0, 4, 0, 0, 2, 2, 0, 0, 0, 22, 0, 
    0, 0, 2, 0, 0, 12, 1, 0, 6, 0, 0, 6, 38, 0, 0, 
    
    -- channel=16
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 6, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 5, 0, 0, 0, 0, 0, 0, 
    7, 27, 0, 0, 27, 20, 0, 0, 0, 6, 0, 0, 5, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 0, 0, 0, 6, 14, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 9, 3, 
    6, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 0, 1, 0, 14, 1, 0, 0, 0, 17, 0, 0, 
    1, 0, 0, 49, 45, 55, 48, 0, 5, 6, 34, 61, 44, 9, 4, 
    15, 2, 9, 35, 0, 0, 0, 0, 20, 41, 50, 50, 55, 52, 51, 
    63, 20, 12, 0, 0, 46, 47, 43, 45, 54, 61, 66, 57, 56, 70, 
    60, 57, 34, 0, 27, 49, 48, 47, 51, 57, 57, 51, 53, 77, 49, 
    62, 62, 45, 0, 30, 38, 40, 49, 61, 59, 55, 55, 79, 73, 54, 
    
    -- channel=17
    26, 35, 27, 33, 31, 28, 31, 35, 36, 32, 23, 15, 18, 24, 29, 
    26, 32, 28, 37, 25, 36, 37, 39, 28, 0, 5, 6, 0, 6, 26, 
    50, 0, 31, 35, 31, 49, 38, 7, 0, 0, 18, 0, 17, 0, 8, 
    57, 0, 30, 28, 50, 0, 28, 3, 0, 0, 36, 7, 13, 2, 0, 
    24, 0, 36, 0, 37, 2, 40, 21, 16, 0, 16, 25, 0, 12, 0, 
    3, 11, 37, 30, 8, 0, 50, 19, 41, 0, 45, 24, 0, 3, 0, 
    0, 57, 4, 65, 0, 0, 50, 20, 43, 0, 42, 18, 0, 0, 8, 
    0, 35, 0, 34, 0, 7, 52, 17, 20, 0, 33, 28, 0, 4, 4, 
    23, 9, 34, 0, 14, 0, 16, 25, 0, 30, 18, 27, 0, 0, 16, 
    24, 9, 60, 0, 31, 0, 0, 37, 2, 21, 24, 0, 0, 1, 28, 
    0, 10, 55, 0, 51, 8, 0, 28, 22, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 105, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 78, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 91, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=18
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 39, 8, 0, 0, 0, 13, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 0, 0, 0, 3, 0, 12, 0, 0, 0, 7, 0, 0, 0, 0, 
    41, 12, 9, 0, 74, 30, 9, 0, 0, 0, 11, 10, 0, 1, 0, 
    0, 0, 18, 0, 0, 0, 36, 5, 10, 0, 6, 0, 0, 0, 5, 
    16, 0, 0, 2, 0, 1, 0, 17, 2, 0, 10, 0, 0, 0, 0, 
    21, 17, 13, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 30, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 0, 117, 38, 0, 0, 8, 0, 0, 0, 0, 0, 0, 
    0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=19
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 9, 0, 0, 0, 13, 0, 0, 0, 0, 
    21, 16, 0, 0, 50, 35, 26, 3, 0, 0, 17, 6, 0, 0, 0, 
    25, 26, 4, 7, 16, 25, 40, 4, 0, 0, 36, 0, 0, 0, 0, 
    27, 41, 0, 0, 0, 22, 36, 19, 2, 1, 26, 1, 0, 0, 0, 
    44, 37, 4, 0, 0, 30, 30, 3, 0, 0, 21, 0, 0, 0, 0, 
    56, 42, 30, 4, 10, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 
    42, 40, 35, 5, 16, 0, 0, 31, 5, 0, 0, 0, 0, 0, 0, 
    24, 39, 30, 20, 78, 33, 30, 30, 13, 0, 0, 0, 0, 0, 0, 
    0, 21, 28, 57, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 11, 75, 13, 0, 0, 0, 0, 0, 0, 0, 1, 0, 5, 
    0, 0, 0, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 4, 23, 0, 
    
    -- channel=20
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 1, 0, 2, 25, 0, 0, 0, 5, 0, 0, 7, 2, 0, 
    0, 10, 0, 0, 1, 30, 0, 0, 0, 41, 0, 0, 0, 8, 11, 
    0, 61, 0, 6, 0, 6, 0, 0, 0, 48, 0, 0, 0, 0, 41, 
    0, 48, 0, 36, 10, 0, 0, 0, 0, 46, 0, 0, 1, 0, 18, 
    0, 14, 0, 0, 48, 0, 0, 0, 0, 118, 0, 0, 9, 0, 0, 
    0, 0, 0, 0, 64, 22, 0, 0, 0, 109, 0, 0, 0, 7, 0, 
    0, 0, 0, 0, 30, 60, 0, 0, 0, 72, 0, 0, 13, 0, 0, 
    0, 0, 0, 17, 0, 0, 0, 0, 14, 0, 14, 0, 8, 11, 8, 
    0, 0, 0, 45, 0, 0, 10, 0, 0, 0, 0, 0, 29, 31, 0, 
    48, 0, 0, 105, 0, 0, 31, 0, 0, 0, 4, 7, 13, 13, 0, 
    56, 7, 0, 90, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 45, 23, 1, 0, 0, 0, 0, 0, 0, 3, 5, 0, 0, 5, 
    0, 0, 76, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 
    0, 0, 0, 2, 0, 4, 0, 0, 0, 0, 0, 0, 23, 0, 0, 
    
    -- channel=21
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 
    0, 0, 0, 0, 0, 4, 22, 0, 0, 0, 29, 22, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 17, 13, 3, 0, 9, 7, 34, 0, 0, 
    80, 0, 5, 0, 10, 0, 21, 15, 7, 0, 28, 0, 18, 21, 0, 
    60, 0, 29, 0, 22, 16, 27, 27, 13, 0, 16, 43, 5, 37, 0, 
    20, 0, 33, 0, 0, 0, 33, 28, 58, 0, 25, 32, 0, 18, 33, 
    24, 18, 0, 34, 0, 0, 0, 25, 44, 0, 38, 34, 2, 0, 23, 
    15, 18, 27, 36, 0, 0, 19, 0, 18, 0, 12, 33, 0, 0, 2, 
    17, 0, 61, 0, 19, 0, 11, 13, 0, 30, 0, 17, 0, 0, 0, 
    0, 0, 65, 0, 22, 0, 0, 31, 7, 0, 18, 3, 0, 0, 2, 
    0, 0, 56, 0, 92, 39, 0, 0, 30, 37, 19, 12, 0, 0, 16, 
    0, 0, 9, 0, 28, 9, 0, 0, 4, 0, 0, 0, 0, 0, 3, 
    19, 0, 0, 0, 43, 1, 4, 1, 4, 1, 0, 0, 0, 0, 0, 
    17, 3, 0, 14, 12, 0, 16, 3, 0, 0, 0, 0, 3, 0, 0, 
    23, 0, 0, 0, 5, 0, 0, 0, 0, 7, 11, 0, 0, 18, 39, 
    
    -- channel=22
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 2, 23, 13, 0, 0, 0, 0, 12, 2, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 4, 13, 15, 0, 
    7, 0, 10, 0, 0, 0, 5, 3, 14, 0, 0, 8, 0, 5, 2, 
    24, 0, 16, 3, 0, 12, 0, 0, 6, 0, 17, 34, 0, 0, 0, 
    9, 0, 13, 8, 0, 0, 0, 0, 17, 0, 27, 3, 0, 0, 0, 
    0, 0, 6, 0, 0, 0, 50, 18, 7, 0, 9, 15, 0, 0, 5, 
    0, 0, 33, 0, 0, 26, 3, 0, 0, 8, 0, 55, 0, 0, 0, 
    0, 0, 26, 0, 7, 4, 0, 0, 0, 20, 52, 8, 0, 0, 0, 
    0, 0, 31, 0, 0, 0, 0, 14, 35, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 76, 57, 13, 12, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 78, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 41, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    2, 0, 0, 16, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
    
    -- channel=23
    23, 17, 21, 16, 19, 19, 20, 23, 17, 15, 22, 26, 20, 18, 17, 
    18, 19, 24, 15, 22, 0, 3, 12, 26, 10, 0, 0, 26, 27, 14, 
    4, 51, 22, 18, 24, 27, 0, 19, 15, 6, 0, 0, 0, 32, 20, 
    0, 33, 12, 22, 0, 24, 0, 0, 0, 37, 0, 0, 0, 0, 51, 
    0, 0, 0, 53, 0, 0, 0, 0, 0, 54, 0, 0, 0, 0, 45, 
    0, 0, 0, 31, 9, 0, 0, 0, 0, 50, 0, 0, 1, 0, 0, 
    0, 0, 11, 0, 35, 0, 0, 0, 0, 33, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 32, 0, 0, 0, 0, 23, 0, 0, 7, 0, 2, 
    0, 0, 0, 0, 0, 27, 0, 0, 5, 0, 0, 0, 24, 8, 6, 
    0, 0, 0, 5, 0, 22, 14, 0, 0, 0, 0, 13, 12, 14, 9, 
    0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 11, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=24
    0, 4, 2, 1, 0, 2, 3, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 4, 3, 1, 17, 1, 2, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 1, 3, 28, 0, 0, 0, 6, 14, 0, 0, 0, 0, 
    0, 0, 0, 2, 5, 0, 5, 0, 0, 16, 13, 5, 0, 0, 0, 
    0, 23, 0, 2, 33, 28, 25, 0, 0, 0, 17, 0, 0, 0, 0, 
    20, 41, 6, 21, 61, 35, 33, 2, 0, 22, 34, 0, 0, 0, 0, 
    15, 47, 0, 0, 24, 33, 50, 15, 0, 38, 21, 0, 0, 0, 0, 
    34, 38, 0, 0, 4, 61, 32, 19, 0, 37, 23, 0, 0, 9, 0, 
    47, 50, 12, 18, 7, 17, 6, 7, 0, 4, 17, 0, 0, 0, 1, 
    54, 53, 19, 21, 14, 0, 5, 25, 12, 11, 0, 0, 0, 7, 2, 
    47, 49, 21, 46, 36, 12, 42, 44, 5, 0, 0, 0, 0, 0, 0, 
    30, 39, 26, 86, 73, 5, 5, 1, 0, 0, 0, 0, 0, 4, 1, 
    0, 23, 32, 90, 5, 0, 0, 0, 0, 0, 0, 0, 6, 2, 2, 
    0, 0, 38, 51, 0, 0, 0, 0, 0, 0, 1, 3, 0, 5, 16, 
    2, 0, 2, 5, 0, 0, 0, 0, 0, 1, 0, 0, 7, 19, 0, 
    
    -- channel=25
    0, 3, 6, 7, 7, 5, 2, 2, 7, 0, 0, 0, 7, 4, 6, 
    8, 8, 7, 6, 10, 59, 8, 3, 0, 16, 29, 4, 0, 0, 10, 
    0, 0, 5, 5, 0, 0, 0, 0, 7, 31, 5, 18, 13, 0, 8, 
    26, 28, 2, 10, 13, 20, 35, 13, 9, 0, 8, 0, 0, 0, 0, 
    36, 49, 4, 27, 103, 44, 5, 6, 0, 9, 22, 13, 17, 22, 0, 
    0, 7, 0, 0, 0, 0, 30, 16, 23, 37, 0, 0, 3, 18, 22, 
    0, 2, 0, 11, 0, 21, 5, 19, 10, 22, 0, 2, 3, 17, 9, 
    0, 26, 3, 29, 13, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 7, 0, 17, 0, 0, 0, 14, 16, 0, 0, 0, 0, 5, 14, 
    0, 0, 7, 16, 0, 0, 19, 51, 0, 0, 0, 0, 24, 21, 3, 
    10, 0, 0, 50, 103, 54, 26, 0, 7, 21, 27, 46, 22, 8, 7, 
    0, 0, 20, 41, 0, 0, 0, 0, 0, 3, 7, 3, 9, 2, 2, 
    3, 0, 0, 0, 0, 6, 2, 2, 4, 9, 15, 16, 3, 3, 26, 
    1, 2, 0, 0, 0, 6, 10, 1, 5, 7, 0, 0, 1, 14, 0, 
    2, 2, 0, 0, 0, 0, 0, 7, 19, 19, 1, 3, 34, 21, 4, 
    
    -- channel=26
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 40, 0, 0, 42, 14, 0, 0, 0, 0, 10, 0, 0, 0, 0, 
    0, 13, 0, 0, 0, 0, 4, 0, 0, 17, 0, 0, 0, 0, 0, 
    0, 13, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 
    3, 30, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 18, 3, 23, 0, 0, 0, 32, 0, 0, 0, 0, 0, 0, 0, 
    17, 13, 0, 57, 70, 49, 19, 0, 0, 0, 15, 28, 23, 4, 0, 
    16, 6, 22, 57, 0, 0, 0, 0, 8, 18, 28, 32, 42, 42, 36, 
    47, 12, 10, 19, 0, 29, 28, 25, 26, 34, 45, 52, 42, 37, 64, 
    48, 42, 14, 0, 3, 35, 35, 31, 29, 38, 38, 37, 39, 60, 31, 
    48, 47, 27, 10, 8, 14, 15, 28, 41, 50, 41, 40, 69, 75, 46, 
    
    -- channel=27
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 16, 10, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 6, 7, 0, 12, 3, 10, 3, 0, 
    32, 0, 0, 0, 0, 3, 11, 8, 8, 0, 10, 11, 4, 9, 0, 
    39, 14, 0, 0, 0, 5, 6, 12, 12, 0, 21, 18, 6, 13, 7, 
    40, 21, 0, 0, 0, 0, 10, 14, 16, 0, 27, 15, 9, 7, 9, 
    31, 32, 17, 0, 0, 0, 29, 10, 9, 0, 14, 17, 6, 4, 0, 
    37, 29, 34, 1, 0, 9, 7, 2, 5, 1, 0, 14, 1, 0, 0, 
    25, 30, 36, 15, 17, 6, 7, 13, 14, 0, 13, 7, 0, 0, 0, 
    13, 26, 37, 5, 40, 24, 13, 30, 31, 23, 23, 24, 33, 25, 23, 
    44, 33, 35, 8, 50, 52, 43, 44, 45, 44, 49, 53, 56, 59, 60, 
    71, 42, 27, 26, 65, 49, 50, 49, 51, 53, 59, 60, 61, 63, 67, 
    77, 61, 32, 49, 48, 53, 55, 50, 51, 56, 63, 65, 68, 65, 71, 
    76, 66, 54, 55, 52, 49, 52, 53, 51, 58, 62, 62, 60, 76, 77, 
    
    -- channel=28
    10, 4, 9, 11, 13, 4, 8, 10, 13, 9, 6, 3, 6, 13, 16, 
    14, 3, 7, 10, 8, 5, 19, 4, 2, 6, 20, 18, 8, 4, 13, 
    8, 0, 9, 10, 10, 0, 19, 15, 16, 0, 18, 23, 31, 12, 1, 
    36, 8, 10, 7, 13, 5, 12, 27, 24, 0, 25, 13, 25, 32, 0, 
    36, 2, 26, 0, 0, 17, 14, 28, 23, 0, 12, 33, 19, 33, 19, 
    34, 0, 27, 14, 0, 1, 14, 23, 37, 0, 24, 31, 10, 26, 33, 
    38, 8, 7, 17, 0, 0, 0, 23, 26, 0, 25, 31, 21, 14, 30, 
    28, 6, 36, 12, 0, 0, 26, 9, 19, 0, 20, 29, 8, 8, 24, 
    21, 0, 48, 0, 27, 0, 15, 17, 8, 22, 0, 28, 10, 10, 14, 
    1, 2, 36, 0, 14, 25, 6, 9, 27, 4, 25, 18, 6, 6, 15, 
    0, 2, 30, 0, 46, 28, 0, 0, 27, 33, 25, 25, 22, 9, 17, 
    0, 0, 13, 0, 14, 24, 10, 12, 23, 23, 25, 23, 25, 28, 29, 
    42, 0, 0, 0, 41, 25, 25, 27, 30, 30, 28, 28, 25, 23, 26, 
    39, 28, 0, 4, 32, 25, 33, 26, 24, 25, 28, 24, 32, 24, 25, 
    41, 27, 27, 4, 31, 20, 20, 27, 25, 30, 32, 30, 21, 34, 45, 
    
    -- channel=29
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 18, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 10, 10, 7, 7, 0, 0, 0, 3, 14, 9, 1, 0, 
    6, 0, 0, 26, 0, 0, 0, 0, 0, 7, 14, 14, 17, 18, 13, 
    22, 3, 0, 6, 0, 9, 10, 10, 11, 16, 20, 22, 18, 13, 23, 
    18, 18, 0, 0, 0, 12, 12, 12, 11, 16, 18, 15, 15, 26, 20, 
    19, 20, 13, 0, 4, 6, 5, 9, 17, 21, 17, 15, 28, 34, 16, 
    
    -- channel=30
    47, 43, 48, 47, 49, 40, 49, 57, 52, 36, 30, 33, 37, 41, 45, 
    49, 46, 48, 47, 48, 15, 40, 33, 33, 12, 0, 1, 16, 31, 38, 
    17, 42, 51, 52, 52, 24, 35, 24, 8, 0, 0, 0, 0, 11, 25, 
    0, 4, 41, 50, 34, 32, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 36, 37, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 12, 
    0, 0, 35, 45, 0, 9, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 22, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 
    0, 0, 0, 0, 8, 9, 2, 0, 0, 14, 0, 11, 3, 8, 21, 
    0, 0, 0, 0, 0, 12, 3, 0, 0, 0, 4, 0, 0, 8, 32, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=31
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=32
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 76, 0, 0, 0, 13, 15, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 18, 0, 0, 0, 37, 0, 0, 0, 0, 19, 
    18, 24, 0, 0, 13, 0, 38, 0, 0, 0, 2, 0, 0, 0, 2, 
    0, 55, 0, 0, 74, 0, 0, 0, 7, 0, 10, 0, 17, 8, 0, 
    0, 36, 0, 0, 62, 0, 49, 0, 37, 39, 0, 0, 1, 0, 0, 
    0, 69, 0, 23, 43, 14, 31, 0, 11, 62, 0, 0, 0, 14, 0, 
    0, 43, 0, 27, 0, 42, 0, 0, 0, 38, 0, 0, 0, 0, 0, 
    0, 9, 0, 39, 0, 0, 0, 42, 0, 4, 20, 0, 0, 14, 0, 
    5, 0, 0, 27, 0, 0, 0, 73, 0, 0, 0, 0, 19, 20, 0, 
    82, 0, 0, 41, 30, 0, 0, 0, 0, 0, 8, 12, 0, 1, 0, 
    0, 0, 0, 71, 0, 0, 0, 0, 0, 0, 3, 2, 9, 2, 0, 
    0, 0, 0, 67, 0, 0, 0, 0, 0, 4, 6, 7, 0, 0, 8, 
    0, 0, 0, 78, 0, 0, 0, 0, 0, 1, 0, 1, 0, 14, 0, 
    0, 8, 0, 25, 0, 0, 0, 0, 6, 13, 0, 0, 16, 22, 0, 
    
    -- channel=33
    4, 8, 4, 6, 3, 2, 9, 7, 0, 0, 0, 0, 0, 0, 0, 
    1, 5, 7, 8, 4, 22, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 6, 5, 38, 0, 0, 0, 7, 20, 4, 0, 0, 2, 
    4, 0, 10, 2, 2, 0, 13, 0, 0, 11, 20, 1, 0, 0, 0, 
    13, 42, 12, 0, 53, 11, 28, 0, 0, 0, 25, 0, 0, 0, 0, 
    0, 57, 15, 0, 59, 16, 46, 12, 4, 0, 35, 0, 2, 0, 0, 
    0, 70, 6, 5, 26, 14, 72, 14, 19, 31, 29, 0, 0, 0, 1, 
    4, 61, 0, 12, 0, 68, 36, 21, 7, 34, 26, 3, 0, 13, 3, 
    33, 56, 0, 29, 0, 11, 10, 9, 2, 9, 16, 0, 0, 7, 10, 
    52, 53, 34, 17, 25, 0, 0, 48, 0, 11, 0, 0, 0, 13, 4, 
    56, 42, 37, 27, 56, 14, 32, 54, 13, 0, 0, 0, 0, 0, 0, 
    39, 40, 37, 85, 85, 0, 0, 0, 0, 0, 0, 0, 2, 7, 2, 
    4, 18, 7, 103, 5, 0, 0, 0, 0, 0, 0, 3, 12, 4, 8, 
    7, 0, 8, 95, 0, 0, 0, 0, 0, 0, 2, 10, 1, 4, 28, 
    10, 3, 0, 35, 0, 0, 4, 0, 2, 6, 6, 0, 8, 33, 8, 
    
    -- channel=34
    0, 0, 0, 1, 2, 4, 0, 0, 5, 0, 0, 0, 0, 0, 2, 
    7, 5, 0, 0, 5, 45, 0, 0, 0, 27, 28, 9, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 12, 18, 18, 0, 6, 0, 0, 0, 
    15, 32, 0, 8, 3, 27, 20, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 21, 0, 30, 44, 1, 0, 0, 0, 32, 25, 1, 9, 8, 0, 
    0, 0, 0, 0, 0, 0, 19, 14, 7, 31, 0, 0, 0, 5, 16, 
    10, 0, 0, 0, 0, 25, 0, 1, 0, 2, 0, 8, 10, 21, 0, 
    4, 16, 5, 18, 6, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 16, 0, 0, 15, 15, 17, 0, 0, 0, 0, 14, 2, 
    0, 0, 0, 27, 0, 0, 27, 30, 0, 0, 0, 4, 10, 0, 0, 
    7, 0, 0, 56, 55, 20, 0, 0, 0, 8, 34, 24, 2, 0, 4, 
    0, 0, 9, 1, 0, 0, 0, 0, 1, 0, 0, 0, 7, 2, 2, 
    0, 0, 15, 0, 0, 2, 0, 0, 3, 7, 11, 8, 0, 0, 20, 
    0, 0, 0, 0, 0, 1, 7, 0, 0, 0, 0, 0, 0, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 13, 0, 6, 31, 0, 0, 
    
    -- channel=35
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 3, 0, 0, 
    16, 3, 0, 0, 0, 18, 4, 0, 0, 0, 12, 0, 3, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 9, 21, 3, 17, 8, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 15, 0, 0, 0, 0, 0, 13, 
    23, 15, 0, 25, 36, 9, 0, 0, 0, 1, 16, 9, 8, 0, 0, 
    6, 21, 6, 0, 13, 0, 15, 0, 1, 12, 9, 4, 5, 1, 5, 
    11, 0, 1, 0, 2, 26, 24, 23, 7, 19, 13, 9, 11, 19, 0, 
    12, 11, 19, 2, 11, 22, 4, 4, 0, 0, 32, 20, 15, 0, 0, 
    21, 20, 8, 0, 13, 11, 0, 0, 20, 30, 17, 3, 0, 0, 0, 
    18, 14, 10, 0, 0, 0, 26, 29, 15, 0, 0, 0, 15, 18, 18, 
    62, 28, 0, 13, 64, 46, 37, 34, 30, 26, 28, 28, 26, 31, 31, 
    39, 56, 15, 44, 36, 23, 25, 24, 25, 26, 24, 26, 36, 34, 21, 
    38, 31, 59, 45, 31, 24, 21, 26, 26, 28, 36, 42, 33, 36, 62, 
    37, 34, 40, 39, 38, 43, 41, 26, 21, 20, 32, 29, 17, 31, 31, 
    
    -- channel=36
    28, 32, 31, 29, 29, 30, 33, 34, 29, 24, 19, 26, 26, 24, 25, 
    32, 35, 34, 30, 33, 46, 8, 25, 14, 21, 3, 6, 19, 31, 28, 
    15, 43, 33, 32, 35, 46, 0, 1, 5, 35, 0, 0, 0, 16, 40, 
    0, 54, 31, 35, 24, 22, 13, 0, 0, 36, 0, 0, 0, 0, 52, 
    0, 38, 0, 32, 21, 0, 0, 0, 0, 31, 0, 0, 8, 0, 14, 
    0, 14, 0, 3, 51, 0, 0, 0, 0, 78, 0, 0, 12, 0, 0, 
    0, 2, 3, 10, 59, 19, 5, 0, 0, 77, 0, 0, 3, 10, 0, 
    0, 0, 0, 15, 26, 46, 0, 0, 0, 54, 0, 0, 12, 7, 0, 
    0, 0, 0, 28, 0, 0, 0, 9, 13, 6, 23, 0, 14, 27, 29, 
    0, 0, 0, 29, 0, 0, 4, 9, 0, 0, 0, 2, 32, 42, 15, 
    43, 0, 0, 55, 0, 0, 9, 0, 0, 0, 0, 0, 0, 5, 0, 
    20, 0, 0, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=37
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 34, 10, 0, 0, 0, 15, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 7, 0, 9, 0, 0, 
    14, 25, 0, 0, 0, 0, 29, 14, 0, 0, 0, 0, 0, 0, 0, 
    13, 61, 3, 13, 83, 68, 0, 0, 0, 0, 16, 16, 4, 9, 0, 
    0, 0, 0, 0, 0, 0, 4, 9, 12, 45, 0, 0, 0, 3, 20, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 21, 0, 0, 0, 8, 11, 
    0, 0, 17, 1, 22, 12, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 0, 0, 4, 0, 0, 0, 0, 0, 0, 20, 
    0, 0, 0, 2, 0, 0, 0, 41, 7, 0, 0, 0, 18, 22, 0, 
    0, 0, 0, 48, 87, 89, 34, 0, 0, 0, 19, 45, 18, 0, 0, 
    0, 0, 0, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 3, 7, 14, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 14, 12, 2, 0, 30, 26, 0, 
    
    -- channel=38
    32, 30, 28, 27, 28, 27, 31, 35, 26, 22, 21, 24, 18, 23, 23, 
    27, 29, 30, 28, 27, 0, 9, 21, 18, 0, 0, 0, 23, 23, 21, 
    23, 39, 31, 30, 37, 62, 0, 9, 0, 0, 0, 0, 0, 27, 23, 
    0, 27, 27, 28, 13, 5, 0, 0, 0, 32, 0, 4, 0, 0, 41, 
    0, 0, 3, 13, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 34, 
    0, 0, 0, 45, 40, 0, 0, 0, 0, 28, 0, 0, 0, 0, 0, 
    0, 0, 10, 0, 43, 0, 0, 0, 0, 36, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 14, 11, 0, 3, 0, 44, 0, 0, 3, 10, 5, 
    0, 0, 0, 0, 0, 23, 0, 0, 0, 11, 25, 0, 21, 11, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 0, 0, 0, 18, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=39
    5, 4, 6, 0, 0, 5, 5, 4, 0, 0, 7, 15, 7, 0, 0, 
    4, 5, 7, 0, 6, 0, 0, 1, 2, 6, 0, 0, 16, 18, 0, 
    0, 43, 5, 1, 6, 22, 0, 0, 2, 25, 0, 0, 0, 17, 21, 
    0, 44, 0, 8, 0, 8, 0, 0, 0, 50, 0, 0, 0, 0, 54, 
    0, 4, 0, 36, 0, 0, 0, 0, 0, 58, 0, 0, 0, 0, 26, 
    0, 1, 0, 3, 63, 0, 0, 0, 0, 98, 0, 0, 6, 0, 0, 
    0, 0, 4, 0, 55, 20, 0, 0, 0, 82, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 22, 36, 0, 0, 0, 52, 0, 0, 13, 2, 0, 
    0, 0, 0, 17, 0, 17, 0, 0, 12, 0, 13, 0, 19, 13, 2, 
    0, 0, 0, 27, 0, 1, 17, 0, 0, 1, 0, 1, 27, 23, 0, 
    33, 0, 0, 69, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 
    48, 21, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 41, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 79, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=40
    6, 6, 0, 2, 4, 0, 5, 9, 8, 16, 21, 12, 3, 4, 8, 
    0, 0, 0, 6, 0, 0, 9, 14, 47, 0, 0, 0, 7, 5, 3, 
    32, 14, 3, 6, 3, 44, 48, 32, 0, 0, 0, 0, 6, 1, 0, 
    28, 0, 5, 0, 11, 0, 0, 0, 0, 0, 18, 6, 20, 5, 0, 
    8, 0, 16, 0, 0, 0, 14, 3, 16, 0, 0, 4, 0, 0, 0, 
    16, 0, 19, 18, 9, 12, 0, 0, 11, 0, 22, 37, 0, 0, 0, 
    0, 14, 21, 37, 0, 0, 10, 0, 25, 0, 40, 6, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 54, 27, 16, 0, 22, 25, 0, 0, 2, 
    0, 0, 27, 0, 0, 39, 21, 0, 0, 28, 11, 61, 0, 0, 0, 
    0, 0, 36, 0, 9, 0, 0, 0, 0, 27, 55, 5, 0, 0, 15, 
    0, 0, 48, 0, 0, 0, 0, 23, 28, 11, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 117, 78, 28, 27, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 99, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 88, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 43, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    
    -- channel=41
    39, 39, 41, 40, 42, 39, 42, 49, 46, 37, 31, 33, 34, 32, 34, 
    44, 43, 43, 42, 44, 28, 32, 37, 34, 20, 0, 0, 16, 35, 33, 
    19, 53, 43, 46, 44, 35, 22, 19, 0, 0, 0, 0, 0, 10, 31, 
    0, 15, 41, 48, 33, 36, 0, 0, 0, 0, 0, 0, 0, 0, 29, 
    0, 0, 23, 51, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 16, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 25, 22, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 22, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 0, 0, 0, 4, 16, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 16, 31, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=42
    4, 0, 0, 0, 0, 0, 0, 0, 0, 2, 11, 10, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 13, 13, 0, 
    0, 42, 0, 0, 2, 48, 0, 18, 3, 0, 0, 0, 0, 27, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 61, 0, 14, 0, 0, 42, 
    0, 0, 0, 41, 0, 0, 0, 0, 0, 48, 0, 0, 0, 0, 30, 
    10, 0, 0, 28, 80, 37, 0, 0, 0, 38, 0, 0, 10, 0, 0, 
    1, 0, 22, 0, 46, 0, 0, 0, 0, 35, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 30, 19, 0, 24, 0, 35, 0, 0, 20, 10, 4, 
    0, 0, 0, 0, 0, 69, 2, 0, 6, 0, 39, 15, 33, 6, 0, 
    0, 1, 0, 11, 0, 16, 12, 0, 0, 31, 5, 17, 0, 0, 0, 
    5, 0, 0, 14, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 
    81, 31, 0, 0, 0, 46, 43, 42, 13, 5, 0, 4, 0, 0, 0, 
    0, 71, 52, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 
    0, 0, 106, 0, 0, 1, 0, 0, 4, 0, 4, 13, 2, 0, 12, 
    0, 0, 11, 40, 13, 30, 25, 1, 0, 0, 0, 6, 0, 0, 0, 
    
    -- channel=43
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 41, 16, 0, 0, 0, 30, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 10, 10, 22, 0, 0, 
    52, 7, 0, 0, 12, 0, 32, 17, 6, 0, 15, 0, 0, 7, 0, 
    42, 26, 14, 0, 65, 49, 17, 23, 0, 0, 22, 34, 10, 27, 0, 
    3, 0, 13, 0, 0, 0, 36, 23, 45, 0, 11, 2, 0, 15, 32, 
    18, 7, 0, 17, 0, 0, 0, 21, 20, 0, 7, 22, 3, 7, 19, 
    20, 12, 21, 19, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 
    20, 0, 38, 0, 26, 0, 0, 20, 0, 13, 0, 0, 0, 0, 11, 
    0, 0, 36, 0, 2, 0, 0, 44, 9, 0, 0, 0, 0, 0, 0, 
    0, 0, 19, 0, 117, 66, 0, 0, 0, 22, 24, 33, 7, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 
    12, 0, 0, 0, 0, 2, 0, 0, 1, 5, 7, 11, 0, 0, 12, 
    5, 0, 0, 0, 0, 0, 14, 1, 0, 0, 0, 0, 0, 4, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 9, 18, 8, 0, 14, 28, 15, 
    
    -- channel=44
    0, 0, 4, 0, 2, 5, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    3, 6, 8, 0, 12, 35, 0, 0, 0, 14, 11, 0, 0, 0, 0, 
    0, 0, 2, 0, 6, 0, 0, 0, 15, 53, 0, 0, 0, 0, 2, 
    0, 65, 0, 11, 0, 26, 12, 0, 0, 43, 0, 0, 0, 0, 29, 
    0, 55, 0, 77, 44, 44, 0, 0, 0, 75, 7, 0, 4, 0, 15, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 136, 0, 0, 6, 0, 2, 
    0, 0, 0, 0, 43, 44, 0, 0, 0, 105, 0, 0, 8, 21, 0, 
    0, 0, 2, 0, 60, 42, 0, 0, 0, 57, 0, 0, 13, 0, 0, 
    0, 4, 0, 13, 1, 0, 0, 0, 23, 0, 0, 0, 0, 9, 19, 
    0, 0, 0, 59, 0, 2, 35, 9, 0, 0, 0, 0, 32, 30, 0, 
    27, 1, 0, 130, 0, 31, 44, 0, 0, 0, 22, 39, 26, 10, 0, 
    6, 0, 0, 101, 0, 0, 0, 0, 0, 0, 1, 5, 6, 4, 0, 
    0, 13, 47, 0, 0, 0, 0, 0, 0, 7, 14, 14, 0, 1, 20, 
    0, 2, 61, 0, 0, 7, 0, 0, 3, 5, 0, 0, 0, 23, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 16, 11, 0, 5, 48, 0, 0, 
    
    -- channel=45
    0, 2, 6, 6, 6, 2, 6, 4, 1, 0, 0, 0, 5, 7, 4, 
    7, 5, 4, 7, 3, 32, 17, 1, 0, 0, 14, 0, 0, 0, 7, 
    0, 0, 6, 4, 1, 0, 0, 0, 0, 0, 9, 10, 18, 0, 0, 
    24, 6, 5, 1, 9, 0, 20, 20, 13, 0, 20, 0, 0, 6, 0, 
    35, 24, 25, 0, 61, 59, 14, 18, 0, 0, 7, 30, 5, 22, 0, 
    14, 0, 33, 9, 0, 0, 28, 11, 28, 0, 24, 5, 0, 13, 27, 
    25, 6, 0, 15, 0, 6, 0, 31, 9, 0, 8, 12, 0, 1, 21, 
    31, 1, 21, 13, 0, 0, 16, 0, 1, 0, 5, 0, 0, 0, 6, 
    24, 0, 42, 0, 33, 0, 0, 3, 0, 3, 0, 0, 0, 0, 15, 
    0, 0, 29, 0, 0, 19, 0, 26, 12, 0, 0, 0, 4, 11, 1, 
    0, 0, 10, 0, 106, 53, 20, 0, 21, 13, 1, 26, 1, 0, 0, 
    0, 0, 13, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 6, 6, 0, 0, 2, 13, 7, 
    
    -- channel=46
    55, 58, 58, 58, 57, 52, 63, 73, 58, 32, 21, 29, 37, 48, 48, 
    57, 65, 62, 61, 57, 27, 40, 34, 19, 0, 0, 0, 0, 25, 40, 
    10, 35, 63, 66, 66, 44, 10, 0, 0, 0, 0, 0, 0, 0, 27, 
    0, 0, 52, 59, 32, 8, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 33, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 29, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 32, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 28, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=47
    0, 0, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 3, 3, 0, 6, 58, 5, 0, 0, 5, 21, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 23, 0, 9, 0, 0, 2, 
    2, 48, 3, 4, 2, 9, 26, 5, 0, 0, 0, 0, 0, 0, 0, 
    17, 58, 4, 26, 92, 42, 0, 0, 0, 20, 16, 4, 9, 10, 0, 
    0, 3, 2, 0, 0, 0, 17, 5, 7, 60, 0, 0, 0, 5, 22, 
    0, 0, 0, 0, 0, 26, 0, 6, 0, 21, 0, 0, 0, 15, 8, 
    0, 6, 10, 17, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 1, 0, 0, 4, 18, 0, 0, 0, 0, 8, 19, 
    0, 0, 0, 9, 0, 0, 15, 37, 0, 0, 0, 0, 25, 23, 0, 
    0, 0, 0, 74, 95, 60, 13, 0, 0, 0, 24, 42, 13, 0, 0, 
    0, 0, 11, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 5, 10, 0, 0, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 0, 0, 34, 7, 0, 
    
    -- channel=48
    69, 71, 71, 72, 70, 68, 76, 80, 71, 55, 44, 50, 59, 66, 65, 
    70, 80, 76, 74, 72, 71, 65, 57, 41, 29, 22, 25, 31, 50, 61, 
    36, 50, 75, 77, 75, 64, 36, 30, 23, 25, 16, 14, 17, 24, 54, 
    30, 34, 73, 74, 59, 45, 40, 14, 11, 20, 20, 19, 14, 13, 43, 
    11, 35, 58, 51, 50, 30, 28, 17, 13, 17, 32, 21, 20, 18, 18, 
    0, 15, 54, 42, 28, 20, 36, 29, 24, 21, 11, 9, 18, 14, 17, 
    0, 18, 37, 67, 41, 26, 27, 17, 24, 22, 13, 15, 14, 18, 21, 
    0, 22, 6, 49, 38, 26, 2, 13, 23, 34, 15, 17, 13, 19, 39, 
    0, 7, 0, 20, 17, 19, 28, 24, 19, 38, 27, 7, 17, 42, 60, 
    6, 5, 6, 15, 15, 2, 17, 36, 7, 11, 4, 11, 22, 53, 53, 
    10, 8, 9, 17, 14, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=49
    4, 0, 3, 0, 0, 2, 1, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 3, 6, 0, 8, 1, 0, 0, 0, 3, 0, 0, 7, 10, 0, 
    0, 33, 2, 0, 5, 19, 0, 0, 3, 46, 0, 0, 0, 17, 16, 
    0, 64, 0, 5, 0, 15, 0, 0, 0, 71, 0, 0, 0, 0, 60, 
    0, 37, 0, 66, 0, 0, 0, 0, 0, 82, 0, 0, 0, 0, 29, 
    0, 10, 0, 0, 48, 0, 0, 0, 0, 138, 0, 0, 14, 0, 0, 
    0, 0, 0, 0, 64, 29, 0, 0, 0, 118, 0, 0, 4, 9, 0, 
    0, 0, 0, 0, 48, 57, 0, 0, 0, 79, 0, 0, 20, 6, 0, 
    0, 4, 0, 20, 0, 16, 0, 0, 29, 0, 2, 0, 20, 24, 13, 
    0, 4, 0, 56, 0, 7, 35, 0, 0, 0, 0, 0, 34, 32, 0, 
    43, 0, 0, 124, 0, 0, 38, 0, 0, 0, 0, 5, 13, 9, 0, 
    66, 31, 0, 88, 0, 0, 0, 0, 0, 0, 0, 5, 1, 2, 0, 
    0, 59, 71, 0, 0, 0, 0, 0, 0, 0, 6, 5, 0, 2, 10, 
    0, 1, 111, 0, 0, 7, 0, 0, 3, 3, 0, 0, 0, 15, 0, 
    0, 0, 3, 0, 0, 10, 3, 0, 7, 0, 0, 6, 33, 0, 0, 
    
    -- channel=50
    94, 98, 98, 98, 96, 93, 102, 107, 99, 84, 75, 78, 84, 86, 86, 
    97, 103, 102, 101, 100, 86, 88, 88, 73, 47, 28, 29, 45, 76, 84, 
    65, 88, 102, 104, 102, 79, 62, 40, 34, 24, 18, 20, 18, 38, 75, 
    27, 40, 95, 101, 83, 67, 44, 25, 19, 31, 28, 25, 21, 19, 57, 
    23, 28, 81, 88, 60, 37, 31, 22, 15, 29, 31, 25, 21, 20, 25, 
    6, 23, 80, 62, 42, 46, 37, 29, 14, 29, 23, 23, 22, 20, 19, 
    12, 9, 66, 84, 42, 43, 38, 31, 23, 20, 24, 17, 15, 21, 24, 
    12, 17, 21, 61, 50, 41, 22, 25, 34, 31, 29, 17, 19, 26, 52, 
    8, 8, 4, 31, 33, 29, 34, 22, 33, 31, 36, 21, 20, 49, 74, 
    20, 10, 10, 7, 26, 21, 30, 26, 10, 39, 21, 17, 28, 66, 81, 
    14, 16, 9, 18, 18, 10, 7, 12, 11, 1, 0, 0, 0, 0, 0, 
    0, 4, 23, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=51
    63, 65, 65, 65, 64, 62, 68, 68, 65, 58, 49, 50, 52, 53, 51, 
    63, 65, 69, 67, 69, 75, 65, 60, 46, 41, 33, 28, 34, 49, 51, 
    45, 57, 65, 67, 68, 76, 47, 29, 25, 48, 43, 37, 27, 29, 50, 
    25, 41, 66, 70, 60, 52, 50, 28, 25, 56, 43, 36, 22, 12, 45, 
    46, 65, 63, 84, 87, 62, 52, 28, 18, 43, 59, 32, 29, 17, 18, 
    45, 72, 62, 46, 85, 71, 65, 44, 17, 67, 58, 30, 36, 27, 14, 
    48, 63, 59, 48, 62, 73, 85, 49, 34, 72, 54, 29, 27, 37, 29, 
    58, 69, 46, 50, 60, 95, 51, 51, 33, 67, 55, 30, 35, 37, 41, 
    68, 78, 30, 62, 38, 50, 47, 40, 49, 43, 50, 18, 18, 45, 60, 
    76, 77, 44, 57, 52, 28, 53, 62, 34, 46, 18, 11, 30, 60, 62, 
    78, 74, 45, 87, 75, 53, 65, 67, 35, 14, 12, 15, 24, 38, 32, 
    51, 68, 68, 112, 73, 22, 21, 21, 17, 14, 14, 14, 16, 20, 16, 
    10, 39, 71, 94, 25, 16, 14, 13, 11, 11, 15, 18, 20, 20, 23, 
    11, 12, 54, 63, 19, 18, 14, 13, 14, 15, 13, 17, 13, 19, 16, 
    9, 11, 14, 32, 8, 13, 18, 15, 19, 19, 14, 14, 30, 27, 7, 
    
    -- channel=52
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 
    0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 2, 5, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 7, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 6, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 13, 4, 0, 7, 0, 0, 6, 22, 2, 
    0, 0, 0, 14, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 5, 10, 0, 0, 
    
    -- channel=53
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 15, 0, 28, 0, 0, 0, 0, 0, 0, 
    21, 0, 0, 0, 0, 0, 60, 26, 0, 0, 8, 8, 29, 0, 0, 
    91, 0, 0, 0, 3, 0, 0, 7, 0, 0, 55, 0, 44, 23, 0, 
    80, 0, 39, 0, 0, 0, 43, 36, 28, 0, 0, 45, 0, 36, 0, 
    54, 0, 59, 0, 0, 12, 33, 28, 59, 0, 58, 83, 0, 16, 5, 
    43, 20, 18, 63, 0, 0, 7, 30, 75, 0, 90, 40, 0, 0, 17, 
    14, 27, 5, 24, 0, 0, 106, 22, 54, 0, 51, 60, 0, 0, 26, 
    25, 0, 95, 0, 0, 8, 34, 0, 0, 19, 0, 97, 0, 0, 0, 
    2, 0, 116, 0, 43, 0, 0, 0, 0, 25, 84, 5, 0, 0, 6, 
    0, 0, 113, 0, 50, 0, 0, 23, 80, 31, 0, 0, 0, 0, 1, 
    0, 0, 20, 0, 151, 107, 6, 11, 19, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 187, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 0, 0, 130, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 
    31, 0, 0, 35, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 
    
    -- channel=54
    78, 83, 82, 83, 84, 80, 85, 92, 89, 75, 65, 66, 69, 72, 73, 
    82, 88, 87, 86, 86, 77, 76, 79, 65, 43, 24, 26, 39, 61, 70, 
    61, 70, 86, 89, 87, 80, 54, 39, 25, 20, 9, 12, 13, 28, 60, 
    24, 33, 78, 90, 79, 62, 37, 16, 10, 22, 19, 17, 11, 9, 45, 
    11, 19, 63, 82, 51, 30, 23, 13, 9, 20, 24, 14, 14, 11, 20, 
    0, 14, 56, 56, 37, 30, 27, 21, 9, 23, 16, 13, 15, 12, 8, 
    0, 8, 44, 71, 43, 34, 32, 20, 15, 21, 14, 9, 9, 12, 10, 
    0, 12, 14, 48, 44, 34, 14, 18, 17, 29, 18, 10, 12, 13, 34, 
    1, 4, 0, 22, 22, 23, 24, 19, 22, 33, 28, 14, 10, 32, 58, 
    12, 5, 0, 8, 11, 15, 25, 20, 4, 27, 14, 10, 14, 53, 69, 
    11, 10, 1, 14, 5, 1, 4, 6, 0, 2, 0, 0, 0, 0, 3, 
    0, 0, 6, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=55
    49, 42, 45, 45, 50, 39, 50, 55, 47, 33, 25, 27, 30, 42, 42, 
    49, 45, 47, 47, 44, 9, 47, 29, 23, 3, 0, 19, 28, 28, 36, 
    21, 28, 50, 50, 55, 50, 24, 29, 4, 0, 0, 0, 6, 30, 24, 
    0, 30, 51, 46, 32, 19, 0, 0, 0, 5, 0, 9, 0, 14, 28, 
    0, 0, 47, 19, 0, 3, 0, 0, 6, 10, 0, 0, 0, 0, 40, 
    0, 0, 37, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 28, 23, 12, 0, 0, 0, 0, 0, 0, 0, 8, 0, 4, 
    0, 0, 20, 7, 17, 0, 0, 4, 0, 17, 0, 8, 0, 6, 27, 
    0, 0, 0, 0, 18, 25, 11, 0, 0, 49, 3, 7, 16, 18, 35, 
    0, 0, 0, 0, 0, 8, 0, 0, 22, 0, 0, 0, 0, 22, 30, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=56
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 3, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    6, 13, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    9, 12, 0, 20, 0, 0, 2, 0, 0, 0, 5, 5, 0, 0, 0, 
    21, 2, 0, 15, 0, 0, 27, 25, 15, 7, 11, 27, 32, 21, 13, 
    61, 44, 12, 9, 9, 39, 40, 40, 42, 48, 54, 59, 60, 59, 58, 
    68, 56, 42, 0, 29, 51, 52, 50, 50, 54, 62, 59, 64, 72, 67, 
    73, 66, 59, 26, 44, 54, 49, 48, 58, 59, 68, 70, 73, 70, 77, 
    70, 73, 65, 44, 49, 57, 62, 58, 57, 55, 57, 66, 68, 62, 68, 
    
    -- channel=57
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 19, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 
    0, 16, 0, 0, 0, 3, 2, 0, 0, 27, 0, 0, 0, 0, 0, 
    6, 4, 0, 0, 0, 20, 0, 0, 0, 9, 0, 0, 0, 0, 0, 
    11, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 15, 0, 14, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 
    21, 13, 0, 34, 16, 17, 30, 4, 0, 0, 0, 9, 12, 0, 0, 
    24, 11, 0, 51, 6, 0, 3, 0, 0, 5, 12, 15, 18, 20, 17, 
    22, 22, 10, 35, 0, 12, 13, 10, 9, 13, 18, 23, 22, 18, 26, 
    18, 21, 35, 0, 0, 14, 13, 13, 14, 18, 21, 19, 16, 32, 27, 
    21, 23, 23, 0, 3, 10, 8, 9, 19, 21, 19, 15, 30, 36, 11, 
    
    -- channel=58
    3, 4, 10, 11, 9, 7, 10, 13, 11, 0, 0, 0, 0, 4, 2, 
    13, 16, 13, 10, 13, 38, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 12, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 8, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 18, 0, 18, 33, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 
    0, 0, 0, 18, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=59
    0, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 1, 5, 
    0, 0, 0, 2, 0, 6, 2, 0, 7, 0, 7, 0, 0, 0, 4, 
    0, 0, 0, 3, 0, 0, 29, 4, 0, 0, 1, 14, 19, 0, 1, 
    57, 0, 0, 0, 5, 0, 7, 0, 1, 0, 38, 0, 26, 5, 0, 
    62, 0, 16, 0, 23, 0, 25, 18, 10, 0, 6, 22, 1, 30, 0, 
    0, 0, 30, 0, 0, 0, 46, 20, 44, 0, 19, 37, 0, 16, 11, 
    0, 21, 3, 40, 0, 0, 11, 26, 47, 0, 46, 18, 0, 0, 10, 
    0, 44, 0, 35, 0, 0, 42, 0, 34, 0, 32, 24, 0, 0, 19, 
    10, 0, 30, 0, 0, 0, 18, 1, 0, 5, 0, 38, 0, 0, 0, 
    7, 0, 70, 0, 11, 0, 0, 28, 0, 0, 41, 3, 0, 0, 3, 
    0, 0, 64, 0, 85, 0, 0, 11, 45, 24, 0, 0, 0, 0, 0, 
    0, 0, 23, 0, 41, 31, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 73, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 83, 16, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 
    
    -- channel=60
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 15, 23, 19, 0, 0, 
    0, 0, 0, 0, 0, 0, 8, 32, 8, 0, 0, 0, 0, 10, 0, 
    3, 21, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 1, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 4, 7, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 12, 0, 0, 25, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 16, 0, 0, 25, 31, 
    0, 0, 0, 0, 0, 26, 31, 27, 9, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=61
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 
    0, 0, 0, 0, 0, 0, 24, 0, 10, 0, 5, 7, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 29, 10, 0, 0, 8, 7, 28, 0, 0, 
    63, 0, 4, 0, 8, 0, 0, 11, 2, 0, 35, 0, 20, 16, 0, 
    55, 0, 39, 0, 0, 9, 33, 26, 14, 0, 2, 39, 0, 26, 0, 
    40, 0, 49, 0, 0, 3, 26, 22, 44, 0, 45, 47, 0, 13, 17, 
    37, 20, 8, 36, 0, 0, 0, 27, 44, 0, 54, 28, 0, 0, 18, 
    24, 17, 27, 22, 0, 0, 63, 4, 22, 0, 25, 34, 0, 0, 11, 
    26, 0, 71, 0, 15, 0, 12, 0, 0, 27, 0, 45, 0, 0, 0, 
    0, 0, 73, 0, 27, 2, 0, 6, 9, 0, 42, 0, 0, 0, 8, 
    0, 0, 68, 0, 67, 13, 0, 7, 50, 30, 0, 0, 0, 0, 4, 
    0, 0, 15, 0, 81, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 85, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 52, 13, 0, 4, 0, 0, 0, 0, 0, 0, 0, 8, 
    21, 0, 0, 0, 3, 0, 0, 0, 0, 0, 1, 0, 0, 3, 36, 
    
    -- channel=62
    0, 0, 2, 5, 4, 0, 2, 3, 3, 0, 0, 0, 4, 7, 8, 
    6, 3, 0, 5, 0, 41, 17, 0, 0, 0, 24, 8, 0, 0, 8, 
    0, 0, 3, 6, 0, 0, 17, 0, 0, 0, 11, 15, 26, 0, 0, 
    63, 0, 5, 0, 18, 0, 26, 14, 11, 0, 42, 0, 19, 14, 0, 
    58, 3, 28, 0, 56, 24, 30, 35, 12, 0, 16, 40, 10, 38, 0, 
    8, 0, 43, 0, 0, 0, 59, 24, 60, 0, 32, 30, 0, 20, 32, 
    21, 25, 0, 42, 0, 0, 0, 40, 38, 0, 36, 32, 0, 0, 26, 
    23, 30, 8, 36, 0, 0, 33, 0, 24, 0, 24, 26, 0, 0, 13, 
    30, 0, 63, 0, 23, 0, 4, 18, 0, 15, 0, 15, 0, 0, 3, 
    1, 0, 73, 0, 9, 0, 0, 42, 0, 0, 16, 0, 0, 0, 4, 
    0, 0, 54, 0, 133, 35, 0, 0, 36, 30, 7, 13, 0, 0, 0, 
    0, 0, 14, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    9, 0, 0, 31, 12, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 0, 0, 0, 0, 0, 0, 0, 0, 8, 2, 0, 0, 17, 28, 
    
    -- channel=63
    30, 33, 29, 30, 29, 29, 33, 38, 34, 31, 33, 31, 28, 29, 29, 
    28, 32, 30, 32, 27, 0, 31, 34, 47, 5, 0, 2, 15, 23, 24, 
    33, 29, 31, 35, 31, 37, 45, 28, 2, 0, 0, 0, 0, 9, 15, 
    9, 0, 27, 30, 27, 12, 0, 0, 0, 0, 12, 9, 13, 7, 1, 
    2, 0, 28, 4, 0, 0, 12, 8, 7, 0, 0, 6, 0, 0, 3, 
    15, 0, 35, 42, 12, 33, 0, 1, 0, 0, 12, 27, 0, 0, 0, 
    12, 0, 30, 44, 0, 0, 0, 3, 10, 0, 21, 5, 0, 0, 0, 
    3, 0, 0, 6, 0, 0, 30, 17, 13, 0, 15, 14, 0, 0, 18, 
    0, 0, 17, 0, 6, 30, 18, 0, 0, 10, 12, 41, 2, 0, 3, 
    0, 0, 11, 0, 7, 8, 0, 0, 0, 27, 31, 8, 0, 0, 28, 
    0, 0, 15, 0, 0, 0, 0, 2, 11, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 39, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end ifmap_package;
