-- https://docs.xilinx.com/r/en-US/ug953-vivado-7series-libraries/BRAM_SINGLE_MACRO

library UNISIM;
use UNISIM.vcomponents.all;
library UNIMACRO;
use unimacro.Vcomponents.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use IEEE.std_logic_arith.all;

-- BRAM_SINGLE_MACRO: Single Port RAM
--                    7 Series
-- Xilinx HDL Language Template, version 2021.2

-- Note -  This Unimacro model assumes the port directions to be "downto".
--         Simulation of this model with "to" in the port directions could lead to erroneous results.

---------------------------------------------------------------------
--  READ_WIDTH | BRAM_SIZE | READ Depth  | ADDR Width |            --
-- WRITE_WIDTH |           | WRITE Depth |            |  WE Width  --
-- ============|===========|=============|============|============--
--    37-72    |  "36Kb"   |      512    |    9-bit   |    8-bit   --
--    19-36    |  "36Kb"   |     1024    |   10-bit   |    4-bit   --
--    19-36    |  "18Kb"   |      512    |    9-bit   |    4-bit   --
--    10-18    |  "36Kb"   |     2048    |   11-bit   |    2-bit   --
--    10-18    |  "18Kb"   |     1024    |   10-bit   |    2-bit   --
--     5-9     |  "36Kb"   |     4096    |   12-bit   |    1-bit   --
--     5-9     |  "18Kb"   |     2048    |   11-bit   |    1-bit   --
--     3-4     |  "36Kb"   |     8192    |   13-bit   |    1-bit   --
--     3-4     |  "18Kb"   |     4096    |   12-bit   |    1-bit   --
--       2     |  "36Kb"   |    16384    |   14-bit   |    1-bit   --
--       2     |  "18Kb"   |     8192    |   13-bit   |    1-bit   --
--       1     |  "36Kb"   |    32768    |   15-bit   |    1-bit   --
--       1     |  "18Kb"   |    16384    |   14-bit   |    1-bit   --
---------------------------------------------------------------------

entity bram_single is
    generic (
        DEVICE     : string := "7SERIES";
        BRAM_NAME  : string := "default"
        );

    port (
        RST  : in std_logic;
        CLK  : in std_logic;
        EN   : in std_logic;
        WE   : in std_logic;
        DI   : in std_logic_vector(36-1 downto 0);
        ADDR : in std_logic_vector(9-1 downto 0);
        DO   : out std_logic_vector(36-1 downto 0)
    );
 end bram_single;

  architecture a1 of bram_single is
    signal bram_wr_en    : std_logic_vector(4-1 downto 0);
    signal bram_addr     : std_logic_vector(9-1 downto 0);

    begin
    bram_wr_en <= (others => '1') when WE = '1' else (others => '0');
    bram_addr <= ADDR(9-1 downto 0);
          

    MEM_IWGHT_LAYER0_INSTANCE0 : if BRAM_NAME = "iwght_layer0_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000018690000112a000008a40000001d00000894fffffa57000004fefffff05b",
            INIT_01 => X"00001da3ffffcfa000000a4b0000188d000013d2fffffebaffffdeecfffffcf0",
            INIT_02 => X"0000000400000000ffffffe5ffffffcafffffff70000000a000000220000001f",
            INIT_03 => X"00000018ffffffddffffffff00000038ffffffd30000002e0000002c00000003",
            INIT_04 => X"ffffffedffffffc3ffffffccffffffc900000018000000200000002100000035",
            INIT_05 => X"ffffffc0ffffffd30000001f0000001bffffffe60000000bffffffdaffffffc6",
            INIT_06 => X"0000000f000000250000001800000017fffffff500000010ffffffe2ffffffc6",
            INIT_07 => X"fffffff3000000320000000700000007ffffffd3fffffff6ffffffd8ffffffd8",
            INIT_08 => X"00000013ffffffcf0000000c00000006ffffffd8000000330000001d00000026",
            INIT_09 => X"ffffffeb0000000bfffffffbffffffff000000240000000500000020fffffff3",
            INIT_0A => X"ffffffdb0000000effffffecfffffff4ffffffdcffffffc1fffffffaffffffdf",
            INIT_0B => X"000000180000002d0000003700000006ffffffe1000000270000000900000032",
            INIT_0C => X"00000016ffffffee0000002d00000021ffffffe6000000020000001200000024",
            INIT_0D => X"ffffffd2fffffffc00000037ffffffc2fffffffbfffffff8ffffffc6ffffffe7",
            INIT_0E => X"0000001000000034000000000000001f00000040ffffffc20000001effffffe6",
            INIT_0F => X"fffffff6ffffffe6ffffffc6ffffffe5ffffffcc0000001e00000052fffffff5",
            INIT_10 => X"fffffffcffffffafffffffbefffffffa0000002b0000004dffffffeb0000002b",
            INIT_11 => X"ffffffc2ffffffe10000003900000044000000220000002bfffffffdffffffcd",
            INIT_12 => X"0000002cfffffff9fffffffa000000330000000b0000003900000001ffffffe1",
            INIT_13 => X"fffffffa0000002f000000450000003b0000002f0000001f0000002600000028",
            INIT_14 => X"fffffff800000021ffffffe400000018ffffffe6fffffff0ffffffef0000001b",
            INIT_15 => X"fffffff4ffffffc6ffffffcaffffffe500000004ffffffd2ffffffd6ffffffd5",
            INIT_16 => X"0000003300000030000000040000001c0000000000000019ffffffd6ffffffe9",
            INIT_17 => X"ffffffc1ffffffb300000005fffffffcffffffbe000000440000000dffffffd6",
            INIT_18 => X"ffffffbc0000001cffffffe400000009fffffff5ffffffd0fffffff000000022",
            INIT_19 => X"0000001100000040000000260000000e000000000000000f0000002500000010",
            INIT_1A => X"ffffffcdfffffff000000000000000340000001fffffffea0000002d00000033",
            INIT_1B => X"00000021ffffffd3ffffffbbffffffc4ffffffc900000009fffffff5fffffff6",
            INIT_1C => X"00000028ffffffc6fffffff200000000ffffffbaffffffc70000000a0000001c",
            INIT_1D => X"ffffffcbfffffff7000000330000003c00000034ffffffff0000002d00000015",
            INIT_1E => X"ffffffd100000017fffffff7fffffff8ffffffde000000030000002fffffffc7",
            INIT_1F => X"0000001c000000390000000bfffffffc0000000afffffff8ffffffc5ffffffc9",
            INIT_20 => X"fffffff8fffffffafffffffb0000000200000003fffffff9ffffffd5fffffff7",
            INIT_21 => X"0000001dffffffdf0000001e0000002bfffffff0ffffffc5ffffffc100000016",
            INIT_22 => X"000000280000003b00000020fffffff30000002d00000031000000170000001b",
            INIT_23 => X"0000003d00000014000000270000002cfffffff70000000600000029ffffffe9",
            INIT_24 => X"0000001dffffffc8ffffffd8fffffff1ffffffd2fffffff50000002500000025",
            INIT_25 => X"ffffffaeffffffbf0000002100000012ffffffe40000001e0000003100000010",
            INIT_26 => X"0000001000000035ffffffdaffffffdcfffffff3000000450000001dffffffe6",
            INIT_27 => X"ffffffd5ffffffe6fffffff7ffffffd00000001cffffffddffffffedffffffcb",
            INIT_28 => X"fffffff9ffffffe2ffffffe300000026fffffffdffffffd9ffffffe0ffffffec",
            INIT_29 => X"0000002cffffffea00000033000000160000002f0000001f0000000100000015",
            INIT_2A => X"ffffffe00000003effffffdbffffffc500000033fffffffbffffffe500000033",
            INIT_2B => X"0000002600000005ffffffd7fffffff800000028ffffffd70000001bfffffff9",
            INIT_2C => X"fffffffeffffffd8000000300000003afffffff30000004b0000000a00000003",
            INIT_2D => X"ffffffddfffffffaffffffebffffffd7ffffffff00000029ffffffc7fffffff9",
            INIT_2E => X"fffffffe0000004dfffffff900000034ffffffe4ffffffdfffffffd9ffffffc9",
            INIT_2F => X"000000030000003d0000001300000019ffffffecffffffbfffffffffffffffd6",
            INIT_30 => X"00000036ffffffff00000007ffffffe9ffffffbcfffffff2ffffffdb0000001b",
            INIT_31 => X"0000000a00000012000000240000000f00000038fffffffb0000003effffffe8",
            INIT_32 => X"0000002900000015fffffffa00000010ffffffe40000000a0000002d00000023",
            INIT_33 => X"0000001900000009ffffffe0ffffffdfffffffd1fffffffdfffffff7ffffffd1",
            INIT_34 => X"ffffffdd0000000dfffffff5ffffffeb0000001afffffff700000010ffffffda",
            INIT_35 => X"0000003100000002ffffffd2ffffffe400000013ffffffefffffffe100000018",
            INIT_36 => X"ffffffdbfffffff50000002b00000042fffffff0000000260000004600000014",
            INIT_37 => X"ffffffccfffffff200000023ffffffdaffffffe4fffffff7fffffff8ffffffcf",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER0_INSTANCE0;


    MEM_IWGHT_LAYER1_INSTANCE0 : if BRAM_NAME = "iwght_layer1_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffa160000101700004a57fffff88dfffffb98fffff23efffff546ffffd97f",
            INIT_01 => X"00001a10fffff2beffffda5300000277000041710000218500000a3200000ea5",
            INIT_02 => X"ffffed1b00000aed00002f1d0000130500000d1ffffff3ef000044f2000041b4",
            INIT_03 => X"00002a6efffff25e00001b8cfffffa92fffff844ffffd00f00002f06fffffb1b",
            INIT_04 => X"000005d9ffffd5f500001e3d000022b7000017290000265700004eda00001aee",
            INIT_05 => X"fffff0af00001eeffffff538ffffd2aa0000091dffffe84800001361ffffed40",
            INIT_06 => X"fffff967fffffec700002c6e00001756fffffaef0000227f00002c7a00000be8",
            INIT_07 => X"00002be400001e3cffffe1000000380e0000257100002da4000018cc00000ac3",
            INIT_08 => X"ffffffff0000001900000000ffffffeb00000006fffffff40000000affffffed",
            INIT_09 => X"ffffffe60000001d0000000bfffffffb0000001ffffffff0fffffff300000010",
            INIT_0A => X"000000340000008f000000280000002d0000002a00000027ffffffe0fffffffa",
            INIT_0B => X"0000000bfffffff6fffffffe0000003800000014000000230000006400000028",
            INIT_0C => X"00000054000000430000003f00000011ffffffd6ffffffd600000006fffffff9",
            INIT_0D => X"ffffffe60000001a0000000000000007000000600000003a000000450000008d",
            INIT_0E => X"00000000fffffffe000000110000001f00000024000000000000000f00000019",
            INIT_0F => X"00000000fffffffeffffffecffffffd800000021fffffffcffffffd30000001b",
            INIT_10 => X"fffffff2ffffffdffffffff7ffffffd8fffffff0ffffffddffffffecfffffffe",
            INIT_11 => X"ffffffee000000020000003b00000012fffffffd000000180000000300000020",
            INIT_12 => X"fffffff800000004fffffffefffffffc000000090000001afffffff4fffffff4",
            INIT_13 => X"fffffffc0000000dfffffffc0000001100000026ffffffe500000005fffffffa",
            INIT_14 => X"fffffffa00000007ffffffdcfffffffb00000008ffffffeaffffffd8ffffffe8",
            INIT_15 => X"0000000700000002000000110000000f0000000300000009ffffffc8ffffffdc",
            INIT_16 => X"000000250000000f00000010000000220000000e0000000bfffffffdffffffef",
            INIT_17 => X"fffffff80000000000000004fffffffa0000000000000015fffffff7ffffffe3",
            INIT_18 => X"000000100000000a0000002400000002000000100000001500000010ffffffcb",
            INIT_19 => X"fffffff1ffffffe900000001fffffff0ffffffcffffffff7ffffffd900000003",
            INIT_1A => X"fffffff0000000010000003700000011fffffff50000000e0000000900000011",
            INIT_1B => X"ffffffe50000000cfffffff3fffffffd000000130000002000000007ffffffdf",
            INIT_1C => X"ffffffd7ffffffb7ffffffffffffffc6ffffffd2ffffffbd00000000ffffffe7",
            INIT_1D => X"00000001fffffff4fffffff900000008ffffffeeffffffdfffffff91ffffffd4",
            INIT_1E => X"fffffff4ffffffd8fffffff7ffffffe5000000120000000000000022fffffffa",
            INIT_1F => X"ffffffe4fffffff600000009fffffffcfffffff000000002fffffff2ffffffde",
            INIT_20 => X"00000005fffffff8000000180000000100000010fffffff6ffffffff00000011",
            INIT_21 => X"00000001ffffffefffffffeb0000000200000002fffffff0fffffff0fffffff5",
            INIT_22 => X"0000001affffffe3fffffff80000002c000000070000000c00000002fffffff7",
            INIT_23 => X"ffffffe600000013ffffffc7000000060000000dffffffed0000001000000007",
            INIT_24 => X"fffffff60000001100000012fffffffb000000300000000e0000000dffffff98",
            INIT_25 => X"0000001afffffffe0000001d00000022ffffffee000000030000000400000008",
            INIT_26 => X"00000000ffffffe800000016fffffffc0000000affffffdcffffffe3ffffffff",
            INIT_27 => X"0000001000000002000000190000001900000021ffffffee000000080000001b",
            INIT_28 => X"00000014ffffffe00000001cffffffdbffffffedffffffd50000001200000015",
            INIT_29 => X"00000004ffffffebfffffffb0000000effffffe7fffffffafffffffcfffffff5",
            INIT_2A => X"ffffffff0000001900000014ffffffff0000001600000003ffffffe900000002",
            INIT_2B => X"ffffffe8ffffffccfffffffd000000040000001d0000000600000010ffffffeb",
            INIT_2C => X"000000000000002300000002fffffff00000001e000000120000000100000000",
            INIT_2D => X"000000250000000500000000ffffffd7ffffffdeffffffc6ffffffddfffffffd",
            INIT_2E => X"ffffffeb0000002600000024ffffffceffffffe2000000110000002c0000006e",
            INIT_2F => X"ffffff9b00000009ffffffaffffffff6fffffff6000000430000002a00000069",
            INIT_30 => X"0000001400000007fffffff1fffffff70000003b0000001cfffffff300000000",
            INIT_31 => X"ffffffe500000007fffffff100000022000000460000003f0000003e00000039",
            INIT_32 => X"0000002100000002ffffffedffffffbeffffffbbfffffffe00000051fffffff5",
            INIT_33 => X"00000010ffffffeaffffffb4ffffffb2ffffffddfffffffdffffffea00000033",
            INIT_34 => X"000000110000000c00000019ffffffbfffffffc6ffffffd00000000300000002",
            INIT_35 => X"00000020000000000000001400000012fffffff8fffffff2fffffffeffffffec",
            INIT_36 => X"0000001800000008000000220000001300000004000000220000003400000014",
            INIT_37 => X"000000200000002900000012fffffff200000009ffffffedffffffd7fffffff5",
            INIT_38 => X"0000003600000054ffffffe200000003ffffffffffffffdc000000210000001f",
            INIT_39 => X"00000006ffffffdafffffffc00000011fffffffaffffffe100000023ffffffda",
            INIT_3A => X"0000000e0000004300000039ffffffc1ffffffcfffffffbaffffffd000000003",
            INIT_3B => X"ffffffefffffffdc000000380000002500000012ffffffe4ffffffddffffffd9",
            INIT_3C => X"00000019ffffffc6ffffffcdffffffcc000000180000003e00000025ffffffd5",
            INIT_3D => X"ffffff8effffff97ffffffd9fffffffe0000000400000005000000180000001f",
            INIT_3E => X"0000002a00000005fffffff40000000cffffffef000000420000003100000034",
            INIT_3F => X"ffffffe2000000050000001e000000230000000d000000330000003000000017",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE0;


    MEM_IWGHT_LAYER1_INSTANCE1 : if BRAM_NAME = "iwght_layer1_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000100000004d00000007ffffffe7000000230000000400000005fffffffd",
            INIT_01 => X"00000022fffffff9fffffffc0000000400000005fffffff70000001dfffffffa",
            INIT_02 => X"0000001d000000030000001afffffffeffffffe5ffffffe0fffffff2fffffffd",
            INIT_03 => X"00000010000000040000001bffffffe0fffffff7000000000000000d00000008",
            INIT_04 => X"fffffffe00000007ffffffe3ffffffd2ffffffe6000000000000001f00000009",
            INIT_05 => X"ffffffdaffffffddfffffff0ffffffd4000000070000000dfffffff7fffffff0",
            INIT_06 => X"ffffffd8ffffffdcffffffe700000023000000490000003100000000fffffffe",
            INIT_07 => X"ffffffd30000004dffffffc7ffffffad00000028fffffff1ffffffb6ffffffde",
            INIT_08 => X"00000014ffffffefffffffceffffffe0fffffff6ffffffdeffffffeaffffffcc",
            INIT_09 => X"000000200000002a000000130000001600000038000000300000003100000024",
            INIT_0A => X"00000024ffffffcefffffff600000015ffffffeeffffffc3fffffff300000011",
            INIT_0B => X"fffffff1ffffffbb00000004fffffffbffffffeeffffffbb0000000000000014",
            INIT_0C => X"0000000500000000ffffffff0000003b000000260000000e00000001ffffffed",
            INIT_0D => X"fffffff300000003ffffffd9ffffffdafffffffaffffffc20000001affffffb7",
            INIT_0E => X"0000003200000018ffffffe9ffffffe1ffffffeeffffffe400000008ffffffe4",
            INIT_0F => X"ffffffddffffffe6ffffffe6fffffffb00000013ffffffeffffffff700000013",
            INIT_10 => X"00000000fffffff900000007ffffffeefffffff2000000140000002200000011",
            INIT_11 => X"0000001cffffffb3ffffffdffffffff500000008fffffff600000002fffffff8",
            INIT_12 => X"ffffffefffffffd9ffffffc7fffffffdffffffeeffffffe9ffffffe500000019",
            INIT_13 => X"0000001f000000590000001d0000001f0000000d0000000b0000000ffffffffc",
            INIT_14 => X"ffffffeeffffffd9ffffffd3ffffffc500000019000000350000000e0000003c",
            INIT_15 => X"0000000d0000000afffffffc00000025fffffff30000000600000001ffffffc4",
            INIT_16 => X"fffffffffffffffd0000001e0000000cfffffff40000000a0000002600000006",
            INIT_17 => X"00000035ffffffeaffffffdcffffffdd0000000400000006ffffffd9fffffff5",
            INIT_18 => X"ffffffeffffffff10000000fffffffcaffffffe400000000000000180000001a",
            INIT_19 => X"0000001000000037fffffffb000000000000000dffffffd200000022ffffffe7",
            INIT_1A => X"ffffffcf0000002e00000019ffffffd60000003800000031ffffffffffffffe0",
            INIT_1B => X"ffffffe30000001e0000001ffffffffbfffffffc0000001c00000028ffffffe2",
            INIT_1C => X"00000026fffffffc0000000ffffffff800000019ffffffe3fffffffcfffffffd",
            INIT_1D => X"ffffffea00000013ffffffe8fffffff30000002c00000024ffffffe900000011",
            INIT_1E => X"00000038000000070000001d000000160000000cffffffe70000000f00000002",
            INIT_1F => X"fffffffd0000000f00000002fffffffc0000001bffffffd8ffffffd8ffffffd6",
            INIT_20 => X"ffffffd200000005fffffff4ffffffceffffffeafffffffe00000008ffffffd4",
            INIT_21 => X"0000002cffffffceffffffc80000003800000004ffffffcf00000036ffffffec",
            INIT_22 => X"0000000700000031ffffffcfffffffd400000023fffffff6fffffff00000002d",
            INIT_23 => X"ffffffc60000002800000008ffffffe50000003c000000010000000afffffff0",
            INIT_24 => X"0000001f000000000000001fffffffddffffffc90000000600000024ffffffe5",
            INIT_25 => X"0000001100000018ffffffe6ffffffff00000001fffffff8ffffffe6fffffff4",
            INIT_26 => X"0000000fffffffe9ffffffe60000001f00000009fffffffbfffffff600000000",
            INIT_27 => X"ffffffe8fffffffe00000024fffffffa000000040000000b0000000d00000010",
            INIT_28 => X"0000001dfffffff30000000200000000fffffff200000007fffffff600000023",
            INIT_29 => X"000000000000001fffffffccffffffc900000022fffffffaffffffd800000031",
            INIT_2A => X"ffffffcb00000003fffffff8ffffffee0000001400000016ffffffb7fffffff3",
            INIT_2B => X"000000360000002600000022000000270000001b0000000d00000032ffffffeb",
            INIT_2C => X"00000037ffffffb7ffffffe8fffffffdffffffe0ffffffeb0000000300000030",
            INIT_2D => X"00000023ffffffd9ffffffc300000023ffffffffffffffdcffffffe30000001d",
            INIT_2E => X"fffffffcffffffe90000002d0000002effffffe400000020ffffffedffffffbe",
            INIT_2F => X"0000000f0000001f00000017000000020000002cffffffe8ffffffe500000030",
            INIT_30 => X"0000001c00000013fffffff80000002c0000004400000025000000490000003e",
            INIT_31 => X"fffffffc00000005fffffffcffffffe3ffffffd8000000350000000fffffffdc",
            INIT_32 => X"ffffffeb000000060000001b000000120000001a0000001300000030ffffffca",
            INIT_33 => X"0000003e00000003ffffffc00000000effffffffffffffbf00000029fffffff4",
            INIT_34 => X"ffffffee0000000cfffffffbfffffffd000000030000000000000000fffffffd",
            INIT_35 => X"fffffff6fffffff3fffffff8ffffffea0000000affffffe4fffffff000000008",
            INIT_36 => X"fffffff6fffffff4ffffffe70000000bffffffed00000006fffffff3ffffffea",
            INIT_37 => X"ffffffe8fffffff0fffffff500000008fffffff0000000000000000efffffff6",
            INIT_38 => X"000000000000000500000000ffffffecfffffffd00000005ffffffeb0000000d",
            INIT_39 => X"fffffff400000007fffffff1ffffffedffffffee00000003fffffff6fffffffa",
            INIT_3A => X"fffffff4fffffffbfffffff6000000060000001100000002fffffffb00000000",
            INIT_3B => X"0000000dfffffffdfffffffd00000006fffffff3fffffff7fffffff0fffffff3",
            INIT_3C => X"00000000ffffffddffffffeb00000000ffffffee00000007000000050000000a",
            INIT_3D => X"ffffffecfffffff900000007000000040000000900000002ffffffe70000000c",
            INIT_3E => X"fffffff9fffffff70000000200000002ffffffff00000008ffffffedfffffffc",
            INIT_3F => X"000000100000000000000003fffffff20000000fffffffebfffffffffffffffc",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE1;


    MEM_IWGHT_LAYER1_INSTANCE2 : if BRAM_NAME = "iwght_layer1_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000007fffffff800000011fffffff8ffffffebffffffdffffffffaffffffea",
            INIT_01 => X"fffffff400000005fffffff80000000500000008fffffffcfffffff200000004",
            INIT_02 => X"ffffffe2fffffffdffffffe1fffffffcfffffff400000002ffffffeb00000000",
            INIT_03 => X"ffffffee0000000100000000fffffffd00000000fffffff20000000b0000000a",
            INIT_04 => X"fffffff8fffffff50000000b000000070000001200000008ffffffeefffffff9",
            INIT_05 => X"fffffff5fffffffbfffffffbfffffff20000000500000003fffffff1ffffffec",
            INIT_06 => X"00000000fffffffbffffffffffffffe8fffffff700000000fffffff00000000b",
            INIT_07 => X"ffffffe7ffffffe9ffffffefffffffebffffffec00000006ffffffffffffffed",
            INIT_08 => X"fffffff20000000afffffff6fffffffe00000000fffffff4fffffffafffffffd",
            INIT_09 => X"00000000fffffff1fffffffe0000000cffffffeafffffff8fffffff4fffffff5",
            INIT_0A => X"fffffff9ffffffed0000000fffffffecffffffebfffffff4ffffffe7fffffff0",
            INIT_0B => X"0000000400000003fffffff4ffffffedfffffff3fffffffbffffffebfffffffb",
            INIT_0C => X"0000000cfffffffefffffff20000000bffffffee00000007fffffffa00000001",
            INIT_0D => X"00000004fffffffcffffffe7fffffff8ffffffeb00000000ffffffe900000005",
            INIT_0E => X"ffffffedfffffff200000003fffffff800000000ffffffeafffffffc00000003",
            INIT_0F => X"00000000fffffffc00000005ffffffe8ffffffeaffffffff00000005ffffffea",
            INIT_10 => X"fffffff0fffffff600000009fffffff300000001fffffff0ffffffeeffffffe0",
            INIT_11 => X"0000000100000000000000110000000400000002fffffffbffffffed00000009",
            INIT_12 => X"0000000800000010ffffffea0000000b0000000bffffffec0000000500000000",
            INIT_13 => X"fffffff0fffffffefffffff2ffffffeaffffffe8fffffff600000002ffffffec",
            INIT_14 => X"0000000700000007fffffff600000009fffffff5fffffff1fffffff1fffffff9",
            INIT_15 => X"fffffff600000009fffffff1fffffffa000000010000000b0000000bffffffed",
            INIT_16 => X"fffffff3fffffff4fffffffb000000090000000d00000008fffffffa00000006",
            INIT_17 => X"fffffff000000008fffffff7fffffff30000001200000004ffffffe3ffffffef",
            INIT_18 => X"000000010000000c00000001fffffff6fffffffb000000170000001b00000009",
            INIT_19 => X"ffffffe6fffffffa0000003e00000012ffffffe3ffffffd5ffffffe3fffffffc",
            INIT_1A => X"ffffffd9fffffff70000000cffffffeaffffffd6ffffffb6fffffff3ffffffee",
            INIT_1B => X"ffffffbeffffffe400000032ffffffceffffffe6000000070000001e00000011",
            INIT_1C => X"0000000affffffcdffffffceffffffd0ffffffc2ffffffe4ffffffdfffffffd5",
            INIT_1D => X"ffffffd3ffffffc3ffffffc3ffffffe5ffffffd6fffffff8ffffffd0ffffffd1",
            INIT_1E => X"00000025000000230000001600000016fffffffeffffffe9ffffffeaffffffbf",
            INIT_1F => X"ffffffff000000360000001c00000008fffffffb0000000f0000001b00000031",
            INIT_20 => X"fffffff20000001f0000000effffffedfffffff7ffffffe10000001800000016",
            INIT_21 => X"0000000e00000003fffffff1000000110000002bfffffff60000000800000007",
            INIT_22 => X"ffffffd7ffffffabffffffcfffffffb6fffffff0ffffffc3fffffff900000024",
            INIT_23 => X"0000000e0000003a000000280000000000000003000000090000000fffffffde",
            INIT_24 => X"00000024fffffff40000000100000014ffffffe90000001d0000000ffffffffa",
            INIT_25 => X"fffffff4fffffff70000001a00000016ffffffdcffffffeefffffffdfffffff0",
            INIT_26 => X"0000001c00000038fffffff3ffffffdfffffffe0fffffff500000000ffffffde",
            INIT_27 => X"00000000ffffffeaffffffe2ffffffebffffffb2ffffffaaffffffcfffffffb5",
            INIT_28 => X"0000000f0000000c0000000300000016fffffff2fffffffaffffffff00000000",
            INIT_29 => X"ffffffc8ffffffe5fffffffc00000000ffffffe0ffffffef00000000fffffffa",
            INIT_2A => X"000000350000001200000060000000410000002affffffe80000000d00000027",
            INIT_2B => X"fffffff9000000220000003fffffffed000000170000001a0000000f0000001d",
            INIT_2C => X"0000000c0000002c00000006fffffff800000000000000060000003700000046",
            INIT_2D => X"000000010000000d0000000afffffffd00000016ffffffd400000000ffffffe4",
            INIT_2E => X"0000000d0000001f000000180000002b00000002fffffffe0000000400000002",
            INIT_2F => X"0000000effffffe60000000200000004fffffffb000000130000001600000013",
            INIT_30 => X"0000001bffffffda0000000dfffffffa0000001400000015ffffffdf00000010",
            INIT_31 => X"fffffff500000002ffffffecfffffff7ffffffe3ffffffeeffffffcefffffff0",
            INIT_32 => X"00000011000000120000001a000000320000003f00000022fffffffffffffff2",
            INIT_33 => X"ffffffec00000023ffffffd6fffffff50000002effffffe7ffffffce00000017",
            INIT_34 => X"fffffff1ffffffd60000002effffffe7ffffffdaffffffdaffffffedffffffbe",
            INIT_35 => X"ffffffeeffffffe9ffffffd4ffffffe5ffffffe0ffffffcc0000000800000005",
            INIT_36 => X"ffffffe900000006ffffffd5fffffff80000000b000000280000000600000008",
            INIT_37 => X"ffffffd900000015ffffffb6ffffffa7fffffffdfffffff70000001cffffffe9",
            INIT_38 => X"ffffffd9fffffffc0000000dfffffff3ffffffd7ffffffbcffffffd1ffffffc7",
            INIT_39 => X"0000000500000029000000110000000600000014fffffff10000000300000024",
            INIT_3A => X"fffffff6fffffff00000000f00000011ffffffe9fffffff70000000c00000014",
            INIT_3B => X"fffffff6ffffffecffffffdbffffffe90000000affffffe5ffffffecffffffeb",
            INIT_3C => X"fffffff5fffffff80000001cfffffff0fffffffffffffffdffffffec0000000f",
            INIT_3D => X"fffffff3ffffffe9fffffff10000000c000000050000002600000038fffffff9",
            INIT_3E => X"ffffffadffffff9fffffffcbffffff92ffffffadfffffffa0000002c0000000e",
            INIT_3F => X"ffffffe5ffffffd0ffffffc4ffffff8dfffffffbffffffd5ffffffe700000036",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE2;


    MEM_IWGHT_LAYER1_INSTANCE3 : if BRAM_NAME = "iwght_layer1_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff0ffffffecffffffb7fffffff2fffffffeffffffdb00000004ffffffcb",
            INIT_01 => X"000000220000003500000023ffffffebfffffff7ffffffd1ffffffc6ffffff9e",
            INIT_02 => X"ffffffd8ffffffe0ffffffedfffffffd00000000000000310000001a00000012",
            INIT_03 => X"0000001bfffffffcfffffff200000008ffffffd8fffffffdfffffff3ffffffde",
            INIT_04 => X"00000019ffffffeeffffffe30000001cffffffef00000007000000120000000a",
            INIT_05 => X"fffffff1ffffffd3ffffffe0ffffffb7ffffffbafffffff4ffffffd4fffffffe",
            INIT_06 => X"00000015fffffff1000000180000002d0000000d00000024fffffffa0000000c",
            INIT_07 => X"ffffffe0ffffffe4ffffffefffffffdfffffffd7fffffffa0000000000000018",
            INIT_08 => X"0000000000000007ffffffe0ffffffdcffffffe800000058000000160000000e",
            INIT_09 => X"00000000000000100000000dfffffffcffffffbeffffffe200000010ffffffbd",
            INIT_0A => X"00000000000000140000001000000006ffffffee0000000100000007fffffffd",
            INIT_0B => X"0000000800000019000000100000000b0000001a000000160000001200000019",
            INIT_0C => X"00000004fffffff9ffffffeeffffffe3ffffffeffffffffeffffffe40000001a",
            INIT_0D => X"ffffffd5000000000000000efffffff8000000110000000f0000001200000020",
            INIT_0E => X"ffffffedffffffd700000001ffffffbcffffffe9ffffffddffffffd1ffffffe5",
            INIT_0F => X"00000014fffffff80000000f0000003e0000001600000003fffffffd00000002",
            INIT_10 => X"fffffffa0000000afffffffeffffffc400000007fffffff9ffffffd3fffffffd",
            INIT_11 => X"0000000d00000002000000110000001200000000ffffffe20000002200000015",
            INIT_12 => X"000000230000002100000025000000140000000a00000007ffffffdb00000023",
            INIT_13 => X"0000002f000000050000000c0000000d00000005ffffffe7000000340000001c",
            INIT_14 => X"0000000bfffffff4ffffffff00000005fffffffd0000003c0000002700000009",
            INIT_15 => X"ffffffedffffffc800000006ffffffedffffffe90000001600000005ffffffe5",
            INIT_16 => X"0000002b000000130000000f0000000afffffffaffffffd2fffffff8ffffffe5",
            INIT_17 => X"fffffff900000033fffffff1fffffff8fffffffbffffffdeffffffb30000001c",
            INIT_18 => X"00000015000000050000000e00000007ffffffeefffffff20000001bffffffe2",
            INIT_19 => X"ffffffd20000000a0000002efffffff70000002100000022000000310000001a",
            INIT_1A => X"00000007ffffffc3fffffff9fffffff1fffffff7ffffffec0000000400000044",
            INIT_1B => X"ffffffd4ffffffbdffffff78ffffffbe0000000200000000ffffffff00000005",
            INIT_1C => X"000000150000000b0000000fffffffd3ffffffd5fffffff0ffffffcdffffffb8",
            INIT_1D => X"0000001d0000000bfffffff8ffffffea0000001e0000003000000021fffffffc",
            INIT_1E => X"000000170000002ffffffffbfffffffc0000001a000000190000000400000010",
            INIT_1F => X"ffffffc60000000c00000025fffffff800000017000000370000001e00000019",
            INIT_20 => X"fffffff2fffffff9fffffffbffffffeafffffff1fffffff1ffffffe5ffffffd8",
            INIT_21 => X"fffffff7000000150000002500000032000000290000002a00000026ffffffeb",
            INIT_22 => X"00000026ffffffeaffffffe2fffffffd0000000e00000000ffffffb8ffffffbb",
            INIT_23 => X"ffffffdaffffffd60000003100000012fffffff60000001afffffff5ffffffe5",
            INIT_24 => X"0000002effffffea0000001cffffffda00000023ffffffedffffffe80000000d",
            INIT_25 => X"000000050000000800000004000000070000001afffffff00000001600000035",
            INIT_26 => X"00000002000000380000003300000031000000270000001c0000003600000015",
            INIT_27 => X"fffffff2ffffffd3ffffffcdfffffff2ffffffedfffffff90000001900000024",
            INIT_28 => X"ffffffcbffffffceffffffdfffffffabffffffa1ffffffb5fffffff1fffffff1",
            INIT_29 => X"000000030000000e000000370000003f00000053000000220000002600000028",
            INIT_2A => X"000000140000000b000000010000000afffffff6fffffff2fffffffbfffffff0",
            INIT_2B => X"0000000b0000000a0000001b00000017fffffffe000000050000000cfffffff0",
            INIT_2C => X"000000000000000200000021ffffffef0000000bffffffddfffffff1ffffffde",
            INIT_2D => X"ffffffe500000020000000210000002100000030fffffffdfffffffc00000040",
            INIT_2E => X"ffffffe7ffffffc4ffffffdefffffff2fffffff5ffffffe80000001300000019",
            INIT_2F => X"000000250000000affffffd2ffffffddffffffeeffffffcaffffffc1ffffffcc",
            INIT_30 => X"0000001800000013fffffff300000006000000230000003a000000220000002c",
            INIT_31 => X"0000002c0000001affffffe40000000efffffffefffffffffffffff7fffffff0",
            INIT_32 => X"ffffff95ffffffaeffffffedffffffb3ffffffabfffffff50000000200000011",
            INIT_33 => X"fffffff50000002f000000160000002200000013000000050000001affffffa3",
            INIT_34 => X"00000031fffffffaffffffd5000000160000000cffffffd30000000600000008",
            INIT_35 => X"00000016fffffff60000001d00000032000000340000001100000034ffffffec",
            INIT_36 => X"ffffffce00000004ffffffee00000004fffffff1fffffff5fffffff0ffffffef",
            INIT_37 => X"0000001a00000027000000250000001500000004fffffffcffffffe9fffffffd",
            INIT_38 => X"0000002d0000002900000011000000150000001ffffffffb000000160000000e",
            INIT_39 => X"0000000bffffffe3ffffffd0ffffffe50000000f00000002000000170000001f",
            INIT_3A => X"fffffffbffffffebffffffe5fffffffe0000000affffffe9ffffffff00000012",
            INIT_3B => X"ffffffefffffffbbffffffacffffffdcffffffe8ffffffcefffffffa0000002b",
            INIT_3C => X"ffffffc6ffffffb6ffffffacffffffb0000000130000000200000007ffffffcd",
            INIT_3D => X"00000024fffffffeffffffec000000030000001100000019ffffffabffffffb6",
            INIT_3E => X"fffffff80000000bffffffec0000000a0000001a00000003ffffffffffffffe0",
            INIT_3F => X"ffffffcdfffffffefffffff8fffffffcffffffb7ffffffbaffffffb6ffffffba",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE3;


    MEM_IWGHT_LAYER1_INSTANCE4 : if BRAM_NAME = "iwght_layer1_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffdeffffffe2000000090000002e0000004efffffff40000002f00000010",
            INIT_01 => X"00000005fffffff6ffffffc3ffffffc3ffffffe4ffffffb3ffffffd3fffffff0",
            INIT_02 => X"fffffff9fffffffefffffff80000001000000000ffffffefffffffd300000006",
            INIT_03 => X"0000001e00000010fffffffe00000016ffffffef000000130000001ffffffff5",
            INIT_04 => X"000000120000000c0000000e0000000bfffffff50000000c0000000ffffffffd",
            INIT_05 => X"ffffffe5fffffff4fffffffb0000000cffffffecfffffffefffffff2fffffffb",
            INIT_06 => X"00000000fffffff300000001fffffffc0000000100000009ffffffe7fffffffa",
            INIT_07 => X"00000000fffffff5ffffffea00000001ffffffe6fffffffa00000002fffffff8",
            INIT_08 => X"ffffffe500000003ffffffeefffffff400000000fffffff6ffffffff00000005",
            INIT_09 => X"ffffffe9ffffffec0000000100000006ffffffebffffffeefffffffafffffff6",
            INIT_0A => X"fffffffe0000000500000001fffffff4fffffff400000000000000090000000a",
            INIT_0B => X"ffffffeffffffff9ffffffedfffffff5ffffffeb00000011fffffffffffffffb",
            INIT_0C => X"00000004fffffff50000000700000005ffffffe80000000400000006fffffff6",
            INIT_0D => X"ffffffe3ffffffff0000000500000005fffffffbfffffff6fffffff1ffffffe0",
            INIT_0E => X"00000014ffffffef0000000bfffffffc00000006fffffff00000000000000005",
            INIT_0F => X"00000000ffffffe3ffffffe5fffffffcfffffff1ffffffe300000006ffffffed",
            INIT_10 => X"fffffffd0000000dfffffff4fffffffc00000003ffffffe700000000ffffffe5",
            INIT_11 => X"000000070000001300000013000000060000000cfffffffafffffff200000008",
            INIT_12 => X"fffffff9fffffff3fffffffa00000013fffffff80000000dffffffebffffffee",
            INIT_13 => X"00000000000000030000000000000007fffffff20000000000000004fffffff8",
            INIT_14 => X"ffffffe4ffffffff0000000dfffffff80000000efffffff7ffffffeafffffffd",
            INIT_15 => X"fffffffdfffffff0fffffff20000000bffffffed0000000800000004fffffff8",
            INIT_16 => X"fffffffd0000000cfffffffefffffff70000000000000001ffffffeafffffff0",
            INIT_17 => X"00000005fffffff2ffffffecfffffffdfffffff7fffffffbfffffff8fffffff0",
            INIT_18 => X"ffffffedffffffeefffffffefffffffb00000003ffffffe700000004fffffff0",
            INIT_19 => X"00000009ffffffe7ffffffe900000000fffffff8fffffff40000000900000007",
            INIT_1A => X"ffffffeafffffffffffffff2fffffff5ffffffe9fffffff30000000100000006",
            INIT_1B => X"fffffff8ffffffeffffffffc00000008ffffffeffffffff9fffffff1ffffffe3",
            INIT_1C => X"00000009fffffff900000005fffffff1fffffffc00000002ffffffe70000000a",
            INIT_1D => X"fffffff8fffffff50000000effffffeefffffff1000000110000000efffffffc",
            INIT_1E => X"ffffffeafffffffafffffff0fffffff9ffffffe6fffffff6fffffff9fffffffb",
            INIT_1F => X"ffffffec00000004ffffffe1fffffffdfffffff70000000b00000001fffffff5",
            INIT_20 => X"ffffffdafffffff1fffffff1fffffff100000003ffffffe6fffffffcffffffea",
            INIT_21 => X"000000070000000200000011fffffff3fffffff500000010ffffffec00000000",
            INIT_22 => X"ffffffed000000030000000afffffffa0000000fffffffef0000000700000014",
            INIT_23 => X"fffffff70000000dffffffffffffffe8ffffffedfffffffe0000000100000004",
            INIT_24 => X"0000000200000001fffffffc000000000000000a00000000fffffff2fffffff1",
            INIT_25 => X"000000060000000400000005fffffff500000001fffffff8fffffffffffffffd",
            INIT_26 => X"fffffffcfffffffc00000008fffffff60000000600000005fffffffe00000001",
            INIT_27 => X"000000000000000bffffffebffffffec00000000fffffff000000003ffffffe9",
            INIT_28 => X"fffffffdfffffff7fffffffd00000003ffffffeb0000000ffffffff900000000",
            INIT_29 => X"ffffffdcffffffdb0000001500000002fffffffc00000004fffffff10000000a",
            INIT_2A => X"000000210000001000000019fffffff7ffffffee00000022ffffffd9ffffffb8",
            INIT_2B => X"00000030fffffff40000000a0000002f0000001c00000005000000050000002e",
            INIT_2C => X"fffffff600000028ffffffedffffffe60000002200000048000000020000002e",
            INIT_2D => X"000000110000001dfffffff70000001900000042000000360000001e00000014",
            INIT_2E => X"0000000fffffffdd000000340000003b00000027ffffffed000000480000002b",
            INIT_2F => X"0000002400000029fffffff4ffffffd5fffffffeffffffc9ffffffdc0000000a",
            INIT_30 => X"000000160000000cffffffe6fffffffdffffffdafffffffffffffff10000000d",
            INIT_31 => X"ffffffea0000001c0000001affffffeeffffffe300000003fffffffeffffffe8",
            INIT_32 => X"0000000600000000ffffffd1ffffffed0000002f00000010ffffffdc00000010",
            INIT_33 => X"ffffffffffffffdfffffffbe00000002ffffffebffffffec00000001fffffff0",
            INIT_34 => X"fffffffaffffffef00000006fffffffcfffffffaffffffe2ffffffc7ffffffb9",
            INIT_35 => X"fffffffbffffffdeffffffebfffffff500000015fffffff4ffffffe80000000f",
            INIT_36 => X"ffffffce0000000afffffff0fffffff3ffffffefffffffd900000017fffffffc",
            INIT_37 => X"fffffff7ffffffebfffffff8ffffffd9ffffffbf00000003ffffffee00000000",
            INIT_38 => X"fffffffd0000000000000002fffffff90000000f0000000dfffffff000000013",
            INIT_39 => X"ffffffdeffffffc9ffffffdfffffffe0ffffffea00000006ffffffe7ffffffd1",
            INIT_3A => X"ffffffdeffffffaaffffffd600000024ffffffbd00000015fffffff900000018",
            INIT_3B => X"ffffffc000000000ffffffd9ffffffc10000002e00000013ffffffef0000000a",
            INIT_3C => X"0000002e000000310000001100000007fffffff400000012fffffff0ffffffef",
            INIT_3D => X"00000004fffffffc00000000ffffffe7ffffffeafffffffb0000002e0000000e",
            INIT_3E => X"fffffff0000000220000000400000001ffffffef0000000500000002fffffffa",
            INIT_3F => X"fffffffa00000009ffffffdffffffff1fffffffafffffffe00000002fffffff5",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE4;


    MEM_IWGHT_LAYER1_INSTANCE5 : if BRAM_NAME = "iwght_layer1_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff2ffffffb3fffffff0ffffffeafffffffc00000004fffffffb0000000f",
            INIT_01 => X"ffffffcbfffffffbffffffdcfffffff400000005fffffff7ffffffda00000023",
            INIT_02 => X"00000016ffffffe0ffffffa20000000fffffffe6ffffffb100000018fffffffa",
            INIT_03 => X"ffffffe50000000800000024000000020000001e0000004dffffffd5ffffffc4",
            INIT_04 => X"ffffffbcffffffe3ffffffeeffffffd1ffffffd9ffffffecfffffffffffffff0",
            INIT_05 => X"00000024ffffffe20000000c0000000c00000009ffffffe800000012fffffffc",
            INIT_06 => X"00000008ffffffde0000001afffffff8ffffffeb0000000affffffcffffffff8",
            INIT_07 => X"0000002a0000001d0000002a00000014ffffffe4ffffffcdffffffdf00000005",
            INIT_08 => X"0000000400000025ffffffe90000003800000069000000560000002a00000016",
            INIT_09 => X"000000030000001afffffff6ffffff9bffffffd6fffffff5fffffffbffffffcb",
            INIT_0A => X"0000000a0000002800000005ffffffd6fffffffefffffff6ffffffe900000015",
            INIT_0B => X"0000000e000000180000001f0000001700000006fffffffc00000007fffffffd",
            INIT_0C => X"0000000f00000001000000020000001efffffff7ffffffe9ffffffeb00000005",
            INIT_0D => X"00000019000000220000002f0000002cfffffff0fffffffe0000001efffffff0",
            INIT_0E => X"0000001200000011fffffff9ffffffe5ffffffd4ffffffe40000000000000016",
            INIT_0F => X"0000003700000005ffffffe5fffffff300000027000000100000001afffffff8",
            INIT_10 => X"00000010ffffffecffffffd0ffffffef00000006000000350000002500000006",
            INIT_11 => X"00000022fffffffdfffffff4ffffffea0000004600000000ffffffda00000000",
            INIT_12 => X"fffffff5fffffffc0000001a000000000000000600000008fffffff900000026",
            INIT_13 => X"00000020000000180000000800000026000000050000000d0000001dffffffdf",
            INIT_14 => X"fffffff300000009fffffffbffffffeb0000001300000028fffffff300000000",
            INIT_15 => X"fffffff1ffffffecfffffff20000001100000011ffffffd0ffffffe7ffffffef",
            INIT_16 => X"ffffffe800000018ffffffebffffffc10000002200000008ffffffd9ffffffd0",
            INIT_17 => X"000000140000000d00000031fffffff7000000140000002d00000020ffffffd1",
            INIT_18 => X"ffffffe4ffffffc800000008ffffffe1ffffffd7ffffffeafffffffd00000013",
            INIT_19 => X"fffffffd000000110000001afffffff8fffffffbffffffdfffffffcf0000000d",
            INIT_1A => X"fffffffb0000001f0000000d00000004000000000000000d0000000efffffffc",
            INIT_1B => X"fffffff6ffffffffffffffeffffffff1ffffffc900000000fffffff7fffffff0",
            INIT_1C => X"ffffffc0ffffffcffffffff900000019ffffffcfffffffd2fffffffc00000016",
            INIT_1D => X"0000004900000002ffffffd900000047ffffffe4ffffffe900000012fffffffd",
            INIT_1E => X"ffffffef000000140000001300000008000000180000000dfffffffc00000002",
            INIT_1F => X"ffffffd900000030ffffffe3ffffffc0ffffffe5ffffffd2ffffffe600000004",
            INIT_20 => X"00000035fffffffdffffffdffffffff400000006ffffffd300000010fffffff0",
            INIT_21 => X"000000110000001c00000013000000170000000c0000000fffffffedfffffffb",
            INIT_22 => X"00000016fffffffc000000120000001b00000016000000020000002effffffff",
            INIT_23 => X"0000001200000002fffffff2fffffff3ffffffda000000040000000affffffe2",
            INIT_24 => X"0000001bfffffff100000002fffffff7ffffffe90000000bfffffff300000019",
            INIT_25 => X"ffffffeb00000008ffffffee0000000a0000002dfffffff4ffffffe900000000",
            INIT_26 => X"ffffffd6fffffff400000023ffffffcc0000000a00000030ffffffefffffffe9",
            INIT_27 => X"0000005300000025000000460000004800000013ffffffed0000001d00000021",
            INIT_28 => X"000000200000000a0000003b00000021ffffffe900000010000000380000004f",
            INIT_29 => X"0000002dffffffcbffffff9800000021ffffffeaffffffd5ffffffe100000018",
            INIT_2A => X"fffffffd0000002c00000014ffffffe1000000020000001efffffffbffffffde",
            INIT_2B => X"fffffff2ffffffeaffffffdefffffffcfffffff80000001a0000003cffffffe0",
            INIT_2C => X"0000002dfffffff9ffffffda000000210000004e00000045fffffff30000002b",
            INIT_2D => X"0000003400000017ffffffd8ffffffd000000009fffffff8ffffffe100000000",
            INIT_2E => X"ffffffaeffffffd9ffffffd60000000affffffdd00000001000000290000000c",
            INIT_2F => X"0000004f00000011ffffffd900000017ffffffd0ffffff9b00000024ffffffe5",
            INIT_30 => X"0000000a000000080000000000000003fffffffefffffff9fffffffefffffffc",
            INIT_31 => X"00000017ffffffafffffffb000000013ffffffaeffffffb700000002ffffffff",
            INIT_32 => X"000000500000002affffffdc0000004300000028ffffffddfffffff1ffffffff",
            INIT_33 => X"00000014fffffff5fffffffb00000001ffffffe60000001dfffffffb00000006",
            INIT_34 => X"0000000dfffffffa0000002cffffffe9000000300000002dffffffe50000002a",
            INIT_35 => X"00000018ffffffedffffffe900000016fffffff9ffffffe3000000450000006e",
            INIT_36 => X"ffffffe00000000000000005fffffffcffffffe60000002c00000009ffffffe5",
            INIT_37 => X"00000006000000030000001e00000027fffffff800000006fffffff1ffffffd4",
            INIT_38 => X"ffffffe0ffffffe20000000500000002ffffffe900000005ffffffdbfffffffb",
            INIT_39 => X"ffffffe80000001700000004fffffff2fffffff900000027ffffffdbfffffffa",
            INIT_3A => X"00000004ffffffbbffffffd000000021ffffffa5ffffffe3fffffff20000000b",
            INIT_3B => X"0000000affffffd60000000700000016ffffffd2ffffffe9ffffffc8ffffffd2",
            INIT_3C => X"ffffffeeffffffde000000160000000dfffffff3fffffffb000000090000000a",
            INIT_3D => X"000000090000001e0000001effffffe2ffffffddfffffffbffffffe100000008",
            INIT_3E => X"ffffffbbffffffd700000012000000120000002b000000160000000d00000007",
            INIT_3F => X"ffffffe6ffffffd0ffffffbdffffffe800000033ffffffc30000000000000064",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE5;


    MEM_IWGHT_LAYER1_INSTANCE6 : if BRAM_NAME = "iwght_layer1_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff2ffffffdfffffffd9ffffffdf000000030000000cffffffe600000029",
            INIT_01 => X"0000000a000000030000001300000026000000360000000f0000000a00000007",
            INIT_02 => X"ffffffb9fffffff4ffffffa2ffffff9afffffffaffffff7cffffffcd0000002a",
            INIT_03 => X"00000027ffffffd7fffffff100000040ffffffe4fffffff200000018ffffffcf",
            INIT_04 => X"ffffffee00000019ffffffea0000000d0000000bfffffff0ffffffddfffffff0",
            INIT_05 => X"fffffffe00000001000000340000002bfffffff3000000000000001bfffffff8",
            INIT_06 => X"00000011000000040000001e0000001c0000000e00000014000000050000001d",
            INIT_07 => X"000000100000000000000013ffffffea0000001ffffffffaffffffee00000009",
            INIT_08 => X"fffffff7ffffffee00000000fffffffc00000000000000260000001200000007",
            INIT_09 => X"00000007000000180000001c00000000ffffffe80000000ffffffff3fffffffc",
            INIT_0A => X"fffffff50000000effffffef0000002a00000003ffffffea0000002700000011",
            INIT_0B => X"ffffffe3fffffff30000005300000014ffffffcb000000580000002affffffc9",
            INIT_0C => X"0000000bfffffff1fffffffc00000015ffffffdaffffffd70000000600000028",
            INIT_0D => X"fffffffbfffffff900000033ffffffd6000000070000000ffffffff2fffffffd",
            INIT_0E => X"00000001ffffffeeffffffecffffffe100000000ffffffc3ffffffe600000009",
            INIT_0F => X"fffffff90000001700000026000000180000001afffffff8fffffff9fffffffc",
            INIT_10 => X"fffffff800000013fffffff300000009fffffff8ffffffd8fffffffa00000007",
            INIT_11 => X"0000001ffffffff4ffffffe7ffffffe7ffffffe60000000affffffec00000018",
            INIT_12 => X"fffffff7ffffffed0000001600000009ffffffecfffffffe0000000d0000000a",
            INIT_13 => X"ffffffe900000007000000200000000f000000080000002600000003fffffff9",
            INIT_14 => X"ffffffdafffffffffffffff600000009fffffff4000000070000001000000004",
            INIT_15 => X"ffffffa4ffffffa9ffffff74ffffff8affffffa8ffffffbeffffff99fffffff8",
            INIT_16 => X"000000150000003700000010000000220000002100000012ffffffccffffffa0",
            INIT_17 => X"0000000000000022fffffffeffffffe3000000240000001afffffffb0000002b",
            INIT_18 => X"0000005f0000002c0000002900000046ffffffe4fffffffcfffffff6ffffffe4",
            INIT_19 => X"fffffff8000000040000000dfffffff100000029000000510000000400000015",
            INIT_1A => X"ffffffffffffffe2ffffffeeffffffe600000002000000060000001d00000000",
            INIT_1B => X"fffffff1fffffff6fffffffd000000190000000bfffffff3fffffffcffffffeb",
            INIT_1C => X"fffffff70000003c000000280000000b0000000a000000170000001f00000024",
            INIT_1D => X"ffffffc8ffffffc3ffffffd7ffffffa1ffffffcf00000003fffffffdfffffffd",
            INIT_1E => X"fffffff9ffffffedfffffff0ffffffedffffffffffffffe9fffffff500000016",
            INIT_1F => X"ffffffcfffffffa0ffffffd2ffffffe5ffffffe2ffffffd200000025fffffff7",
            INIT_20 => X"0000000400000018ffffffdfffffffd8ffffffdcfffffff9ffffffc9fffffff0",
            INIT_21 => X"0000000cffffffefffffffe5ffffffe8ffffffebffffffea00000009ffffffe5",
            INIT_22 => X"000000020000001b0000000d000000100000001d0000001bffffffea00000009",
            INIT_23 => X"fffffffffffffffefffffffc0000000e0000001500000013fffffff5fffffffa",
            INIT_24 => X"ffffffe8fffffff2ffffffe1fffffff80000000200000007ffffffe8ffffffe4",
            INIT_25 => X"0000000c000000180000002bffffffe8ffffffe800000014ffffffd9fffffff5",
            INIT_26 => X"ffffffeeffffffe0fffffff0ffffffd7ffffffb1ffffffefffffffd3ffffffb0",
            INIT_27 => X"0000000d00000003ffffffecfffffff8ffffffd6ffffffd9fffffff90000000f",
            INIT_28 => X"fffffff60000000bfffffff60000001900000029fffffff000000006fffffffe",
            INIT_29 => X"0000001700000005fffffffe0000000a00000005ffffffe4ffffffebfffffff4",
            INIT_2A => X"0000001400000007fffffffcfffffff8000000050000001e0000000ffffffffa",
            INIT_2B => X"fffffffcfffffff2ffffffe9ffffffdefffffffd0000001cffffffed00000006",
            INIT_2C => X"ffffffe5ffffffef0000000afffffffb00000012ffffffecfffffff6ffffffe9",
            INIT_2D => X"0000002700000014fffffff6fffffff300000008fffffff9ffffffe4fffffff4",
            INIT_2E => X"0000000400000008fffffff000000012fffffff6ffffffeb0000001200000005",
            INIT_2F => X"00000010ffffffd00000002afffffff1000000000000000ffffffffffffffffe",
            INIT_30 => X"00000008000000090000001b0000000800000020000000140000001d00000031",
            INIT_31 => X"00000006000000060000001e00000014fffffffefffffff7fffffff1ffffffed",
            INIT_32 => X"ffffffe70000000300000005ffffffeafffffffd0000003a0000000100000000",
            INIT_33 => X"0000000300000011000000290000003400000000fffffffc000000140000001f",
            INIT_34 => X"0000001500000009ffffffdb0000000c00000021000000090000000300000031",
            INIT_35 => X"0000001100000003000000000000000cfffffff50000002e00000002ffffffe1",
            INIT_36 => X"00000017ffffffddfffffff600000002fffffff70000000d0000000d0000000f",
            INIT_37 => X"0000000a000000180000002d0000001e000000170000001a0000001500000000",
            INIT_38 => X"fffffff8000000070000000affffffebfffffff7ffffffdf0000000100000008",
            INIT_39 => X"00000005ffffffed0000002d00000023fffffff30000000a0000000400000000",
            INIT_3A => X"fffffff3000000060000001e000000560000002e0000000bffffffaeffffffce",
            INIT_3B => X"0000000cffffffc6000000000000001500000004ffffffefffffffe4ffffffed",
            INIT_3C => X"fffffff3000000220000001b0000003700000013fffffff2ffffffba0000002a",
            INIT_3D => X"ffffffe1ffffffb3ffffffd9ffffffd0ffffffd7fffffff1ffffffd800000006",
            INIT_3E => X"fffffff3000000190000004400000029000000290000000fffffffb10000000c",
            INIT_3F => X"0000000bffffffe1ffffffe3fffffff400000017ffffffeaffffffdf00000012",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE6;


    MEM_IWGHT_LAYER1_INSTANCE7 : if BRAM_NAME = "iwght_layer1_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffeaffffffef00000002ffffffff0000001ffffffff10000001300000005",
            INIT_01 => X"ffffffd5ffffffe200000021fffffffe000000280000001a00000011ffffffed",
            INIT_02 => X"fffffff5ffffffd7ffffffe3ffffffeefffffff0ffffffe8ffffffd5ffffffe5",
            INIT_03 => X"ffffffedfffffffe00000033ffffffe40000000000000011fffffffbffffffe0",
            INIT_04 => X"ffffffdefffffff7fffffff2fffffff200000017ffffffddffffffeffffffff9",
            INIT_05 => X"00000012ffffffd6ffffffd8fffffffafffffff8ffffffe8fffffffbffffffe9",
            INIT_06 => X"000000310000000500000005000000310000001e000000080000000800000004",
            INIT_07 => X"ffffffad00000003ffffffea00000003ffffffe700000009000000150000001e",
            INIT_08 => X"000000000000003d0000001d0000003600000009ffffffcc00000044ffffffae",
            INIT_09 => X"00000018ffffffe50000000300000015000000110000000c000000190000000c",
            INIT_0A => X"ffffffdc0000001effffffbf0000000c00000003ffffffdbffffffe90000000d",
            INIT_0B => X"ffffffe2fffffff9fffffff6ffffffc500000002fffffff6ffffffd7ffffffd6",
            INIT_0C => X"0000004d0000004d000000100000002500000034fffffffc00000026ffffffda",
            INIT_0D => X"ffffffd800000010ffffffebffffffdf00000001ffffffedffffffff0000001c",
            INIT_0E => X"ffffffec0000000bffffffee0000002400000018ffffffff0000002600000025",
            INIT_0F => X"00000016ffffffe8ffffffedfffffffdffffffec0000000000000000ffffffdc",
            INIT_10 => X"fffffffeffffffca0000001f000000070000000c00000020ffffffe2fffffff1",
            INIT_11 => X"fffffff40000000cfffffff5ffffffec00000000fffffffaffffffdffffffff4",
            INIT_12 => X"00000028000000110000002b0000001b000000100000000cffffffebffffffbc",
            INIT_13 => X"ffffffe5ffffffdcfffffff90000003b00000026000000310000006d00000010",
            INIT_14 => X"fffffff0fffffff100000004fffffffb0000002800000013fffffff8ffffffe5",
            INIT_15 => X"0000001afffffff20000001700000009fffffffffffffff6ffffffbfffffffec",
            INIT_16 => X"0000000e00000005ffffffe0ffffffdb0000000b00000006fffffff9ffffffed",
            INIT_17 => X"fffffffd000000350000001300000018fffffff70000000600000010fffffff3",
            INIT_18 => X"ffffffdeffffffda00000002fffffffffffffff9fffffff10000000a0000000f",
            INIT_19 => X"ffffffde00000006fffffff7fffffff7ffffffecffffffe20000001900000008",
            INIT_1A => X"fffffffa00000011000000050000000200000000ffffffe500000006fffffffa",
            INIT_1B => X"00000028000000180000001f0000001d0000001bfffffffe0000000b00000001",
            INIT_1C => X"fffffff900000014000000000000001dfffffff700000001fffffffb00000008",
            INIT_1D => X"ffffffeefffffff8fffffff7fffffffafffffff800000010fffffff1fffffffe",
            INIT_1E => X"000000170000002afffffff7ffffffcafffffff8ffffffe000000023fffffff5",
            INIT_1F => X"ffffffe6ffffffdb000000080000000b0000001c000000590000006000000051",
            INIT_20 => X"00000025ffffffb1ffffffd9fffffff8ffffffdbfffffff200000019fffffff5",
            INIT_21 => X"00000013000000150000000700000014000000270000004fffffffd40000000d",
            INIT_22 => X"0000000affffffee00000001ffffffe60000000a00000003ffffffddffffffec",
            INIT_23 => X"fffffff9fffffff4fffffff20000000b00000008ffffffe1ffffffe300000019",
            INIT_24 => X"0000001e000000160000000c0000000000000002ffffffed0000001fffffffd8",
            INIT_25 => X"ffffffed0000001cffffffd90000001600000014ffffffbbffffffd800000004",
            INIT_26 => X"0000000ffffffff30000002f00000027fffffffefffffffaffffffec00000000",
            INIT_27 => X"fffffff80000000700000006ffffffc4fffffff2ffffffe2ffffffdb0000000b",
            INIT_28 => X"fffffffeffffffee0000001dfffffff1ffffffeffffffffefffffff0ffffffda",
            INIT_29 => X"fffffffa000000020000000effffffeffffffffe0000002c0000000100000032",
            INIT_2A => X"0000002d000000080000000afffffff9ffffffdcffffffd100000014fffffff5",
            INIT_2B => X"0000000e0000001500000006000000130000000cffffffdf000000180000000b",
            INIT_2C => X"ffffffe400000010ffffffe20000001200000000000000020000000100000010",
            INIT_2D => X"ffffffd30000000000000012fffffff6fffffffdffffffed0000000affffffd5",
            INIT_2E => X"fffffffc00000023000000600000004a000000710000002d0000002f00000025",
            INIT_2F => X"000000120000000c0000001500000005000000050000000dffffffe50000001f",
            INIT_30 => X"fffffff3ffffffd600000002fffffff200000001ffffffffffffffed00000007",
            INIT_31 => X"ffffffc7fffffff900000024ffffffe2fffffff7fffffff0ffffffdbffffffdb",
            INIT_32 => X"fffffff20000002a0000001300000006fffffffbfffffff1fffffff7ffffffd0",
            INIT_33 => X"0000001ffffffffdfffffff4000000040000000400000001ffffffe1ffffffca",
            INIT_34 => X"fffffff8fffffff3fffffffefffffffb00000017ffffffe3fffffff9ffffffcd",
            INIT_35 => X"00000000ffffffef0000000300000015fffffff30000000c00000024fffffff0",
            INIT_36 => X"fffffff0ffffffc1ffffffea00000024fffffff7000000030000001cffffffeb",
            INIT_37 => X"0000000200000014ffffffddffffffeefffffff5ffffffe30000001000000009",
            INIT_38 => X"0000001300000003ffffffeb000000080000000000000000ffffffff00000000",
            INIT_39 => X"fffffff70000002a0000000effffffe10000000ffffffffc0000001500000026",
            INIT_3A => X"ffffffeefffffff300000007ffffffe7ffffffd8ffffffd3ffffffec00000003",
            INIT_3B => X"fffffff9fffffffcfffffff5ffffffc2000000270000001d00000014fffffff2",
            INIT_3C => X"0000002d00000032fffffffeffffffe5fffffff300000023fffffffbfffffff6",
            INIT_3D => X"000000000000003200000014fffffffbffffffe900000042fffffff3fffffffa",
            INIT_3E => X"ffffffeffffffff6fffffff3fffffff9fffffff2ffffffd7fffffffa00000027",
            INIT_3F => X"fffffff0fffffffd0000000a000000140000001dfffffff8fffffff900000019",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE7;


    MEM_IWGHT_LAYER1_INSTANCE8 : if BRAM_NAME = "iwght_layer1_instance8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001c0000002a0000000b00000014000000090000001effffffecffffffef",
            INIT_01 => X"ffffffd60000000c000000060000002cfffffffd00000013000000270000001c",
            INIT_02 => X"00000034000000520000001400000011fffffffe0000000e0000000dffffffd4",
            INIT_03 => X"0000003d0000002b0000001f000000380000002c000000270000002100000041",
            INIT_04 => X"00000034ffffffe0fffffffc0000002dffffffdefffffffc000000020000000e",
            INIT_05 => X"000000320000000cfffffff3ffffffe7fffffff700000005ffffffe300000050",
            INIT_06 => X"ffffffdd000000020000001d0000000f0000002f0000000ffffffff7ffffffff",
            INIT_07 => X"fffffffcfffffff40000000f00000006ffffffbaffffffd6ffffffd6fffffff9",
            INIT_08 => X"000000030000001e0000001c0000000a000000260000000b00000002ffffffe7",
            INIT_09 => X"ffffffe0ffffffe4fffffff400000002fffffffefffffff0000000240000002c",
            INIT_0A => X"0000000000000000ffffffdfffffffda000000230000001e0000000800000004",
            INIT_0B => X"ffffffe5fffffff000000002ffffffe6fffffff300000025fffffffdfffffff3",
            INIT_0C => X"00000009ffffffdd00000002ffffffdf0000000fffffffe9ffffffd6fffffff8",
            INIT_0D => X"ffffffc80000000700000005ffffffd2ffffffeaffffffdc00000018fffffff3",
            INIT_0E => X"fffffff2ffffffcefffffff60000000400000007ffffffe6fffffff7ffffffe3",
            INIT_0F => X"0000001bfffffffd0000001e000000150000001c000000050000000100000029",
            INIT_10 => X"ffffffc50000001a0000003d000000420000001700000001ffffffe000000001",
            INIT_11 => X"ffffffef0000000dffffffe100000010ffffffc8ffffffa30000000afffffff3",
            INIT_12 => X"ffffffffffffffebffffffc2ffffffeb0000000afffffff6ffffffd100000043",
            INIT_13 => X"0000002200000001fffffff7000000090000001cfffffff9ffffffe200000026",
            INIT_14 => X"ffffffdfffffffe3ffffffbe0000001effffffe1ffffffd3000000020000000c",
            INIT_15 => X"fffffff3ffffffddfffffff300000005fffffff500000004fffffff900000020",
            INIT_16 => X"ffffffd70000001ffffffff100000023fffffff1ffffffe80000001c00000011",
            INIT_17 => X"000000230000002a0000000100000010fffffff5ffffffea00000018ffffffe0",
            INIT_18 => X"fffffff7fffffff800000006000000110000000b00000016fffffffdffffffe3",
            INIT_19 => X"0000003a0000002400000034fffffff00000001efffffff4ffffffcc0000000a",
            INIT_1A => X"ffffffddffffffe700000001ffffffc5ffffffd600000001fffffff8fffffff8",
            INIT_1B => X"fffffff5ffffffed0000002000000032000000250000004b00000029fffffff2",
            INIT_1C => X"ffffffeeffffffea000000120000001effffffe0ffffffe5fffffffcfffffffb",
            INIT_1D => X"00000028ffffffedfffffffc00000032ffffffecfffffffe00000000fffffff5",
            INIT_1E => X"00000004ffffffe60000000cfffffff6ffffffdf000000050000001d00000014",
            INIT_1F => X"0000001500000003000000580000001700000011ffffffea0000000c00000017",
            INIT_20 => X"0000000dffffff99ffffffc0ffffffd00000001c00000019ffffffe70000005c",
            INIT_21 => X"fffffff800000005fffffff600000015fffffffefffffff6ffffffe3ffffffe7",
            INIT_22 => X"0000000000000029000000060000000a0000000200000000fffffff40000000d",
            INIT_23 => X"fffffffefffffffe0000000400000020fffffffafffffff2000000130000000f",
            INIT_24 => X"0000000b0000000c0000001700000013000000020000000900000009fffffff4",
            INIT_25 => X"0000000e0000001000000000fffffff4000000360000001b0000002a0000000d",
            INIT_26 => X"ffffffff0000001900000042000000250000000a000000390000001d00000021",
            INIT_27 => X"ffffffcdffffffd000000013ffffffe1ffffffdc000000170000001800000015",
            INIT_28 => X"000000100000002c000000210000001bffffffc5ffffffb9ffffffbfffffffe1",
            INIT_29 => X"0000000f0000000cfffffff600000005fffffffaffffffe80000004000000043",
            INIT_2A => X"00000018fffffffdfffffffafffffff60000001e0000000000000015ffffffdb",
            INIT_2B => X"00000000ffffffeaffffffe6fffffffefffffffb000000180000000200000032",
            INIT_2C => X"000000180000000affffffe8000000000000000700000013ffffffeaffffffff",
            INIT_2D => X"fffffffb00000028fffffff00000000a0000001efffffff5ffffffd00000000d",
            INIT_2E => X"ffffffefffffffeb00000003fffffffc000000000000001a0000000500000000",
            INIT_2F => X"0000001b00000015fffffffa0000000cfffffff0000000150000000cfffffff0",
            INIT_30 => X"0000000dffffffc700000027000000130000001f0000001a000000170000001b",
            INIT_31 => X"000000000000002c0000000effffffffffffffe60000002d00000003fffffff2",
            INIT_32 => X"000000060000000dfffffff7ffffffd1ffffffe1ffffffe10000000cffffffe7",
            INIT_33 => X"00000015000000170000001100000015ffffffdd00000009000000190000000f",
            INIT_34 => X"0000000cfffffff900000011fffffffffffffff3ffffffeaffffffca00000034",
            INIT_35 => X"ffffffe900000000fffffff4000000090000000d000000050000003300000022",
            INIT_36 => X"00000022ffffffff0000002f00000006fffffff4ffffffe50000003400000002",
            INIT_37 => X"ffffffd6fffffff60000001afffffff10000001c0000001b0000002500000012",
            INIT_38 => X"ffffffccfffffff0ffffffc7ffffffccffffffccffffff9bffffffea00000001",
            INIT_39 => X"fffffffbfffffff80000000efffffffb00000000ffffffd600000015ffffffd3",
            INIT_3A => X"ffffffdaffffffda00000000ffffffeefffffff2000000080000000b00000006",
            INIT_3B => X"fffffff80000001b00000016000000080000000cffffffecfffffff1ffffffd6",
            INIT_3C => X"000000240000001b0000000efffffff90000001dffffffe5ffffffedffffffe5",
            INIT_3D => X"ffffffdbffffffebffffffde000000050000001fffffffebfffffffd00000035",
            INIT_3E => X"ffffffe10000002000000010ffffffe70000000dffffffdc0000000e00000012",
            INIT_3F => X"fffffff00000001dffffffcdffffffe900000007ffffffd5ffffffc2fffffff3",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE8;


    MEM_IWGHT_LAYER1_INSTANCE9 : if BRAM_NAME = "iwght_layer1_instance9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffebfffffffd0000000d0000001bffffffcbffffffeefffffff800000019",
            INIT_01 => X"ffffffe7fffffff400000019fffffff90000002500000019fffffff60000000e",
            INIT_02 => X"ffffffe1fffffffafffffffefffffff2fffffff5ffffffe00000000afffffff1",
            INIT_03 => X"ffffffc000000010ffffffdbffffffdaffffffd5ffffffda00000002fffffff2",
            INIT_04 => X"fffffff3ffffffe7ffffffe6ffffffc4ffffffd4ffffffddffffffeaffffffbb",
            INIT_05 => X"ffffffe5ffffffe9ffffffeb0000000100000003ffffffddfffffff2fffffff1",
            INIT_06 => X"00000025ffffffee0000000ffffffff1ffffffd1ffffffdbffffffd9ffffffc5",
            INIT_07 => X"ffffffd4ffffffdcffffffec00000000000000000000000e0000004300000039",
            INIT_08 => X"ffffffff0000000500000015fffffff9fffffff1000000160000000dfffffff0",
            INIT_09 => X"0000001f0000002700000001fffffffaffffffe9ffffffe2ffffffdffffffffb",
            INIT_0A => X"ffffffa6ffffffb3ffffffc6ffffffe1ffffffc70000000e0000001400000005",
            INIT_0B => X"ffffffc5fffffff2ffffffb3ffffffb60000001bffffffa9ffffffa9ffffffe4",
            INIT_0C => X"ffffffa0ffffffc6ffffffa8ffffffdaffffff940000001e00000019ffffffa7",
            INIT_0D => X"ffffffeaffffffd4ffffffc1ffffffa8fffffff4ffffffc4ffffff9bffffffc5",
            INIT_0E => X"fffffff2fffffff4000000100000000bfffffffb00000015fffffff0ffffffda",
            INIT_0F => X"00000029ffffffca000000000000000affffffe10000000bfffffff3ffffffdb",
            INIT_10 => X"ffffffdb0000000a000000270000000c0000002600000031fffffff10000001d",
            INIT_11 => X"00000017fffffffc0000001500000017ffffffe6000000220000000000000001",
            INIT_12 => X"fffffff000000027ffffffd4fffffffe00000036ffffffecffffffe90000000a",
            INIT_13 => X"ffffffff00000007fffffff20000001600000008fffffff60000004700000021",
            INIT_14 => X"ffffff7affffffd1ffffffbdffffff9cffffff8600000001fffffff8fffffffd",
            INIT_15 => X"00000003ffffffd1fffffff2ffffffe2ffffffe8fffffff500000015ffffffbe",
            INIT_16 => X"ffffffe80000000000000007fffffff5fffffffefffffff2fffffff400000000",
            INIT_17 => X"ffffffccffffffad00000000ffffffe400000017ffffffecfffffff2fffffffe",
            INIT_18 => X"ffffffd9ffffffd6ffffffe3ffffffd0ffffffdfffffffaeffffffd4ffffffe3",
            INIT_19 => X"0000001700000013000000080000002f0000001600000011fffffff5ffffffeb",
            INIT_1A => X"0000000c000000020000000c0000000200000012000000100000002600000033",
            INIT_1B => X"fffffffafffffff6ffffffe4fffffff4ffffffd8ffffffeefffffff1ffffffde",
            INIT_1C => X"ffffffdaffffffd8ffffffee000000100000001c00000011fffffffbffffffe9",
            INIT_1D => X"000000240000002e0000001a00000034fffffffbffffffc0ffffffbaffffffb0",
            INIT_1E => X"fffffff9fffffff0ffffffebffffffe7fffffffa0000002d0000001d0000001e",
            INIT_1F => X"0000000500000000fffffff0fffffffcfffffffa00000000ffffffef00000015",
            INIT_20 => X"000000000000000600000000000000280000000c00000017fffffff8fffffffc",
            INIT_21 => X"000000050000001a000000040000000b0000002a0000000c00000013ffffffee",
            INIT_22 => X"fffffff50000001efffffff700000003fffffffb00000011fffffff400000029",
            INIT_23 => X"000000540000007a0000002f0000006d0000004f000000330000001a00000006",
            INIT_24 => X"0000000dfffffff40000000300000032fffffffb000000130000002a00000064",
            INIT_25 => X"0000001efffffff9ffffffed00000023fffffff7fffffff8ffffffd500000010",
            INIT_26 => X"0000000d0000001b00000013fffffff2fffffff80000003affffffff00000003",
            INIT_27 => X"ffffffb1fffffff6ffffffbbfffffff8fffffff30000000bfffffffdfffffff1",
            INIT_28 => X"000000060000001500000018ffffffafffffffd2ffffffeaffffffb9ffffffa3",
            INIT_29 => X"0000002000000027fffffffffffffff80000001500000000ffffffe8ffffffdd",
            INIT_2A => X"ffffffdfffffffd3fffffff6fffffff5000000010000002100000012fffffffc",
            INIT_2B => X"0000003700000015000000140000001affffffeefffffff500000006fffffff1",
            INIT_2C => X"fffffff00000000a0000000ffffffffafffffffefffffff9fffffff900000000",
            INIT_2D => X"fffffff6ffffffcfffffff86ffffffacffffff99ffffff8bffffffb600000006",
            INIT_2E => X"0000001400000007000000020000004200000047ffffffdcffffffd6ffffffca",
            INIT_2F => X"00000009fffffff10000004400000016fffffffbffffffd7ffffffe8ffffffe8",
            INIT_30 => X"0000001c000000210000003000000030ffffffcfffffffe000000001ffffffe3",
            INIT_31 => X"0000001e0000003e000000190000000ffffffffe000000110000004d00000006",
            INIT_32 => X"ffffffd7ffffffdc0000001300000018000000070000001f0000001f0000001f",
            INIT_33 => X"fffffffa00000003ffffffebffffffd1ffffffe5ffffffd7fffffff0ffffffc2",
            INIT_34 => X"000000090000001900000024000000050000001e000000160000001000000019",
            INIT_35 => X"ffffffd1ffffffd9ffffffefffffffcbffffffddfffffff8ffffffe4fffffffa",
            INIT_36 => X"ffffffe500000004fffffffbffffffc1ffffffefffffffe4ffffffa200000000",
            INIT_37 => X"ffffffddffffffcdfffffffbffffffcbffffffbcffffffe7ffffffdf00000009",
            INIT_38 => X"ffffffe3ffffffeb00000013ffffffd0ffffffc9ffffffe6ffffffdf0000000d",
            INIT_39 => X"fffffff500000011fffffff400000000ffffffddffffffd600000012ffffffe1",
            INIT_3A => X"ffffffd4ffffffd3ffffffcf0000001800000011fffffff90000000f00000001",
            INIT_3B => X"ffffffebfffffffb00000006ffffffeeffffffc9ffffffe1ffffffd2fffffff4",
            INIT_3C => X"ffffffc3ffffffd600000000fffffff3ffffffebfffffffefffffff300000012",
            INIT_3D => X"0000002400000039fffffff4000000060000000affffffd6fffffff6ffffffe7",
            INIT_3E => X"ffffffbfffffffc7ffffffbeffffffc5ffffffa6ffffffa7ffffffeaffffffd5",
            INIT_3F => X"0000001cffffffe3ffffffef00000001ffffffdcffffffbfffffffdeffffffb7",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE9;


    MEM_IWGHT_LAYER1_INSTANCE10 : if BRAM_NAME = "iwght_layer1_instance10" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000007ffffffe9ffffffe8000000270000000e0000001effffffe600000000",
            INIT_01 => X"000000270000000f00000006fffffffe00000008ffffffef00000000ffffffaa",
            INIT_02 => X"ffffffef000000200000000fffffffeb0000002f00000017fffffff900000022",
            INIT_03 => X"fffffffffffffffcfffffff80000001900000016fffffff90000000300000010",
            INIT_04 => X"ffffffdaffffffc2000000160000001a000000010000000c000000080000000a",
            INIT_05 => X"00000018fffffffdffffffeb0000000cffffffe4fffffff5ffffffccffffffc5",
            INIT_06 => X"fffffffa0000000cfffffff6ffffffef0000001500000019000000110000000a",
            INIT_07 => X"ffffffdeffffffa400000005fffffff2ffffffb7ffffffff0000002bffffffed",
            INIT_08 => X"fffffff500000005fffffff2ffffffff000000250000002a0000001000000006",
            INIT_09 => X"fffffffafffffff3fffffff00000000ffffffffbffffffe700000005ffffffe6",
            INIT_0A => X"00000008ffffffe5ffffffe0ffffffc8ffffffebfffffff800000009fffffff3",
            INIT_0B => X"0000000800000037000000130000001c0000000400000000ffffffbefffffff6",
            INIT_0C => X"ffffffd900000005fffffffa00000012ffffffadffffffe3fffffff200000000",
            INIT_0D => X"0000003200000019ffffffcb00000002ffffffe1ffffffdffffffff2ffffffd6",
            INIT_0E => X"00000000000000170000001afffffff8000000110000001ffffffff80000000c",
            INIT_0F => X"00000004fffffffd0000002afffffffd000000160000001200000000ffffffeb",
            INIT_10 => X"ffffffe9000000000000000a000000030000000d00000014ffffffeeffffffee",
            INIT_11 => X"fffffff50000000a0000001c000000050000003e0000000f0000001600000017",
            INIT_12 => X"0000000e0000001bfffffffc0000000100000000ffffffe90000000300000000",
            INIT_13 => X"00000006000000320000000fffffffe3ffffffce0000001c0000000afffffff4",
            INIT_14 => X"0000000b00000002fffffffcffffffee000000000000000b0000002fffffffe7",
            INIT_15 => X"0000000300000018fffffff700000007fffffffc0000002200000008fffffffb",
            INIT_16 => X"0000001b000000000000002200000004ffffffef00000009ffffffeeffffffed",
            INIT_17 => X"ffffffea0000000fffffffffffffffee0000001800000001000000030000000f",
            INIT_18 => X"0000005000000018000000480000003100000017ffffffe50000002500000000",
            INIT_19 => X"0000000100000028ffffffdc000000340000001bffffffc7ffffffdd0000001e",
            INIT_1A => X"ffffffa9ffffffd8fffffffeffffffedfffffff20000002200000011fffffff7",
            INIT_1B => X"ffffffe50000000dfffffff900000011000000000000001bffffffd0ffffffe2",
            INIT_1C => X"ffffffcaffffffd30000002cfffffff00000000dfffffff200000009ffffffe6",
            INIT_1D => X"ffffffe7000000240000002600000023ffffffebffffffd4ffffffc4ffffffc8",
            INIT_1E => X"000000200000002b0000001400000013fffffff9fffffff900000008ffffffe1",
            INIT_1F => X"ffffffddfffffff200000043fffffff700000011000000190000001bfffffff7",
            INIT_20 => X"0000004a0000003e0000003d0000002cffffffdfffffffe5ffffffecffffffde",
            INIT_21 => X"ffffffc6ffffffc2ffffffbe00000000fffffff8ffffffe40000002100000046",
            INIT_22 => X"ffffffefffffffd10000000c0000001cffffffecffffffb4ffffffd1ffffffc7",
            INIT_23 => X"ffffffb6fffffff6fffffffeffffffe20000000f0000002500000021ffffffdf",
            INIT_24 => X"fffffff80000003100000002ffffffd3ffffffdeffffffe100000003fffffffa",
            INIT_25 => X"fffffffaffffffe9fffffff5ffffffff0000000dffffffcdffffffe9ffffffba",
            INIT_26 => X"000000130000000e0000000a000000000000001effffffe5fffffff0ffffffea",
            INIT_27 => X"000000160000001e0000002100000004ffffffedfffffffb0000002e00000011",
            INIT_28 => X"0000002d0000005200000003ffffffdc0000000e00000013fffffff1fffffff5",
            INIT_29 => X"ffffffccfffffff6fffffff1fffffff6ffffffce00000000000000000000001a",
            INIT_2A => X"0000001200000012ffffffeafffffff8ffffffe2ffffffe9ffffffd0ffffffac",
            INIT_2B => X"ffffffd4fffffff5ffffffe1ffffffeffffffff4ffffffafffffffa5ffffffd8",
            INIT_2C => X"0000002a0000000c000000340000000efffffff7ffffffd7ffffffb2ffffffbc",
            INIT_2D => X"ffffffdbfffffff5ffffffd0fffffffc0000000efffffffefffffffdfffffff7",
            INIT_2E => X"00000012000000000000000f000000000000000f0000000fffffffebffffffb2",
            INIT_2F => X"0000001dffffffcafffffff1fffffff000000037fffffff2ffffffe300000014",
            INIT_30 => X"fffffff20000000700000018ffffffcc000000000000000fffffffcdfffffffa",
            INIT_31 => X"ffffffe8ffffffd60000003cfffffff2000000010000003b00000015fffffffe",
            INIT_32 => X"000000100000000b0000001e0000001b00000022000000230000001bfffffffc",
            INIT_33 => X"ffffffe8ffffffeeffffffcc0000000b00000000ffffffe30000001c00000029",
            INIT_34 => X"0000000200000015fffffffcfffffff40000000e0000001a000000060000000c",
            INIT_35 => X"000000420000003e00000040000000430000002a0000004b00000033fffffff9",
            INIT_36 => X"ffffffbcffffff8affffffbcfffffff5ffffffbafffffff00000003a00000038",
            INIT_37 => X"ffffffc0ffffffdeffffffe3ffffffdfffffffdeffffffdaffffff94ffffffbe",
            INIT_38 => X"ffffffc4ffffffe6ffffffe2fffffff7ffffffe5ffffffe4ffffffa2ffffffef",
            INIT_39 => X"ffffffd9ffffffe9fffffffaffffffe1ffffffbeffffff860000000cffffffbb",
            INIT_3A => X"00000042fffffffe000000420000002f00000037ffffffff000000000000000c",
            INIT_3B => X"0000000effffffefffffffe0ffffffdc0000000dffffffebfffffff700000027",
            INIT_3C => X"000000080000001500000027000000050000002100000010fffffffb00000001",
            INIT_3D => X"000000100000000c0000000afffffff10000001e00000022000000150000000a",
            INIT_3E => X"ffffffcb0000000200000005ffffffdb0000001b0000000b0000001400000038",
            INIT_3F => X"00000029fffffff5000000220000000d000000100000002100000003ffffffdb",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE10;


    MEM_IWGHT_LAYER1_INSTANCE11 : if BRAM_NAME = "iwght_layer1_instance11" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff7fffffff0ffffffd8fffffff0fffffff800000017fffffffdffffffee",
            INIT_01 => X"ffffffefffffffebffffffe90000000b0000000a0000001effffffe4ffffffe7",
            INIT_02 => X"000000160000002100000013fffffff20000000cfffffffffffffff1fffffff3",
            INIT_03 => X"ffffffe90000000c0000000900000007ffffffed000000320000003100000014",
            INIT_04 => X"ffffffe400000006000000100000001efffffffb00000000ffffffedfffffffe",
            INIT_05 => X"0000000900000010fffffffa0000000300000000ffffffdaffffffe9fffffffc",
            INIT_06 => X"00000013000000200000003a00000048fffffff90000005e0000005d00000033",
            INIT_07 => X"fffffff700000000000000050000000afffffffd0000001e0000000e00000025",
            INIT_08 => X"ffffffe60000000dffffffe3ffffffe800000000ffffffea0000000d0000000e",
            INIT_09 => X"fffffff6000000010000001f0000000f0000001dffffffe4fffffff8ffffffe8",
            INIT_0A => X"0000000fffffffeafffffff5ffffffd200000019000000140000001400000008",
            INIT_0B => X"00000003000000190000001100000007000000020000001affffffe700000018",
            INIT_0C => X"000000120000001c00000011000000070000000bffffffe60000000ffffffffc",
            INIT_0D => X"0000000300000003fffffff6fffffff40000001c000000110000000300000029",
            INIT_0E => X"fffffff300000004ffffffd3000000060000000dfffffff900000004fffffff1",
            INIT_0F => X"ffffff70ffffff97ffffffc3ffffff94ffffffb7fffffff7ffffffdeffffffbb",
            INIT_10 => X"00000004000000230000000f0000001000000024000000210000000affffffc0",
            INIT_11 => X"000000090000002dffffffd80000002100000013000000030000001900000011",
            INIT_12 => X"fffffffb0000000a000000090000001800000032000000060000000affffffe6",
            INIT_13 => X"ffffffd2fffffff4ffffffd4fffffff6ffffffec0000001000000025ffffffed",
            INIT_14 => X"00000001ffffffe9ffffffef00000008ffffffe7ffffffc800000009ffffffd5",
            INIT_15 => X"ffffffe8fffffff1ffffffdfffffffea00000004ffffffea0000000800000009",
            INIT_16 => X"fffffff000000000000000150000000d000000030000001200000018ffffffe6",
            INIT_17 => X"0000000900000000fffffffb000000030000000e00000003fffffffc0000000f",
            INIT_18 => X"0000000a00000003000000030000000bffffffea00000000ffffffeaffffffeb",
            INIT_19 => X"ffffffd4ffffffe2ffffffc7ffffffeffffffffc00000004000000110000000a",
            INIT_1A => X"ffffffedffffff9affffffabffffffccffffffc1ffffffc2ffffffdeffffffd8",
            INIT_1B => X"0000000300000029ffffffd6fffffff70000000900000015fffffffb0000000b",
            INIT_1C => X"ffffffb2ffffffb3ffffffc1ffffff96fffffffe0000003500000036ffffffe5",
            INIT_1D => X"00000033000000420000001a000000050000002400000005ffffffe9ffffffd6",
            INIT_1E => X"ffffffe9ffffffd8ffffffd6fffffff1ffffffcf000000270000001600000000",
            INIT_1F => X"0000001b0000002cffffffeb00000009ffffffe5ffffffdeffffffa3ffffffbf",
            INIT_20 => X"000000340000000a0000001c0000001e00000000fffffff70000000f0000000e",
            INIT_21 => X"ffffffe7ffffffcbfffffff6ffffffcaffffffdafffffff9fffffffdfffffffa",
            INIT_22 => X"fffffff800000007ffffffed00000001fffffffc0000001400000010ffffffee",
            INIT_23 => X"ffffffedfffffff3ffffffd8fffffff500000007fffffff2ffffffee0000000a",
            INIT_24 => X"0000000c00000008000000070000001d000000140000002400000029fffffff3",
            INIT_25 => X"000000020000001800000003fffffffcffffffc60000001efffffffafffffff2",
            INIT_26 => X"ffffffd3ffffffd6ffffffdbffffffda000000010000000000000005fffffff9",
            INIT_27 => X"000000360000000e0000003b000000300000004dfffffff2fffffff900000003",
            INIT_28 => X"ffffffe9ffffffe3ffffffedffffffc4ffffffec0000000effffffe700000018",
            INIT_29 => X"00000000ffffffedffffffd8ffffffebfffffffdfffffffdfffffff100000001",
            INIT_2A => X"000000360000001700000034000000100000000bffffffd50000000700000004",
            INIT_2B => X"00000008fffffffffffffff10000001b00000006fffffff5fffffff400000016",
            INIT_2C => X"ffffffff00000005fffffff0ffffffd2fffffff9ffffffd60000000b00000014",
            INIT_2D => X"00000015ffffffed0000001b0000000cfffffffbffffffe40000000a0000002a",
            INIT_2E => X"0000001ffffffff40000000d0000000c0000001300000005ffffffeffffffff6",
            INIT_2F => X"ffffffff0000001000000031ffffffeb00000004fffffff7fffffff60000001c",
            INIT_30 => X"0000001afffffffd00000014ffffffeeffffffd2ffffffe70000000efffffffa",
            INIT_31 => X"00000003fffffff700000006ffffffeb0000002800000015000000020000000c",
            INIT_32 => X"000000110000001a0000000dffffffecfffffff600000006000000120000000f",
            INIT_33 => X"0000000effffffc60000005000000034ffffffcf0000002d0000001dffffffc4",
            INIT_34 => X"0000002affffffe600000000ffffffe2ffffffcbffffffcdffffffc90000008d",
            INIT_35 => X"fffffff3ffffffeffffffff400000004fffffff3000000010000002e0000003a",
            INIT_36 => X"fffffff1ffffffe50000000a00000008ffffffe4000000010000002000000031",
            INIT_37 => X"0000002affffffd9fffffff4fffffff00000001600000015ffffffbffffffff9",
            INIT_38 => X"000000160000002e00000011ffffffeb0000003600000037ffffffe700000009",
            INIT_39 => X"0000000e000000220000001dffffffe9ffffffd80000000d00000006ffffffea",
            INIT_3A => X"00000025fffffff8000000100000001bfffffffd0000001e00000025fffffff3",
            INIT_3B => X"fffffffa000000220000001cffffffd900000016000000360000002800000017",
            INIT_3C => X"00000017000000040000001a0000000a000000060000000c00000008fffffffe",
            INIT_3D => X"00000005000000180000000600000003fffffff300000004fffffff7fffffff5",
            INIT_3E => X"ffffffe9ffffffeafffffff0fffffff3fffffffa0000000fffffffed00000030",
            INIT_3F => X"ffffffea00000006ffffffd1ffffffe2fffffff7fffffffbffffffd900000015",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE11;


    MEM_IWGHT_LAYER1_INSTANCE12 : if BRAM_NAME = "iwght_layer1_instance12" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffdefffffffaffffffbfffffffe20000004d0000001a000000020000002c",
            INIT_01 => X"0000000fffffffecfffffff4ffffffaaffffffa3fffffffeffffffffffffffd2",
            INIT_02 => X"0000002500000021fffffff1ffffffe2ffffffecfffffffbfffffff300000000",
            INIT_03 => X"ffffffec00000000ffffffc5ffffffc5ffffffd6ffffffa8ffffffa2fffffff1",
            INIT_04 => X"0000002e0000000effffffe00000000afffffff0ffffffca000000070000001b",
            INIT_05 => X"fffffff3fffffffbffffffea0000000600000004000000110000001500000022",
            INIT_06 => X"00000011ffffffd50000000600000016ffffffc9ffffffe50000000affffffe9",
            INIT_07 => X"ffffffe4000000220000001d0000001f000000160000000affffffacfffffff2",
            INIT_08 => X"0000000800000007fffffff9fffffff600000000ffffffd5ffffffecffffffea",
            INIT_09 => X"ffffffd8ffffffe4ffffffe9ffffffe1000000090000000a00000022ffffffef",
            INIT_0A => X"fffffff500000023000000180000000600000002ffffffe100000001fffffff9",
            INIT_0B => X"000000050000000b0000000e00000006000000160000000b0000001dfffffffd",
            INIT_0C => X"fffffff8ffffffd1ffffffabffffffc6ffffffee000000150000000600000001",
            INIT_0D => X"fffffff400000003fffffff5fffffff2fffffffc00000028ffffffedfffffffd",
            INIT_0E => X"0000000d0000000c000000020000003b00000047000000210000002600000036",
            INIT_0F => X"fffffff9fffffff80000002100000005000000000000000ffffffff700000002",
            INIT_10 => X"fffffff500000026ffffffdffffffffb000000270000002300000006ffffffe2",
            INIT_11 => X"ffffffedfffffff1000000140000000d0000000effffffc7fffffff3ffffffb5",
            INIT_12 => X"ffffffe10000001c0000002f00000033ffffffffffffffd1ffffffbb00000007",
            INIT_13 => X"000000210000001d0000003300000002ffffffdeffffffc200000015ffffffcf",
            INIT_14 => X"ffffffd9ffffffec00000023ffffffcbffffffe00000000dfffffff80000000e",
            INIT_15 => X"fffffffdffffffff0000000900000010ffffffd90000000700000006ffffffff",
            INIT_16 => X"ffffffdaffffffc3ffffff9d0000000f000000100000000c0000002000000024",
            INIT_17 => X"ffffffc20000002400000006ffffffb100000028fffffff7ffffffe800000036",
            INIT_18 => X"ffffffee0000000ffffffff400000009000000050000000300000004ffffffd8",
            INIT_19 => X"fffffff20000002a0000000ffffffff100000026000000220000001900000001",
            INIT_1A => X"fffffff6fffffffbffffffd0ffffffe4ffffffe7ffffffcc000000240000000b",
            INIT_1B => X"ffffffe1ffffffe9ffffffd800000006fffffff9ffffffd4ffffffeaffffffed",
            INIT_1C => X"fffffff2fffffffbffffffee00000034000000030000000700000012ffffffef",
            INIT_1D => X"0000000b0000001dffffffe8ffffffde0000000cfffffff8ffffffecffffffe9",
            INIT_1E => X"0000000a00000027ffffffd4ffffffadfffffffcffffffffffffffd900000002",
            INIT_1F => X"fffffffb0000001d00000029fffffff30000002c00000022ffffffe000000013",
            INIT_20 => X"0000000a000000160000000dfffffff600000013000000040000001800000001",
            INIT_21 => X"000000100000003500000028000000130000001bfffffffa0000000000000001",
            INIT_22 => X"000000120000002d0000001ffffffff4000000210000003bffffffef00000031",
            INIT_23 => X"ffffffe3ffffffc9ffffffeffffffff800000013fffffff900000001ffffffd9",
            INIT_24 => X"00000000000000130000000600000028fffffff1ffffffd600000004ffffffed",
            INIT_25 => X"fffffff8ffffffd4ffffffe6ffffffff0000000d000000070000000400000023",
            INIT_26 => X"fffffff6ffffffe4ffffffd5ffffffb9fffffff3ffffffd9ffffffbeffffffe2",
            INIT_27 => X"fffffffd0000000900000011ffffffe20000000c0000001ffffffff800000009",
            INIT_28 => X"000000290000001fffffffe40000000e000000200000000400000000fffffff6",
            INIT_29 => X"fffffff3ffffffe00000000affffffedfffffff9fffffff6fffffff600000011",
            INIT_2A => X"fffffffeffffffeb000000060000002dfffffffffffffffcfffffffe0000000e",
            INIT_2B => X"0000001000000020000000190000001a0000002000000027ffffffd7fffffff6",
            INIT_2C => X"fffffffeffffffc40000001800000003000000050000001efffffff7fffffffa",
            INIT_2D => X"ffffffe40000000e0000001c00000006ffffffe0ffffffd4fffffff700000000",
            INIT_2E => X"ffffffe7ffffffd9ffffffedffffffd8fffffff600000006fffffff6fffffff8",
            INIT_2F => X"ffffffd2fffffff0ffffffe700000004fffffffd0000000c0000001dffffffe8",
            INIT_30 => X"00000011fffffff4ffffffcefffffff2ffffffe9ffffffbdffffffe8fffffff0",
            INIT_31 => X"ffffffd8fffffffd00000032fffffff0ffffffdd000000250000000a00000008",
            INIT_32 => X"00000018ffffffdaffffffce00000017ffffffcb0000001000000030fffffff3",
            INIT_33 => X"ffffffd80000002f00000012fffffffefffffff80000002c0000001d00000001",
            INIT_34 => X"fffffff90000002b000000360000001effffffe600000012ffffffe900000017",
            INIT_35 => X"ffffffd1fffffffd0000000b0000001000000012ffffffe1ffffffd900000039",
            INIT_36 => X"000000120000000e0000001000000008fffffffaffffffe2fffffffc00000000",
            INIT_37 => X"0000000a000000110000000bffffffe6ffffffdeffffffebfffffff6ffffffe7",
            INIT_38 => X"fffffff1ffffffdefffffff4ffffffe9000000050000000dffffffd4fffffff4",
            INIT_39 => X"00000020fffffff4fffffff3000000080000000dfffffff8fffffffa00000015",
            INIT_3A => X"00000033fffffffbfffffff10000000dfffffff0fffffffe0000000c00000000",
            INIT_3B => X"000000010000001afffffff80000000400000009fffffff7ffffffd600000011",
            INIT_3C => X"ffffffd7000000290000003c000000110000000c000000220000001000000003",
            INIT_3D => X"00000000000000080000000f0000000000000002fffffffa0000001d00000029",
            INIT_3E => X"00000006ffffffc80000001dfffffff600000003ffffffd60000000500000045",
            INIT_3F => X"ffffffd100000001ffffffecfffffff2ffffffd1fffffffcfffffff1ffffffe7",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE12;


    MEM_IWGHT_LAYER1_INSTANCE13 : if BRAM_NAME = "iwght_layer1_instance13" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000ffffffe5fffffff8ffffffd5ffffffa9ffffffe7ffffffdcffffffbe",
            INIT_01 => X"0000000000000004ffffffd80000002b00000003ffffffc1ffffffcdffffffe1",
            INIT_02 => X"000000050000000900000002ffffffee00000001fffffffdfffffff7fffffffa",
            INIT_03 => X"ffffffe0fffffff10000001c00000019fffffffb00000020000000050000000e",
            INIT_04 => X"fffffff00000000afffffff2fffffffe0000000a00000010fffffff6fffffff6",
            INIT_05 => X"00000028ffffffc4ffffffeb00000025ffffffdbffffffc9ffffffdefffffff5",
            INIT_06 => X"0000000dfffffff0ffffffe6ffffffd6ffffffc7ffffffe3ffffffec00000004",
            INIT_07 => X"fffffffbffffffe6ffffffd8ffffffb8fffffff4000000290000000affffffdb",
            INIT_08 => X"ffffffeeffffffc8ffffffb7ffffffea00000033fffffff0ffffffe800000028",
            INIT_09 => X"ffffffeefffffffbffffffda0000004d00000054fffffff200000010ffffffea",
            INIT_0A => X"000000170000001b0000002f0000002900000029ffffffe60000000effffffe2",
            INIT_0B => X"00000028ffffffc2ffffffc7ffffffd90000001a000000310000001effffffff",
            INIT_0C => X"00000011ffffffedfffffff0000000180000003a0000003f0000001300000018",
            INIT_0D => X"000000490000002effffffeefffffffafffffff1ffffffecfffffff5ffffffcf",
            INIT_0E => X"ffffffc80000003a0000002000000028000000240000001a0000001800000010",
            INIT_0F => X"0000000300000007fffffff9ffffffd9ffffffddffffffcffffffff5ffffffd7",
            INIT_10 => X"0000002800000000fffffff4ffffffdcffffffdc00000000000000210000000c",
            INIT_11 => X"00000006ffffffedfffffffb00000009000000350000000cffffffe40000000a",
            INIT_12 => X"000000250000000e0000004200000012fffffff7fffffff9fffffff800000015",
            INIT_13 => X"ffffffe5ffffffa2fffffff0ffffffc3ffffffee00000019000000280000006e",
            INIT_14 => X"000000050000000d0000003f00000023000000090000003c00000000ffffffbc",
            INIT_15 => X"ffffffedffffffdb0000000dfffffff5ffffffe5ffffffedfffffffa00000014",
            INIT_16 => X"000000350000001500000046000000300000005100000031000000300000002c",
            INIT_17 => X"ffffffdcfffffffc00000000fffffffffffffff2fffffffd000000050000000e",
            INIT_18 => X"00000001ffffffeeffffffe10000000d00000004fffffff1ffffffeeffffffcd",
            INIT_19 => X"ffffffff00000000ffffffc0ffffffecffffffd2ffffffd500000006ffffffd7",
            INIT_1A => X"00000017ffffffccffffffe0ffffffdc000000020000003500000019ffffffdf",
            INIT_1B => X"ffffffbefffffff9ffffffebfffffff90000003b0000003bfffffff70000001a",
            INIT_1C => X"0000000700000024000000030000003500000042ffffffdefffffffa0000000f",
            INIT_1D => X"ffffffcbffffffeeffffffcbffffffdc00000001fffffffb0000001300000012",
            INIT_1E => X"ffffffcf0000000c0000000affffffed0000002d00000001ffffffecffffffd5",
            INIT_1F => X"00000018ffffffcc0000001800000040ffffffd80000000000000034ffffffb9",
            INIT_20 => X"fffffffc000000040000000500000045ffffffe2ffffffc9000000230000004b",
            INIT_21 => X"0000003cfffffffafffffff30000001a0000002dfffffff8ffffffe1ffffffe5",
            INIT_22 => X"00000023000000140000002d000000440000001efffffffaffffffbeffffffe1",
            INIT_23 => X"0000000d0000000affffffd5ffffffeffffffff100000008ffffffef0000001c",
            INIT_24 => X"00000048000000430000000c0000003afffffffdfffffff100000013ffffffda",
            INIT_25 => X"ffffffe800000002ffffffd5ffffffd7ffffffbd0000002f0000001d0000000d",
            INIT_26 => X"00000003fffffff70000000d0000002a000000100000002a00000022ffffffec",
            INIT_27 => X"00000001ffffffefffffffea00000013ffffffe7fffffffd0000002c00000018",
            INIT_28 => X"00000007fffffff7fffffff20000000a0000000800000000fffffffa00000000",
            INIT_29 => X"fffffff5fffffff5fffffff600000002fffffff400000013ffffffed00000012",
            INIT_2A => X"fffffff0fffffff3fffffff90000000a00000007fffffffcfffffffafffffff3",
            INIT_2B => X"ffffffff00000000fffffff50000000e00000000fffffffbfffffff900000010",
            INIT_2C => X"00000000ffffffe6ffffffedfffffffd0000000bfffffff40000000700000002",
            INIT_2D => X"000000030000000000000005fffffff9ffffffffffffffee00000000fffffffc",
            INIT_2E => X"fffffff6fffffffefffffff1fffffffcffffffebfffffff4fffffff4fffffff7",
            INIT_2F => X"fffffff3fffffff6000000040000000000000000ffffffecfffffffd00000010",
            INIT_30 => X"fffffffa000000030000001000000004ffffffe9000000010000000dfffffff4",
            INIT_31 => X"00000000fffffffcfffffffbfffffff0fffffffdffffffef00000009fffffff1",
            INIT_32 => X"0000000300000011000000030000000a0000000a000000000000000afffffffb",
            INIT_33 => X"00000004fffffffe00000002fffffffb00000013fffffffdfffffff5fffffff6",
            INIT_34 => X"fffffff50000000c0000000700000006fffffff9fffffffdfffffff100000017",
            INIT_35 => X"fffffff700000002ffffffec0000000f000000070000000000000000fffffff3",
            INIT_36 => X"0000000bffffffeb00000006fffffffd0000000d000000000000000100000003",
            INIT_37 => X"0000000efffffffdfffffffbfffffff7fffffff5fffffff000000002ffffffef",
            INIT_38 => X"00000003fffffff4ffffffecfffffff10000000bfffffff90000000000000000",
            INIT_39 => X"ffffffea00000011ffffffecffffffff00000006ffffffeaffffffea00000000",
            INIT_3A => X"00000005fffffff50000000f0000000cfffffff0ffffffee0000001100000010",
            INIT_3B => X"0000000400000007fffffff500000000fffffff6fffffff8ffffffeb0000000e",
            INIT_3C => X"fffffffb00000007fffffff30000000200000011000000150000000afffffff1",
            INIT_3D => X"0000000cfffffff3ffffffed0000000e00000003fffffff0fffffff9fffffffa",
            INIT_3E => X"00000004ffffffe8fffffffffffffff900000002ffffffff0000000efffffff3",
            INIT_3F => X"fffffff40000000b00000006fffffffd00000003fffffff5000000020000000d",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE13;


    MEM_IWGHT_LAYER1_INSTANCE14 : if BRAM_NAME = "iwght_layer1_instance14" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000dfffffff00000000affffffeb000000090000000afffffff4ffffffe9",
            INIT_01 => X"fffffffdfffffff900000012ffffffeeffffffe900000005fffffffafffffffc",
            INIT_02 => X"ffffffeaffffffedfffffff300000004fffffff0fffffff2fffffff4fffffff1",
            INIT_03 => X"fffffffe000000050000000afffffffe00000003fffffff6fffffff8fffffff0",
            INIT_04 => X"00000003fffffff9fffffff300000004ffffffe8fffffffefffffff4ffffffe8",
            INIT_05 => X"fffffff60000000f000000050000000bfffffff6fffffffe00000000fffffffe",
            INIT_06 => X"fffffffbffffffeffffffff500000009fffffff60000000d0000000700000011",
            INIT_07 => X"fffffff80000000400000000fffffff6ffffffee00000004ffffffebfffffffa",
            INIT_08 => X"fffffff2fffffff800000000fffffff500000003fffffff6fffffff500000001",
            INIT_09 => X"00000009ffffffeaffffffec0000000700000000fffffffcfffffff9ffffffeb",
            INIT_0A => X"0000000600000003fffffffbfffffff7fffffff900000000ffffffeefffffff3",
            INIT_0B => X"ffffffe9fffffff4fffffff3ffffffeefffffffbfffffff9ffffffff00000008",
            INIT_0C => X"ffffffe900000006ffffffe700000008fffffff8fffffffefffffffafffffff8",
            INIT_0D => X"fffffffaffffffd5ffffffe9fffffffd0000000200000015fffffffdffffffee",
            INIT_0E => X"0000001f00000014fffffffcffffffdffffffffcffffffddfffffff3ffffffe4",
            INIT_0F => X"000000180000003a00000040000000480000001d00000028000000430000002e",
            INIT_10 => X"00000030ffffffdafffffff2fffffff9ffffffe6000000020000000b0000001e",
            INIT_11 => X"fffffff7ffffffe0fffffffb00000033000000310000002cfffffff00000000b",
            INIT_12 => X"0000000affffffeaffffffe100000017ffffffe9ffffffeefffffffdffffffe0",
            INIT_13 => X"00000005ffffffe9fffffff6fffffff4fffffff7ffffffd7fffffffefffffffe",
            INIT_14 => X"0000000000000027000000200000002600000022000000130000000400000018",
            INIT_15 => X"ffffffe90000000d00000001fffffff40000001b000000190000001c00000016",
            INIT_16 => X"00000022ffffffe5ffffffc3ffffffdbffffffe8ffffff9affffffb200000006",
            INIT_17 => X"ffffffefffffffdbfffffff2000000020000002f000000080000002400000000",
            INIT_18 => X"ffffffc4ffffffd2ffffffe6ffffffc1ffffffc9ffffffe0ffffffe80000000c",
            INIT_19 => X"fffffffcffffffe5ffffffce00000001ffffffcfffffffbfffffffeeffffffd5",
            INIT_1A => X"000000020000000cffffffed000000100000002100000013fffffff500000003",
            INIT_1B => X"ffffffee000000160000002e0000000d00000017fffffffe0000000500000002",
            INIT_1C => X"ffffffeaffffffeffffffff90000000100000015fffffff200000010fffffff6",
            INIT_1D => X"0000001e0000000900000007fffffff9fffffff2ffffffddfffffff2ffffffd1",
            INIT_1E => X"ffffffe0ffffffe5ffffffddffffffaeffffffafffffffefffffffc6ffffffcf",
            INIT_1F => X"fffffffd00000009ffffffc300000000fffffffffffffff7ffffffc7ffffffcd",
            INIT_20 => X"ffffffb1ffffffb1ffffffb8fffffff40000001b0000000100000007fffffff8",
            INIT_21 => X"0000002c00000026ffffffec0000000900000028ffffffc7ffffffa3ffffffba",
            INIT_22 => X"00000013fffffff400000001000000150000001f000000130000002500000006",
            INIT_23 => X"ffffffec0000000b00000027fffffff5ffffffecffffffdefffffff1ffffffeb",
            INIT_24 => X"ffffffebffffffd500000009fffffffa0000000900000004000000130000002b",
            INIT_25 => X"fffffffe0000001c0000000a0000001600000006ffffffd1fffffff2fffffff6",
            INIT_26 => X"ffffffff00000007fffffff900000004fffffffffffffff30000001400000007",
            INIT_27 => X"fffffffb00000000fffffffd000000290000002c000000190000003000000020",
            INIT_28 => X"000000230000002400000007000000230000002000000042000000240000000b",
            INIT_29 => X"00000007fffffffcffffffc7fffffff7ffffffbdffffffb70000001700000001",
            INIT_2A => X"00000028fffffffcfffffffbffffffe200000017000000200000000bfffffffd",
            INIT_2B => X"00000024000000240000002e0000004100000013000000060000000a0000001f",
            INIT_2C => X"0000000cffffffcaffffffdcfffffff0ffffffee0000000b0000001400000014",
            INIT_2D => X"000000100000000f00000001000000080000000d00000003ffffffda00000004",
            INIT_2E => X"ffffffedfffffff2ffffffeffffffff50000001d0000000b0000002800000013",
            INIT_2F => X"00000022000000140000000b00000010ffffffdcffffffbe00000002ffffffb8",
            INIT_30 => X"00000006fffffffdfffffff7fffffff60000000700000015fffffff900000000",
            INIT_31 => X"0000000300000023fffffff900000003000000280000001300000035ffffffe9",
            INIT_32 => X"000000150000002e0000002d0000003cfffffffc0000002a0000000200000000",
            INIT_33 => X"ffffffdffffffff7ffffffe9fffffff1ffffffc800000016000000300000002c",
            INIT_34 => X"00000037ffffffcc00000019ffffffefffffffcf0000000c00000012ffffffee",
            INIT_35 => X"ffffffd8ffffffddffffffdb000000020000001d000000140000001400000035",
            INIT_36 => X"000000380000004d000000070000001e0000000e00000023000000270000000e",
            INIT_37 => X"0000001cffffffc3ffffffc7fffffff5000000200000001c0000000e00000033",
            INIT_38 => X"fffffffbffffffc9ffffffe8ffffffd3fffffff7ffffffe90000001600000033",
            INIT_39 => X"0000001b000000120000002a0000002c0000000100000007fffffff80000002e",
            INIT_3A => X"00000026ffffffe7ffffffdf0000002bfffffffe000000110000002c00000017",
            INIT_3B => X"0000003300000000ffffffdd00000006ffffffeb00000001ffffffef00000000",
            INIT_3C => X"0000001fffffffe20000000e0000002dfffffff6fffffff3fffffff2ffffffe9",
            INIT_3D => X"0000000a00000004000000040000001bffffffe0ffffffdc000000070000001e",
            INIT_3E => X"000000350000001200000030ffffffe3fffffff800000006ffffffdf00000011",
            INIT_3F => X"0000000d0000000cffffffe9ffffffe5fffffff2ffffffddffffffe200000002",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE14;


    MEM_IWGHT_LAYER1_INSTANCE15 : if BRAM_NAME = "iwght_layer1_instance15" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000006000000180000003e00000010000000210000003f00000010ffffffed",
            INIT_01 => X"00000001ffffffe7fffffff6ffffffe5fffffffa0000001d0000000300000008",
            INIT_02 => X"ffffffd6ffffffd100000029ffffffef0000000b00000013fffffffbffffffe4",
            INIT_03 => X"fffffff600000027fffffff40000000500000028000000100000001afffffff9",
            INIT_04 => X"000000090000000400000018fffffff500000006fffffff6ffffffe9ffffffde",
            INIT_05 => X"0000003500000008fffffff4fffffffd0000000efffffff10000000700000024",
            INIT_06 => X"0000000afffffff4fffffff2fffffffdfffffff600000008fffffff200000000",
            INIT_07 => X"ffffffe90000000100000000000000060000000efffffff6ffffffde00000003",
            INIT_08 => X"0000002a0000004a0000000f0000000b0000001c00000010000000130000000f",
            INIT_09 => X"ffffffe3fffffff7ffffffef00000028000000170000000b0000001500000028",
            INIT_0A => X"ffffffe0fffffffb0000000dfffffff50000000a00000005ffffffd7fffffff2",
            INIT_0B => X"00000001ffffffdc0000003ffffffff80000001200000000ffffffcf00000001",
            INIT_0C => X"ffffffbcffffffdcffffffe7ffffffeffffffffa0000000bfffffffe00000022",
            INIT_0D => X"00000001ffffffe100000011fffffffffffffffd00000013ffffffb5ffffffc7",
            INIT_0E => X"00000003000000190000001e0000001300000048fffffffeffffffd800000019",
            INIT_0F => X"00000001fffffff4fffffff6fffffff1fffffff3fffffff4fffffffe00000011",
            INIT_10 => X"000000190000002500000020fffffff10000003a0000001a0000001f00000004",
            INIT_11 => X"fffffffaffffffe100000013ffffffdbfffffffbfffffff8000000020000001b",
            INIT_12 => X"0000001effffffeb00000001ffffffe9fffffff1fffffff5fffffff7ffffffdd",
            INIT_13 => X"ffffffed0000000100000019fffffff6ffffffd7fffffff5fffffffb00000010",
            INIT_14 => X"0000000a00000015000000080000000300000014ffffffebffffffee0000000a",
            INIT_15 => X"00000008fffffffeffffffea00000001ffffffeffffffff0ffffffe700000000",
            INIT_16 => X"00000008fffffff5ffffffed000000050000000a000000020000000000000002",
            INIT_17 => X"000000040000000dfffffff40000000bffffffe8ffffffedffffffebfffffffd",
            INIT_18 => X"00000007fffffff6fffffffd00000002fffffffd0000000200000011fffffff3",
            INIT_19 => X"fffffffcfffffff8fffffffe000000020000000a0000000cfffffff600000015",
            INIT_1A => X"000000070000000b00000003ffffffff00000005ffffffe60000000bfffffffe",
            INIT_1B => X"0000000700000006ffffffe5fffffff1fffffff4fffffff400000000ffffffff",
            INIT_1C => X"00000001fffffff6fffffffbfffffff8ffffffeafffffffc00000001ffffffeb",
            INIT_1D => X"fffffff2fffffff5ffffffe7fffffff0ffffffef0000000500000009fffffff1",
            INIT_1E => X"ffffffe8ffffffe70000000000000009ffffffebfffffff10000000cffffffed",
            INIT_1F => X"ffffffee0000000a000000010000000900000005ffffffe7fffffff9ffffffe5",
            INIT_20 => X"fffffff50000000ffffffffdfffffff90000000affffffeefffffff9fffffffd",
            INIT_21 => X"fffffff1fffffffcffffffebffffffecfffffffd0000000000000000fffffff9",
            INIT_22 => X"fffffff400000009ffffffeffffffffffffffffa000000090000000bffffffe5",
            INIT_23 => X"fffffff5ffffffe6ffffffe600000000fffffffcfffffffe00000002fffffff5",
            INIT_24 => X"fffffff0000000020000000400000004fffffff10000000000000001ffffffe9",
            INIT_25 => X"00000001fffffff9fffffff1fffffff10000000f0000000f0000000700000004",
            INIT_26 => X"00000007fffffff1000000000000000b00000000fffffff5fffffff3fffffffc",
            INIT_27 => X"ffffffeafffffff900000002ffffffeb000000010000000b00000003fffffffc",
            INIT_28 => X"0000000000000002ffffffec000000080000000dfffffff5ffffffee00000009",
            INIT_29 => X"fffffff3fffffffffffffff2fffffffc000000070000000f0000000fffffffec",
            INIT_2A => X"ffffffec0000000bfffffff9fffffff2fffffff6ffffffe3fffffffefffffff6",
            INIT_2B => X"000000050000000effffffeb00000000fffffff0ffffffe3ffffffedfffffff8",
            INIT_2C => X"0000000d00000000ffffffec0000000effffffeefffffff60000000d00000007",
            INIT_2D => X"fffffff000000007ffffffedfffffff4fffffff8ffffffef00000004ffffffff",
            INIT_2E => X"00000005ffffffee00000007fffffff9ffffffeafffffff00000000000000004",
            INIT_2F => X"0000000b00000007ffffffe400000004fffffff2ffffffe70000000200000000",
            INIT_30 => X"fffffff4ffffffdeffffffdfffffffe60000000300000000ffffffe1ffffffed",
            INIT_31 => X"fffffffdfffffff3fffffff60000001300000006fffffff8ffffffefffffffe0",
            INIT_32 => X"fffffff8fffffffa00000001fffffff3ffffffe9fffffff000000000fffffff6",
            INIT_33 => X"fffffffdffffffe600000007fffffff4ffffffe700000005ffffffecffffffeb",
            INIT_34 => X"0000000bffffffecffffffffffffffe30000000500000013fffffff200000007",
            INIT_35 => X"ffffffe7fffffffbfffffffcffffffe5fffffff300000005fffffff400000010",
            INIT_36 => X"fffffff4fffffffd00000006ffffffebfffffffefffffff2fffffff500000000",
            INIT_37 => X"00000005ffffffe80000000f00000006ffffffecfffffff9fffffffdfffffff4",
            INIT_38 => X"00000006fffffffdfffffffe00000014ffffffed00000012fffffffdfffffff6",
            INIT_39 => X"000000030000000a0000000300000009ffffffebfffffffd00000004ffffffef",
            INIT_3A => X"000000110000000400000005fffffffdfffffff7ffffffed00000000ffffffff",
            INIT_3B => X"fffffff7ffffffefffffffecffffffeb00000000ffffffe90000000500000001",
            INIT_3C => X"fffffffc00000003fffffff3ffffffeefffffff2fffffff700000009ffffffec",
            INIT_3D => X"00000002ffffffe4ffffffe9ffffffeefffffff4fffffff00000000600000009",
            INIT_3E => X"ffffffe8fffffff4fffffff40000000b00000009ffffffe2ffffffefffffffe4",
            INIT_3F => X"ffffffeafffffffeffffffecfffffffa0000000200000002fffffff5fffffffe",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE15;


    MEM_IWGHT_LAYER1_INSTANCE16 : if BRAM_NAME = "iwght_layer1_instance16" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffecffffffe7fffffff5fffffff1fffffff600000005fffffff9fffffff3",
            INIT_01 => X"0000000b00000000fffffffe0000000000000000ffffffe7ffffffef00000007",
            INIT_02 => X"0000000800000008fffffffeffffffedfffffff6fffffff00000000600000003",
            INIT_03 => X"00000005ffffffe3fffffffcfffffffc00000005000000000000000500000008",
            INIT_04 => X"ffffffe9ffffffea0000000bfffffff9ffffffeb00000000fffffff7fffffff5",
            INIT_05 => X"00000005fffffffa0000000f0000000800000003ffffffe9fffffffc0000000e",
            INIT_06 => X"0000000c0000000400000002000000040000000b0000000f0000000800000009",
            INIT_07 => X"0000000affffffe9fffffffffffffff60000000affffffecfffffffdffffffe9",
            INIT_08 => X"fffffffaffffffeb00000006000000080000000000000006fffffff2fffffffe",
            INIT_09 => X"fffffffcfffffff7fffffff300000001fffffff800000000fffffff60000000e",
            INIT_0A => X"ffffffed00000000fffffff1fffffffefffffff60000000c000000120000000e",
            INIT_0B => X"00000008ffffffedffffffeafffffffdfffffff400000006fffffff800000004",
            INIT_0C => X"fffffffb00000005fffffff60000000a00000005fffffffcfffffff7fffffffc",
            INIT_0D => X"fffffff9fffffffcfffffff9ffffffea0000000dfffffffaffffffef00000013",
            INIT_0E => X"ffffffff0000000affffffec00000002ffffffe50000000affffffe9fffffff1",
            INIT_0F => X"00000007fffffff400000002ffffffeffffffff200000003fffffff5fffffff0",
            INIT_10 => X"fffffffbffffffeffffffff2ffffffebffffffecfffffff200000005fffffff9",
            INIT_11 => X"00000006ffffffed00000000fffffff1fffffff6fffffffe00000000ffffffec",
            INIT_12 => X"fffffffafffffff9ffffffe7fffffffaffffffff000000040000000b00000005",
            INIT_13 => X"ffffffebfffffffaffffffe60000000ffffffff60000000a00000009fffffff4",
            INIT_14 => X"ffffffeefffffff8ffffffe9ffffffeb00000003fffffff2ffffffeb0000000c",
            INIT_15 => X"fffffff5ffffffeafffffff0000000000000000ffffffff9fffffff300000004",
            INIT_16 => X"ffffffeaffffffec0000001000000005ffffffe9fffffffcffffffe4fffffff8",
            INIT_17 => X"fffffff500000007fffffffbffffffeaffffffeefffffff5fffffffafffffff1",
            INIT_18 => X"fffffff5ffffffe5ffffffeefffffffafffffff9fffffff500000009ffffffef",
            INIT_19 => X"fffffffaffffffec00000003fffffff10000000e0000000200000003ffffffeb",
            INIT_1A => X"ffffffeeffffffeefffffff3fffffffa00000000fffffff500000005fffffffa",
            INIT_1B => X"fffffff7ffffffee0000000dfffffff9fffffffffffffffeffffffff00000006",
            INIT_1C => X"ffffffedfffffffafffffff700000008ffffffe9000000110000000800000000",
            INIT_1D => X"00000016fffffff6ffffffeeffffffdc0000001e0000002d0000000200000000",
            INIT_1E => X"fffffff40000002600000032000000050000002e00000022000000000000000c",
            INIT_1F => X"ffffffc9fffffff2ffffffd4ffffffe9fffffffdfffffff90000003100000035",
            INIT_20 => X"0000003effffffd9fffffffb0000001effffffb3ffffffa700000012ffffffa9",
            INIT_21 => X"fffffff20000000b0000000b0000000a0000000a00000038fffffffc0000000b",
            INIT_22 => X"000000220000002affffffe2ffffffe8ffffffe9000000170000002900000016",
            INIT_23 => X"ffffffe1ffffffb7ffffffecffffffe4ffffffea00000003fffffffa0000000f",
            INIT_24 => X"0000002d000000150000003afffffff300000010ffffffdf00000018ffffffff",
            INIT_25 => X"0000000f00000003fffffff0ffffffe100000007fffffff20000001a00000035",
            INIT_26 => X"0000001600000026fffffffcffffffe900000022ffffffd50000000d0000000e",
            INIT_27 => X"ffffffe4ffffffbeffffffd3000000010000002e000000040000002afffffff8",
            INIT_28 => X"ffffffe0000000180000000e00000026fffffffb0000000cfffffff700000013",
            INIT_29 => X"fffffffdffffffddffffffea0000000100000006ffffffc900000012fffffff5",
            INIT_2A => X"0000001300000000ffffffdc0000001300000008000000150000001800000007",
            INIT_2B => X"0000000c00000038fffffff500000015fffffffa00000006ffffffffffffffd6",
            INIT_2C => X"ffffffecffffffe7fffffff3fffffffcfffffffe00000018ffffffff00000004",
            INIT_2D => X"0000002000000005ffffffd10000002afffffff1ffffffe40000001500000003",
            INIT_2E => X"0000000efffffff4ffffffd9ffffffd2ffffffbd00000014fffffff2ffffffc6",
            INIT_2F => X"000000000000001affffffe9000000020000002300000001fffffffeffffffcb",
            INIT_30 => X"0000003ffffffffc0000000a00000012fffffff7ffffffc6000000050000000c",
            INIT_31 => X"000000090000001d0000001a0000002e00000016ffffffe5ffffffdcffffffce",
            INIT_32 => X"fffffff00000002a0000001bffffffe3fffffff10000000dfffffff90000000b",
            INIT_33 => X"0000000a0000002d00000031000000190000001cffffffed0000001300000000",
            INIT_34 => X"0000002600000018fffffff70000000effffffec000000030000000d00000005",
            INIT_35 => X"00000034fffffffc0000001c0000000cfffffffdffffffff000000170000000a",
            INIT_36 => X"ffffffeefffffff4ffffffeffffffffc0000000800000006ffffffe600000014",
            INIT_37 => X"ffffffe4ffffffaafffffff4ffffffdbffffffe90000001e0000002d00000016",
            INIT_38 => X"00000005ffffffeb0000000dfffffffe0000001300000003fffffff2ffffffd3",
            INIT_39 => X"0000003500000008fffffff900000018ffffffe6fffffff6ffffffe3fffffff8",
            INIT_3A => X"0000001000000017fffffff10000001d0000001f00000019fffffffffffffff9",
            INIT_3B => X"fffffff8ffffffaffffffff8fffffff8ffffffed0000001dffffffe90000000d",
            INIT_3C => X"0000000000000006fffffff8ffffffbfffffffcfffffffdaffffffcdfffffff0",
            INIT_3D => X"00000003ffffffcfffffffefffffffff000000090000002b0000000dffffffeb",
            INIT_3E => X"000000010000000c0000000800000015ffffffda00000000ffffffe8fffffff9",
            INIT_3F => X"0000000700000001ffffffe100000017fffffff30000000e0000001cffffffd7",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE16;


    MEM_IWGHT_LAYER1_INSTANCE17 : if BRAM_NAME = "iwght_layer1_instance17" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff40000000cffffffef0000000d00000007fffffff9fffffffe0000000c",
            INIT_01 => X"ffffffe1ffffffedfffffffeffffffdcffffffe4ffffffe3000000020000000e",
            INIT_02 => X"ffffffedfffffff7ffffffe8ffffffdf00000002ffffffeffffffff00000000a",
            INIT_03 => X"00000009fffffff9fffffffdffffffe900000004fffffff9ffffffee0000000d",
            INIT_04 => X"fffffff5fffffff0fffffff4ffffffe4ffffffebffffffd4ffffffedfffffff7",
            INIT_05 => X"fffffff90000000fffffffed0000000000000003fffffffefffffffa0000000c",
            INIT_06 => X"00000002ffffffedffffffe90000000100000000fffffff40000000400000001",
            INIT_07 => X"fffffff7fffffff200000000ffffffebffffffeefffffffbffffffe500000003",
            INIT_08 => X"fffffffd00000007ffffffe9fffffff400000006ffffffebfffffff000000002",
            INIT_09 => X"00000008ffffffe9ffffffecfffffffdffffffeb0000000a00000000fffffff6",
            INIT_0A => X"0000000dffffffe8fffffff800000007fffffff20000000300000009fffffff1",
            INIT_0B => X"fffffff3fffffff1fffffffe0000000dfffffff5fffffff500000016ffffffff",
            INIT_0C => X"fffffff8ffffffe900000013000000120000000000000004ffffffe8ffffffea",
            INIT_0D => X"fffffff6ffffffea0000000f0000000600000005ffffffe9fffffffdffffffe6",
            INIT_0E => X"fffffff1ffffffe400000005fffffff1fffffffefffffffeffffffedffffffe4",
            INIT_0F => X"000000110000000b0000000afffffff70000000100000000ffffffe800000002",
            INIT_10 => X"ffffffeefffffffdffffffe5fffffff4ffffffebfffffff3ffffffe9ffffffee",
            INIT_11 => X"fffffff8000000000000000cfffffff9fffffff7ffffffed00000003fffffff9",
            INIT_12 => X"00000020000000080000000cfffffffefffffff7fffffffb0000001000000016",
            INIT_13 => X"00000001fffffffd00000000000000110000001400000019fffffffd00000000",
            INIT_14 => X"fffffffafffffff9fffffffd00000011fffffff50000000500000004fffffff6",
            INIT_15 => X"ffffffe6fffffff1ffffffeb00000000ffffffe80000000000000002fffffff6",
            INIT_16 => X"ffffffefffffffefffffffecffffffe000000002fffffff7ffffffe8ffffffff",
            INIT_17 => X"00000000ffffffe0fffffff5ffffffe3ffffffec00000000fffffff4ffffffe0",
            INIT_18 => X"ffffffe6ffffffe00000000800000002fffffffdfffffff2ffffffebfffffff7",
            INIT_19 => X"0000000bfffffff300000020fffffffd0000000cfffffff90000000ffffffff7",
            INIT_1A => X"00000008ffffffed0000000600000000000000000000000900000012fffffffa",
            INIT_1B => X"0000000c00000000ffffffe6ffffffe8ffffffe9ffffffdcfffffff4fffffff1",
            INIT_1C => X"ffffffebffffffeafffffff0ffffffe6ffffffd9fffffffc0000000bffffffdb",
            INIT_1D => X"fffffffc0000000f0000001200000011fffffffafffffff3ffffffedffffffed",
            INIT_1E => X"ffffffe3fffffff8fffffff00000000800000004ffffffe60000000effffffe5",
            INIT_1F => X"fffffff7fffffff400000002ffffffe8fffffff0fffffffefffffff8fffffffa",
            INIT_20 => X"fffffff100000000fffffff6fffffff5ffffffec0000000300000001fffffffa",
            INIT_21 => X"000000070000000afffffff0fffffff1ffffffea00000009ffffffffffffffea",
            INIT_22 => X"ffffffe3fffffffefffffff9fffffff2fffffffa00000008ffffffebfffffff0",
            INIT_23 => X"ffffffffffffffe9ffffffebfffffff9fffffffc0000000efffffff9fffffffa",
            INIT_24 => X"0000001a000000180000000e0000000700000004ffffffee0000001a00000019",
            INIT_25 => X"000000570000003a000000620000004a000000420000003c0000001c00000005",
            INIT_26 => X"ffffffaeffffffb6ffffffc0fffffff7ffffffef00000000ffffffc600000006",
            INIT_27 => X"fffffff4ffffffe500000012fffffff5ffffffe5ffffff74ffffffb8ffffff83",
            INIT_28 => X"ffffffdcfffffffd00000006fffffffd000000630000000f0000001b0000001c",
            INIT_29 => X"fffffffa000000180000001affffffbeffffff63ffffffebffffffc4ffffffbc",
            INIT_2A => X"0000000afffffff600000054000000340000002affffffedffffffe000000004",
            INIT_2B => X"0000000900000000ffffffe500000000000000000000000800000012fffffff4",
            INIT_2C => X"000000070000002d0000001600000006fffffff4fffffffcfffffffa00000011",
            INIT_2D => X"000000090000002c000000140000003a00000019000000300000001400000016",
            INIT_2E => X"00000007ffffffb0ffffffe0fffffff5ffffffc3fffffff1ffffffe5ffffffbb",
            INIT_2F => X"ffffffff0000002a00000047000000020000002400000025fffffff1fffffff5",
            INIT_30 => X"ffffff84ffffffc9ffffffb5fffffff5fffffffdffffff6effffff9e00000023",
            INIT_31 => X"000000040000000effffffeeffffffddffffffdfffffffc1fffffffeffffffcb",
            INIT_32 => X"ffffffdc000000230000000f00000065000000310000001dfffffff9ffffffed",
            INIT_33 => X"ffffffd600000012fffffff9fffffffbfffffffdfffffff90000001f00000031",
            INIT_34 => X"fffffffc000000310000001f0000000affffffa8ffffffe4fffffff0ffffffd7",
            INIT_35 => X"000000220000001600000003ffffffe7ffffffde00000014ffffffd6ffffffe1",
            INIT_36 => X"00000002fffffff6ffffffed000000070000002c00000014000000490000000a",
            INIT_37 => X"000000010000001700000021000000220000000b0000000f00000028ffffffea",
            INIT_38 => X"ffffffe800000016ffffffe10000000effffffda0000000200000015fffffffc",
            INIT_39 => X"00000002fffffff9000000150000000e0000001bfffffffb00000018fffffff6",
            INIT_3A => X"ffffffdcfffffffdfffffff90000000e00000013000000130000000900000002",
            INIT_3B => X"fffffffd000000000000001d00000001fffffff6fffffff8fffffff6ffffffea",
            INIT_3C => X"0000000cffffffe800000009fffffffbfffffff80000000a00000000fffffff1",
            INIT_3D => X"000000210000000000000009fffffff3ffffffee0000000ffffffffd0000000f",
            INIT_3E => X"ffffffc7ffffffcdffffffebffffffe4ffffffe60000001efffffff300000001",
            INIT_3F => X"ffffffb5fffffff5ffffff9bffffffd6ffffffb8ffffffffffffffb8ffffffe6",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE17;


    MEM_IWGHT_LAYER1_INSTANCE18 : if BRAM_NAME = "iwght_layer1_instance18" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000c000000070000002a0000002000000032000000240000002fffffffa2",
            INIT_01 => X"ffffffdefffffffbfffffffaffffffecfffffff90000002effffffe9fffffff4",
            INIT_02 => X"fffffff80000000effffffeafffffffefffffff30000000ffffffffffffffff7",
            INIT_03 => X"ffffffe40000001dffffffd0fffffff00000000e0000000f0000000cfffffff0",
            INIT_04 => X"ffffffd3ffffffd2ffffffe00000000e000000190000003bfffffffafffffff3",
            INIT_05 => X"0000000ffffffff1000000140000000b00000013ffffffcfffffffc0ffffffbb",
            INIT_06 => X"0000000e0000001a0000000b0000000900000017ffffffe6fffffff900000001",
            INIT_07 => X"0000001b0000001afffffffdfffffffeffffffff00000005fffffff6ffffffe5",
            INIT_08 => X"000000100000000e00000008fffffffc000000040000001400000018fffffffc",
            INIT_09 => X"ffffffefffffffeffffffff700000017fffffffd000000210000001200000002",
            INIT_0A => X"ffffffc4ffffffd2ffffffeeffffffccffffffedfffffff90000000cffffffd0",
            INIT_0B => X"000000190000002f00000007000000000000001affffffcbffffffd500000003",
            INIT_0C => X"ffffffe5ffffffe0ffffff96fffffff3fffffff0000000210000003b0000002c",
            INIT_0D => X"ffffffc4fffffff2ffffffcaffffffe6ffffffeaffffffd9ffffffcfffffff94",
            INIT_0E => X"00000000000000160000003100000040ffffffdffffffff500000009ffffffe9",
            INIT_0F => X"ffffffdbffffffeeffffffedffffffe20000001dffffffee0000000900000013",
            INIT_10 => X"0000001ffffffffc0000000f0000002900000013fffffff600000005ffffffd3",
            INIT_11 => X"fffffffffffffff9ffffffea000000050000004d0000000f000000320000004d",
            INIT_12 => X"ffffffe9ffffffdafffffff40000000afffffff5ffffffea00000002fffffff6",
            INIT_13 => X"ffffffe0ffffffd700000024ffffffff0000002100000025ffffffe3fffffff6",
            INIT_14 => X"0000001dfffffffeffffffecffffffeb00000000ffffffe100000000fffffff5",
            INIT_15 => X"fffffff3fffffffbffffffdffffffff3fffffffefffffffbfffffff200000002",
            INIT_16 => X"ffffffdeffffffe7ffffffde0000001700000018000000150000002900000016",
            INIT_17 => X"ffffffef0000001100000001fffffff900000022000000370000000500000015",
            INIT_18 => X"000000010000000800000012fffffff40000000bfffffff6ffffffe4ffffffd8",
            INIT_19 => X"000000120000000d000000010000001900000019ffffffe9ffffffe0ffffffda",
            INIT_1A => X"00000006fffffff400000026000000280000002e00000026000000390000005f",
            INIT_1B => X"0000000800000026fffffffc00000012000000110000000b0000000900000024",
            INIT_1C => X"fffffff0fffffff8ffffffecffffffb4ffffffd0fffffff6ffffffe8ffffffeb",
            INIT_1D => X"ffffffe10000000effffffe5ffffffee0000000000000019ffffffeeffffffea",
            INIT_1E => X"ffffffbfffffffd8ffffffe7ffffffe70000002e00000022ffffffe5fffffffd",
            INIT_1F => X"ffffffdeffffffeffffffff60000002a0000001cffffffd8ffffffe8ffffffe6",
            INIT_20 => X"ffffffeafffffffe0000004200000040fffffff8ffffffd8ffffffdcffffffc1",
            INIT_21 => X"00000040fffffff7ffffffeaffffffd300000004ffffffeefffffff2ffffffd1",
            INIT_22 => X"fffffff6fffffff6fffffffefffffffdffffffe5000000170000000a00000019",
            INIT_23 => X"0000001e00000000ffffffd2fffffffe0000004cffffffbfffffffdbfffffffa",
            INIT_24 => X"00000001000000080000000dfffffff0fffffff1ffffffe50000000500000017",
            INIT_25 => X"000000050000000500000022000000130000000effffffff0000000a00000005",
            INIT_26 => X"ffffffeefffffffaffffffcdffffffd8ffffffddfffffff3fffffff800000007",
            INIT_27 => X"0000003000000021000000190000000600000004fffffff4ffffffeb00000009",
            INIT_28 => X"fffffff6fffffffcfffffff3ffffffde000000010000001f0000000f00000008",
            INIT_29 => X"ffffffeeffffffdb00000012ffffffe7fffffff6ffffffe60000000dfffffff4",
            INIT_2A => X"ffffffe3000000180000000cfffffff4fffffff4ffffffe5ffffffb0ffffffd4",
            INIT_2B => X"00000012fffffff9000000180000002f00000011fffffffb0000001700000002",
            INIT_2C => X"ffffffe8ffffffe30000000afffffff6ffffffdfffffffed00000001fffffff7",
            INIT_2D => X"ffffff78ffffffb9ffffff9affffff9bffffffebfffffff60000001affffffe8",
            INIT_2E => X"fffffffc00000006ffffffe0ffffffea0000001900000018ffffffc6ffffff87",
            INIT_2F => X"ffffffc10000000affffffdcffffffb3000000020000000e0000001b00000026",
            INIT_30 => X"0000002700000000ffffffee0000000affffffd6ffffffe900000011ffffffcc",
            INIT_31 => X"ffffffff00000022000000290000000a0000002c0000002bffffffef00000014",
            INIT_32 => X"00000008ffffffeffffffff6000000170000000cfffffff60000002700000039",
            INIT_33 => X"0000000cfffffff3fffffff2fffffffdffffffe0fffffff5fffffff9ffffffeb",
            INIT_34 => X"000000190000001a00000026000000380000001bfffffff40000000100000020",
            INIT_35 => X"fffffff0ffffffcaffffffeeffffffc9ffffffb8fffffff6ffffffe4fffffff4",
            INIT_36 => X"0000000cffffffe9fffffff7ffffffff00000005000000110000000100000003",
            INIT_37 => X"ffffffc7ffffffc3ffffffdcfffffffd0000000900000001fffffffefffffff9",
            INIT_38 => X"ffffffd00000001effffffed0000000b0000000a0000000efffffff1ffffffda",
            INIT_39 => X"00000005ffffffe1fffffff4fffffffaffffffe3ffffffd80000002fffffffdd",
            INIT_3A => X"00000028000000220000000dffffffc80000001000000020fffffff1fffffffd",
            INIT_3B => X"fffffff200000003000000020000000300000006fffffffffffffffaffffffe3",
            INIT_3C => X"fffffff0fffffff00000001200000013fffffff20000000e0000003fffffffe9",
            INIT_3D => X"fffffffa0000000e00000019fffffff10000001b0000000f0000000dfffffff5",
            INIT_3E => X"ffffffb000000004ffffffbbffffffe0ffffffb4ffffffc4ffffffe2ffffffcc",
            INIT_3F => X"00000002ffffffe4000000110000000000000011000000140000001effffffc2",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE18;


    MEM_IWGHT_LAYER1_INSTANCE19 : if BRAM_NAME = "iwght_layer1_instance19" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffedffffffda000000070000004c0000004a0000002cffffffcefffffffa",
            INIT_01 => X"0000000d0000001700000000ffffffe7fffffffbffffffdaffffffbbfffffffc",
            INIT_02 => X"000000220000001cfffffff80000000400000019000000230000000f0000000b",
            INIT_03 => X"fffffff9fffffff70000000700000000fffffff2fffffff9fffffff800000004",
            INIT_04 => X"fffffff7000000000000001a0000000800000007000000000000000b00000019",
            INIT_05 => X"00000020ffffffef0000002200000000fffffff50000000700000005fffffffc",
            INIT_06 => X"0000000b0000001900000020000000080000000d00000013fffffffdfffffff7",
            INIT_07 => X"00000021fffffff10000003000000003ffffffebffffffd900000010fffffff3",
            INIT_08 => X"00000017ffffffe1fffffff5ffffffdb0000000d000000110000000000000042",
            INIT_09 => X"ffffffef0000000e000000000000002900000026fffffffa0000000effffffed",
            INIT_0A => X"00000000ffffffe8ffffffccffffffebfffffffcffffffe3fffffff600000026",
            INIT_0B => X"00000019ffffffe6000000000000001d00000005000000210000000600000009",
            INIT_0C => X"ffffffcc00000021fffffff4ffffffe80000003afffffffbffffffd900000008",
            INIT_0D => X"ffffffe6ffffffffffffffecfffffffb00000029ffffffff0000002c00000007",
            INIT_0E => X"000000210000000c00000006000000140000000effffffec0000000e00000001",
            INIT_0F => X"ffffffce0000002300000010000000020000001b0000000e000000320000001b",
            INIT_10 => X"fffffffa000000010000000e00000010fffffffcffffffe3fffffff5ffffffed",
            INIT_11 => X"0000000e0000003200000016000000360000000e00000015fffffffdfffffff0",
            INIT_12 => X"0000000c00000011ffffffdd0000001a000000110000002f0000002000000020",
            INIT_13 => X"0000003b000000180000000700000015ffffffe8000000420000001c00000015",
            INIT_14 => X"0000001000000015ffffffda0000001c0000000bffffffeaffffffd600000007",
            INIT_15 => X"ffffffebffffffd8ffffffcd0000002700000008ffffffe8000000290000000f",
            INIT_16 => X"fffffff9ffffffeaffffffe7ffffffc7ffffffb8ffffffeeffffffe4ffffffe7",
            INIT_17 => X"00000022fffffffcfffffff2fffffffeffffffb5ffffffb9ffffffafffffffd5",
            INIT_18 => X"00000015fffffff900000011ffffffe5fffffff100000012fffffff50000003a",
            INIT_19 => X"00000001ffffffc80000001100000009ffffffe800000002fffffffbffffffec",
            INIT_1A => X"0000000600000002fffffff700000009000000180000000bffffffee0000003e",
            INIT_1B => X"0000001afffffffe000000090000001a0000000dffffffe90000000d0000000b",
            INIT_1C => X"fffffff1ffffffb70000000effffffa8ffffffe5000000130000002900000003",
            INIT_1D => X"ffffffc9fffffffbfffffff4ffffffeaffffffcfffffffe2ffffffc0ffffffe7",
            INIT_1E => X"ffffffd5fffffffaffffffdeffffffbbffffffc2fffffffa0000000ffffffff2",
            INIT_1F => X"ffffffbfffffffdfffffffec00000012fffffffdffffffe3ffffffccffffffd8",
            INIT_20 => X"fffffff0ffffffc9ffffffa5ffffff97fffffffbffffff9affffffc0fffffff0",
            INIT_21 => X"ffffffbfffffffd7fffffff200000001ffffffeaffffffea0000001e00000000",
            INIT_22 => X"ffffff82ffffffcaffffffa9ffffffabffffffbbffffffe7ffffffeaffffffcc",
            INIT_23 => X"ffffffd9ffffffe1ffffffabfffffff00000001a00000000ffffffd1ffffffd7",
            INIT_24 => X"0000000000000000ffffffe100000024fffffffcffffffffffffffe6fffffffd",
            INIT_25 => X"00000014000000020000001b000000180000000e0000001cffffffcfffffffdd",
            INIT_26 => X"0000001700000030000000450000000fffffffd7ffffffdf0000001300000003",
            INIT_27 => X"00000033000000330000000effffffedffffffe3fffffffa0000003e00000036",
            INIT_28 => X"ffffffefffffffe2ffffffedffffffedffffffe0000000140000003500000011",
            INIT_29 => X"ffffffef0000000e00000001ffffffeb000000070000000bffffffe900000002",
            INIT_2A => X"ffffffe5ffffffcaffffffdd00000015ffffffe3ffffffe20000001bfffffff7",
            INIT_2B => X"0000001a00000031000000160000003200000024ffffffec0000001d00000008",
            INIT_2C => X"00000005000000060000001600000000ffffffe7000000130000002bfffffff3",
            INIT_2D => X"000000430000002100000000000000390000001500000000fffffff0fffffff3",
            INIT_2E => X"ffffffb0ffffffeeffffffdeffffffd2ffffffdb000000380000001afffffff8",
            INIT_2F => X"000000300000002c0000000000000008ffffff9effffffb60000002fffffffd1",
            INIT_30 => X"ffffffc3ffffff95ffffff97000000110000000d0000000c0000003100000004",
            INIT_31 => X"0000001500000008ffffffcd0000000400000022ffffff76ffffff90ffffffc5",
            INIT_32 => X"fffffff4ffffffcfffffffe3000000040000000d000000310000001500000032",
            INIT_33 => X"0000001ffffffff4fffffffb0000001a0000002b00000011000000440000000c",
            INIT_34 => X"0000000000000001fffffff300000002ffffffe1ffffffef0000001300000013",
            INIT_35 => X"ffffffeaffffffa7ffffffbcffffffd0ffffff9affffffceffffffe600000000",
            INIT_36 => X"00000003ffffffde0000000bffffffcaffffffea00000004fffffff6ffffffe0",
            INIT_37 => X"00000011ffffffe4fffffff1fffffffbffffffeeffffffe1fffffffe00000002",
            INIT_38 => X"00000004ffffffc9ffffffd8fffffff1fffffffa00000005ffffffe200000016",
            INIT_39 => X"0000002e0000002d0000000fffffffe5ffffffdaffffffd6ffffffe5fffffff0",
            INIT_3A => X"ffffffdd00000014fffffffdfffffffc00000025000000200000001c0000001f",
            INIT_3B => X"fffffffb00000014fffffffb0000002200000005ffffffec0000000effffffca",
            INIT_3C => X"ffffffe30000000e00000012000000180000000f00000029ffffffdf00000017",
            INIT_3D => X"ffffffeeffffffe9fffffff7ffffffdf00000000fffffffaffffffe400000019",
            INIT_3E => X"0000001100000002ffffffffffffffedfffffff3ffffffe0ffffffed0000000c",
            INIT_3F => X"fffffff9fffffff10000001cffffffcbffffffe9000000130000001500000024",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE19;


    MEM_IWGHT_LAYER1_INSTANCE20 : if BRAM_NAME = "iwght_layer1_instance20" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001c0000001700000037fffffff9000000050000001a0000000c00000004",
            INIT_01 => X"fffffff80000002e00000009ffffffe3000000040000000a0000001f00000026",
            INIT_02 => X"ffffffccfffffff1fffffffe0000000900000004fffffff90000001e00000001",
            INIT_03 => X"0000002a00000019fffffff20000000affffffd6ffffffdfffffffc7ffffffec",
            INIT_04 => X"ffffffeaffffffda0000000700000024000000080000001c0000002100000021",
            INIT_05 => X"0000000afffffffdffffffe100000000ffffffe6ffffffda00000010ffffffd6",
            INIT_06 => X"fffffff3ffffffe1ffffffc4ffffffd6fffffffbffffffd7ffffffcaffffffe6",
            INIT_07 => X"0000000d0000001300000000000000190000000dffffffeafffffffeffffffda",
            INIT_08 => X"0000000400000004ffffffd10000002c00000004000000330000001700000038",
            INIT_09 => X"0000001c00000011000000120000001dfffffffb0000004700000000fffffff4",
            INIT_0A => X"0000001100000004000000110000001effffffecfffffffc0000002900000006",
            INIT_0B => X"00000015000000160000000e0000000d0000001900000011fffffff700000012",
            INIT_0C => X"fffffff1fffffff700000009fffffff2fffffffd0000000b00000004fffffff5",
            INIT_0D => X"00000009000000150000001b000000110000001a000000080000000cfffffff0",
            INIT_0E => X"ffffffdbffffffe500000021fffffffdfffffff500000018fffffff10000001e",
            INIT_0F => X"000000220000005b000000690000004c0000002d000000470000003d00000063",
            INIT_10 => X"00000004ffffffdcffffffbfffffffeeffffffbdffffffd9fffffffa00000011",
            INIT_11 => X"0000001c0000001600000005fffffff300000005fffffff6fffffff9ffffffde",
            INIT_12 => X"fffffff900000022fffffffefffffffb00000001000000240000003c00000014",
            INIT_13 => X"00000002000000140000000b000000110000000c000000280000002ffffffffa",
            INIT_14 => X"fffffff9000000000000000700000023fffffff2ffffffde0000001a00000001",
            INIT_15 => X"0000001400000014000000030000002100000041000000150000002600000011",
            INIT_16 => X"ffffffeffffffffafffffff00000000dffffffea0000000e0000001200000011",
            INIT_17 => X"0000001a00000027000000060000000fffffffed0000000000000006fffffff5",
            INIT_18 => X"0000001600000014fffffff30000000efffffff3fffffff000000008ffffffff",
            INIT_19 => X"ffffffddffffffebfffffff6ffffffceffffffd7fffffffe00000008fffffffe",
            INIT_1A => X"0000000c0000004700000034000000190000004bffffffffffffffc0ffffffc0",
            INIT_1B => X"ffffffda000000090000001ffffffff1fffffffc000000000000000700000020",
            INIT_1C => X"fffffffe0000003d000000240000002c00000026000000050000002dffffffea",
            INIT_1D => X"00000006000000000000000c0000003c000000050000004affffffe6fffffff5",
            INIT_1E => X"ffffffe7ffffffd4ffffffd1fffffffb00000000ffffffea0000001d00000032",
            INIT_1F => X"ffffffe8fffffffdfffffff6ffffffc30000001600000002ffffffd8fffffff3",
            INIT_20 => X"0000001f0000000d00000002ffffffecffffffd1fffffffa0000000b00000011",
            INIT_21 => X"fffffffa000000020000002400000000000000010000000a000000140000001b",
            INIT_22 => X"ffffffd9fffffffe000000370000001fffffffe4fffffff5ffffffdf0000001a",
            INIT_23 => X"0000001e00000006fffffffbfffffff7ffffffec000000110000000afffffffa",
            INIT_24 => X"ffffffcf0000001700000007fffffff2ffffffdf0000001f0000001cfffffff4",
            INIT_25 => X"ffffffceffffffddffffffc4ffffffa2ffffffe1ffffffc9ffffffe20000000f",
            INIT_26 => X"fffffff00000000400000002ffffffd5ffffffdffffffffaffffffc7ffffffca",
            INIT_27 => X"ffffffd700000000ffffffd6fffffff0ffffffd8fffffff2ffffffe600000012",
            INIT_28 => X"ffffff91ffffffeaffffffe8fffffff9ffffffecfffffffbffffffe9ffffffff",
            INIT_29 => X"ffffffff0000000300000012ffffffdaffffffc6ffffffbfffffffd7ffffff95",
            INIT_2A => X"0000000300000016000000160000000effffffe2ffffff9dffffffb9ffffffdd",
            INIT_2B => X"ffffffe500000013ffffffdffffffff2ffffffcdffffffedffffffbcffffffdf",
            INIT_2C => X"0000000cffffffff000000370000002a0000001b000000260000000c00000015",
            INIT_2D => X"fffffffaffffffffffffffffffffffe5ffffffec00000029fffffff800000024",
            INIT_2E => X"0000000dfffffff2000000050000000900000017fffffff2fffffff3fffffffc",
            INIT_2F => X"fffffffeffffffe8ffffffe90000001d000000010000000f00000009fffffffa",
            INIT_30 => X"ffffffc4ffffffa5fffffffeffffffebffffffef0000000c0000000a00000007",
            INIT_31 => X"fffffff2fffffffcffffffe8fffffffbffffffd9ffffffdffffffff3ffffffdc",
            INIT_32 => X"00000029000000070000000c000000190000001100000016ffffffffffffffe9",
            INIT_33 => X"00000024ffffffdbffffffd2ffffffeaffffffc6ffffffff0000001cffffffe2",
            INIT_34 => X"0000002000000033000000250000001400000000000000030000002900000010",
            INIT_35 => X"ffffffddfffffffd00000018ffffffecfffffff7ffffffff0000001e00000031",
            INIT_36 => X"ffffffe7ffffffc6ffffffd1fffffff4ffffffb900000001ffffffe9fffffffd",
            INIT_37 => X"00000011000000250000002e00000027ffffffdc00000017ffffffb2fffffff1",
            INIT_38 => X"ffffffb1ffffffd2ffffffe9000000040000001c0000002ffffffff9fffffff2",
            INIT_39 => X"0000000300000011000000170000000bffffffe400000013ffffffefffffffe8",
            INIT_3A => X"0000000c00000015000000190000000d0000001b000000020000001900000005",
            INIT_3B => X"ffffffeefffffff1ffffffdcffffffcdffffffaafffffff3ffffffe2ffffffee",
            INIT_3C => X"00000010fffffffcfffffff70000000500000002fffffff4fffffff1fffffff5",
            INIT_3D => X"ffffffe1ffffffe600000009ffffffe9ffffffe7000000010000000f0000000d",
            INIT_3E => X"0000002a0000002d00000005000000360000001a0000000fffffffe5fffffff2",
            INIT_3F => X"0000001500000017ffffffe5000000120000005f000000160000003600000011",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE20;


    MEM_IWGHT_LAYER1_INSTANCE21 : if BRAM_NAME = "iwght_layer1_instance21" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001e00000005000000250000002b000000140000000dffffffe6ffffffe8",
            INIT_01 => X"00000002ffffffacffffffb100000010fffffff900000001fffffff400000031",
            INIT_02 => X"ffffffcbffffffeafffffff6ffffffe7ffffffc90000001affffffe8ffffffd0",
            INIT_03 => X"fffffff5000000270000000c000000250000000bffffffeaffffffe4ffffffd1",
            INIT_04 => X"0000000d0000000a0000002c0000003a00000009000000360000000000000019",
            INIT_05 => X"fffffff6ffffffcdffffffeffffffff9ffffffa9ffffffd600000008ffffffde",
            INIT_06 => X"00000008ffffffdbffffffeaffffffeeffffffdeffffffccffffffbefffffff4",
            INIT_07 => X"00000013fffffffaffffffd600000011ffffffe3ffffffeeffffffe6fffffff1",
            INIT_08 => X"ffffffbbfffffff20000001dfffffff5fffffff4fffffff7ffffffdffffffff6",
            INIT_09 => X"fffffff7fffffff3ffffffeaffffffd1ffffffd0ffffffd3ffffffcafffffffb",
            INIT_0A => X"ffffffeb000000110000001c0000002000000011fffffffa0000000300000016",
            INIT_0B => X"ffffffdbffffffaafffffff2fffffffb0000002f0000000d0000001f00000059",
            INIT_0C => X"fffffff7ffffffdfffffffdc0000000200000002fffffffdffffffc7ffffffe6",
            INIT_0D => X"0000000200000023000000010000001100000007fffffff1000000000000000a",
            INIT_0E => X"ffffffbf00000016ffffffc5fffffff90000004800000003fffffff500000042",
            INIT_0F => X"0000000700000010ffffffecffffffeffffffff2ffffffe4ffffffd6fffffffa",
            INIT_10 => X"ffffffc7ffffffebfffffff5ffffffd1ffffffc0ffffffdf0000002400000011",
            INIT_11 => X"00000002fffffff0000000150000000cffffffed0000000bffffffe300000011",
            INIT_12 => X"fffffffe00000003fffffffefffffff100000021000000020000000100000010",
            INIT_13 => X"0000000400000023fffffffbffffffe600000007fffffffdfffffff9fffffff9",
            INIT_14 => X"fffffffbffffffecffffffe8ffffffeefffffffc0000001b00000020fffffffe",
            INIT_15 => X"ffffffee00000036000000130000000700000013ffffffe6ffffffff00000013",
            INIT_16 => X"0000002d0000000e0000000efffffff500000000fffffff200000018ffffffd7",
            INIT_17 => X"ffffffccffffffd90000002f00000014ffffffd40000002c00000034fffffff9",
            INIT_18 => X"0000002e00000006000000130000002f000000120000002000000037ffffffe9",
            INIT_19 => X"fffffffc000000250000002efffffff3fffffffbffffffed0000000400000006",
            INIT_1A => X"ffffffe700000004ffffffd1ffffffdcffffffc4000000070000000cfffffff9",
            INIT_1B => X"0000000dffffffd3ffffffe000000012000000200000001e0000000000000016",
            INIT_1C => X"0000001affffffd3ffffffbaffffffe900000020ffffffe0ffffffcefffffffd",
            INIT_1D => X"00000014ffffffeb00000033fffffff500000004fffffffaffffffe7ffffffe7",
            INIT_1E => X"fffffff000000004000000010000000a00000012000000070000001100000019",
            INIT_1F => X"fffffffc000000230000001900000013000000160000000cfffffffc0000000c",
            INIT_20 => X"00000010fffffff9ffffffdffffffff6ffffffebffffffe9fffffff6ffffffec",
            INIT_21 => X"ffffffb20000001d00000003fffffff600000015fffffff6fffffff400000003",
            INIT_22 => X"00000009fffffffa00000017ffffffebffffffedffffffdf0000001000000002",
            INIT_23 => X"0000000900000001000000280000001ffffffffe0000001800000037ffffffff",
            INIT_24 => X"00000009ffffffd4ffffffcfffffffd4ffffffd2fffffff80000000dffffffe9",
            INIT_25 => X"fffffffdfffffffe00000000000000000000004d00000024000000060000002c",
            INIT_26 => X"0000000f00000003fffffff40000001e00000034ffffffdd0000001000000023",
            INIT_27 => X"ffffffe10000000e00000000000000090000000900000012fffffff000000023",
            INIT_28 => X"00000003000000070000001a0000000cfffffff0fffffff20000002000000002",
            INIT_29 => X"0000000000000012000000020000002500000035fffffff30000002400000013",
            INIT_2A => X"ffffffae0000003100000036ffffffb30000001600000014ffffffaeffffffd9",
            INIT_2B => X"ffffffed0000000600000021fffffff40000001300000003000000460000000a",
            INIT_2C => X"fffffffbffffffc900000000fffffffcffffffe3ffffffdafffffff1fffffffa",
            INIT_2D => X"ffffffe8fffffff80000000900000000000000000000001dfffffff60000000b",
            INIT_2E => X"0000001500000019ffffffbbffffffdeffffffd100000015fffffff6fffffff7",
            INIT_2F => X"00000007000000040000003900000005ffffff9b0000000600000020ffffffc1",
            INIT_30 => X"00000000ffffffef000000390000002bfffffffa0000000b00000036ffffffdb",
            INIT_31 => X"00000012fffffffc0000000d0000002000000009fffffff20000001cfffffff5",
            INIT_32 => X"fffffffbffffffc20000005200000045000000190000004a0000004afffffffa",
            INIT_33 => X"ffffffda0000001d00000026ffffffdf0000002dfffffff4ffffffc600000016",
            INIT_34 => X"00000014ffffffceffffffffffffffe900000005000000390000001700000017",
            INIT_35 => X"fffffff20000002cffffffdaffffffe200000027000000170000000a00000005",
            INIT_36 => X"0000002cffffffdbffffffef00000037ffffffd4000000000000002affffffd2",
            INIT_37 => X"ffffffd0ffffffcf0000002fffffffd9000000000000003fffffffd1fffffff1",
            INIT_38 => X"00000018ffffffeeffffffe5fffffff50000002cffffffc9fffffff600000010",
            INIT_39 => X"000000020000002bffffffe8ffffffe10000002d0000000effffffcc00000006",
            INIT_3A => X"ffffffac000000030000001cffffffdc0000000200000030ffffffccffffffe2",
            INIT_3B => X"fffffff100000019000000070000001a0000001500000001000000310000003f",
            INIT_3C => X"ffffffdefffffff4000000150000000afffffffd0000000dffffffd40000000d",
            INIT_3D => X"0000004b00000023ffffffd000000033fffffff2ffffff9f00000001fffffffb",
            INIT_3E => X"fffffff8ffffffe9fffffff7fffffff3fffffffa0000003f0000000cffffffb6",
            INIT_3F => X"0000000ffffffffe0000001cffffffe900000012fffffff50000001400000005",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE21;


    MEM_IWGHT_LAYER1_INSTANCE22 : if BRAM_NAME = "iwght_layer1_instance22" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000bfffffff6ffffffcdffffffe3fffffff8fffffff30000001500000016",
            INIT_01 => X"fffffff50000002b0000001affffffefffffffe80000001cfffffffcffffffcb",
            INIT_02 => X"ffffffdcffffffcc0000000a00000050ffffffddffffffe900000023ffffffeb",
            INIT_03 => X"00000015fffffff6ffffffc10000002e00000000ffffffc80000003bffffffff",
            INIT_04 => X"fffffff100000005ffffffe800000001ffffffe4fffffff60000000200000014",
            INIT_05 => X"00000003ffffffedfffffffc0000002f000000270000000a00000023ffffffea",
            INIT_06 => X"ffffffd2ffffffc60000000dfffffff7fffffff0ffffffe9ffffffcaffffffe4",
            INIT_07 => X"ffffffc90000002000000016ffffffcdffffffcffffffff90000001600000033",
            INIT_08 => X"00000015ffffffaeffffffc7fffffff3ffffffeeffffffcb0000002dffffffbb",
            INIT_09 => X"ffffffe8fffffffb00000033fffffff3000000250000005fffffffc0ffffffc7",
            INIT_0A => X"0000000800000037ffffffd6fffffff3ffffffe7ffffffeffffffff600000010",
            INIT_0B => X"ffffffe8ffffffec0000000700000005ffffffea000000000000000dfffffff2",
            INIT_0C => X"0000001bffffffedffffffce00000011fffffff0ffffffc90000005200000011",
            INIT_0D => X"ffffffff00000004ffffffd3fffffffb0000001fffffffed0000001c0000000e",
            INIT_0E => X"00000015fffffff5fffffffc00000028ffffffd6ffffffc00000000effffffd4",
            INIT_0F => X"00000000ffffffeffffffffc0000000a000000010000000fffffffc1fffffffd",
            INIT_10 => X"ffffffdbffffffe10000002affffffebffffffedfffffffe0000000bffffffeb",
            INIT_11 => X"0000000b00000009ffffffe300000031ffffffd9ffffffbeffffffe9fffffff3",
            INIT_12 => X"00000026ffffffe900000002ffffffcdffffffe1ffffffe4ffffffceffffffe8",
            INIT_13 => X"0000000500000003ffffffed0000000a0000001f00000008000000130000004c",
            INIT_14 => X"00000031ffffffc6ffffffddffffffd2ffffffe0ffffffe00000000400000007",
            INIT_15 => X"0000000d0000002700000021fffffff7000000030000002bfffffffbfffffff3",
            INIT_16 => X"000000140000003d0000004b00000051000000430000000f0000002900000008",
            INIT_17 => X"00000008ffffffdd0000000b0000001200000009fffffff000000010fffffff9",
            INIT_18 => X"000000060000000500000008ffffffe5ffffffe1ffffffccffffffc7fffffffb",
            INIT_19 => X"fffffffcfffffff60000000a0000000300000001fffffff1000000210000000c",
            INIT_1A => X"ffffffed00000018fffffffefffffff6000000080000000bfffffff400000002",
            INIT_1B => X"0000000300000011fffffff90000001500000006fffffff50000000f00000017",
            INIT_1C => X"0000000200000022000000110000003e0000000c00000013ffffffe8fffffffe",
            INIT_1D => X"00000014ffffffc4fffffffbfffffff4ffffffdcfffffffb00000036ffffffd2",
            INIT_1E => X"000000160000000400000008ffffffff0000000100000000ffffffc7ffffffd9",
            INIT_1F => X"00000015ffffffee0000003e0000004a0000000f0000004d000000700000004b",
            INIT_20 => X"0000002700000019fffffffc00000026000000020000000bffffffec00000033",
            INIT_21 => X"fffffffa000000070000002effffffdbffffffd30000001b0000001e00000007",
            INIT_22 => X"0000000000000006fffffffb0000002d0000000cffffffd8fffffff80000002e",
            INIT_23 => X"fffffff2fffffff6ffffffb1ffffffe0ffffffd600000000ffffffe600000004",
            INIT_24 => X"0000000e0000000e00000017ffffffe2fffffff800000039ffffffb3ffffffd8",
            INIT_25 => X"ffffffe0fffffff1ffffffc4ffffffe8ffffffd10000001dfffffff8ffffffdf",
            INIT_26 => X"0000001e00000001ffffffdfffffffbf00000016fffffff7ffffffe60000000f",
            INIT_27 => X"ffffffec0000003100000011ffffffe7fffffffe00000033ffffffe7ffffffe1",
            INIT_28 => X"0000001c0000001c0000001f00000014fffffffbfffffffb00000019ffffffff",
            INIT_29 => X"0000000800000029ffffffeeffffffc900000039ffffffc0ffffffbd0000000f",
            INIT_2A => X"ffffff9fffffffaaffffffbdffffffcbffffffa3ffffffa8fffffff600000008",
            INIT_2B => X"000000200000000f00000041000000310000001100000008ffffffe200000003",
            INIT_2C => X"ffffff9cffffffb0ffffff7dffffffda0000000e0000001f000000150000000c",
            INIT_2D => X"0000001b0000003300000041fffffffffffffffefffffff4ffffffeeffffffbe",
            INIT_2E => X"ffffffe9fffffff400000005ffffffe800000007000000100000001f00000018",
            INIT_2F => X"fffffff60000001e00000018fffffffd00000000fffffff9fffffff4fffffff9",
            INIT_30 => X"ffffffeb00000009ffffffe3ffffffe3ffffffd9000000090000000100000003",
            INIT_31 => X"fffffff9ffffffdf0000002000000000ffffffe10000003dffffffdeffffffdd",
            INIT_32 => X"ffffffeb0000000cfffffffeffffffe900000015fffffffafffffff10000000d",
            INIT_33 => X"00000012fffffff0fffffff9fffffff8ffffffd7ffffffcf0000002200000015",
            INIT_34 => X"0000000b00000004ffffffff000000090000001000000008fffffffb00000011",
            INIT_35 => X"00000017000000080000000c0000002dfffffff0fffffff800000008ffffffc5",
            INIT_36 => X"0000001effffffe6ffffffbf0000001d0000000d0000000b000000210000001f",
            INIT_37 => X"0000002c000000330000000b00000013ffffffe30000001700000003ffffffd1",
            INIT_38 => X"000000160000000ffffffff900000018fffffff4000000280000001100000015",
            INIT_39 => X"0000000c0000002800000003fffffff900000024ffffffe50000000b0000000c",
            INIT_3A => X"0000005500000017000000480000003400000002000000440000002bffffffc7",
            INIT_3B => X"0000001e00000003ffffffef00000000fffffffcffffffdaffffffde00000039",
            INIT_3C => X"fffffffa00000022fffffffafffffff30000002dfffffffc0000002400000003",
            INIT_3D => X"0000000e00000014fffffff6000000240000001efffffff10000001bfffffff2",
            INIT_3E => X"0000001cffffffdf0000001a000000030000001c0000000b000000190000000c",
            INIT_3F => X"ffffffee0000000000000004ffffffd90000000ffffffff1ffffffe3fffffffb",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE22;


    MEM_IWGHT_LAYER1_INSTANCE23 : if BRAM_NAME = "iwght_layer1_instance23" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff40000000bfffffff80000000300000007fffffff5000000180000002a",
            INIT_01 => X"0000000b000000070000001efffffff00000000300000026ffffffe40000002d",
            INIT_02 => X"00000015fffffff40000001a00000003000000110000000cffffffdb00000004",
            INIT_03 => X"00000029ffffffecffffffd9fffffff8ffffffef0000000bffffffb20000000a",
            INIT_04 => X"0000003a00000034ffffffeffffffff900000016ffffffd6ffffffc600000001",
            INIT_05 => X"0000001500000006ffffffd50000001700000012ffffffe00000000900000029",
            INIT_06 => X"0000001c0000000d0000001400000011ffffffff0000002500000007ffffffe7",
            INIT_07 => X"000000060000001affffffe8fffffff100000001fffffff8fffffff900000015",
            INIT_08 => X"0000000600000009ffffffef0000002b0000000b0000000f0000000c0000000c",
            INIT_09 => X"0000001600000000fffffffd00000002ffffffee0000000bfffffff7fffffffa",
            INIT_0A => X"fffffff2ffffffecfffffff800000014fffffff40000000400000017ffffffe0",
            INIT_0B => X"0000000400000000ffffffe60000001100000010ffffffe500000002fffffff0",
            INIT_0C => X"ffffffefffffffe9ffffffe9ffffffe700000006fffffff9fffffff60000000f",
            INIT_0D => X"0000001f0000001600000012fffffffb00000032fffffffcffffffdffffffff9",
            INIT_0E => X"00000009ffffffd1ffffffe6ffffffe1ffffffe8ffffffccfffffff00000003c",
            INIT_0F => X"00000052000000130000001200000035ffffffeefffffffaffffffbdffffffe0",
            INIT_10 => X"fffffff5ffffffff00000022ffffffd9000000380000001e0000003200000053",
            INIT_11 => X"fffffff50000001e00000010ffffffe8fffffff7ffffffdd0000003900000002",
            INIT_12 => X"ffffffefffffffe9fffffff4fffffff5ffffffdafffffff50000000000000015",
            INIT_13 => X"fffffff900000045ffffffff000000050000002c000000210000001600000020",
            INIT_14 => X"00000007ffffffde0000000fffffffeeffffffefffffffe70000002a00000015",
            INIT_15 => X"00000036ffffffc50000002800000019ffffffa400000015ffffffe8ffffffc0",
            INIT_16 => X"ffffffffffffffbdffffffe200000013ffffffebffffffee00000022ffffffe1",
            INIT_17 => X"0000002500000009ffffffab00000033ffffffdeffffffc5ffffffee00000003",
            INIT_18 => X"ffffffb1ffffffbcffffffd7ffffffddfffffff3ffffffd1ffffffe1ffffffee",
            INIT_19 => X"000000000000000b000000010000001cffffff97ffffffaefffffff0ffffffb2",
            INIT_1A => X"fffffff2fffffff7000000010000000c000000180000001effffffe2fffffff4",
            INIT_1B => X"00000005ffffffedfffffffefffffff800000027ffffffdf000000110000001d",
            INIT_1C => X"00000023fffffff9ffffffcdffffffec00000002ffffffddffffffe7fffffffe",
            INIT_1D => X"ffffffee000000090000000dffffffefffffffe700000020ffffffe3fffffff7",
            INIT_1E => X"0000000b000000100000003400000002fffffff2ffffffd4ffffffe9ffffffe4",
            INIT_1F => X"00000028000000170000000800000014fffffffcffffffedfffffff700000013",
            INIT_20 => X"000000170000003c0000002b0000000b00000034000000250000000800000004",
            INIT_21 => X"fffffffc00000012000000250000002000000025ffffffd3000000030000002f",
            INIT_22 => X"fffffff9ffffffdf00000013000000160000002700000012ffffffea0000000e",
            INIT_23 => X"0000001b0000001600000002ffffffe7ffffffe3ffffffd1fffffffcffffffed",
            INIT_24 => X"00000007000000010000000b0000000a000000130000000f0000000b00000012",
            INIT_25 => X"ffffffb90000000e0000002e0000001a000000060000001b0000002600000021",
            INIT_26 => X"0000002e00000003fffffff30000000b00000015ffffffd700000018fffffff7",
            INIT_27 => X"ffffffabffffffaeffffffeffffffff0ffffffc3fffffff2ffffffc4ffffffd3",
            INIT_28 => X"000000100000002700000030000000030000002800000009ffffffc7ffffffc7",
            INIT_29 => X"ffffffca000000070000002dffffffd8ffffffea00000025fffffffd0000001d",
            INIT_2A => X"fffffffe00000009fffffffdfffffff600000010ffffffed000000000000000f",
            INIT_2B => X"00000016fffffffafffffffd00000003ffffffec00000008fffffffbffffffe1",
            INIT_2C => X"ffffffe0ffffffd70000000b0000002b00000015000000000000004800000060",
            INIT_2D => X"0000001500000008ffffffeeffffffd6ffffffe5ffffffbcffffffb800000004",
            INIT_2E => X"00000009fffffff000000006ffffffea0000000900000006ffffffd4fffffff8",
            INIT_2F => X"fffffff10000000700000022fffffffb000000020000001a0000000300000012",
            INIT_30 => X"0000001300000000fffffff8ffffffec00000008ffffffe800000009ffffffff",
            INIT_31 => X"00000036ffffffe4ffffffbeffffffe9000000010000002affffffeb00000019",
            INIT_32 => X"0000004d0000004700000013000000420000003700000017ffffffeb0000001e",
            INIT_33 => X"0000001800000045ffffffe80000000e00000028000000280000004100000011",
            INIT_34 => X"0000004a0000001a0000004b000000380000002200000017fffffff900000008",
            INIT_35 => X"0000002c000000260000001f0000002e0000002e000000170000003e00000037",
            INIT_36 => X"000000160000002ffffffffffffffffcffffffe7000000350000003e00000021",
            INIT_37 => X"fffffff00000000b00000004fffffff5ffffffe6fffffffcffffffc900000010",
            INIT_38 => X"fffffff0fffffff3fffffff0ffffffc7ffffffdaffffffc80000000b0000000b",
            INIT_39 => X"000000030000001200000000ffffffdfffffffd900000000000000090000000a",
            INIT_3A => X"ffffffeafffffff700000013fffffff2000000180000002e0000002300000019",
            INIT_3B => X"ffffffeafffffff0fffffff1ffffffd100000026000000000000000afffffff9",
            INIT_3C => X"0000000600000021ffffffd5ffffffe40000001d0000000e0000001b00000008",
            INIT_3D => X"fffffff0fffffffbfffffff600000022fffffffbfffffff900000027ffffffe9",
            INIT_3E => X"fffffff4fffffff8ffffffd8fffffff1ffffffe1ffffffdfffffffec00000000",
            INIT_3F => X"00000024fffffffc000000290000002afffffffcffffffc9ffffffbbffffffba",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE23;


    MEM_IWGHT_LAYER1_INSTANCE24 : if BRAM_NAME = "iwght_layer1_instance24" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000034ffffffe2ffffffc7ffffffdb0000000b0000002300000007fffffff1",
            INIT_01 => X"ffffffc300000000ffffffef000000060000000d00000022fffffff500000011",
            INIT_02 => X"0000002b00000017fffffff40000000afffffff1000000290000000800000000",
            INIT_03 => X"0000000a00000000fffffffefffffff5ffffffebfffffff600000019fffffffe",
            INIT_04 => X"0000000effffffc400000012fffffff7ffffffdcfffffff5ffffffda00000007",
            INIT_05 => X"ffffffed00000011ffffffe000000007fffffffd00000004fffffffbfffffffd",
            INIT_06 => X"00000006fffffff0ffffffdbffffffebffffffefffffffe0ffffffd200000000",
            INIT_07 => X"fffffffbfffffff800000024ffffffdcffffffefffffffe700000018ffffffee",
            INIT_08 => X"0000002300000033ffffffccffffffddffffffe40000000d000000170000000e",
            INIT_09 => X"fffffff9ffffffe1fffffff3ffffffcbfffffff1fffffffcfffffffd0000000c",
            INIT_0A => X"0000002c0000000bfffffff9ffffffe9fffffff90000000effffffccffffffd4",
            INIT_0B => X"ffffffecffffffe500000049000000530000001200000012000000400000003d",
            INIT_0C => X"ffffffe3ffffffd7ffffffd8ffffffd8ffffffeb00000018ffffffdc0000002f",
            INIT_0D => X"ffffffe2fffffffdfffffffffffffff60000000c00000003fffffffd0000000c",
            INIT_0E => X"0000001affffffdaffffffdd0000003100000024fffffff1ffffffebffffffdf",
            INIT_0F => X"00000039fffffff80000001a00000039fffffff8fffffff1fffffff3ffffffea",
            INIT_10 => X"ffffffc6ffffffcaffffffe0ffffffe700000029ffffffe40000001500000057",
            INIT_11 => X"ffffffd5fffffff6ffffffdbffffffdaffffffe6ffffffd5fffffffeffffffdc",
            INIT_12 => X"0000001b00000004ffffffff00000006ffffffee0000000000000005fffffff1",
            INIT_13 => X"ffffffee0000000000000009ffffffee0000000affffffff00000012fffffffa",
            INIT_14 => X"000000130000000d000000090000001000000022000000240000001300000004",
            INIT_15 => X"00000036000000220000001300000014fffffffeffffffd4fffffff8fffffff9",
            INIT_16 => X"000000270000004c00000029fffffff400000021000000000000003d00000036",
            INIT_17 => X"fffffff900000012fffffff7ffffffddffffffff000000510000006500000056",
            INIT_18 => X"00000052fffffff900000014fffffffc00000018fffffffdffffffc3ffffffd6",
            INIT_19 => X"00000042000000480000002f000000570000004000000044000000330000006c",
            INIT_1A => X"0000001600000008ffffffb9ffffff98ffffff830000000000000011ffffffdd",
            INIT_1B => X"fffffffbffffffe0ffffffc5ffffffc2ffffffafffffffca0000000000000014",
            INIT_1C => X"00000010000000100000000cfffffff3ffffffd60000002cffffffe5ffffffe1",
            INIT_1D => X"000000190000000300000013fffffff9ffffffeb0000000e000000170000000a",
            INIT_1E => X"fffffffb0000000cfffffff800000001fffffff800000005fffffff600000020",
            INIT_1F => X"0000001e0000000d0000000d00000023000000090000001bffffffdafffffff8",
            INIT_20 => X"fffffff4fffffffd000000270000002000000012000000010000000400000014",
            INIT_21 => X"ffffffee00000017000000290000000effffffe300000000ffffffc3ffffffdf",
            INIT_22 => X"ffffffe300000003ffffffffffffffe700000004ffffffcbffffffdb0000001e",
            INIT_23 => X"000000270000001f0000001300000016fffffff1fffffff0ffffffc6fffffff0",
            INIT_24 => X"fffffff7ffffffd4ffffffbaffffff8cfffffffbffffffceffffffca00000023",
            INIT_25 => X"fffffff2ffffffeaffffffef0000000b00000013ffffffe00000001a0000000d",
            INIT_26 => X"00000000fffffffd00000009000000280000000b000000400000004700000036",
            INIT_27 => X"ffffffe6ffffffe7fffffffefffffffa000000060000001c00000032ffffffde",
            INIT_28 => X"fffffff500000006fffffffb0000004b00000042000000380000000d00000006",
            INIT_29 => X"00000018fffffff6000000230000003000000011ffffffe5ffffffa1ffffffb8",
            INIT_2A => X"fffffff20000001c0000001400000010ffffffc8ffffffbfffffffe900000013",
            INIT_2B => X"00000018000000390000002affffffdeffffffa1ffffffd5fffffffcfffffffb",
            INIT_2C => X"00000004ffffffffffffffe7ffffffd7ffffffbd0000001800000012fffffff5",
            INIT_2D => X"00000027ffffffe8fffffffefffffff6fffffffafffffff6fffffffc00000014",
            INIT_2E => X"ffffffc1ffffff96ffffff9d000000000000000ffffffff00000004400000033",
            INIT_2F => X"000000060000001200000000ffffffd6ffffffdcffffffccffffffebffffffee",
            INIT_30 => X"000000030000001bffffffeb0000001afffffffdfffffff0000000000000000f",
            INIT_31 => X"fffffff200000001ffffffe7fffffff60000000a0000000efffffff2ffffffee",
            INIT_32 => X"fffffff4ffffffdd0000000cfffffff700000001ffffffe1fffffff400000004",
            INIT_33 => X"fffffff6ffffffc7ffffffdcffffffeaffffffeeffffffe7fffffff900000012",
            INIT_34 => X"fffffffa000000050000000100000021ffffffe6ffffffc6ffffffe000000001",
            INIT_35 => X"000000160000000ffffffff20000001b0000000bffffffd3fffffffcffffffcc",
            INIT_36 => X"0000001cffffffcdffffffcaffffffc7ffffffe3ffffffeeffffffea00000020",
            INIT_37 => X"ffffffec00000014fffffff10000000500000011fffffff20000002100000025",
            INIT_38 => X"0000000e00000012000000010000000efffffffe0000000500000003ffffffef",
            INIT_39 => X"fffffff7ffffffeaffffffdbffffffe5ffffffeeffffffecffffffe50000001a",
            INIT_3A => X"0000007000000051000000140000003d0000004500000000ffffffd3ffffffe3",
            INIT_3B => X"00000047ffffffe6fffffffe00000011fffffffe00000015fffffff3fffffff7",
            INIT_3C => X"00000020fffffffc0000003b0000003e0000001300000029ffffffd900000029",
            INIT_3D => X"000000020000000100000007ffffffff00000021ffffffdb0000004500000044",
            INIT_3E => X"0000000effffffe6000000120000001e0000002900000013000000030000000c",
            INIT_3F => X"000000010000000c00000005fffffff1ffffffdd00000008fffffff7ffffffe7",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE24;


    MEM_IWGHT_LAYER1_INSTANCE25 : if BRAM_NAME = "iwght_layer1_instance25" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000190000000c0000000bfffffff6fffffff9ffffffebfffffff800000000",
            INIT_01 => X"ffffffdbfffffffa00000001fffffff60000000a000000210000003100000010",
            INIT_02 => X"0000002500000001fffffff600000010fffffff5ffffffe2fffffff000000008",
            INIT_03 => X"0000000a00000000000000070000001a0000000affffffebfffffffaffffffee",
            INIT_04 => X"0000002500000014000000190000000200000005ffffffccffffffb8ffffffc9",
            INIT_05 => X"00000017fffffff4fffffff2fffffff4ffffffce0000001dfffffff700000007",
            INIT_06 => X"ffffffebffffffe20000000b000000070000002a00000020ffffffdffffffffa",
            INIT_07 => X"0000000f00000000fffffffbfffffffe00000028000000110000000500000006",
            INIT_08 => X"00000018fffffffd000000310000000e000000260000001a0000002e00000020",
            INIT_09 => X"00000034000000360000004fffffffd7ffffffd700000019ffffffd5ffffffce",
            INIT_0A => X"000000240000004cffffffd9ffffffe6ffffffe3ffffffd7fffffffafffffff2",
            INIT_0B => X"00000005fffffff7ffffffe5ffffffe6ffffffd2ffffffdcffffffdc0000002b",
            INIT_0C => X"000000160000001a000000280000000b000000160000000c0000000300000024",
            INIT_0D => X"fffffffe00000010ffffffebfffffff1ffffffe8000000160000003300000009",
            INIT_0E => X"ffffffe400000004ffffffdf000000090000001a0000000000000003ffffffde",
            INIT_0F => X"fffffff7ffffffe4fffffff8fffffff10000001f0000001effffffd1ffffffeb",
            INIT_10 => X"ffffffccffffffd9fffffffd0000001700000000ffffffe9fffffffd00000008",
            INIT_11 => X"0000000c0000002b0000003100000028000000190000000000000008ffffffe6",
            INIT_12 => X"00000003ffffffec00000001ffffffeb0000000500000005ffffffec00000023",
            INIT_13 => X"ffffffd8ffffffe2000000470000002f0000001200000058000000430000000b",
            INIT_14 => X"000000150000000d00000004fffffffffffffff7ffffffe40000000a00000011",
            INIT_15 => X"ffffffffffffffe5fffffffffffffffeffffffe6fffffffc0000001000000009",
            INIT_16 => X"00000004fffffff5ffffffcfffffffd9ffffffe40000001d0000000d0000002a",
            INIT_17 => X"fffffff5fffffffb0000002e00000029000000220000001b0000002900000007",
            INIT_18 => X"00000012fffffffbfffffff1000000170000001effffffda0000003e00000051",
            INIT_19 => X"000000000000000d0000002a000000090000001a0000000a00000004fffffff1",
            INIT_1A => X"ffffffe7000000160000002600000023ffffffe4ffffffeeffffffe6ffffffec",
            INIT_1B => X"00000005000000240000001e00000000ffffffe500000003ffffffebffffffdd",
            INIT_1C => X"fffffff000000008fffffffbfffffff6ffffffec00000008fffffffffffffffb",
            INIT_1D => X"00000000ffffffe0fffffff00000000000000006fffffffbfffffffa0000000f",
            INIT_1E => X"ffffffec00000000ffffffeffffffff700000006ffffffe80000000400000004",
            INIT_1F => X"0000000d00000012fffffffcfffffff2ffffffeb00000010fffffffffffffff7",
            INIT_20 => X"0000001e00000006000000020000000cffffffe8ffffffe8fffffff60000001a",
            INIT_21 => X"0000000b000000000000001afffffff9ffffffef0000000cfffffffbfffffffd",
            INIT_22 => X"ffffffe9fffffff5ffffffedfffffff1fffffffefffffff800000007fffffff5",
            INIT_23 => X"ffffffe4ffffffe9ffffffebffffffe4ffffffecffffffe5ffffffda00000007",
            INIT_24 => X"000000000000000b000000080000000c00000000000000070000000dffffffe5",
            INIT_25 => X"ffffffdffffffffbffffffffffffffe8fffffff6ffffffeafffffff2ffffffed",
            INIT_26 => X"ffffffed0000000bffffffebffffffebffffffe5ffffffe30000000600000014",
            INIT_27 => X"00000004fffffffbffffffeaffffffe700000008ffffffeefffffff0ffffffed",
            INIT_28 => X"ffffffe8fffffffaffffffedfffffff3ffffffe800000000ffffffecfffffff8",
            INIT_29 => X"ffffffe600000004fffffff5ffffffedffffffebfffffff3fffffff2fffffff3",
            INIT_2A => X"ffffffdfffffffe1ffffffefffffffeeffffffe2ffffffedffffffee0000000a",
            INIT_2B => X"ffffffe50000000100000005ffffffecfffffff0000000090000000600000000",
            INIT_2C => X"ffffffebfffffffbfffffff8fffffff00000000affffffdcffffffeb00000008",
            INIT_2D => X"fffffff00000000100000000ffffffe800000004ffffffe30000000a00000001",
            INIT_2E => X"0000000d00000005fffffff6fffffff4fffffffaffffffeefffffffbffffffe6",
            INIT_2F => X"0000000c0000000000000001fffffffefffffff4ffffffd9ffffffddfffffffd",
            INIT_30 => X"fffffff1fffffff0fffffff100000003fffffffcfffffff5fffffff8ffffffe5",
            INIT_31 => X"00000000fffffffeffffffffffffffe1ffffffe5000000000000000c0000000b",
            INIT_32 => X"fffffff500000008ffffffe70000000ffffffff000000003ffffffeeffffffec",
            INIT_33 => X"00000007fffffffa0000000a0000000dffffffe400000000ffffffec00000006",
            INIT_34 => X"ffffffe2fffffffaffffffeeffffffe8ffffffeaffffffe9ffffffe1ffffffe3",
            INIT_35 => X"ffffffe4fffffff5fffffffcfffffff00000000500000005ffffffdf00000001",
            INIT_36 => X"ffffffeaffffffe7ffffffff0000000affffffe5ffffffec0000000300000003",
            INIT_37 => X"0000000dffffffe6fffffff4ffffffe9ffffffe9ffffffffffffffe6fffffff6",
            INIT_38 => X"ffffffefffffffe90000000000000008fffffff5ffffffedffffffe7fffffff8",
            INIT_39 => X"fffffffcffffffee00000004ffffffe7ffffffe9ffffffec00000007fffffffb",
            INIT_3A => X"fffffffc000000070000000affffffe9fffffffffffffffcffffffed00000001",
            INIT_3B => X"000000020000000efffffff5fffffff3fffffff70000000200000002ffffffe2",
            INIT_3C => X"fffffff800000000fffffffbffffffe2000000080000000100000002ffffffe7",
            INIT_3D => X"0000000affffffeafffffff2fffffffa00000000fffffff7ffffffef00000005",
            INIT_3E => X"0000000afffffffb0000000900000009ffffffecffffffed0000000000000002",
            INIT_3F => X"0000000800000016fffffffffffffff1fffffff900000008fffffffcfffffff2",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE25;


    MEM_IWGHT_LAYER1_INSTANCE26 : if BRAM_NAME = "iwght_layer1_instance26" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000b0000000a00000007ffffffe80000000800000000ffffffecfffffff6",
            INIT_01 => X"00000015ffffffedfffffff800000014ffffffd3fffffff2ffffffefffffffeb",
            INIT_02 => X"00000010000000310000003c0000000a0000000a00000018ffffffdb00000001",
            INIT_03 => X"ffffffe5ffffffc1ffffffd80000000bffffffdb0000002b000000370000002f",
            INIT_04 => X"0000001a0000001cfffffff9fffffffcffffffc7ffffffb6ffffffd8ffffffb8",
            INIT_05 => X"0000001700000022fffffffa0000003000000055000000230000004d0000003b",
            INIT_06 => X"0000001b00000021fffffffdffffffdefffffff0fffffffb0000000affffffea",
            INIT_07 => X"fffffffcffffffe6ffffffcbffffffe2fffffff1ffffffd2ffffffd800000017",
            INIT_08 => X"000000050000000b0000000bfffffff8ffffffff00000016ffffffedffffffe7",
            INIT_09 => X"ffffff95ffffffb9fffffff20000001afffffff3000000230000000d0000002a",
            INIT_0A => X"fffffff40000000000000017ffffffc9000000140000000000000002ffffffb0",
            INIT_0B => X"ffffffdfffffffdafffffff600000008ffffffe2fffffff400000003fffffffe",
            INIT_0C => X"0000000cfffffffb0000000000000010fffffff7ffffffceffffffcbffffffd1",
            INIT_0D => X"ffffffe9fffffff10000000f000000130000001dffffffeaffffffc4fffffff9",
            INIT_0E => X"fffffffc00000006ffffffcc0000001400000002ffffffe30000000e00000010",
            INIT_0F => X"000000110000001b0000002200000016000000150000000f0000000ffffffffb",
            INIT_10 => X"fffffff2ffffffd0ffffffabffffffa80000000000000001ffffffd900000019",
            INIT_11 => X"0000003500000044000000210000000c0000003000000010ffffffd00000000b",
            INIT_12 => X"00000021000000020000001a00000007fffffff90000000d00000001ffffffe9",
            INIT_13 => X"ffffffb7fffffff4ffffffefffffffef0000001f000000190000000600000014",
            INIT_14 => X"ffffffc1ffffffb6ffffffc1ffffffbdffffffedffffffd6ffffffe9ffffffdf",
            INIT_15 => X"fffffff000000004000000050000000e0000000effffffe200000002ffffffd5",
            INIT_16 => X"00000027ffffffd6ffffffeeffffffe30000000e000000190000000500000008",
            INIT_17 => X"ffffffe6fffffff0fffffffcfffffff8000000190000003bffffffdcfffffff5",
            INIT_18 => X"0000002200000010000000060000001900000023ffffffeb0000001500000015",
            INIT_19 => X"0000001dffffffddffffffccffffffd40000000a00000005ffffffee00000015",
            INIT_1A => X"ffffffe5ffffffbdffffff9d00000007fffffffcffffffda0000002700000016",
            INIT_1B => X"ffffff9afffffffbffffffd9ffffffccffffffd0ffffffee00000032ffffffec",
            INIT_1C => X"00000027fffffffd0000001e00000020000000180000000500000015ffffffce",
            INIT_1D => X"00000015fffffffdfffffff20000002300000001ffffffe7000000070000001f",
            INIT_1E => X"ffffffeeffffffe300000003000000090000000a0000001700000015fffffff8",
            INIT_1F => X"ffffffc100000009ffffffffffffffe6fffffffbffffffe00000000e0000000c",
            INIT_20 => X"00000017fffffff2ffffffdeffffffecffffffc9ffffffc5ffffffccffffffb8",
            INIT_21 => X"0000000b00000007fffffffbffffffd5ffffffbe00000001fffffff7ffffffeb",
            INIT_22 => X"fffffff3000000120000003500000039ffffffed000000210000001900000005",
            INIT_23 => X"fffffff7fffffffcffffffd80000002f00000017000000040000001a0000000b",
            INIT_24 => X"ffffffff0000002400000012000000010000000d0000000f0000000cfffffffe",
            INIT_25 => X"ffffffb9ffffffd0ffffff98ffffffc9fffffff5ffffffe9fffffff7fffffffb",
            INIT_26 => X"0000004e00000035000000330000000c00000009fffffff0ffffffdeffffff8a",
            INIT_27 => X"0000004300000034000000260000005900000026000000260000005500000043",
            INIT_28 => X"0000002affffffe2ffffffecfffffffd00000008000000180000002c00000031",
            INIT_29 => X"ffffffe6000000080000000afffffffa0000001800000031ffffffe600000026",
            INIT_2A => X"ffffffe4ffffffef00000022000000280000002c0000000f0000001b0000001b",
            INIT_2B => X"ffffffdfffffffff0000000000000025ffffffedfffffff7fffffffeffffffcd",
            INIT_2C => X"fffffff0ffffffd9ffffffc7ffffffedfffffffdffffffeeffffffe000000000",
            INIT_2D => X"fffffff6fffffffbfffffffcfffffff40000001affffffff0000000a00000039",
            INIT_2E => X"0000001effffffebfffffff600000023ffffffeeffffffdeffffffe800000000",
            INIT_2F => X"ffffffe1ffffffed0000001b000000100000000600000016fffffffdfffffffc",
            INIT_30 => X"00000023fffffff900000020fffffffcfffffff0fffffff1fffffff1ffffffec",
            INIT_31 => X"0000001800000000fffffff7ffffffed00000022000000060000002c0000001b",
            INIT_32 => X"ffffffe7ffffffccfffffffc000000030000002800000015000000130000000b",
            INIT_33 => X"fffffffd0000000effffffe1ffffffcfffffffebffffffe1ffffffcf0000001a",
            INIT_34 => X"fffffffffffffff900000034000000170000000000000022000000040000000a",
            INIT_35 => X"0000000a000000060000000b000000120000001800000012ffffffe5fffffffe",
            INIT_36 => X"ffffffd3ffffffe2ffffffdbffffffab0000002affffffedffffffe300000006",
            INIT_37 => X"0000001affffffd70000000900000051ffffffe3fffffff500000018ffffffd2",
            INIT_38 => X"fffffffaffffffdcffffffe5ffffffbbffffffccffffffd1ffffffd2fffffff3",
            INIT_39 => X"ffffffeaffffffdd00000014fffffff1ffffffdcfffffff5fffffff0ffffffea",
            INIT_3A => X"ffffffe70000000c0000000dffffffe000000016fffffff5fffffff000000017",
            INIT_3B => X"00000006ffffffe1ffffffc900000007ffffffe8ffffffdb0000002200000009",
            INIT_3C => X"00000000ffffffee0000002200000000ffffffe90000001d0000000affffffe9",
            INIT_3D => X"00000011fffffff10000000500000035ffffffe0000000020000003400000005",
            INIT_3E => X"000000040000000300000016fffffff500000016fffffff8fffffff9fffffff1",
            INIT_3F => X"000000450000005a0000001d0000006f0000003f000000200000004500000036",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE26;


    MEM_IWGHT_LAYER1_INSTANCE27 : if BRAM_NAME = "iwght_layer1_instance27" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffd2fffffffbffffffe5ffffffe1fffffff2ffffffe20000000100000035",
            INIT_01 => X"ffffffd5fffffffa00000031fffffff4fffffffc00000008ffffffd3ffffffae",
            INIT_02 => X"ffffffe0ffffffdb00000014ffffffe7ffffffdaffffffe0fffffff900000034",
            INIT_03 => X"0000007b0000001700000049000000350000001bfffffff2ffffffe1fffffffe",
            INIT_04 => X"00000011ffffffdcffffffd6000000360000002700000069000000380000005b",
            INIT_05 => X"ffffffefffffffe60000000fffffffe6ffffffe5ffffffe800000005fffffffe",
            INIT_06 => X"fffffff700000016fffffff1ffffffec000000220000001cffffffe700000012",
            INIT_07 => X"ffffffc8fffffffb00000035fffffff1ffffffe50000001efffffff100000000",
            INIT_08 => X"00000000ffffffe100000000fffffff90000001600000004fffffff700000014",
            INIT_09 => X"fffffff000000026fffffff9ffffffd7ffffffbd0000001e0000003f00000008",
            INIT_0A => X"000000210000000a0000000affffffd8000000010000001afffffff9ffffffd8",
            INIT_0B => X"fffffff0ffffffd100000001ffffffdfffffffd400000009ffffffecffffffef",
            INIT_0C => X"0000000f000000280000000c0000001afffffff0fffffff6ffffffca00000010",
            INIT_0D => X"0000000b00000019ffffffe9ffffffd800000006fffffffe00000028fffffffc",
            INIT_0E => X"ffffffd6ffffffb0000000150000002300000018000000140000000efffffff7",
            INIT_0F => X"ffffffccffffffd5fffffff8fffffff0ffffffd4ffffffe6ffffffd700000003",
            INIT_10 => X"00000006ffffffd1ffffffeaffffffe200000002ffffffd8ffffffc2ffffffcb",
            INIT_11 => X"fffffff8ffffffd900000033fffffff7ffffffdf000000350000003300000031",
            INIT_12 => X"fffffffcffffffc1fffffff2ffffffd0ffffffd3fffffff9ffffffe500000023",
            INIT_13 => X"00000044ffffffddffffffc50000000d000000160000000ffffffff9fffffff4",
            INIT_14 => X"ffffffc2fffffff0fffffff1ffffffebffffffdb00000020ffffffe3ffffffd9",
            INIT_15 => X"ffffffddffffffeaffffffceffffffd7fffffff0ffffffdd0000001000000001",
            INIT_16 => X"fffffff9ffffffccffffffe2ffffffc5ffffffcb00000003fffffffeffffff9f",
            INIT_17 => X"00000022ffffffbe00000002fffffffaffffffe8fffffffaffffffdf00000001",
            INIT_18 => X"ffffffd2ffffffe4ffffffddfffffff800000003ffffffdfffffffd900000048",
            INIT_19 => X"ffffffcd0000001600000017ffffff9cffffffdafffffffaffffffd7fffffff4",
            INIT_1A => X"0000000bffffffd00000003000000005ffffffc4fffffff80000003600000007",
            INIT_1B => X"fffffffc00000028fffffff2ffffffb40000000b0000000efffffff30000002b",
            INIT_1C => X"0000003c0000004e00000069000000390000003800000006fffffff7fffffff1",
            INIT_1D => X"ffffffc4ffffffda00000000fffffffaffffffe0000000230000006600000055",
            INIT_1E => X"fffffffcfffffff9ffffffd6ffffffdfffffffaaffffffcaffffffdbffffffb1",
            INIT_1F => X"fffffffc0000000d00000004ffffffd0fffffffdfffffffaffffffb4fffffff2",
            INIT_20 => X"ffffffeffffffff1ffffffdb00000018fffffffbffffffe4ffffffeafffffff7",
            INIT_21 => X"00000001ffffffe40000004700000013ffffffebffffffdcffffffe5fffffff2",
            INIT_22 => X"0000001cffffffdbffffffd500000023ffffffeeffffffd00000003d0000002e",
            INIT_23 => X"ffffffd600000007000000270000000bffffffdefffffff20000000bfffffff0",
            INIT_24 => X"ffffffdf0000000afffffff9ffffffe90000000cffffffe90000002100000003",
            INIT_25 => X"ffffffe6fffffff5fffffff7fffffffbfffffff2ffffffe900000015ffffffe1",
            INIT_26 => X"ffffffe3ffffffd6fffffffcffffffe7ffffffd10000003200000007ffffffed",
            INIT_27 => X"fffffff80000002800000014ffffffd6ffffffd70000000effffffdcfffffffb",
            INIT_28 => X"ffffffecffffffcbffffffd80000002900000011000000030000003a0000000e",
            INIT_29 => X"ffffffccffffffdc0000004300000017ffffffef00000007fffffff4ffffffea",
            INIT_2A => X"00000014ffffffd2ffffffef0000000cffffffe2ffffffe10000000400000005",
            INIT_2B => X"000000230000001a0000002100000011fffffff90000000a0000001200000024",
            INIT_2C => X"fffffff2fffffff0fffffff0000000140000000cfffffffcfffffffc00000012",
            INIT_2D => X"fffffff2000000090000001300000003fffffff1000000370000003600000019",
            INIT_2E => X"fffffffb00000041fffffffc0000000a00000015ffffffce0000000ffffffffc",
            INIT_2F => X"0000002c00000010ffffffd2fffffff8ffffffd600000009fffffffbffffffe6",
            INIT_30 => X"0000001e00000031fffffffeffffffd50000003a000000230000000c00000011",
            INIT_31 => X"0000000c0000001900000006fffffff6ffffffc900000034fffffffcffffffdc",
            INIT_32 => X"00000010fffffffaffffffda00000001fffffff3fffffff90000000800000000",
            INIT_33 => X"ffffffebffffffe0fffffffffffffffa000000060000000e00000000ffffffc4",
            INIT_34 => X"000000130000000dfffffff40000001f00000007fffffff500000000ffffffe0",
            INIT_35 => X"00000006fffffff9fffffff700000015fffffff1000000070000002a0000000a",
            INIT_36 => X"fffffff0ffffffb7ffffffc4ffffffffffffffecfffffff00000000a00000036",
            INIT_37 => X"00000017000000070000001dffffffeb0000001cfffffff1ffffffedffffffe5",
            INIT_38 => X"ffffffddfffffffdfffffff1ffffffd2fffffffc00000024fffffff60000001c",
            INIT_39 => X"fffffff800000010ffffffea00000000ffffffa8ffffffdbffffffc4ffffffe7",
            INIT_3A => X"ffffffdd00000007fffffff3ffffffd3ffffffd9ffffffd0ffffffebffffffe5",
            INIT_3B => X"ffffffd4fffffffb00000019000000060000000100000000fffffff40000000b",
            INIT_3C => X"00000007ffffffb7ffffffcdffffffccffffffddfffffff000000007ffffffef",
            INIT_3D => X"fffffff1ffffffebffffffe4ffffffc4ffffffe3ffffffe1ffffffd9ffffffda",
            INIT_3E => X"00000006ffffffdfffffffe0ffffffc8ffffff93ffffffbdffffffa4ffffffcd",
            INIT_3F => X"00000010fffffffa000000040000002dffffffe7000000110000001fffffffdb",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE27;


    MEM_IWGHT_LAYER1_INSTANCE28 : if BRAM_NAME = "iwght_layer1_instance28" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000005b000000660000000d000000480000004a000000100000000a0000000a",
            INIT_01 => X"ffffffe0ffffffd900000007fffffff3ffffffee000000380000009000000053",
            INIT_02 => X"ffffffe7fffffffdfffffff1ffffffdbfffffff3ffffffcaffffffdefffffffc",
            INIT_03 => X"ffffffedfffffffbfffffff9ffffffeffffffffbfffffff400000010fffffff0",
            INIT_04 => X"000000000000001dffffffddffffffedffffffecfffffffe00000009ffffffd0",
            INIT_05 => X"00000008ffffffedfffffffefffffff6fffffffefffffff900000023ffffffe2",
            INIT_06 => X"ffffffffffffffc8ffffffdaffffffcfffffffd20000000fffffffcdffffffca",
            INIT_07 => X"ffffffe9fffffffefffffffb0000003b00000018000000120000003e00000009",
            INIT_08 => X"ffffffed0000000b00000006ffffffeb0000000700000000fffffffc0000000d",
            INIT_09 => X"ffffffc6000000010000000bffffffe2000000000000003b000000450000000f",
            INIT_0A => X"ffffffffffffffe6ffffffff0000003afffffff7ffffffd9ffffffdaffffffe7",
            INIT_0B => X"00000025fffffff100000012fffffff4ffffffdfffffffceffffffddffffffca",
            INIT_0C => X"00000013fffffff5000000020000003e000000340000002a000000180000004e",
            INIT_0D => X"fffffffaffffffc6ffffffe3fffffff3ffffffe3ffffffbf00000006fffffff7",
            INIT_0E => X"000000370000000700000012fffffff000000010fffffff6ffffffda00000008",
            INIT_0F => X"fffffff20000000afffffffcffffffda0000000d0000001effffffec0000000e",
            INIT_10 => X"fffffffeffffffe00000001b000000040000001200000024fffffffdfffffff8",
            INIT_11 => X"0000000c00000022fffffff0fffffffd000000000000000a00000011fffffff5",
            INIT_12 => X"ffffffccffffffcfffffffd6ffffffdaffffffbcffffffc40000001600000017",
            INIT_13 => X"00000025ffffffa10000001c00000012ffffffc5ffffffeeffffffddfffffff8",
            INIT_14 => X"ffffffa5ffffffe1ffffffa0ffffff760000001000000016fffffff000000000",
            INIT_15 => X"0000001f0000000d0000000f00000001ffffffc1000000030000000bffffff7b",
            INIT_16 => X"00000021000000040000002c0000002200000001000000160000002800000000",
            INIT_17 => X"00000039fffffff7ffffffbeffffffaa00000025ffffffe8ffffffe200000011",
            INIT_18 => X"0000001e0000001a00000020fffffff20000002900000028fffffff200000006",
            INIT_19 => X"ffffffcfffffffdbffffffeeffffffdeffffffe8fffffff9ffffffe500000037",
            INIT_1A => X"ffffffe80000001000000021ffffffed000000280000001c00000027ffffffd6",
            INIT_1B => X"0000000ffffffff800000000fffffff90000001a00000012fffffffbfffffff9",
            INIT_1C => X"00000017ffffffd60000002d0000002c0000000dffffffd8ffffffe50000001a",
            INIT_1D => X"ffffffea000000190000000f000000100000000d00000013ffffffe700000015",
            INIT_1E => X"00000002000000100000001b000000200000000b000000000000001100000020",
            INIT_1F => X"0000002afffffff80000002500000006ffffffdffffffffc00000023ffffffff",
            INIT_20 => X"ffffffe00000000bffffffecffffffe300000020fffffffeffffffe80000002e",
            INIT_21 => X"000000230000000c000000120000000300000006ffffffe00000000ffffffff2",
            INIT_22 => X"00000039ffffffc4ffffffdaffffffc3ffffffc9fffffff6ffffffdeffffffb6",
            INIT_23 => X"ffffffc100000023fffffff3fffffffd0000003800000028fffffffc00000003",
            INIT_24 => X"00000019ffffffd6fffffff7ffffffe7fffffff00000001c00000005ffffffff",
            INIT_25 => X"ffffffe100000016ffffffecffffffc3ffffffe0ffffffee00000011fffffff7",
            INIT_26 => X"00000035ffffffdaffffffc7fffffff900000005fffffffb00000033ffffffe7",
            INIT_27 => X"ffffffe1ffffffe3ffffffeeffffffec0000001c00000059ffffffb7fffffffa",
            INIT_28 => X"00000002fffffffbffffffe3000000010000003bffffffe8ffffffdf00000022",
            INIT_29 => X"ffffffdf00000019fffffff4ffffffd3fffffffa0000000dfffffffd00000027",
            INIT_2A => X"fffffff2ffffffe9ffffffe800000016ffffffebffffffe00000001bfffffff3",
            INIT_2B => X"0000002a00000023ffffffcf0000002a00000016ffffffd5ffffffdfffffffc0",
            INIT_2C => X"0000003a000000040000001200000006ffffffe300000003ffffffe400000000",
            INIT_2D => X"000000130000000cffffffc5000000160000000cffffffeb0000001600000017",
            INIT_2E => X"fffffff1fffffff20000000afffffff4fffffff400000008fffffff4ffffffb8",
            INIT_2F => X"ffffffa8fffffffeffffffe2fffffffe00000025ffffffc7fffffff80000000e",
            INIT_30 => X"0000002700000020ffffffe50000001bfffffffeffffffc1ffffffecfffffff3",
            INIT_31 => X"fffffff700000002000000000000000dfffffffa00000009000000250000000c",
            INIT_32 => X"fffffff0ffffffef000000160000004dffffffdcfffffff00000002dffffffed",
            INIT_33 => X"0000001cfffffffdffffffd40000000d0000000effffffad0000002600000013",
            INIT_34 => X"00000012fffffffefffffffb000000060000001200000004fffffff800000000",
            INIT_35 => X"00000005ffffffeafffffff9fffffff9fffffff900000007fffffff2fffffff7",
            INIT_36 => X"fffffff000000001fffffffefffffff6fffffff8fffffff100000003ffffffee",
            INIT_37 => X"0000000000000006ffffffff00000000fffffff4fffffff60000000b00000006",
            INIT_38 => X"fffffffe0000000dffffffff00000006fffffff300000005ffffffe800000000",
            INIT_39 => X"fffffff6fffffff200000006fffffffdffffffe9fffffff60000000efffffff2",
            INIT_3A => X"0000000afffffffc00000006ffffffffffffffefffffffeaffffffea00000007",
            INIT_3B => X"fffffffafffffffbffffffe9fffffff5fffffffa0000000c0000000cfffffff1",
            INIT_3C => X"000000000000000000000006fffffff400000006fffffff2ffffffe700000004",
            INIT_3D => X"ffffffe700000009fffffff700000002ffffffef0000000bfffffff9fffffffe",
            INIT_3E => X"000000080000000afffffff4ffffffec0000001200000002fffffffbfffffff2",
            INIT_3F => X"0000000000000000fffffff100000001fffffff2ffffffed00000000fffffff9",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE28;


    MEM_IWGHT_LAYER1_INSTANCE29 : if BRAM_NAME = "iwght_layer1_instance29" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000a0000000affffffec00000000ffffffec0000000dffffffe70000000e",
            INIT_01 => X"0000000ffffffff3fffffff50000000fffffffed00000010fffffffbffffffec",
            INIT_02 => X"fffffff2fffffffffffffffb00000011fffffff00000000dfffffff40000000a",
            INIT_03 => X"00000001fffffff800000000ffffffe60000000100000000ffffffeefffffffc",
            INIT_04 => X"00000006fffffff800000007fffffffdfffffff7ffffffeafffffff1fffffff0",
            INIT_05 => X"ffffffeeffffffefffffffefffffffedffffffebfffffffbfffffff9fffffffd",
            INIT_06 => X"ffffffeffffffff1ffffffeefffffff4fffffffcfffffff800000002fffffffd",
            INIT_07 => X"ffffffecfffffffb0000000efffffff20000000fffffffea0000000b00000009",
            INIT_08 => X"00000009fffffff40000000d0000000f0000000700000012fffffff3ffffffeb",
            INIT_09 => X"0000000000000006ffffffe9ffffffebffffffe8fffffff9000000010000000d",
            INIT_0A => X"fffffff0fffffff30000000effffffed0000000c00000008ffffffe5ffffffe7",
            INIT_0B => X"fffffff80000000500000006ffffffe90000000affffffe7ffffffecfffffff3",
            INIT_0C => X"ffffffecfffffff9000000060000000100000004fffffff90000000b00000003",
            INIT_0D => X"0000000500000001fffffff00000000dffffffeefffffff7fffffff6ffffffed",
            INIT_0E => X"00000006fffffffcffffffe9fffffff300000000ffffffeffffffff4ffffffec",
            INIT_0F => X"ffffffeafffffffdffffffecffffffef0000000afffffffc00000005ffffffec",
            INIT_10 => X"00000009fffffff80000000afffffff3fffffffdffffffe9fffffffdfffffffe",
            INIT_11 => X"ffffffea00000001fffffffe00000007ffffffe70000000100000000ffffffe2",
            INIT_12 => X"0000000d00000003fffffff000000008ffffffeefffffffbfffffff5fffffff4",
            INIT_13 => X"0000000e0000000cfffffff00000000500000007ffffffeffffffffe0000000f",
            INIT_14 => X"0000000b0000000cfffffff0ffffffe4fffffffbfffffff3ffffffed00000015",
            INIT_15 => X"ffffffedfffffffbfffffff4ffffffe90000000d0000001200000005fffffff1",
            INIT_16 => X"fffffff00000000a0000000d0000000fffffffebffffffe80000000bfffffff0",
            INIT_17 => X"0000000d00000004fffffff3fffffffc000000070000000c0000000200000007",
            INIT_18 => X"000000150000000c000000040000001100000010ffffffea00000000fffffff0",
            INIT_19 => X"ffffffff0000000affffffe6fffffffcfffffff5ffffffe4fffffffdfffffff7",
            INIT_1A => X"fffffffb00000026000000050000000b000000320000001d00000019fffffffe",
            INIT_1B => X"fffffff900000000fffffffaffffffd5ffffffdf00000002000000240000001a",
            INIT_1C => X"fffffffcfffffff900000015fffffff3fffffffa000000080000001400000011",
            INIT_1D => X"0000000ffffffffeffffffe60000000a0000000f00000003000000130000002d",
            INIT_1E => X"ffffffe1fffffff7fffffff4ffffffc7fffffff1fffffffd00000001ffffffce",
            INIT_1F => X"fffffffdffffffcdffffffd300000000fffffffc0000000200000004ffffffed",
            INIT_20 => X"ffffffe7000000180000002500000005000000130000002bffffffe6fffffff5",
            INIT_21 => X"0000000700000005000000250000000fffffffec0000000b0000000600000000",
            INIT_22 => X"fffffffaffffffa2ffffffc200000009fffffffdffffffbfffffffe6fffffffb",
            INIT_23 => X"00000014fffffff80000000d0000001c0000001800000007fffffff7fffffff3",
            INIT_24 => X"fffffffffffffff2fffffff20000000a0000001f0000002d00000014fffffff6",
            INIT_25 => X"000000040000001a000000160000000100000000fffffff4ffffffde00000003",
            INIT_26 => X"ffffffc6ffffffc30000000d0000000f0000000c0000000f0000000b00000001",
            INIT_27 => X"00000008ffffffe900000004fffffff3fffffff4ffffffc2ffffffc00000000f",
            INIT_28 => X"0000000f0000000effffffe9ffffffc500000006fffffffbffffffd800000005",
            INIT_29 => X"ffffffcafffffff400000033fffffffa000000050000000b0000000000000006",
            INIT_2A => X"ffffffb4ffffffe7ffffffafffffffc500000000fffffffcffffffe000000013",
            INIT_2B => X"fffffffeffffffc6ffffffe300000020fffffff0fffffffafffffff1fffffff0",
            INIT_2C => X"ffffffd2ffffffe4fffffff3000000000000003b00000025ffffffcfffffffca",
            INIT_2D => X"00000009ffffffdc0000001d0000000bfffffff0ffffffc8ffffffc8fffffff7",
            INIT_2E => X"fffffffa0000001100000000ffffffd60000000800000000ffffffeffffffffe",
            INIT_2F => X"0000000c00000010fffffff0fffffff4ffffffe9ffffffd7ffffffe5fffffffa",
            INIT_30 => X"00000004ffffffeffffffffffffffff4fffffff300000006fffffffcffffffe4",
            INIT_31 => X"0000000affffffe8ffffffbc00000029ffffffeeffffffdc0000000bffffffe5",
            INIT_32 => X"fffffff80000000dffffffff000000170000000b0000000400000026fffffffa",
            INIT_33 => X"000000530000003400000001000000120000004d0000001900000017fffffff6",
            INIT_34 => X"0000000b00000000ffffffff0000000e00000000ffffffe700000010ffffffff",
            INIT_35 => X"ffffffe9ffffffdd0000003bfffffff7ffffffe7fffffff30000002bfffffff5",
            INIT_36 => X"fffffffa00000006ffffffe6ffffffebfffffff6ffffffe4ffffffe70000000e",
            INIT_37 => X"ffffffffffffffecffffffd0ffffffe4ffffffd4ffffffedffffffef0000000c",
            INIT_38 => X"000000310000002000000009fffffff6fffffffd00000012fffffff0ffffffdb",
            INIT_39 => X"00000012ffffffd2fffffff00000000cffffffe8ffffffe2ffffffe300000018",
            INIT_3A => X"00000029000000240000001efffffff00000001800000003fffffff100000023",
            INIT_3B => X"ffffffc6fffffff50000001cffffffb8fffffff500000028ffffffe300000000",
            INIT_3C => X"fffffffe00000000fffffff300000001000000080000000600000000ffffffff",
            INIT_3D => X"ffffffdc00000029000000380000000e00000013000000060000002300000007",
            INIT_3E => X"ffffffd9ffffffd1fffffffd00000019fffffffdfffffff80000001000000007",
            INIT_3F => X"ffffff99ffffffb7ffffffd8ffffffd0ffffffb9ffffffafffffffbefffffff2",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE29;


    MEM_IWGHT_LAYER1_INSTANCE30 : if BRAM_NAME = "iwght_layer1_instance30" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffb70000002600000046ffffffe7ffffff9dffffff86ffffffafffffffc5",
            INIT_01 => X"00000013000000280000003d00000001ffffffc0fffffff5fffffffbffffffef",
            INIT_02 => X"fffffff6fffffffc000000230000001000000034000000230000000000000000",
            INIT_03 => X"fffffff8fffffffd00000000fffffff8000000000000000500000003fffffffe",
            INIT_04 => X"0000001c0000000f00000022000000220000001f0000001e0000000f00000014",
            INIT_05 => X"0000000afffffff0ffffffd000000012ffffffdffffffffcffffffebffffffdc",
            INIT_06 => X"ffffffed0000000afffffffcfffffff3ffffffedffffffeb0000000affffffef",
            INIT_07 => X"fffffff2ffffffec0000000affffffe2fffffff1ffffffeafffffff9fffffff5",
            INIT_08 => X"00000001fffffffd00000001fffffffcfffffff800000001000000080000000c",
            INIT_09 => X"fffffffb00000012000000000000000bfffffff3000000020000001400000004",
            INIT_0A => X"00000009000000020000000a00000012000000140000001b00000015ffffffef",
            INIT_0B => X"0000001400000025000000180000001200000000000000370000004700000012",
            INIT_0C => X"000000100000002a000000270000002100000016000000150000000700000033",
            INIT_0D => X"0000001400000005ffffffedfffffffc00000003ffffffe5fffffff90000000c",
            INIT_0E => X"00000024ffffffe60000001000000028ffffffec000000180000000cffffffd3",
            INIT_0F => X"fffffffc000000050000000e0000000900000005fffffffefffffffefffffff5",
            INIT_10 => X"ffffffecffffffce00000014ffffffe7ffffffea00000018fffffffa00000016",
            INIT_11 => X"ffffffecfffffff3000000010000000dfffffff7fffffff90000001dfffffff9",
            INIT_12 => X"fffffff2fffffff8ffffffffffffffe4000000080000001300000026fffffffb",
            INIT_13 => X"0000000800000009fffffff900000014fffffff800000000fffffff6ffffffed",
            INIT_14 => X"fffffffefffffff90000001ffffffffffffffffffffffffbfffffff2fffffff1",
            INIT_15 => X"fffffffcfffffffc000000050000000fffffffe60000001b0000000effffffe8",
            INIT_16 => X"fffffff1000000080000001900000005ffffffdcfffffff1fffffffdffffffe1",
            INIT_17 => X"ffffffa3ffffffdeffffff94ffffff6effffff6dffffff95ffffffe1ffffff84",
            INIT_18 => X"0000000e0000003400000032000000080000001d000000310000000fffffff84",
            INIT_19 => X"0000001200000011fffffff8000000010000001dfffffffafffffff2fffffff8",
            INIT_1A => X"000000080000001afffffff0ffffffeefffffffafffffff1000000020000000c",
            INIT_1B => X"ffffffb5ffffffdcffffffe4ffffffd3000000290000002d0000002b00000024",
            INIT_1C => X"0000000dfffffffb00000000ffffffa9ffffffa1ffffffaaffffffa7ffffffa5",
            INIT_1D => X"ffffffe7ffffffe90000002e0000002700000030000000110000001700000006",
            INIT_1E => X"0000001c0000001cffffffff00000023fffffffdfffffff1fffffff3ffffffec",
            INIT_1F => X"fffffff3fffffffafffffff0fffffffe0000000cffffffeb000000140000001b",
            INIT_20 => X"0000001500000003000000150000001700000000ffffffff0000001800000009",
            INIT_21 => X"ffffffe900000015ffffffed0000000a0000000900000022000000150000000e",
            INIT_22 => X"0000004800000057000000270000000800000018000000190000000e00000002",
            INIT_23 => X"ffffffe6000000150000000e0000000100000022000000490000000b00000035",
            INIT_24 => X"00000023ffffffedfffffff100000018ffffffc7ffffffe4ffffffeb00000008",
            INIT_25 => X"fffffff2ffffffe4ffffffe20000002c0000000c0000001a0000004000000029",
            INIT_26 => X"000000320000000afffffff9000000260000003c0000000400000013fffffff6",
            INIT_27 => X"fffffff9ffffffd1ffffffc9ffffffd3fffffff200000008fffffff10000001f",
            INIT_28 => X"0000001bfffffff3ffffffe8ffffffeb00000004ffffffe40000000fffffffff",
            INIT_29 => X"00000002000000170000000600000021000000370000000a0000002b00000033",
            INIT_2A => X"00000001ffffffdf0000001dfffffffbfffffffd000000270000000800000006",
            INIT_2B => X"000000090000001500000006000000090000003600000014ffffffd500000004",
            INIT_2C => X"000000040000000a00000021fffffff1ffffffe100000018fffffff700000017",
            INIT_2D => X"ffffffd700000016fffffffeffffffdbffffffe60000000b0000000700000024",
            INIT_2E => X"0000002c00000038fffffffcffffffc9fffffff1ffffffeaffffffdcffffffe2",
            INIT_2F => X"ffffffe0ffffffe60000001200000012ffffffe3ffffffe300000006ffffffd1",
            INIT_30 => X"ffffffda00000016000000060000004300000007fffffff60000001efffffff9",
            INIT_31 => X"0000000700000004ffffffce00000014ffffffe5ffffffbe000000320000000d",
            INIT_32 => X"fffffff4ffffffc7ffffff81fffffff0fffffffdffffffd10000003a00000013",
            INIT_33 => X"00000008fffffff0fffffff1000000030000003c0000003700000018ffffffda",
            INIT_34 => X"fffffff7ffffffedffffffbffffffff3fffffff7ffffffe4ffffffc0ffffffdf",
            INIT_35 => X"ffffffebffffffe200000008fffffff0fffffff1ffffffc900000003ffffffd4",
            INIT_36 => X"ffffffd90000001100000000fffffffffffffffdffffffe70000000ffffffff3",
            INIT_37 => X"0000002dfffffff7fffffff80000002c00000009ffffffe00000002100000006",
            INIT_38 => X"00000019fffffff60000002400000002fffffff30000002f00000018ffffffed",
            INIT_39 => X"00000017ffffffc5ffffffe8fffffff70000000900000009ffffffe800000023",
            INIT_3A => X"fffffff10000000600000018000000080000000f00000008ffffffe50000000b",
            INIT_3B => X"ffffffd0fffffff500000014ffffffb3ffffffd0ffffffd0ffffffb5fffffff7",
            INIT_3C => X"fffffff3ffffffe3ffffffe8ffffffeaffffffe60000001500000011ffffffe0",
            INIT_3D => X"fffffff1fffffffcffffffea0000000b0000002e000000030000000c00000011",
            INIT_3E => X"fffffff8ffffffd00000001bfffffff0fffffff7000000070000001300000004",
            INIT_3F => X"fffffff70000002d0000001dfffffffefffffff2ffffffd100000013ffffffc1",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE30;


    MEM_IWGHT_LAYER1_INSTANCE31 : if BRAM_NAME = "iwght_layer1_instance31" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffffcffffffe2ffffffdc00000011ffffffe8fffffffb0000001600000015",
            INIT_01 => X"fffffffb00000001fffffff3fffffff4ffffffe5ffffffbaffffffeaffffffa8",
            INIT_02 => X"000000080000001300000009fffffff800000021fffffff6ffffffebffffffee",
            INIT_03 => X"fffffffafffffff2ffffffcf0000000200000003ffffffd70000002000000006",
            INIT_04 => X"00000002fffffff6fffffffd000000100000000000000000fffffff2fffffff7",
            INIT_05 => X"00000018fffffff400000023000000490000000f0000001400000026fffffff8",
            INIT_06 => X"fffffffaffffffed0000000000000020000000040000000e0000005900000033",
            INIT_07 => X"000000320000002800000017fffffffb00000013ffffffe9ffffffbf00000006",
            INIT_08 => X"ffffffc90000002d0000002afffffff00000003400000036000000110000003f",
            INIT_09 => X"0000001300000020fffffffcffffffe5ffffffe6ffffffe2fffffffefffffff3",
            INIT_0A => X"0000001efffffff900000000ffffffeaffffffd10000001affffffdbffffffd8",
            INIT_0B => X"fffffff900000013fffffff1fffffffa0000003e00000006ffffffd000000018",
            INIT_0C => X"ffffffe2ffffffeafffffff90000002400000038000000030000003b0000002e",
            INIT_0D => X"0000001f0000000affffffec00000013fffffff7fffffff8ffffffd400000004",
            INIT_0E => X"00000005ffffffe2ffffffc7ffffffd9ffffffffffffffe30000000a0000002a",
            INIT_0F => X"00000010fffffffaffffffd8ffffffeffffffffcffffffefffffffedffffffdb",
            INIT_10 => X"0000000cffffffca000000200000002d000000180000003b00000012ffffffe0",
            INIT_11 => X"ffffffef0000001a000000280000002600000019ffffffe5ffffffbe0000001b",
            INIT_12 => X"00000002000000010000000d000000020000000cffffffff000000040000000b",
            INIT_13 => X"00000025fffffff0fffffff0fffffff200000026ffffffd2ffffffe800000009",
            INIT_14 => X"0000003100000019fffffff0ffffff8800000006ffffffedffffff8400000021",
            INIT_15 => X"ffffffe3fffffff90000001affffffdcffffffe700000016fffffffd0000001d",
            INIT_16 => X"0000001b00000022000000280000005000000008ffffffdcffffffee00000003",
            INIT_17 => X"ffffffe6000000300000000f000000040000000500000017000000290000003e",
            INIT_18 => X"000000170000002e000000130000001afffffffbffffffe10000001b00000013",
            INIT_19 => X"ffffffffffffffdc0000000c00000026fffffffc000000100000001b00000014",
            INIT_1A => X"fffffff2fffffff6ffffffffffffffd9fffffff50000000fffffffd700000038",
            INIT_1B => X"0000000f0000001c0000002afffffff6fffffffbffffffd6000000160000002e",
            INIT_1C => X"fffffff200000017fffffffeffffffedffffffe000000018000000250000001a",
            INIT_1D => X"ffffffddffffffeffffffff1ffffffe600000017ffffffd7ffffffdf00000008",
            INIT_1E => X"0000000e00000024ffffffde0000001f0000001affffffc300000004fffffff6",
            INIT_1F => X"ffffffec0000002900000002ffffffd5ffffffe500000012ffffffdeffffffe8",
            INIT_20 => X"ffffffe3fffffff6fffffffdffffffe3ffffffffffffffeaffffffe9ffffffe2",
            INIT_21 => X"ffffffc9ffffffd800000004ffffffefffffffd0fffffffefffffffeffffffec",
            INIT_22 => X"ffffffccffffffb3000000220000001600000007fffffffb000000000000002f",
            INIT_23 => X"ffffffff00000005fffffff100000002fffffff7ffffffe50000000600000020",
            INIT_24 => X"00000018fffffff9000000090000001900000019000000090000002600000008",
            INIT_25 => X"00000000ffffffd9ffffffd6ffffffda0000002600000011ffffffe4ffffffcd",
            INIT_26 => X"000000120000000b0000000affffffc3000000060000001cffffffdc00000016",
            INIT_27 => X"000000130000000600000033ffffffd7fffffff80000002900000017fffffff7",
            INIT_28 => X"0000000efffffff90000000e000000220000000c000000100000000300000014",
            INIT_29 => X"ffffffe4ffffffdc0000001ffffffff400000002000000000000001700000002",
            INIT_2A => X"fffffffc0000003800000017fffffffb0000002e0000003d00000022ffffffe2",
            INIT_2B => X"000000060000003dfffffff40000001d000000370000000afffffff0fffffffc",
            INIT_2C => X"0000003cffffffe4ffffffe4fffffff1ffffffd60000000700000040ffffffe0",
            INIT_2D => X"0000001700000000ffffffd8fffffffdffffffcf00000043ffffffbbffffffe9",
            INIT_2E => X"0000000400000000000000290000000400000038000000130000000b00000010",
            INIT_2F => X"ffffffd100000009ffffffdd0000001a0000001ffffffff6ffffffed0000002c",
            INIT_30 => X"fffffffbffffffceffffffefffffffcffffffff3ffffffbbffffffcaffffffe6",
            INIT_31 => X"ffffffd900000002fffffff60000000affffffecffffffe9fffffff80000000f",
            INIT_32 => X"00000001000000150000001a0000000b0000000600000000fffffff1ffffffe9",
            INIT_33 => X"0000000d00000016ffffffe90000000a000000070000000c000000130000001c",
            INIT_34 => X"00000003000000000000001a00000009fffffff300000009ffffffe0ffffffcd",
            INIT_35 => X"ffffffdb00000012fffffffbffffffeb000000010000000a0000001700000037",
            INIT_36 => X"fffffffa000000030000001f0000002a0000000a0000001500000006ffffffeb",
            INIT_37 => X"ffffffe4ffffffc6fffffff30000000800000022fffffff90000000fffffffe6",
            INIT_38 => X"ffffffd9fffffff600000017ffffffe90000000400000005fffffff700000018",
            INIT_39 => X"000000090000002000000013fffffffa00000006ffffffe3fffffffcffffffe6",
            INIT_3A => X"ffffffebfffffffcfffffff9000000200000000bfffffff40000000600000000",
            INIT_3B => X"0000000c0000002b0000001b000000010000002e0000000effffffe1ffffffef",
            INIT_3C => X"000000280000000600000050000000100000002a00000047fffffffe0000000d",
            INIT_3D => X"ffffffd8ffffffc8ffffffe9ffffffdbffffffde000000540000006b0000004b",
            INIT_3E => X"ffffffedffffffcc00000012fffffff9fffffff1fffffff2ffffffc7ffffffe6",
            INIT_3F => X"ffffffceffffffd70000000800000009fffffff7ffffffc3ffffffd300000009",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE31;


    MEM_IWGHT_LAYER1_INSTANCE32 : if BRAM_NAME = "iwght_layer1_instance32" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffffe00000007fffffffaffffffe8ffffffe0ffffffd0fffffff0ffffffef",
            INIT_01 => X"ffffffe4fffffff3000000060000001f00000017ffffffecfffffff800000016",
            INIT_02 => X"ffffffe3ffffffe90000001500000010fffffffb00000018000000090000000c",
            INIT_03 => X"00000005ffffffd7ffffffe5000000300000001cffffffe1ffffffe3ffffffeb",
            INIT_04 => X"fffffff3ffffffdd00000024fffffffefffffff6000000020000000e0000000b",
            INIT_05 => X"fffffffe000000160000000d00000003ffffffeeffffffecfffffff9ffffffd1",
            INIT_06 => X"00000005ffffffe800000013ffffffecffffffe20000000b0000002700000031",
            INIT_07 => X"00000033fffffffd000000230000000e0000001d0000001bfffffff7ffffffe9",
            INIT_08 => X"ffffffe900000000ffffffea000000030000001c0000000affffffdbfffffff0",
            INIT_09 => X"ffffffd2fffffffa0000003c0000003700000023000000220000002200000001",
            INIT_0A => X"00000018fffffff7ffffffd6ffffffc1ffffffe000000002ffffffceffffffc2",
            INIT_0B => X"0000002000000016000000410000000400000000fffffffe0000000900000000",
            INIT_0C => X"0000001dfffffff70000000a00000010fffffff7ffffffec0000000dfffffff9",
            INIT_0D => X"00000013000000170000001a00000019000000260000001b0000000d00000018",
            INIT_0E => X"ffffffa4000000280000002dffffffc2ffffffee000000420000002100000011",
            INIT_0F => X"ffffffc0ffffffefffffffd0ffffffe200000004fffffffdffffffff00000028",
            INIT_10 => X"00000036ffffffbfffffffb60000003fffffffaeffffffe6fffffff5ffffff8f",
            INIT_11 => X"0000001dffffffecfffffff7ffffffac0000000900000055ffffffbeffffffb7",
            INIT_12 => X"000000200000000a00000000fffffff2ffffffea000000090000002200000006",
            INIT_13 => X"00000024000000130000000e000000070000000affffffff00000006fffffff2",
            INIT_14 => X"000000050000001e000000190000000d00000009000000230000003500000040",
            INIT_15 => X"ffffffe400000002ffffffcd00000000ffffffedffffffbcffffffeefffffff2",
            INIT_16 => X"fffffff8fffffffc00000027ffffffd4ffffffe800000008ffffffe8ffffffdc",
            INIT_17 => X"fffffffb000000300000001effffffe7ffffffee00000002fffffffb00000003",
            INIT_18 => X"ffffffe1ffffffffffffffe3fffffff9ffffffe7000000120000000e0000000b",
            INIT_19 => X"ffffffec0000000ffffffffb000000000000001100000001ffffffce00000000",
            INIT_1A => X"0000000e00000036ffffffe000000013ffffffeaffffffc10000002cfffffff5",
            INIT_1B => X"0000000cfffffff50000000c00000012fffffffe0000002c0000003b00000001",
            INIT_1C => X"0000000dfffffffc00000003ffffffe100000028fffffffcffffffe1fffffffb",
            INIT_1D => X"fffffff7ffffffeaffffffc20000000b0000001affffffec0000000a0000000e",
            INIT_1E => X"00000004000000030000001e000000420000001e0000003200000028ffffffce",
            INIT_1F => X"fffffff70000001400000029fffffff80000000e00000010ffffffcd00000015",
            INIT_20 => X"0000000b0000000bfffffff8ffffff97ffffffd0ffffffeefffffff100000018",
            INIT_21 => X"0000001bffffffe800000014000000030000001b0000000a00000009ffffffe5",
            INIT_22 => X"0000000000000004000000130000000f0000001500000000ffffffe40000001c",
            INIT_23 => X"0000001300000021000000130000001e00000000fffffff70000003a00000025",
            INIT_24 => X"000000090000002200000006ffffffe3ffffffe5000000140000000600000002",
            INIT_25 => X"ffffffed000000020000000bffffffdcfffffff0ffffffdafffffffeffffffeb",
            INIT_26 => X"0000001600000001ffffffe100000002fffffffefffffff4ffffffdbffffffd2",
            INIT_27 => X"ffffffc400000038ffffff8cffffff9d00000003ffffffaeffffff9900000028",
            INIT_28 => X"fffffffd0000000e000000020000001c000000020000002600000012ffffff77",
            INIT_29 => X"0000000e00000016ffffffff0000000a00000000ffffffed0000001f00000015",
            INIT_2A => X"ffffffeaffffffd300000025fffffff9fffffffc0000000e000000190000001a",
            INIT_2B => X"ffffffc6ffffffbcffffff91ffffffdb00000000fffffff20000001b00000003",
            INIT_2C => X"ffffffedffffffe2ffffffcfffffffb7ffffffcd00000006ffffffb1ffffff9c",
            INIT_2D => X"000000000000001000000003fffffffeffffffecfffffffc0000000affffffc8",
            INIT_2E => X"0000000400000018fffffffeffffffee000000160000002b0000000200000011",
            INIT_2F => X"00000001000000070000000e0000001c0000001000000006ffffffe5ffffffea",
            INIT_30 => X"ffffffee00000009ffffffff00000005fffffff30000000e0000001f0000000c",
            INIT_31 => X"fffffff1fffffff80000002500000047fffffff20000003100000018fffffff9",
            INIT_32 => X"ffffffefffffffa6fffffff3ffffffe2ffffffc2fffffff1000000120000001f",
            INIT_33 => X"0000003100000041000000280000003b00000017ffffffd9ffffffd600000017",
            INIT_34 => X"ffffffd9ffffffdcffffffa7ffffffc9ffffffff00000028000000380000003d",
            INIT_35 => X"fffffff2ffffffcdffffffbdffffffe7fffffff2fffffff0ffffffd9ffffffb3",
            INIT_36 => X"0000001afffffff4ffffffdafffffffe0000002cffffffdaffffffb1fffffff3",
            INIT_37 => X"00000012ffffffdd00000004000000000000002f0000003e0000003a00000045",
            INIT_38 => X"00000015ffffffecffffffd800000015fffffffb00000011000000070000000c",
            INIT_39 => X"000000180000002d000000130000002200000052fffffff700000048fffffffd",
            INIT_3A => X"fffffffbfffffff800000001fffffff5fffffff6ffffffdc00000001fffffff3",
            INIT_3B => X"000000110000000c000000210000001e000000160000000f0000000300000015",
            INIT_3C => X"ffffffbbffffffbbffffffbfffffff96ffffffd600000018000000140000000d",
            INIT_3D => X"00000014fffffffffffffff7000000140000000ffffffff8fffffffa00000000",
            INIT_3E => X"ffffffd20000001200000006fffffff1ffffffedffffffef0000001000000004",
            INIT_3F => X"ffffffbbffffffe3ffffffd3ffffffdbffffffabffffffe50000001500000023",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE32;


    MEM_IWGHT_LAYER1_INSTANCE33 : if BRAM_NAME = "iwght_layer1_instance33" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000041ffffffff000000130000001200000022ffffffe0ffffffd7ffffffde",
            INIT_01 => X"ffffffe6ffffffe600000024fffffff1fffffff00000001a00000004fffffff2",
            INIT_02 => X"0000001bffffffe6ffffffdb00000004fffffffa0000002c0000000500000009",
            INIT_03 => X"0000000c00000002000000110000000700000010000000220000001700000010",
            INIT_04 => X"fffffffd0000001100000046ffffffd700000017000000230000000f00000009",
            INIT_05 => X"0000001200000009000000260000000afffffff4fffffff1fffffff70000001e",
            INIT_06 => X"ffffffe5fffffff7fffffff10000000a00000010fffffffa000000070000000b",
            INIT_07 => X"0000002000000003fffffffc000000300000002e00000002ffffffe9ffffffe8",
            INIT_08 => X"00000011fffffffd0000001a0000000d00000025000000110000001000000004",
            INIT_09 => X"fffffffefffffff600000003000000010000000a000000010000000c00000015",
            INIT_0A => X"ffffffe00000001b0000000b000000290000001e0000001f0000001800000002",
            INIT_0B => X"0000004500000035fffffff50000001f0000002900000027000000160000001d",
            INIT_0C => X"ffffffd8ffffffefffffffeffffffff9ffffffe500000017ffffffeb0000001c",
            INIT_0D => X"ffffffe80000000a00000010ffffffeb000000060000000f00000023ffffffff",
            INIT_0E => X"00000007ffffffe400000009fffffff90000000000000004fffffff80000001a",
            INIT_0F => X"000000240000003c0000000a0000001dfffffffcffffffe9fffffff300000024",
            INIT_10 => X"ffffffceffffffc2ffffffedffffffe10000001100000014fffffffcfffffff1",
            INIT_11 => X"00000006fffffff0ffffffddffffffc9ffffffd7fffffff8ffffffb7ffffffd7",
            INIT_12 => X"0000001dfffffff90000002a000000050000002500000003ffffffdbffffffee",
            INIT_13 => X"0000002d0000001d00000049fffffff90000001a0000002600000015fffffff7",
            INIT_14 => X"00000010000000180000000ffffffff10000000300000017000000080000000b",
            INIT_15 => X"0000002d0000000e0000001c00000025ffffffe20000000600000014fffffff8",
            INIT_16 => X"0000000000000009ffffffeaffffffd90000000c00000003000000190000002a",
            INIT_17 => X"ffffffecffffffe4ffffffafffffffc3ffffffe9ffffffe60000000cffffffe4",
            INIT_18 => X"000000020000000a0000002a0000004fffffffbdffffffbbffffffc6ffffffbe",
            INIT_19 => X"fffffffffffffff3fffffff60000000600000012ffffffe50000000a0000003e",
            INIT_1A => X"0000001400000018ffffffee00000008fffffff00000001400000021fffffff9",
            INIT_1B => X"00000017fffffff9ffffffceffffffc6fffffff1fffffff2fffffffb0000000d",
            INIT_1C => X"000000290000000b0000000400000000fffffff20000000c0000001100000001",
            INIT_1D => X"00000000000000080000001cfffffffa00000005000000050000000500000003",
            INIT_1E => X"ffffff92000000020000001c000000160000001c0000002c0000002800000011",
            INIT_1F => X"0000002a0000000800000020000000080000001b00000015ffffffc6ffffffb7",
            INIT_20 => X"fffffff200000009ffffffcaffffffd400000001ffffffef0000000600000004",
            INIT_21 => X"00000013fffffff5fffffff6fffffff4ffffffb9ffffffd8ffffffefffffffc9",
            INIT_22 => X"00000010000000160000000f00000003ffffffe3ffffffedfffffffdfffffffe",
            INIT_23 => X"fffffffcffffffe7ffffffe4fffffffefffffffbffffffe50000000000000005",
            INIT_24 => X"0000000cffffffeaffffffe5fffffffbfffffff70000000d0000000800000000",
            INIT_25 => X"ffffffd5fffffff5fffffffeffffffff000000150000001fffffffd500000016",
            INIT_26 => X"ffffff8effffffc2ffffffabffffffbbffffffbffffffffeffffffe0ffffffd4",
            INIT_27 => X"ffffffb600000000fffffff00000000f0000001d0000002200000019ffffffab",
            INIT_28 => X"ffffffeefffffffb00000040ffffffef0000003f00000031ffffffc3ffffffb8",
            INIT_29 => X"000000160000001300000001fffffffefffffff60000000a0000002e0000001c",
            INIT_2A => X"0000002efffffff400000002000000010000001000000029fffffffc00000001",
            INIT_2B => X"000000050000000a00000007000000240000000d000000380000000100000022",
            INIT_2C => X"0000003dffffffe90000002a000000050000001e000000180000001f00000012",
            INIT_2D => X"fffffff5ffffff9cffffffcbffffff80ffffffe0ffffffffffffffed00000019",
            INIT_2E => X"0000001affffffd1ffffffd800000012fffffffbffffffeb00000010ffffffff",
            INIT_2F => X"ffffffd0ffffff9affffffb9ffffffbbffffffceffffffebffffffd1ffffffe1",
            INIT_30 => X"00000018000000170000001200000023000000230000002700000019ffffffc2",
            INIT_31 => X"fffffffcfffffff30000001e0000001e00000046000000440000000efffffffd",
            INIT_32 => X"ffffffd3ffffffd3fffffffeffffffe3fffffffaffffffd7ffffffe9ffffffcc",
            INIT_33 => X"ffffffedffffffd6ffffffcc0000001affffffd1ffffffd7ffffffebfffffffa",
            INIT_34 => X"00000021ffffffccffffffdaffffffebffffffbbffffffedffffffefffffffed",
            INIT_35 => X"000000170000000affffffb1ffffff90ffffffd3ffffffa6ffffff7bffffffa5",
            INIT_36 => X"00000016000000090000002500000018000000080000000d0000002300000000",
            INIT_37 => X"ffffffb9ffffffe6ffffffbf0000002900000004fffffff5000000040000003d",
            INIT_38 => X"00000006fffffffdffffffef0000001400000010fffffff4000000040000000d",
            INIT_39 => X"00000006ffffffe40000000300000009000000000000000b000000100000000c",
            INIT_3A => X"00000010000000100000000ffffffffe00000011000000030000002400000018",
            INIT_3B => X"ffffffeaffffffb2ffffffefffffffe0ffffffc5000000200000001d00000011",
            INIT_3C => X"00000022fffffff4fffffff600000006ffffffeaffffffe2ffffffcfffffffde",
            INIT_3D => X"0000000fffffffdc000000040000002d0000004800000001000000180000002b",
            INIT_3E => X"fffffff40000001dffffffe50000001800000008fffffff8fffffffa00000013",
            INIT_3F => X"ffffffecffffffeffffffff2fffffff6ffffffe0fffffff4fffffffefffffffa",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE33;


    MEM_IWGHT_LAYER1_INSTANCE34 : if BRAM_NAME = "iwght_layer1_instance34" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002d0000002b000000070000000bffffffff00000004ffffffedfffffff3",
            INIT_01 => X"fffffffc00000015ffffffdd0000001e00000047000000080000001a0000000c",
            INIT_02 => X"ffffffdc00000021ffffffefffffffdf00000008fffffffb000000160000000c",
            INIT_03 => X"ffffffedffffffed0000000ffffffff900000018fffffffe0000001cffffffd8",
            INIT_04 => X"ffffffcfffffffd5ffffffe1ffffffe8ffffffe7fffffffaffffffed0000002b",
            INIT_05 => X"fffffff900000009fffffff400000004ffffffcdffffffe1ffffffd1fffffff0",
            INIT_06 => X"000000000000001500000007ffffffeafffffffa0000000d00000009fffffffe",
            INIT_07 => X"ffffffeefffffff70000001900000020ffffffeb000000340000001e00000002",
            INIT_08 => X"00000004ffffffcc000000000000001affffffeffffffffa0000000cffffffe6",
            INIT_09 => X"0000001d00000004ffffffed000000130000002b0000001b000000000000001e",
            INIT_0A => X"ffffff97ffffffb9fffffff3ffffffcaffffffe0ffffffbeffffffd3ffffffaf",
            INIT_0B => X"fffffff0ffffffdaffffffdbffffffe50000000600000001fffffff4ffffffa8",
            INIT_0C => X"ffffffdaffffffd0ffffffc60000002300000006fffffffcffffffdeffffffd8",
            INIT_0D => X"0000001d0000001d000000130000001b0000001affffffebffffffdfffffff8d",
            INIT_0E => X"0000001afffffffa0000000a0000000b000000230000002e00000010fffffffc",
            INIT_0F => X"fffffff8000000000000001d00000021ffffffee000000040000002200000012",
            INIT_10 => X"ffffffe5ffffffce0000000a0000000800000019000000000000001000000008",
            INIT_11 => X"00000006ffffffd0ffffffc3ffffffc8ffffffb2ffffffe3ffffffcbffffffec",
            INIT_12 => X"fffffff8fffffff300000006ffffffeafffffff4000000160000002200000013",
            INIT_13 => X"ffffffdd00000006ffffffaeffffffd7ffffffceffffffdafffffff5ffffffcf",
            INIT_14 => X"0000001d0000000f000000160000001b0000002c000000100000000dffffffd9",
            INIT_15 => X"000000090000000ffffffff70000001bfffffffc000000070000001b00000014",
            INIT_16 => X"000000000000001500000009ffffffe80000000800000012ffffffe5ffffffd6",
            INIT_17 => X"ffffffe40000001300000002fffffff900000006000000000000000100000003",
            INIT_18 => X"0000002b0000001b00000000ffffffd800000000fffffff8fffffffdfffffff1",
            INIT_19 => X"fffffffe00000002ffffffddffffffceffffffe2ffffffdaffffffc5ffffffde",
            INIT_1A => X"00000012fffffffbffffffed000000010000000a000000040000000300000016",
            INIT_1B => X"ffffffecffffffdeffffffcafffffffe00000009ffffffe9000000010000000f",
            INIT_1C => X"0000000000000000fffffff9ffffffecfffffff7000000050000000e00000008",
            INIT_1D => X"ffffffbf0000001f00000021ffffffdfffffffdfffffffeb0000001bffffffef",
            INIT_1E => X"00000019000000100000000c00000000fffffffb00000019ffffffebffffffcf",
            INIT_1F => X"fffffffb00000002ffffffffffffffe3ffffffe6ffffffbbfffffff8ffffffd6",
            INIT_20 => X"fffffff8fffffff3fffffff0fffffff400000012fffffffbffffffe500000020",
            INIT_21 => X"fffffffaffffffcfffffffdafffffff4ffffffd60000000dffffffe1fffffffa",
            INIT_22 => X"00000002ffffffeefffffff20000000b00000029fffffffdffffffcd00000006",
            INIT_23 => X"00000000fffffff1fffffffa00000007ffffffc60000001f0000000d0000000b",
            INIT_24 => X"00000037fffffffbfffffff70000002a00000010ffffffe40000001f0000001f",
            INIT_25 => X"ffffffe2ffffffd500000000fffffffefffffff30000000800000011ffffffd9",
            INIT_26 => X"0000002affffffc7ffffffe900000015ffffffc0fffffff100000016ffffffed",
            INIT_27 => X"0000004e00000003ffffffd90000002c00000044fffffff8fffffff7fffffff0",
            INIT_28 => X"00000007000000270000000f000000050000000effffffdcfffffff8ffffffb6",
            INIT_29 => X"00000023ffffffefffffffdb0000001cffffffeb000000120000002900000047",
            INIT_2A => X"ffffffe6000000190000000f0000000c0000002500000036ffffffdbfffffff3",
            INIT_2B => X"fffffff7ffffffcf00000013fffffff6fffffffb000000050000000bffffffd4",
            INIT_2C => X"0000003a00000003000000270000002ffffffff9ffffffdaffffffff00000016",
            INIT_2D => X"00000006fffffffc00000040ffffffd8ffffffe70000003cffffffdcffffffd0",
            INIT_2E => X"ffffffecffffffbefffffff90000002affffffd0ffffffe00000001cfffffff4",
            INIT_2F => X"00000015ffffffd60000001affffffe7ffffffeeffffffeffffffff500000023",
            INIT_30 => X"ffffffcc00000007fffffffdfffffffe00000006000000310000000800000032",
            INIT_31 => X"ffffffeefffffff00000000bffffffd7fffffff400000002fffffff80000002a",
            INIT_32 => X"0000001500000016fffffff8ffffffddffffffed00000001fffffff2fffffffe",
            INIT_33 => X"00000020ffffffefffffffe20000002700000003ffffffeb0000000400000002",
            INIT_34 => X"ffffffe2fffffffafffffffdfffffff8000000100000001dffffffe0ffffffef",
            INIT_35 => X"ffffffe3fffffff70000001900000022ffffffc0ffffffe800000006ffffffbe",
            INIT_36 => X"00000011fffffff5ffffffee00000055ffffffedffffffc10000004000000019",
            INIT_37 => X"0000001e000000060000005e00000052000000500000001b0000002e00000042",
            INIT_38 => X"ffffffc80000001600000013ffffffdaffffffe10000001bffffffe200000023",
            INIT_39 => X"ffffffceffffffed0000000dffffffde000000010000001a0000002800000003",
            INIT_3A => X"ffffffeafffffff5fffffffdffffffe300000000fffffff70000001c0000002d",
            INIT_3B => X"0000001e0000000500000027000000170000001d0000001c0000000affffffe3",
            INIT_3C => X"ffffffe600000008000000050000001d0000001200000018000000210000001f",
            INIT_3D => X"ffffffc3ffffffca000000500000003b00000017000000320000003e00000029",
            INIT_3E => X"00000008fffffffefffffff8ffffffeffffffffaffffffd3ffffffdc00000008",
            INIT_3F => X"000000110000002200000054ffffffd6ffffffef00000036ffffffcaffffffda",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE34;


    MEM_IWGHT_LAYER1_INSTANCE35 : if BRAM_NAME = "iwght_layer1_instance35" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff000000004ffffffe5fffffffefffffffffffffff2fffffffe00000006",
            INIT_01 => X"0000001d0000001d00000005000000250000002e0000002900000004fffffff3",
            INIT_02 => X"ffffff8fffffff89ffffffbbffffffb5ffffffa7ffffffb40000000700000029",
            INIT_03 => X"00000037000000280000002f00000037fffffff8ffffffa1ffffffbeffffff93",
            INIT_04 => X"ffffffb3ffffffaeffffffb7ffffffad000000150000002900000027ffffffff",
            INIT_05 => X"000000180000002700000000ffffffcaffffffafffffffa9ffffffcfffffff96",
            INIT_06 => X"000000280000000e0000001000000012ffffffd7000000340000002b00000002",
            INIT_07 => X"00000026fffffff6ffffffdcffffffc5fffffff3ffffffedffffffec00000032",
            INIT_08 => X"fffffffc000000020000000200000007fffffff50000000dffffffef0000001c",
            INIT_09 => X"fffffff5ffffffe40000001afffffff500000004fffffff4ffffffdaffffffe7",
            INIT_0A => X"00000000fffffff7ffffffd2fffffff700000017ffffffeffffffff0ffffffc7",
            INIT_0B => X"0000001e00000000fffffff9fffffffeffffffe9fffffff90000000000000009",
            INIT_0C => X"0000001c00000004ffffffe5fffffff1ffffffecffffffcaffffffeeffffffdd",
            INIT_0D => X"000000020000001efffffffe0000001d00000014ffffffdafffffff700000009",
            INIT_0E => X"00000007000000060000000f0000000a00000000ffffffec0000002a00000028",
            INIT_0F => X"00000019000000110000001a0000000e0000000ffffffff1ffffffeb0000000e",
            INIT_10 => X"ffffffffffffffeaffffffddffffffe2000000190000001a0000000700000007",
            INIT_11 => X"000000110000000f0000000e0000000a00000012fffffffe0000000000000006",
            INIT_12 => X"0000000e00000021fffffffa000000000000001600000007ffffffe4ffffffe4",
            INIT_13 => X"0000000b0000000f000000050000000c00000027000000160000002600000019",
            INIT_14 => X"ffffffacffffffd80000001effffffd2ffffffee00000015fffffff3fffffff7",
            INIT_15 => X"00000017000000020000002b0000001efffffff6ffffffd6ffffffe30000000d",
            INIT_16 => X"fffffffdfffffff80000000bfffffffe0000000bfffffff9fffffff700000027",
            INIT_17 => X"0000000f000000280000001e0000000000000005ffffffeeffffffebfffffffd",
            INIT_18 => X"00000023000000100000001f0000001a0000001300000017fffffffd0000000f",
            INIT_19 => X"0000001700000000fffffffbfffffff90000000cfffffffd0000000700000029",
            INIT_1A => X"fffffff2ffffffc7ffffffc400000016000000290000000a0000001b00000009",
            INIT_1B => X"ffffffe3ffffffb2ffffffd5ffffffe3ffffffa0ffffff99ffffffc5ffffff77",
            INIT_1C => X"0000001efffffffaffffffe5fffffff90000000900000007fffffff20000000b",
            INIT_1D => X"fffffff3fffffff5fffffff1000000080000000afffffffe0000000800000005",
            INIT_1E => X"00000023fffffff20000000a000000030000001300000013fffffff1fffffffb",
            INIT_1F => X"00000018fffffffc00000017ffffffeb0000000200000006ffffffde00000029",
            INIT_20 => X"fffffffa00000007fffffff5ffffffca0000000bfffffff1ffffffc6fffffff4",
            INIT_21 => X"0000000800000002ffffffecffffffdeffffffedfffffff9ffffffe3fffffffe",
            INIT_22 => X"00000011fffffffdffffffe4ffffffe700000000000000080000000d00000007",
            INIT_23 => X"0000000500000024000000200000001d0000001b000000190000000700000013",
            INIT_24 => X"000000030000000900000012fffffffbffffffecffffffe5fffffff3fffffffd",
            INIT_25 => X"0000004600000018000000260000001c00000000000000180000000f00000005",
            INIT_26 => X"fffffffdffffffc70000000dffffffff00000007000000220000002300000047",
            INIT_27 => X"ffffffe5ffffffe60000000ffffffffcfffffffe00000002ffffffd7ffffffeb",
            INIT_28 => X"ffffff9600000000ffffffe7ffffffff0000000bffffffc7ffffff97fffffffc",
            INIT_29 => X"00000013000000230000000effffffe7ffffffcfffffffa0ffffffd0ffffffbc",
            INIT_2A => X"0000000800000027000000230000002500000041fffffff10000000a0000000e",
            INIT_2B => X"00000006fffffff5ffffffeaffffffcaffffffef00000013ffffffe700000027",
            INIT_2C => X"fffffff00000000affffffecfffffffafffffff2fffffff80000000500000004",
            INIT_2D => X"ffffffee000000090000002400000015ffffffffffffffed00000004ffffffff",
            INIT_2E => X"fffffff9000000170000001300000005000000040000001b0000000a0000001d",
            INIT_2F => X"000000230000000b0000000bfffffffc0000000600000000fffffff300000020",
            INIT_30 => X"ffffffd2fffffff7fffffffcffffffe2ffffffd900000005000000160000000b",
            INIT_31 => X"ffffffe30000000cfffffff3ffffffeffffffff40000000400000006ffffffee",
            INIT_32 => X"fffffffc00000021ffffffdafffffff7ffffffee0000000cffffffe4ffffffe8",
            INIT_33 => X"ffffffed000000030000001b0000003a000000000000000f0000002cfffffff4",
            INIT_34 => X"00000009ffffffff00000004fffffffefffffffdffffffdfffffffeafffffffd",
            INIT_35 => X"0000000c0000000a00000015ffffffeffffffff9ffffffecfffffff5fffffffc",
            INIT_36 => X"0000000efffffff800000045000000460000001b000000390000001e00000009",
            INIT_37 => X"ffffffe4000000010000000b0000000600000017000000230000000b0000003f",
            INIT_38 => X"ffffffb0ffffffd4fffffffcffffffe300000026000000460000000ffffffff9",
            INIT_39 => X"fffffff400000008000000120000000800000039ffffffcaffffffd7ffffffd4",
            INIT_3A => X"fffffffd00000004fffffff60000000cffffffedffffffedffffffee00000003",
            INIT_3B => X"0000000c000000270000001bffffffc7ffffffb8ffffffe8ffffffc1ffffffce",
            INIT_3C => X"0000001e00000004ffffffdcfffffff9ffffffe9ffffffe2ffffffe5fffffff4",
            INIT_3D => X"0000000bffffffd60000000dffffffe6ffffffff0000000effffffe800000014",
            INIT_3E => X"ffffffeafffffffaffffffed0000001000000018fffffff60000001200000010",
            INIT_3F => X"ffffffca0000000bffffffdeffffffacffffffcbffffffc6ffffffc4fffffff4",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE35;


    MEM_IWGHT_LAYER1_INSTANCE36 : if BRAM_NAME = "iwght_layer1_instance36" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffed0000001b000000220000001200000015000000060000001fffffff9d",
            INIT_01 => X"0000001600000028fffffff20000000c00000008fffffff80000001200000014",
            INIT_02 => X"fffffffdfffffff900000005fffffffa000000060000002d00000016ffffffef",
            INIT_03 => X"ffffffd7ffffffec00000002fffffff1ffffffe5ffffffeb00000025fffffff3",
            INIT_04 => X"ffffffe3ffffffd5ffffffe000000016ffffffc4ffffffadffffffe4ffffffd5",
            INIT_05 => X"000000040000002d00000013fffffffe0000001fffffffd3ffffffedffffffef",
            INIT_06 => X"00000002ffffffd5ffffffd4fffffff4ffffffd1ffffffe300000000fffffff7",
            INIT_07 => X"0000001f0000000ffffffff0fffffff90000000cffffffd6000000000000000b",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE36;


    MEM_IWGHT_LAYER2_INSTANCE0 : if BRAM_NAME = "iwght_layer2_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00002a0cffffb7b00000300100000073fffff170fffffe76fffff509fffff8e0",
            INIT_01 => X"000016b300000b7a000015ce00000dc2ffffe731ffffe7ef000006a400000521",
            INIT_02 => X"00000a63fffff8a10000232300000bd500002342fffff083fffffd10fffff645",
            INIT_03 => X"00002a49000018e6ffffee1e000007d6ffffddff000017c20000027000000f0a",
            INIT_04 => X"fffffff7ffffffedfffffffaffffffed00000000fffffff2fffffff500000006",
            INIT_05 => X"ffffffdd00000017fffffffdffffffcfffffffd7ffffffef00000005fffffff2",
            INIT_06 => X"ffffffdcffffffebffffffeb00000005ffffffe4fffffffdffffffe900000010",
            INIT_07 => X"fffffff50000000400000008ffffffd1ffffffe2ffffffdc00000002fffffff5",
            INIT_08 => X"0000000cfffffff7ffffffdeffffffeaffffffdcffffffdfffffffd3fffffffe",
            INIT_09 => X"0000001300000009000000140000001cffffffe800000000fffffffbffffffff",
            INIT_0A => X"fffffff5fffffffc00000015fffffff900000004fffffff6ffffffea00000000",
            INIT_0B => X"ffffffeafffffffafffffffcffffffec0000001300000016fffffffaffffffe4",
            INIT_0C => X"000000040000001afffffff20000001cffffffe4ffffffea00000009fffffff9",
            INIT_0D => X"00000015fffffff5ffffffe2ffffffe4fffffff4fffffff300000007ffffffed",
            INIT_0E => X"ffffffd9ffffffe2fffffff1ffffffdb0000000ffffffff000000000fffffff8",
            INIT_0F => X"ffffffdaffffffefffffffdaffffffe2fffffff5fffffff4ffffffd7ffffffd4",
            INIT_10 => X"0000000cffffffe80000001600000000ffffffe4ffffffd0ffffffe3fffffff8",
            INIT_11 => X"000000030000000efffffff200000005ffffffddffffffd0ffffffe6fffffff9",
            INIT_12 => X"0000000d00000017fffffffaffffffe0ffffffdbffffffe3ffffffedfffffff3",
            INIT_13 => X"ffffffdefffffffbffffffe500000013ffffffe700000000ffffffef00000006",
            INIT_14 => X"0000000d0000000a0000000500000012ffffffeaffffffeaffffffe600000004",
            INIT_15 => X"fffffff5ffffffe0ffffffdaffffffdc00000000fffffffcfffffffafffffff9",
            INIT_16 => X"ffffffeefffffff50000001e0000000a000000090000002c0000001500000014",
            INIT_17 => X"ffffffed00000013fffffffe0000000affffffff00000016000000160000000e",
            INIT_18 => X"ffffffe800000000ffffffeafffffffd0000000b000000080000001400000014",
            INIT_19 => X"0000000f0000000d00000015000000260000003000000000fffffff6ffffffee",
            INIT_1A => X"00000029000000120000003600000027ffffffe2ffffffcbffffffd2fffffff1",
            INIT_1B => X"0000000c000000360000000a0000002e0000003c000000040000004f00000057",
            INIT_1C => X"0000001a00000011ffffffd9ffffffd4ffffffdfffffffecfffffff400000009",
            INIT_1D => X"00000004ffffffe6ffffffc1ffffffaf00000007000000000000000affffffed",
            INIT_1E => X"ffffffd7ffffffc3ffffffe0fffffff0fffffffafffffff8000000310000001d",
            INIT_1F => X"0000000ffffffff000000030000000680000003d000000110000005800000014",
            INIT_20 => X"ffffffd4fffffff700000012ffffffe8000000300000000a0000000fffffffde",
            INIT_21 => X"0000006200000060000000590000004e0000003f0000003affffffdd00000001",
            INIT_22 => X"ffffffe6fffffff60000000b0000001200000017000000370000004900000029",
            INIT_23 => X"00000017fffffff80000001100000010ffffffea00000003ffffffe600000006",
            INIT_24 => X"ffffffbfffffffc7ffffffec0000001afffffffbfffffffa00000005fffffffb",
            INIT_25 => X"0000003d0000002100000004000000120000001e000000210000002bffffffee",
            INIT_26 => X"0000000bffffffe3ffffffe9ffffffd2fffffff8000000090000000d00000035",
            INIT_27 => X"ffffffcaffffffc8ffffffdaffffffde0000000200000006000000220000001c",
            INIT_28 => X"ffffffe40000003200000006ffffffbf0000001effffffefffffffc500000009",
            INIT_29 => X"ffffffcefffffff600000004ffffffe20000000200000017ffffffd200000009",
            INIT_2A => X"fffffff40000001bffffffcafffffff20000001f000000110000002cfffffff6",
            INIT_2B => X"ffffffb20000005f00000019ffffffae0000003b0000000700000008fffffff8",
            INIT_2C => X"00000001ffffffd9ffffffd000000012fffffffeffffffd70000005e00000013",
            INIT_2D => X"0000001affffffee0000001efffffffcfffffffbffffffeaffffffe4fffffff3",
            INIT_2E => X"00000056ffffffa400000005000000030000001f00000000ffffffcffffffff7",
            INIT_2F => X"0000001f0000001d00000046ffffff8a0000000b0000008bffffff6300000017",
            INIT_30 => X"ffffffffffffffd400000016fffffff3ffffffea00000014ffffffdd0000000b",
            INIT_31 => X"ffffffdcfffffff4fffffff7ffffffea0000001bffffffe6fffffff000000014",
            INIT_32 => X"0000002200000014ffffffe1fffffff600000017fffffff7ffffffe2fffffff7",
            INIT_33 => X"ffffffed0000000200000062fffffff0ffffffe500000033ffffffeffffffff5",
            INIT_34 => X"00000050ffffff920000001300000045ffffffdbfffffffe000000230000000f",
            INIT_35 => X"ffffff490000000c00000047ffffff730000001c0000001affffffbb00000005",
            INIT_36 => X"fffffffaffffffd2000000120000000e00000054ffffff680000001b00000057",
            INIT_37 => X"0000000300000008fffffff6fffffffd00000019ffffffe9ffffffd6fffffff2",
            INIT_38 => X"0000004200000001ffffffd500000004fffffffdfffffff80000002200000012",
            INIT_39 => X"ffffffd8fffffffbfffffffa0000000dffffffc90000004500000001ffffffaa",
            INIT_3A => X"00000000ffffffddfffffff4ffffffe300000030fffffff40000001c0000001b",
            INIT_3B => X"ffffffdc00000011ffffffebfffffff30000001efffffff800000016fffffffb",
            INIT_3C => X"0000003b0000000bffffffee0000001effffffe6ffffffae0000003600000016",
            INIT_3D => X"ffffffc4ffffff83ffffffe3ffffffdeffffffb50000002dfffffff300000006",
            INIT_3E => X"fffffff50000002400000000ffffffc500000040ffffffefffffffa70000000a",
            INIT_3F => X"ffffffee0000000e0000000affffffe30000001a000000160000001400000042",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE0;


    MEM_IWGHT_LAYER2_INSTANCE1 : if BRAM_NAME = "iwght_layer2_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002a00000016fffffffbfffffff0ffffffd900000009ffffffe3ffffffe6",
            INIT_01 => X"0000002900000004fffffffe000000470000001c0000001c0000004c00000047",
            INIT_02 => X"fffffff0fffffff9ffffffe1ffffffdbffffffc800000011ffffffe8ffffffdf",
            INIT_03 => X"00000000ffffffac00000008ffffffc1ffffffcdffffffe6ffffffe20000001f",
            INIT_04 => X"ffffffd70000001600000011ffffffef0000002dffffffefffffffdefffffff9",
            INIT_05 => X"0000000dffffffcaffffffceffffffcdffffffce00000000000000300000000f",
            INIT_06 => X"0000000effffffed0000000bfffffff9ffffffd900000002ffffffc8ffffff94",
            INIT_07 => X"000000500000004d00000042000000160000002800000017000000010000003f",
            INIT_08 => X"0000003900000031ffffffcafffffff20000002a000000490000003c0000004f",
            INIT_09 => X"00000012ffffffe2000000210000002a0000003affffffea000000320000000f",
            INIT_0A => X"ffffffe90000000600000029ffffffdb000000190000001bffffffc40000000c",
            INIT_0B => X"ffffffecffffffd2ffffffaaffffffdcffffff9fffffffc0ffffff8cffffffae",
            INIT_0C => X"00000034ffffffecffffffd50000000afffffff6fffffff0000000150000000f",
            INIT_0D => X"fffffffe0000000bffffffe00000000500000006ffffffe700000018ffffffd5",
            INIT_0E => X"00000025ffffffcc0000002c00000005fffffff4fffffff8fffffffcfffffff2",
            INIT_0F => X"00000061ffffffdaffffffd2000000440000000c00000027ffffffc00000002f",
            INIT_10 => X"ffffffcaffffffe5fffffff000000003ffffffc80000004affffffe5ffffffac",
            INIT_11 => X"ffffffee0000000cfffffffd0000000effffffc40000001dffffffd5ffffffcc",
            INIT_12 => X"ffffffbb0000001bffffffc500000019fffffff1ffffffd80000002e0000000c",
            INIT_13 => X"0000002b0000005fffffff6a0000003100000068ffffff380000003900000019",
            INIT_14 => X"ffffffc7000000390000000f0000000500000033ffffffe60000001900000005",
            INIT_15 => X"00000007ffffffccffffffddfffffffbfffffffbfffffff30000000300000000",
            INIT_16 => X"00000029fffffff100000000fffffff8ffffffeefffffff70000000fffffffc4",
            INIT_17 => X"ffffffe10000003effffffcbffffffe90000002cffffffd1ffffffebfffffffc",
            INIT_18 => X"ffffffa50000001e00000023ffffffda0000001dffffffd300000039ffffffbf",
            INIT_19 => X"0000005400000012ffffffd00000001c0000005bffffff780000002a0000002a",
            INIT_1A => X"fffffff300000004000000200000007fffffff67000000590000004effffff86",
            INIT_1B => X"000000160000000dfffffffa000000030000000f00000017ffffffe20000001e",
            INIT_1C => X"ffffffdeffffffe70000000000000031ffffffc40000001cfffffffeffffffe8",
            INIT_1D => X"ffffffac0000004c00000009ffffff8100000060ffffffd3ffffffc900000033",
            INIT_1E => X"0000000400000007ffffffecfffffff1fffffff0fffffff1ffffffef00000013",
            INIT_1F => X"ffffffdbffffffe0ffffffffffffffc600000019fffffff400000010fffffff9",
            INIT_20 => X"0000001100000010ffffffe900000023fffffffa00000011ffffffc5ffffffbe",
            INIT_21 => X"000000080000000a0000000c000000050000002f00000021000000010000000f",
            INIT_22 => X"ffffff69ffffff88ffffff90ffffff91ffffffedfffffffd0000003a00000011",
            INIT_23 => X"fffffff90000000c00000022ffffff94ffffff7dffffff7dffffff8bffffff23",
            INIT_24 => X"000000270000000effffffe10000001700000038ffffffe6fffffffa0000001a",
            INIT_25 => X"0000000dffffffe80000000ffffffffd0000000900000023fffffffd00000012",
            INIT_26 => X"00000009000000120000000f0000001fffffffecffffffef0000001500000016",
            INIT_27 => X"ffffffa5ffffffaeffffffa8ffffffb1ffffffc5ffffffebffffffd600000006",
            INIT_28 => X"fffffffeffffffdbfffffff600000017ffffffe30000000affffffdeffffff9b",
            INIT_29 => X"ffffff84ffffff87ffffffc3fffffff7ffffffb7ffffffe700000015fffffff0",
            INIT_2A => X"fffffffffffffffe0000001fffffffed0000000fffffff8effffff94ffffffbc",
            INIT_2B => X"000000100000000700000023ffffffe30000000b00000001ffffffe700000020",
            INIT_2C => X"ffffffa9ffffff7effffff8f000000020000002f000000140000000700000028",
            INIT_2D => X"00000002fffffff7ffffffe3ffffffc8ffffffadffffffb0ffffff70ffffff71",
            INIT_2E => X"fffffff8000000010000000c0000001cffffffcdffffffe500000012ffffffe2",
            INIT_2F => X"0000002200000019000000130000000a0000001e00000000ffffffee0000000d",
            INIT_30 => X"0000003b00000026fffffff00000001dfffffff7fffffffc0000002800000016",
            INIT_31 => X"ffffffd50000000dfffffff3fffffffdffffffdd0000002f0000001b00000017",
            INIT_32 => X"00000008000000040000002a000000280000001000000032ffffffd3ffffffd9",
            INIT_33 => X"fffffff70000001dffffffea0000002f0000002c0000000c0000000300000014",
            INIT_34 => X"00000030ffffffd700000042fffffffdfffffff000000018fffffffd0000000d",
            INIT_35 => X"fffffff2ffffffe3ffffffc30000000d0000000a0000001b0000002100000030",
            INIT_36 => X"00000006ffffffea0000000b0000003f00000044fffffffffffffffbffffffef",
            INIT_37 => X"ffffffac0000000f00000035000000190000002f000000190000002100000003",
            INIT_38 => X"00000013000000270000001d00000001fffffffcfffffffcffffffaeffffff9b",
            INIT_39 => X"0000003cfffffff1ffffffe600000002fffffff7ffffffddffffffdbffffffec",
            INIT_3A => X"0000001900000000fffffff3fffffffb0000000f000000080000002b00000016",
            INIT_3B => X"ffffffe700000016fffffffa0000002800000025000000330000000dffffffdf",
            INIT_3C => X"0000000f00000005000000060000001000000037ffffffcf0000000dfffffffd",
            INIT_3D => X"000000270000003600000026000000180000000effffffcdffffffcd0000000e",
            INIT_3E => X"ffffffea0000000a00000016ffffffe2ffffffbeffffffe900000006fffffff9",
            INIT_3F => X"00000009ffffffc5ffffffdfffffffd600000002ffffffd8ffffffe50000000f",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE1;


    MEM_IWGHT_LAYER2_INSTANCE2 : if BRAM_NAME = "iwght_layer2_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffd600000029000000180000002d0000001f0000001c00000020fffffff0",
            INIT_01 => X"ffffffc4ffffffdeffffffed00000026ffffffd5ffffffcd0000000900000006",
            INIT_02 => X"0000001f00000002ffffffe9ffffffdefffffff6ffffffc7ffffffdeffffffdd",
            INIT_03 => X"ffffffedffffffecffffffd8ffffffd600000000ffffffd7ffffffee00000016",
            INIT_04 => X"fffffff5fffffffefffffff90000001c00000001fffffff100000002ffffffd3",
            INIT_05 => X"fffffff8fffffff4fffffffbffffffff000000020000000a00000000fffffff7",
            INIT_06 => X"0000003cfffffff60000002a0000002600000006ffffffefffffffdc00000000",
            INIT_07 => X"fffffff70000000afffffff5000000270000004800000044000000130000003b",
            INIT_08 => X"000000260000000000000007000000260000002400000012fffffffffffffff5",
            INIT_09 => X"ffffffcd0000000cfffffff3000000160000002e000000030000001800000030",
            INIT_0A => X"ffffff6bffffffa0ffffff9dffffff82ffffffaeffffffc1ffffffaaffffff92",
            INIT_0B => X"00000006ffffffcfffffffe10000001e00000004fffffff4ffffffda00000023",
            INIT_0C => X"00000015ffffffdffffffff1fffffff80000000bffffffdf00000000ffffffef",
            INIT_0D => X"0000000c0000003d0000002100000001000000200000002bffffffde0000001b",
            INIT_0E => X"fffffffffffffff9000000200000000000000022000000210000001e00000002",
            INIT_0F => X"00000008fffffff100000015fffffffbffffffec00000000ffffffff00000002",
            INIT_10 => X"ffffffe0ffffffd0fffffff20000000efffffff50000000200000020ffffffe2",
            INIT_11 => X"fffffff0ffffffd0ffffffd8ffffffd8ffffffc8ffffffd1ffffffdf00000013",
            INIT_12 => X"000000000000000dfffffff8000000080000000bffffffe2fffffff4ffffffe1",
            INIT_13 => X"fffffffcffffffeaffffffecffffffd0fffffff8fffffffbffffffd4fffffff2",
            INIT_14 => X"ffffffca00000000fffffff5fffffffbfffffff1000000150000000d00000019",
            INIT_15 => X"0000001cfffffff90000000cfffffff80000002b0000001bffffffe8ffffffb6",
            INIT_16 => X"00000020fffffff1fffffff6ffffffe4000000010000000900000025fffffff0",
            INIT_17 => X"00000020000000270000001000000012fffffffc00000015ffffffe7ffffffe5",
            INIT_18 => X"ffffff8dffffffd6ffffffc60000001500000014000000120000000f00000012",
            INIT_19 => X"000000220000000200000023000000040000000fffffffd200000021ffffffb7",
            INIT_1A => X"fffffff90000001affffffe5ffffffecfffffff900000012fffffffe00000006",
            INIT_1B => X"0000001d0000001100000016fffffff30000001d0000001affffffef00000014",
            INIT_1C => X"0000000f0000000e000000150000002000000016000000260000000c0000000c",
            INIT_1D => X"0000002e0000000afffffff90000000e000000050000000c0000002600000027",
            INIT_1E => X"00000003ffffffebffffffd70000000affffffff0000001a0000002c00000000",
            INIT_1F => X"000000210000003d00000049000000180000003ffffffffeffffffd0ffffffe0",
            INIT_20 => X"fffffff8ffffffd3fffffff6ffffffd7ffffffc400000029000000390000003f",
            INIT_21 => X"ffffffeaffffffebffffffde00000031fffffffd00000010fffffff3fffffff3",
            INIT_22 => X"ffffffc4ffffffd30000000d0000001affffffe5fffffff0ffffffd8ffffffaa",
            INIT_23 => X"00000013000000230000002800000029ffffffe4fffffff8fffffff6ffffffd2",
            INIT_24 => X"00000018ffffffdeffffffbdffffffd1fffffff1ffffffe6fffffff4fffffff3",
            INIT_25 => X"fffffff8ffffffcbffffffe4ffffffcefffffff1fffffffdfffffff10000001e",
            INIT_26 => X"00000024fffffff7ffffffe8fffffffbffffffedffffffc5ffffffe80000002e",
            INIT_27 => X"000000380000000a0000001d0000002afffffff500000004fffffff700000004",
            INIT_28 => X"fffffffdffffffebfffffff100000014000000130000001cfffffffdfffffff2",
            INIT_29 => X"0000002500000026fffffff70000000f0000003400000004ffffffed00000002",
            INIT_2A => X"0000006500000002000000060000000c000000070000001c0000001cfffffffb",
            INIT_2B => X"ffffffddfffffff7ffffffe00000000600000017000000350000002a00000038",
            INIT_2C => X"ffffffcbffffffddffffffcafffffff9ffffffe5ffffffc3ffffffddffffffe8",
            INIT_2D => X"00000035ffffff9cffffff96fffffff5ffffff62ffffff78ffffffa7ffffffbc",
            INIT_2E => X"ffffffd7ffffffbfffffffdcffffffe9ffffffbdffffffc7000000050000003b",
            INIT_2F => X"00000023fffffff7ffffffdc0000001d0000000400000010ffffffc70000002e",
            INIT_30 => X"fffffffaffffffe9ffffffe20000001900000000000000080000000afffffff5",
            INIT_31 => X"0000001e0000001200000019fffffff70000001e000000000000000300000011",
            INIT_32 => X"fffffff8fffffffa0000001a0000000efffffff6000000230000001b0000001c",
            INIT_33 => X"fffffff2ffffffc1ffffffa1ffffffb10000000f0000001b0000002bfffffff2",
            INIT_34 => X"ffffffea0000000e00000005ffffffb4ffffffccfffffffaffffffa5ffffffc1",
            INIT_35 => X"00000008ffffffe500000030000000370000000a0000003e0000003c00000040",
            INIT_36 => X"ffffffe7ffffffed00000014ffffffebfffffff7ffffffe9fffffff100000016",
            INIT_37 => X"00000028000000290000002b00000008000000050000002c00000001fffffff8",
            INIT_38 => X"00000018fffffffbfffffffe0000000000000001ffffffeb00000005ffffffe8",
            INIT_39 => X"ffffffe70000004b0000003300000011fffffff4ffffffe400000021fffffffb",
            INIT_3A => X"0000001c0000000a000000240000001d000000110000002900000022fffffff5",
            INIT_3B => X"0000001e0000000500000034ffffffedfffffff9fffffff3ffffffe7ffffffe6",
            INIT_3C => X"00000012000000180000001dfffffffbffffffe1ffffffe6fffffff1ffffffed",
            INIT_3D => X"ffffffe10000000d00000013000000120000001b000000230000001e00000013",
            INIT_3E => X"000000010000003cffffffce0000000d00000013fffffffe0000002400000014",
            INIT_3F => X"00000016000000320000003500000005000000040000003c0000001dffffffe7",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE2;


    MEM_IWGHT_LAYER2_INSTANCE3 : if BRAM_NAME = "iwght_layer2_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000250000001b0000001b0000003e0000003200000042ffffffed00000000",
            INIT_01 => X"0000003a0000002b0000002a00000062000000410000001500000020fffffffc",
            INIT_02 => X"ffffffe800000017fffffffa0000000d00000009fffffffd0000001800000044",
            INIT_03 => X"0000004e0000005200000036000000000000001900000007ffffffcaffffffcc",
            INIT_04 => X"000000230000000000000002fffffffbffffffef000000410000003800000014",
            INIT_05 => X"00000002000000140000001e0000001bfffffff900000011fffffffd0000002a",
            INIT_06 => X"fffffff2fffffff00000000a00000009ffffffe2fffffff8ffffffef00000004",
            INIT_07 => X"00000013fffffff4ffffffc9fffffff200000019ffffffd4ffffffde00000010",
            INIT_08 => X"fffffffafffffffdffffffd3ffffffd9fffffffa0000000afffffff9fffffffc",
            INIT_09 => X"fffffff800000009fffffff7000000000000001efffffffb0000002300000009",
            INIT_0A => X"00000013fffffff70000002b00000008000000040000002100000000ffffffea",
            INIT_0B => X"fffffffb0000001e00000014ffffffe400000017fffffffd0000001f00000003",
            INIT_0C => X"ffffffea00000010ffffffdc000000160000000700000005000000350000002d",
            INIT_0D => X"ffffffdcffffffd50000002a0000001afffffff6fffffffc00000013ffffffe1",
            INIT_0E => X"ffffff4affffffe5ffffffd8ffffffae00000015ffffffbbffffffcefffffff0",
            INIT_0F => X"ffffffe40000000f00000000ffffff65ffffff73ffffff74ffffff63ffffff45",
            INIT_10 => X"0000001300000031ffffffe90000001afffffff600000000000000040000000e",
            INIT_11 => X"fffffff7ffffffda0000001800000037ffffffe7000000220000005bffffffc9",
            INIT_12 => X"000000060000002000000051ffffffd80000000300000028ffffffcbfffffffa",
            INIT_13 => X"0000002d0000004bfffffffa0000001100000002ffffffc5ffffffd7ffffffe2",
            INIT_14 => X"ffffffcb000000320000001effffffdb000000370000002bffffffee0000001d",
            INIT_15 => X"ffffffd3ffffffc9ffffffc9ffffffccffffff7effffffc10000000e00000001",
            INIT_16 => X"000000200000000b000000060000000100000016ffffffebffffffc6ffffffcb",
            INIT_17 => X"0000003f0000000c0000000500000032000000190000002dfffffff500000013",
            INIT_18 => X"000000220000000cfffffffa0000001500000037000000330000001b00000026",
            INIT_19 => X"0000002500000018fffffff3ffffffc3ffffffcbffffffd1ffffff99ffffff82",
            INIT_1A => X"00000002ffffffcdffffffe90000000100000019fffffffb00000018fffffff8",
            INIT_1B => X"0000001a00000019000000180000001900000015fffffff800000027ffffffd9",
            INIT_1C => X"fffffffe00000012ffffffeeffffffddffffffe6fffffffaffffffe0ffffffec",
            INIT_1D => X"fffffff8ffffffd90000000c0000000cffffffdf00000011fffffff000000018",
            INIT_1E => X"0000001100000005fffffffc00000012fffffff400000005ffffffdcfffffffb",
            INIT_1F => X"0000000000000000fffffff900000011ffffffff00000016ffffffe1ffffffee",
            INIT_20 => X"ffffffcdffffffa3ffffff9fffffffceffffffecffffffe2fffffff60000000e",
            INIT_21 => X"0000001f0000000f0000000cffffffffffffffec00000012ffffffbfffffffc8",
            INIT_22 => X"fffffffeffffffee00000018fffffff90000001300000007000000140000000a",
            INIT_23 => X"ffffffaf00000012fffffff1ffffffcfffffffefffffffdbffffffdefffffffc",
            INIT_24 => X"ffffffd6ffffffcaffffffeeffffffddffffffb0ffffffafffffffd2ffffffd0",
            INIT_25 => X"00000013fffffff4ffffffe9ffffffbdffffffefffffff97ffffffa8ffffff96",
            INIT_26 => X"0000001f0000002300000017fffffffe00000001fffffffd00000006fffffff0",
            INIT_27 => X"ffffffc5ffffffb5ffffffc2ffffff95ffffff63ffffffad0000000600000023",
            INIT_28 => X"00000008ffffffe1fffffff80000001400000017ffffffdeffffffe2ffffffc4",
            INIT_29 => X"00000012000000030000001e0000000bfffffff0000000090000000afffffffb",
            INIT_2A => X"ffffffb100000000fffffff1000000110000000e00000017fffffff0fffffff7",
            INIT_2B => X"fffffffbffffffec00000014000000280000001fffffffefffffffcfffffffe8",
            INIT_2C => X"fffffff3ffffffdefffffffbffffffe3000000080000000f0000000dfffffff3",
            INIT_2D => X"fffffff700000028fffffffdffffffcd0000000bffffffefffffffd0ffffffd7",
            INIT_2E => X"00000023000000010000001cfffffffeffffffd9000000010000000dffffffcd",
            INIT_2F => X"0000000affffffecffffffe00000000efffffff9ffffffef000000100000002a",
            INIT_30 => X"fffffff5ffffffdfffffffff00000011fffffff200000003ffffffddfffffffb",
            INIT_31 => X"fffffff2ffffffed000000160000000300000003000000100000000a0000001b",
            INIT_32 => X"0000006a0000002c000000140000003dfffffff1fffffff1fffffffd00000003",
            INIT_33 => X"ffffffb6ffffffc6ffffffbb000000750000004d000000690000005c0000005f",
            INIT_34 => X"ffffffd2ffffffc0000000290000001e00000020fffffffbfffffff8ffffffae",
            INIT_35 => X"ffffff9bffffffe9ffffffcbffffffd3ffffffc6ffffff95ffffffa9ffffffc3",
            INIT_36 => X"00000013000000270000001bffffffb5ffffffb5ffffffbdffffffbdffffffa7",
            INIT_37 => X"0000001effffffe900000014000000440000002cffffffe2000000070000002b",
            INIT_38 => X"0000000000000001fffffff100000000000000110000001efffffff100000002",
            INIT_39 => X"00000009000000070000000200000005000000190000001c0000000fffffffee",
            INIT_3A => X"ffffffec00000007000000190000000300000029ffffffd1fffffff900000010",
            INIT_3B => X"fffffff5000000020000001e0000000cfffffffeffffffd8fffffffd0000000b",
            INIT_3C => X"fffffffdfffffff7fffffffc00000007ffffffe20000000c000000150000000e",
            INIT_3D => X"fffffff2ffffffcf000000320000003b00000060000000280000003a0000004f",
            INIT_3E => X"fffffffa00000038fffffffffffffffbffffffed00000018fffffffbfffffff4",
            INIT_3F => X"0000000800000016fffffff6fffffffbffffffe6fffffff8fffffff6ffffffe3",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE3;


    MEM_IWGHT_LAYER2_INSTANCE4 : if BRAM_NAME = "iwght_layer2_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff0fffffffefffffffa0000000700000018fffffffdfffffff000000006",
            INIT_01 => X"ffffffb600000006fffffffaffffffe10000002e00000000ffffffdffffffff0",
            INIT_02 => X"ffffffecffffffe1ffffffdf0000001ffffffffefffffffdfffffff2ffffffdb",
            INIT_03 => X"000000080000001e0000001f0000000600000019000000010000000900000000",
            INIT_04 => X"fffffef2ffffffe3ffffff56ffffff63ffffffeb00000005fffffffe00000005",
            INIT_05 => X"ffffffed0000002b0000003cffffff2fffffff1effffff33ffffff1bfffffeb6",
            INIT_06 => X"fffffffd0000001900000000000000270000003bfffffff30000001900000029",
            INIT_07 => X"0000001effffffea0000000c00000011fffffff20000000300000039fffffff8",
            INIT_08 => X"0000002a0000001900000051fffffffb000000040000000f00000000fffffff6",
            INIT_09 => X"fffffff5000000130000002cffffffef0000002d00000010ffffffd700000000",
            INIT_0A => X"fffffffd0000001ffffffff5ffffffeb0000000b0000000d00000024fffffff3",
            INIT_0B => X"ffffffdeffffffe3ffffffddffffffeaffffffd3fffffff0ffffffff0000000f",
            INIT_0C => X"fffffffbffffffde00000001fffffffdfffffffefffffffaffffffc7ffffffe6",
            INIT_0D => X"00000017ffffffea0000001e00000024ffffffe4ffffffd7fffffff20000001c",
            INIT_0E => X"0000000effffff7cffffff88fffffff8fffffffc00000006ffffffdcfffffff7",
            INIT_0F => X"000000030000001fffffff84ffffff38ffffff6bffffff5dffffff3affffff12",
            INIT_10 => X"ffffffcdffffffecfffffffeffffffed000000010000002100000011fffffff8",
            INIT_11 => X"00000013ffffffea00000000fffffff9ffffffe5ffffffd1fffffff0fffffff5",
            INIT_12 => X"00000033000000300000001d00000016ffffffe7fffffff60000002e00000033",
            INIT_13 => X"00000016ffffffdf00000001000000290000001afffffff40000002f0000000b",
            INIT_14 => X"ffffffe9ffffffd0fffffffb000000150000000ffffffffafffffff4fffffff4",
            INIT_15 => X"00000003fffffff9fffffffdffffffecffffffffffffffd0ffffffc8fffffff9",
            INIT_16 => X"fffffff6fffffff3ffffffecffffffda00000009ffffffdcffffffe5ffffffed",
            INIT_17 => X"ffffffe0ffffffe3ffffffe600000001ffffffebffffffd100000007ffffffb0",
            INIT_18 => X"ffffffb3ffffffce00000001ffffffe7ffffffe5fffffff2fffffffeffffffee",
            INIT_19 => X"ffffff52ffffffbeffffff8dffffff92ffffffc3ffffffaeffffffc4ffffffab",
            INIT_1A => X"ffffff90ffffff75ffffff94ffffffb4ffffff75ffffff83ffffffd6ffffffa2",
            INIT_1B => X"ffffffc7ffffffc2ffffffd6ffffffe5ffffffcaffffffdfffffffd9ffffffd3",
            INIT_1C => X"000000140000001f0000001f0000002700000001000000250000002bffffffc4",
            INIT_1D => X"ffffffeafffffff9ffffffeb00000010ffffffee000000210000000100000017",
            INIT_1E => X"000000000000000700000027000000140000000b00000007ffffffe4fffffff1",
            INIT_1F => X"000000160000000e0000003ffffffffdffffffff000000230000001c0000000a",
            INIT_20 => X"ffffffc00000001cffffffe90000003f0000003600000028000000280000004a",
            INIT_21 => X"00000008ffffffdb0000000f0000000c0000001900000001ffffffecffffffcb",
            INIT_22 => X"00000026ffffffe5ffffffebffffffcefffffffeffffffdd0000000000000010",
            INIT_23 => X"000000730000007e0000004d0000006900000065000000380000000d0000001d",
            INIT_24 => X"ffffffe3ffffffeafffffffe00000012fffffffc000000070000002b00000028",
            INIT_25 => X"00000036000000240000002000000019ffffffb9ffffff8dffffffbeffffffd5",
            INIT_26 => X"fffffff1fffffff400000016000000070000001900000011000000460000002d",
            INIT_27 => X"0000001e00000008ffffffe8ffffffbbffffffc8fffffff0fffffff4ffffffdc",
            INIT_28 => X"0000000e000000220000001d0000004100000025000000200000001affffffe6",
            INIT_29 => X"000000200000005000000036ffffffcffffffff00000002a0000001b00000017",
            INIT_2A => X"000000480000004fffffffd7ffffffaaffffffd8fffffff8ffffffed00000012",
            INIT_2B => X"00000062ffffffd9ffffffa2ffffffd000000004ffffffe9ffffffec00000023",
            INIT_2C => X"ffffffabffffff8effffffb7fffffffa0000001d000000040000004d0000007d",
            INIT_2D => X"ffffffdaffffffbf0000001a000000170000001d000000260000003200000042",
            INIT_2E => X"0000000f000000150000001600000013fffffff6ffffffdaffffffe0ffffffea",
            INIT_2F => X"ffffffff000000100000000effffffc1ffffffb7ffffffc00000002400000004",
            INIT_30 => X"0000000bfffffff1ffffffb5ffffffa6ffffffdb00000021000000290000002a",
            INIT_31 => X"ffffffe800000011fffffff7fffffffe00000031000000460000004100000007",
            INIT_32 => X"fffffff30000000b00000025ffffffe5ffffffd8fffffff9ffffffe1fffffff5",
            INIT_33 => X"00000004fffffffdfffffffe000000000000002b000000110000001500000016",
            INIT_34 => X"00000019ffffffc3ffffffddffffffe20000001900000010fffffffa00000033",
            INIT_35 => X"ffffffc0ffffffcbffffffdd000000040000000d00000010000000280000002f",
            INIT_36 => X"ffffffe7ffffffcafffffffe00000000fffffff8ffffffefffffffe9fffffffb",
            INIT_37 => X"00000024000000060000003700000014ffffffdffffffff30000000affffffdc",
            INIT_38 => X"0000002efffffff3000000010000003600000023fffffff20000002500000003",
            INIT_39 => X"00000010000000000000001a0000002a00000023fffffff900000002fffffff2",
            INIT_3A => X"00000036fffffffe000000130000002e0000000cfffffffa0000001400000016",
            INIT_3B => X"ffffffe6ffffffe3ffffffdcfffffff500000020000000060000000800000001",
            INIT_3C => X"0000000ffffffffbfffffff8fffffff7fffffff100000003ffffffefffffffec",
            INIT_3D => X"0000000b000000380000001200000027000000130000000a0000000100000010",
            INIT_3E => X"000000490000003a000000420000001f0000005a00000060ffffffe80000001f",
            INIT_3F => X"00000016000000260000002c0000003d00000022fffffff40000001700000021",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE4;


    MEM_IWGHT_LAYER2_INSTANCE5 : if BRAM_NAME = "iwght_layer2_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffe3000000240000000cfffffff50000002800000000ffffffe90000001a",
            INIT_01 => X"ffffffc7000000260000001bffffffe9fffffff700000015000000040000000e",
            INIT_02 => X"0000002b0000001f0000001cfffffffd0000001effffffd8ffffffdbfffffff7",
            INIT_03 => X"fffffff200000023fffffffbffffffd100000030000000130000001d00000028",
            INIT_04 => X"ffffffe500000010fffffff1ffffffe3ffffffd7ffffffdaffffffdcffffffe8",
            INIT_05 => X"0000001dfffffff8fffffffc0000001100000021000000080000000500000028",
            INIT_06 => X"ffffffc6ffffffe7fffffff0ffffffeafffffff3ffffffef0000001affffffea",
            INIT_07 => X"ffffffa8ffffffcaffffffd3ffffffcdffffffd3ffffffb5ffffffb8ffffffbe",
            INIT_08 => X"000000330000001900000020000000360000003d000000110000002d00000031",
            INIT_09 => X"00000063000000000000000f00000043000000520000002d0000004500000021",
            INIT_0A => X"00000057fffffff6000000020000001500000011000000360000001500000025",
            INIT_0B => X"ffffff8bffffffa7ffffff96fffffff2ffffffe4000000370000002a0000000e",
            INIT_0C => X"ffffffbb00000012ffffffe3ffffffcb00000018ffffffa8ffffffbfffffffa6",
            INIT_0D => X"ffffffd70000000dffffffe700000012ffffffffffffffe600000029ffffffe0",
            INIT_0E => X"ffffffbfffffffb70000000bfffffffbffffffcfffffffea00000004ffffffe1",
            INIT_0F => X"ffffffe200000003000000030000000a0000000effffffcaffffffe3ffffffb1",
            INIT_10 => X"0000002100000029ffffffe9000000200000000afffffff4ffffffe7fffffffe",
            INIT_11 => X"0000000affffffdf0000000c00000011fffffff1ffffffe6fffffff4ffffffe5",
            INIT_12 => X"ffffffbeffffffd2ffffffc8ffffffdbffffffcd00000001fffffff000000030",
            INIT_13 => X"00000010fffffffa0000000f000000060000003dffffffcefffffffeffffffe1",
            INIT_14 => X"ffffffd20000000f000000270000001b0000002300000032fffffff5fffffffd",
            INIT_15 => X"0000000400000001000000080000003cfffffffaffffffef000000190000000e",
            INIT_16 => X"0000002bffffffebffffffff0000001a0000003e00000004000000200000002c",
            INIT_17 => X"00000023000000090000002200000031fffffff500000049fffffffaffffffd9",
            INIT_18 => X"000000400000002efffffff8ffffffe100000022000000240000000ffffffff0",
            INIT_19 => X"00000030000000200000002c0000004e000000440000004d0000003f00000056",
            INIT_1A => X"000000200000000bfffffffc000000150000000fffffffe7fffffffa0000001c",
            INIT_1B => X"ffffffcbffffffdcffffffbaffffffa8ffffffc9ffffffc4fffffff9ffffffed",
            INIT_1C => X"00000002000000000000001b0000000effffffe4fffffff2ffffffcdffffffbd",
            INIT_1D => X"0000001f0000001600000003ffffffebfffffff500000009000000000000000b",
            INIT_1E => X"ffffffe8fffffffbfffffffbffffffedfffffff5000000080000002500000000",
            INIT_1F => X"fffffffffffffffd00000019000000350000001bffffffddffffffdeffffffeb",
            INIT_20 => X"0000000ffffffff900000026000000290000001800000009000000030000001c",
            INIT_21 => X"ffffffdeffffffea0000001500000019ffffffe7fffffff30000000bffffffe7",
            INIT_22 => X"ffffffccffffffb6ffffffd6ffffffe8fffffff4ffffffd9ffffffc9fffffff5",
            INIT_23 => X"ffffffe7fffffffd00000007ffffffdbffffffdeffffffff0000000afffffff8",
            INIT_24 => X"00000010ffffffef000000110000001300000012fffffff700000019fffffff7",
            INIT_25 => X"00000009fffffffd0000000ffffffffdffffffe4fffffffb0000001700000007",
            INIT_26 => X"ffffffcefffffffaffffffe0ffffffd7ffffffdd00000007ffffffee00000004",
            INIT_27 => X"00000010fffffff00000001afffffffafffffff7fffffff9ffffffe4ffffffec",
            INIT_28 => X"ffffffc7ffffffc9ffffffc10000001700000024ffffffe1ffffffe80000000a",
            INIT_29 => X"000000160000001cffffffcfffffffbcffffffc600000009ffffffb9ffffffcf",
            INIT_2A => X"ffffffe600000002000000010000001effffffef000000190000001e0000000f",
            INIT_2B => X"ffffffffffffffdffffffff2ffffffef000000040000000affffffe000000006",
            INIT_2C => X"00000035fffffff2000000120000000200000019000000190000001400000005",
            INIT_2D => X"fffffff50000000affffffd7ffffffd30000000300000000ffffffec00000022",
            INIT_2E => X"ffffffd1ffffffdfffffffd2fffffff7ffffffc2ffffffc000000003ffffffeb",
            INIT_2F => X"ffffffe4ffffffe3ffffffd2ffffffefffffffdaffffffe6fffffff600000005",
            INIT_30 => X"fffffff8fffffff80000001500000025fffffff4ffffffe9ffffffe6ffffffec",
            INIT_31 => X"00000014000000210000000d00000002fffffffafffffff600000023fffffff9",
            INIT_32 => X"ffffffe3ffffffed000000100000000800000021fffffff10000000bfffffffc",
            INIT_33 => X"ffffffe9ffffffddfffffff300000012ffffffe9ffffffcaffffffc5ffffffdf",
            INIT_34 => X"ffffffe3ffffffdeffffffedffffffe6ffffffe0ffffffe3ffffffd2fffffff7",
            INIT_35 => X"fffffffb0000001bfffffff1fffffff500000004fffffffb0000000f0000000f",
            INIT_36 => X"fffffff7000000050000000600000006ffffffee0000000300000013ffffffe0",
            INIT_37 => X"0000001a000000190000000e0000000100000023000000080000000200000015",
            INIT_38 => X"ffffffe3fffffff300000008fffffffa00000007000000310000000cfffffffe",
            INIT_39 => X"000000060000003e0000002c00000004ffffffdbffffffdafffffffdffffffd5",
            INIT_3A => X"000000050000000afffffff40000001600000035000000080000003f0000000f",
            INIT_3B => X"ffffffddffffffe60000000bffffffefffffffd000000000ffffffdbfffffff5",
            INIT_3C => X"0000000efffffff8ffffffe70000001d00000008fffffff50000000b0000000e",
            INIT_3D => X"0000001b0000002b00000010000000370000001e000000100000002d00000036",
            INIT_3E => X"fffffff0ffffffff000000190000000800000017000000070000000bffffffe4",
            INIT_3F => X"fffffffeffffffc5ffffffc5ffffffc3ffffffeb00000000000000110000000c",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE5;


    MEM_IWGHT_LAYER2_INSTANCE6 : if BRAM_NAME = "iwght_layer2_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffebfffffff5ffffffd7fffffff7ffffffe70000000effffffdbffffffd1",
            INIT_01 => X"ffffffdb0000000800000001000000140000001bfffffff0ffffffd7ffffffd3",
            INIT_02 => X"ffffffdaffffffefffffffd0ffffffed0000000b0000000cfffffff9ffffffe8",
            INIT_03 => X"0000001cffffffeafffffff20000000bffffffc1ffffffd8ffffffe5fffffff8",
            INIT_04 => X"00000000ffffffe7000000250000000d00000022000000280000001700000015",
            INIT_05 => X"fffffff40000000afffffff400000006ffffffff00000014ffffffe200000004",
            INIT_06 => X"fffffff5ffffffe7ffffffe2ffffffe8fffffff000000006ffffffe6ffffffd4",
            INIT_07 => X"ffffffce000000140000000bffffffecfffffff700000001fffffffc00000035",
            INIT_08 => X"fffffff30000000900000018ffffffef00000006000000110000001cfffffffc",
            INIT_09 => X"fffffff4fffffff6000000280000001b000000090000000effffffec00000008",
            INIT_0A => X"0000000000000000fffffff2fffffff8fffffffbffffffffffffffed0000000d",
            INIT_0B => X"fffffff600000010fffffff000000000ffffffcbffffffc4fffffff8ffffffbe",
            INIT_0C => X"ffffffcfffffffdcffffffd500000007000000280000001800000006fffffff7",
            INIT_0D => X"00000007fffffff1ffffffceffffffc9ffffffcbffffffd0fffffff0ffffffc2",
            INIT_0E => X"ffffffdcffffffd9fffffff8fffffffcfffffff9ffffffdcffffffe500000008",
            INIT_0F => X"0000000d0000001b0000000e0000002cfffffffeffffffed0000000200000008",
            INIT_10 => X"fffffff500000004ffffffff00000017ffffffdeffffffdfffffffe1fffffff9",
            INIT_11 => X"ffffffeaffffffee0000001dfffffff1ffffffe400000006fffffff800000017",
            INIT_12 => X"fffffff30000000c00000009ffffffe20000001f00000037ffffffefffffffe9",
            INIT_13 => X"0000001f0000000c000000200000001a000000390000000c0000001000000000",
            INIT_14 => X"ffffffeffffffff30000000b0000001bfffffffa0000001c00000026fffffffb",
            INIT_15 => X"ffffffdbfffffff1ffffffeefffffff70000000a00000014fffffff4fffffff2",
            INIT_16 => X"ffffffcc000000200000000500000001ffffffe9ffffffd5ffffffc4ffffffdf",
            INIT_17 => X"ffffffceffffffb70000001f00000000ffffffc0ffffffe100000000ffffffd1",
            INIT_18 => X"0000003c000000360000003b00000003ffffffa5ffffffd4ffffffbeffffffb9",
            INIT_19 => X"fffffffefffffff3fffffff1fffffff100000001fffffff1fffffff7ffffffe3",
            INIT_1A => X"ffffffed00000000000000270000000b00000009000000300000001a0000001c",
            INIT_1B => X"fffffff9000000240000003500000026000000100000000afffffff20000000e",
            INIT_1C => X"0000000500000009ffffffe0ffffffec0000000afffffff800000019ffffffe7",
            INIT_1D => X"00000001ffffffde00000001fffffffaffffffe6fffffff8fffffff2ffffffe4",
            INIT_1E => X"ffffffe80000000300000015ffffffe0000000170000000bffffffa7ffffffdb",
            INIT_1F => X"fffffff200000017fffffff2ffffffe700000010fffffffd0000001400000019",
            INIT_20 => X"ffffff9d0000000efffffff00000001fffffffe3fffffff1fffffffd00000001",
            INIT_21 => X"fffffffd00000006ffffffebfffffff000000006ffffffccffffffef00000000",
            INIT_22 => X"000000170000000b0000000b00000013fffffff4ffffffdf00000007ffffffe2",
            INIT_23 => X"0000000e00000002ffffffdcfffffff40000000400000018000000300000000d",
            INIT_24 => X"000000010000002a00000050fffffffe0000000b00000022ffffff8bfffffffa",
            INIT_25 => X"ffffffea0000001afffffff5ffffffeafffffff500000007000000390000003b",
            INIT_26 => X"fffffff0ffffffe400000015ffffffdd00000019000000200000002efffffffc",
            INIT_27 => X"000000290000001300000014000000070000000d00000005fffffffbffffffe0",
            INIT_28 => X"0000002d000000420000003e00000007fffffff6000000560000003c00000008",
            INIT_29 => X"00000014000000570000003e0000003d00000037000000600000004c00000033",
            INIT_2A => X"0000001b0000002b000000110000006b00000041000000450000001500000047",
            INIT_2B => X"fffffff90000001c00000024000000070000001500000039000000240000001f",
            INIT_2C => X"00000006fffffffdffffffe20000000bfffffffffffffff10000001800000015",
            INIT_2D => X"00000001ffffffb7ffffffc7fffffffdffffffe3ffffffdf00000005ffffffe7",
            INIT_2E => X"ffffffdf00000010ffffffe6ffffffd20000000afffffff4ffffffbfffffffe5",
            INIT_2F => X"fffffffeffffffe5ffffffd9ffffffefffffffc90000000e0000003affffffa8",
            INIT_30 => X"ffffffdcffffffdafffffff6ffffffccffffffe6ffffffdcffffffabffffffca",
            INIT_31 => X"0000000500000009fffffffa000000170000001fffffffe700000003ffffffff",
            INIT_32 => X"ffffffbf000000080000000d000000010000002300000020ffffffe000000018",
            INIT_33 => X"ffffffdfffffffccffffffe3ffffffbeffffffcafffffff9ffffffd8ffffffe3",
            INIT_34 => X"fffffff900000013fffffff9ffffffff00000003fffffffcfffffff7ffffffeb",
            INIT_35 => X"00000036ffffffcafffffff10000002a00000016fffffff20000003400000000",
            INIT_36 => X"ffffffedffffffd500000027ffffffb4ffffffca00000006ffffffaa00000003",
            INIT_37 => X"0000002f00000063ffffffc00000001a00000033ffffffeeffffffef0000002e",
            INIT_38 => X"00000019ffffffc90000001b00000034000000020000004e00000040fffffff8",
            INIT_39 => X"ffffffeb000000230000001d0000002e00000024ffffffbb0000000400000006",
            INIT_3A => X"ffffffc5ffffffdf0000002100000000000000090000001500000003ffffffef",
            INIT_3B => X"ffffffedffffffe3ffffffb30000001100000009ffffffa4ffffffea00000048",
            INIT_3C => X"0000000b00000018fffffff30000001d00000002fffffff20000001e0000000a",
            INIT_3D => X"ffffffedffffffe6ffffffe7ffffffdbfffffff500000019ffffffe2ffffffea",
            INIT_3E => X"00000031ffffffb1ffffffe800000043ffffffcaffffffe000000002ffffffe7",
            INIT_3F => X"000000300000001300000010000000210000002600000009ffffffc50000001f",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE6;


    MEM_IWGHT_LAYER2_INSTANCE7 : if BRAM_NAME = "iwght_layer2_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffff9f00000038fffffffdffffffe2ffffffff00000018fffffffaffffffff",
            INIT_01 => X"ffffffb30000000cffffffe3ffffffb9ffffffbefffffff400000056fffffffe",
            INIT_02 => X"ffffffc5ffffffe100000002fffffff8ffffff85fffffff4fffffffcffffff5d",
            INIT_03 => X"ffffffe400000010ffffffec0000000effffffe6ffffffd1ffffffd3fffffff7",
            INIT_04 => X"0000001bffffffe60000001a00000014ffffffde0000001600000009ffffffd6",
            INIT_05 => X"000000590000001fffffffca000000590000002affffffeb000000130000002f",
            INIT_06 => X"fffffffe0000002c00000009000000150000000b0000001dfffffff2ffffffe1",
            INIT_07 => X"00000006fffffff2fffffff400000013ffffffc2ffffffeaffffffc8fffffff4",
            INIT_08 => X"00000000ffffffe80000001300000012ffffffec0000000cffffffd4ffffffdf",
            INIT_09 => X"000000000000000e00000007000000030000000700000007ffffffee00000001",
            INIT_0A => X"0000007400000029000000370000005700000019000000180000000000000016",
            INIT_0B => X"fffffff600000009fffffffa0000002f00000056000000360000007200000083",
            INIT_0C => X"00000013fffffff0fffffffd00000006fffffff3fffffff7fffffff2ffffffee",
            INIT_0D => X"0000000f0000001b0000000a0000000cffffffee00000033ffffffec0000000d",
            INIT_0E => X"ffffffdffffffff9ffffffd1ffffffe900000017ffffffee0000001b00000014",
            INIT_0F => X"fffffff4ffffffecffffffe50000002600000008000000380000002efffffff8",
            INIT_10 => X"00000000fffffff400000001ffffffe8ffffffdd00000008ffffffe5ffffffd6",
            INIT_11 => X"0000003a00000039000000580000002f0000000f000000220000001ffffffffa",
            INIT_12 => X"00000027ffffffdffffffffb0000000e0000000f000000200000001a00000036",
            INIT_13 => X"000000030000000cfffffff800000000ffffffd6fffffffdffffffe7ffffffd3",
            INIT_14 => X"00000031000000340000001e000000260000002b000000010000003000000004",
            INIT_15 => X"ffffffe50000001e0000003f0000002f0000003c000000300000002a00000029",
            INIT_16 => X"0000000700000014fffffff9ffffffe8ffffffefffffffed00000004fffffff4",
            INIT_17 => X"ffffffd3ffffffef0000000b00000000ffffffd10000001200000012ffffffd7",
            INIT_18 => X"ffffffc5ffffffd7ffffffdbffffffe5ffffffcb000000060000000000000007",
            INIT_19 => X"0000004dfffffffc0000001a0000001c0000000400000006fffffff4fffffff1",
            INIT_1A => X"ffffffe3ffffffe000000011fffffffc0000000dffffffe90000001e00000035",
            INIT_1B => X"ffffffff00000014ffffffddffffffe50000001f00000003000000010000001b",
            INIT_1C => X"fffffff70000001c0000002a0000000c00000019000000130000000c00000016",
            INIT_1D => X"0000000300000000ffffffc900000022fffffffc000000210000000800000031",
            INIT_1E => X"00000000fffffff9ffffffa5ffffffd1ffffffafffffffd0ffffffaeffffffc3",
            INIT_1F => X"fffffff1ffffffc0ffffffe2fffffff3ffffffe9ffffffbbffffffdcfffffff9",
            INIT_20 => X"ffffffb1ffffffd2ffffffaafffffff8ffffff9bffffff960000005d00000023",
            INIT_21 => X"00000007ffffffcd00000024ffffffe0ffffffd80000000afffffffeffffffe9",
            INIT_22 => X"000000140000001600000002fffffffcfffffffb0000000f0000000affffffdc",
            INIT_23 => X"0000003a0000000400000005000000080000000a0000001cffffffe9fffffff4",
            INIT_24 => X"ffffffff0000001c000000280000000bfffffffd0000000cffffffdffffffffe",
            INIT_25 => X"fffffffbffffffedfffffff9fffffff500000036000000250000004500000040",
            INIT_26 => X"00000003ffffffff0000001d00000001ffffffd6ffffffefffffffeffffffff8",
            INIT_27 => X"ffffffe9fffffff60000002b0000001c00000004000000190000003300000004",
            INIT_28 => X"ffffffecffffffc4fffffff4ffffffe8ffffffd5ffffffd9ffffffcd0000001b",
            INIT_29 => X"00000000fffffffafffffff40000003300000015fffffff50000001900000015",
            INIT_2A => X"000000220000002bfffffffcfffffff80000001bffffffe8fffffff6fffffff8",
            INIT_2B => X"00000010ffffffe8fffffff50000000dffffffec000000030000000600000037",
            INIT_2C => X"fffffff1ffffffe6fffffffafffffffd0000000900000004000000170000000e",
            INIT_2D => X"000000080000001200000014fffffffe000000260000000fffffffef0000000a",
            INIT_2E => X"fffffff700000023ffffffec00000000fffffff60000001d0000000d00000012",
            INIT_2F => X"ffffffe0fffffff00000001700000045000000320000002f0000001900000009",
            INIT_30 => X"fffffff0fffffff4000000300000003800000037000000070000003f0000003e",
            INIT_31 => X"0000000d0000002dffffffc6ffffffd000000015ffffffc5ffffffe5fffffff7",
            INIT_32 => X"fffffff1ffffffc4ffffffc3ffffffd7ffffffcfffffffe8ffffffbc00000001",
            INIT_33 => X"ffffffebffffffc2ffffffe900000032fffffff1fffffff2fffffff30000002f",
            INIT_34 => X"0000002c00000001fffffff300000031000000090000000effffffecffffffe6",
            INIT_35 => X"ffffffcf00000000ffffffcc00000021ffffffdbffffffe400000023fffffff6",
            INIT_36 => X"ffffffda00000003000000000000000ffffffff3fffffff9ffffffe3ffffffc8",
            INIT_37 => X"ffffffcdffffffeaffffffb0ffffffa800000010ffffffe0fffffffb0000000a",
            INIT_38 => X"0000002d00000018fffffff900000005ffffffe8ffffffc20000000fffffffc3",
            INIT_39 => X"fffffffb0000001a000000370000001600000024fffffff9ffffffe6ffffffed",
            INIT_3A => X"ffffffd00000000a000000030000001c00000007000000040000002100000010",
            INIT_3B => X"ffffffe300000034fffffff0ffffffbcffffffe4ffffffbdffffffeeffffffe4",
            INIT_3C => X"ffffffe200000007ffffffe8ffffffea00000012ffffffdd000000090000000c",
            INIT_3D => X"000000000000003c0000000100000020000000430000000300000014ffffffe4",
            INIT_3E => X"0000002600000003ffffffd50000001fffffffed0000000000000039fffffffb",
            INIT_3F => X"ffffffb10000000effffffd4ffffffe80000002a0000001e00000021fffffffb",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE7;


    MEM_IWGHT_LAYER2_INSTANCE8 : if BRAM_NAME = "iwght_layer2_instance8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffba00000009ffffffdbffffff9a0000001cffffffe2fffffffd0000001d",
            INIT_01 => X"fffffffb0000001efffffffdffffffe2fffffffbfffffff6ffffffe7fffffff4",
            INIT_02 => X"00000023ffffffddfffffff5fffffffbffffffe7ffffffe600000000fffffff1",
            INIT_03 => X"00000016000000340000001f000000160000005300000032ffffffe600000046",
            INIT_04 => X"00000000ffffffec00000016ffffffd1ffffffd500000029fffffff100000018",
            INIT_05 => X"ffffffaaffffffe0ffffffb7ffffffa800000020ffffffb6fffffff90000001d",
            INIT_06 => X"ffffffd600000018ffffffe0ffffffdb00000001ffffffdfffffffe7ffffffa4",
            INIT_07 => X"ffffff8effffffb90000005dffffffa7000000070000002f0000003bffffffe4",
            INIT_08 => X"00000019fffffff90000003700000016ffffffdeffffffc2ffffff8500000021",
            INIT_09 => X"ffffffdd0000001e00000021ffffffd70000002a000000310000000500000028",
            INIT_0A => X"0000003f00000024fffffff30000005400000043fffffff80000005a0000003c",
            INIT_0B => X"ffffffff00000011fffffff90000001dffffffe4000000300000001cffffffee",
            INIT_0C => X"000000130000001700000008ffffffebfffffff7ffffffe0fffffffe00000008",
            INIT_0D => X"ffffffb8ffffffc0fffffffaffffffd0ffffffd700000023ffffffb50000000a",
            INIT_0E => X"00000019ffffffe800000000ffffffe900000002fffffff1ffffffd20000000f",
            INIT_0F => X"00000012fffffff3fffffffc00000027fffffff4ffffffecffffffec0000000a",
            INIT_10 => X"0000001efffffff20000001b0000000dfffffff5ffffffe800000004fffffffd",
            INIT_11 => X"0000001200000010ffffffd8fffffffc0000001d000000240000001700000037",
            INIT_12 => X"fffffffd0000001b00000031000000390000000a000000390000001700000018",
            INIT_13 => X"ffffffec0000001d000000070000004700000052000000230000003c00000040",
            INIT_14 => X"ffffffe2ffffffe400000022000000230000000400000019000000010000001e",
            INIT_15 => X"00000027ffffffb3fffffff2fffffff8ffffffeeffffffd60000001500000010",
            INIT_16 => X"0000001afffffffbfffffff4000000480000000a0000002a000000470000001a",
            INIT_17 => X"ffffff9cffffffb1ffffffb3ffffffbeffffffc30000000dffffffe8ffffffd6",
            INIT_18 => X"0000002afffffff6fffffffc00000021ffffffe1ffffffe8fffffffeffffffe0",
            INIT_19 => X"ffffff84ffffff6bffffff82ffffffc6ffffffe6ffffffc00000001200000031",
            INIT_1A => X"0000000200000001ffffffecffffffe1ffffffe5ffffff6affffff53ffffff67",
            INIT_1B => X"ffffffc600000000ffffffddffffffd800000032000000150000001affffffeb",
            INIT_1C => X"fffffffe000000010000000effffffabffffff9dffffffefffffff8dffffffa4",
            INIT_1D => X"ffffffee0000000e000000350000002f00000018000000230000003d00000005",
            INIT_1E => X"0000000b0000000c0000002200000000fffffff2000000100000002200000006",
            INIT_1F => X"ffffffeeffffffe0ffffffcd000000170000002bffffffccfffffff100000034",
            INIT_20 => X"0000002000000000ffffffe8fffffffefffffff10000000f00000000ffffffee",
            INIT_21 => X"ffffffe3fffffff2fffffff0ffffffd1ffffffa8ffffffdfffffffd20000001a",
            INIT_22 => X"ffffffddffffffeeffffffdbffffffd0ffffffdbffffffd4ffffffeffffffff2",
            INIT_23 => X"ffffffe9ffffffdeffffffddffffffc0ffffffed00000000ffffffedfffffff3",
            INIT_24 => X"000000160000000c00000009fffffffffffffffdffffffeeffffffd8fffffff1",
            INIT_25 => X"0000001a00000009fffffff4000000220000000d0000000b0000000400000000",
            INIT_26 => X"ffffffe2000000110000001d00000021000000070000000dffffffff00000012",
            INIT_27 => X"fffffff800000007000000150000001afffffffb0000000cfffffff5ffffffee",
            INIT_28 => X"ffffffddffffffefffffffdfffffffeafffffff70000000600000019ffffffe2",
            INIT_29 => X"fffffff8ffffffe7fffffff8ffffffeefffffff3ffffffe90000000dfffffff5",
            INIT_2A => X"fffffff6000000200000000600000007ffffffe8ffffffecffffffeeffffffec",
            INIT_2B => X"ffffffe70000000effffffe1ffffffe6fffffffeffffffe00000001300000022",
            INIT_2C => X"ffffffebffffffe6ffffffbdffffffc2ffffffd6fffffffdffffffe7fffffff8",
            INIT_2D => X"0000002c0000000e00000037000000140000000e00000002ffffffc7ffffffff",
            INIT_2E => X"fffffff2fffffff9fffffffe0000000d00000006000000340000001900000028",
            INIT_2F => X"0000000400000005fffffff800000009ffffffd7fffffff9ffffffecffffffeb",
            INIT_30 => X"000000280000000b0000000e0000001cffffffffffffffe90000000dfffffff7",
            INIT_31 => X"fffffff0fffffffc00000022fffffff50000001d000000260000001700000019",
            INIT_32 => X"ffffffb2ffffffcfffffffefffffffe2fffffffbffffffe3ffffffecfffffff9",
            INIT_33 => X"0000003d00000014fffffff400000001fffffff6ffffffeefffffff4ffffffc3",
            INIT_34 => X"00000016ffffffddffffffdc00000017ffffffdf0000000fffffffef00000012",
            INIT_35 => X"ffffffebfffffffc000000110000000f000000150000001b00000006ffffffe5",
            INIT_36 => X"ffffffc3ffffffadffffffeffffffff30000002800000006000000170000000e",
            INIT_37 => X"00000002fffffff9fffffff3ffffffe800000005ffffffe0ffffffd2ffffffee",
            INIT_38 => X"fffffffcffffffd4ffffffbaffffffd2ffffff88fffffffeffffffe9ffffffbd",
            INIT_39 => X"ffffffe2fffffffcffffffccfffffff100000000ffffffcdffffffd200000002",
            INIT_3A => X"ffffffe1ffffffc9ffffffc0ffffffdbffffffbdffffffb10000003900000029",
            INIT_3B => X"ffffffbdffffffccffffffe2ffffffcdffffffc5fffffffaffffffe1ffffffde",
            INIT_3C => X"0000000000000013ffffffed0000001a0000002000000020ffffffeeffffffed",
            INIT_3D => X"fffffffbffffffedffffffe40000001300000006fffffff900000002fffffff1",
            INIT_3E => X"000000010000001700000029ffffffe10000001f0000000b00000000fffffff2",
            INIT_3F => X"0000000900000016fffffff30000000d0000001500000016000000130000002c",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE8;


    MEM_IWGHT_LAYER2_INSTANCE9 : if BRAM_NAME = "iwght_layer2_instance9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffadffffffed0000000500000027000000170000000f000000010000001a",
            INIT_01 => X"0000001600000019000000190000001a00000011fffffff20000000dfffffffd",
            INIT_02 => X"00000023fffffff0fffffff8ffffffbefffffff80000000cffffffd700000024",
            INIT_03 => X"00000013000000030000002c0000003b000000170000002dffffffd30000000f",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE9;


    MEM_IFMAP_LAYER0_INSTANCE0 : if BRAM_NAME = "ifmap_layer0_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000009f000000a20000009c000000a0000000a6000000a50000009f0000009e",
            INIT_01 => X"000000aa000000a9000000a6000000a1000000a0000000a10000009f0000009e",
            INIT_02 => X"0000009400000096000000950000009c000000a0000000a0000000a2000000a7",
            INIT_03 => X"000000740000007e000000890000008f0000008d0000008c0000008f00000095",
            INIT_04 => X"000000a2000000a4000000a0000000a2000000a60000009f0000009700000098",
            INIT_05 => X"000000ab000000ab000000aa000000a30000009f0000009b0000009c000000a3",
            INIT_06 => X"0000008d0000008c0000008b00000091000000970000009a000000a0000000a9",
            INIT_07 => X"000000770000007d000000880000008f0000008e000000910000009300000095",
            INIT_08 => X"000000a5000000a5000000a3000000a0000000a70000009e0000009700000097",
            INIT_09 => X"000000a9000000a7000000a6000000a10000009d0000009e000000a2000000a3",
            INIT_0A => X"0000007200000065000000620000006e00000079000000910000009f000000aa",
            INIT_0B => X"00000078000000820000008b0000008e0000008c0000008f0000008600000078",
            INIT_0C => X"000000a9000000a9000000a7000000a7000000ae000000a00000009b0000009b",
            INIT_0D => X"000000a4000000a20000009d000000b1000000bf000000a7000000a5000000a5",
            INIT_0E => X"0000004a000000500000005c000000620000006700000068000000950000009e",
            INIT_0F => X"0000007f000000880000008c0000008c00000084000000710000005300000056",
            INIT_10 => X"000000a6000000a9000000a3000000a9000000aa000000a10000009c0000009b",
            INIT_11 => X"0000008e0000009200000097000000c3000000f6000000ad000000a4000000a4",
            INIT_12 => X"0000005d000000610000006a0000007000000071000000550000004e0000006f",
            INIT_13 => X"00000081000000850000008a000000800000006900000055000000540000004a",
            INIT_14 => X"000000a7000000a7000000a5000000a100000093000000820000008500000094",
            INIT_15 => X"0000004200000061000000800000009d000000b4000000a3000000a5000000a3",
            INIT_16 => X"0000005e00000072000000770000007a00000076000000590000004200000045",
            INIT_17 => X"000000860000008a0000008c0000006c000000430000003a0000005b00000063",
            INIT_18 => X"000000aa000000a8000000aa00000099000000580000002f0000006d0000007f",
            INIT_19 => X"00000044000000640000007f0000008100000093000000a4000000a6000000a9",
            INIT_1A => X"0000006b000000690000007c000000920000008400000053000000480000004e",
            INIT_1B => X"000000860000008d000000840000004f0000002e0000003f0000005500000073",
            INIT_1C => X"000000a8000000a5000000a70000008f000000460000002a0000006300000083",
            INIT_1D => X"00000058000000740000009000000082000000780000008c000000a1000000ab",
            INIT_1E => X"0000006a0000006600000088000000a30000007c0000004d000000550000005b",
            INIT_1F => X"000000880000008a0000006b0000003900000031000000360000005500000064",
            INIT_20 => X"000000a6000000a3000000a1000000990000007c0000003600000067000000aa",
            INIT_21 => X"00000056000000790000009c0000009d0000007d00000071000000ae000000a5",
            INIT_22 => X"0000005700000071000000920000008a00000051000000500000005400000052",
            INIT_23 => X"00000089000000850000004a0000002800000038000000470000005600000053",
            INIT_24 => X"000000990000009c0000009e000000ae0000009a0000005e00000086000000b4",
            INIT_25 => X"0000005d0000007d00000094000000ae0000009c000000cf000000ed000000cf",
            INIT_26 => X"0000006a000000850000008f000000890000004c0000003b0000004a00000056",
            INIT_27 => X"000000840000005f00000028000000320000004b000000540000005700000056",
            INIT_28 => X"0000007a0000009f0000009b000000b1000000a50000008e0000006c000000b7",
            INIT_29 => X"000000780000007d0000009c000000b7000000a4000000dc000000ed000000d5",
            INIT_2A => X"0000006b0000009b0000009d000000af0000005b0000002d000000500000004e",
            INIT_2B => X"000000680000003b000000290000003b0000004e000000580000006700000057",
            INIT_2C => X"00000086000000ad000000a6000000bb000000aa0000008700000064000000bc",
            INIT_2D => X"0000007500000086000000bd000000b9000000aa000000c7000000c200000075",
            INIT_2E => X"0000005d00000092000000a0000000d20000007d000000260000005400000066",
            INIT_2F => X"0000004c0000003e000000370000004900000055000000680000005e00000053",
            INIT_30 => X"0000009f000000b2000000a6000000ae000000af0000007f0000005a000000bd",
            INIT_31 => X"0000007b000000a0000000d8000000ba00000089000000a8000000a800000061",
            INIT_32 => X"0000005b0000007b0000009b000000c200000096000000320000007300000078",
            INIT_33 => X"000000490000004f0000004900000054000000560000005f0000005400000054",
            INIT_34 => X"000000a7000000ad0000008800000077000000b9000000980000005d000000bd",
            INIT_35 => X"0000008d000000b4000000e2000000bd000000a7000000910000009300000067",
            INIT_36 => X"000000570000007200000095000000ba0000009a00000047000000750000007e",
            INIT_37 => X"0000005e000000610000005a0000006400000063000000500000004800000050",
            INIT_38 => X"000000a70000009c0000006300000069000000ba000000a80000006c000000c2",
            INIT_39 => X"0000009a00000091000000ac000000be000000c60000008a0000007300000064",
            INIT_3A => X"0000006e0000008200000089000000b300000098000000470000006700000092",
            INIT_3B => X"000000750000006100000064000000730000006d0000005f0000005b00000055",
            INIT_3C => X"0000009b0000008c0000004e00000082000000b8000000ac00000084000000c5",
            INIT_3D => X"000000830000008700000091000000f2000000e60000008f0000008200000073",
            INIT_3E => X"000000570000007000000098000000a8000000900000005f0000006c00000079",
            INIT_3F => X"0000008800000079000000670000007800000070000000690000005700000047",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE0;


    MEM_IFMAP_LAYER0_INSTANCE1 : if BRAM_NAME = "ifmap_layer0_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000008a0000007e0000004e000000a8000000bf000000a800000092000000cb",
            INIT_01 => X"00000071000000710000008c000000a2000000ad0000009a000000600000008a",
            INIT_02 => X"0000006d00000087000000940000009c000000ab000000700000006900000065",
            INIT_03 => X"00000090000000970000007d0000006b000000650000005e0000004f0000004e",
            INIT_04 => X"0000009c000000600000005e000000b0000000b7000000a4000000a3000000d6",
            INIT_05 => X"0000007300000066000000740000007200000076000000810000006a00000094",
            INIT_06 => X"0000004b00000085000000800000004400000076000000900000006500000056",
            INIT_07 => X"0000008c000000960000008f0000007400000066000000470000003a0000003c",
            INIT_08 => X"0000008d000000560000007c000000b0000000ad000000a7000000b2000000d4",
            INIT_09 => X"00000093000000810000007c000000860000004d000000680000008700000099",
            INIT_0A => X"000000400000004b0000006b0000007500000084000000960000005c00000055",
            INIT_0B => X"000000970000009a000000a00000009b0000008500000056000000410000002c",
            INIT_0C => X"000000770000005600000090000000b1000000ae000000ab000000bb000000c7",
            INIT_0D => X"000000b8000000910000006c000000810000004600000090000000890000007a",
            INIT_0E => X"0000003400000033000000590000008600000089000000830000004900000074",
            INIT_0F => X"000000950000009e000000a4000000ab000000a3000000790000005a0000002f",
            INIT_10 => X"000000830000006300000098000000b5000000b1000000b3000000c3000000a5",
            INIT_11 => X"000000bf000000b20000007a0000005d000000500000005d00000067000000ab",
            INIT_12 => X"00000018000000260000002e0000003c00000057000000590000006400000096",
            INIT_13 => X"000000780000007f0000008000000090000000900000006c0000003c0000002e",
            INIT_14 => X"00000096000000530000008a000000b5000000b2000000b1000000c300000075",
            INIT_15 => X"000000c2000000be000000b0000000950000008600000085000000db000000f5",
            INIT_16 => X"0000003a0000003100000022000000230000003d0000006e0000007d000000a8",
            INIT_17 => X"000000370000003b000000450000004e00000048000000450000003a0000003d",
            INIT_18 => X"000000d30000006d0000008c000000b1000000b0000000ae000000af0000004f",
            INIT_19 => X"0000007a000000740000007c000000720000007c000000d0000000fc000000fd",
            INIT_1A => X"000000380000003300000032000000340000003c000000440000004400000068",
            INIT_1B => X"0000002a0000002b000000300000003b000000330000002b0000003300000038",
            INIT_1C => X"000000f6000000a5000000a5000000b2000000a8000000900000006000000029",
            INIT_1D => X"000000300000003100000031000000350000003c0000006e000000e3000000fd",
            INIT_1E => X"0000002b0000002e0000002e000000260000002a0000002e0000002a0000002d",
            INIT_1F => X"0000002d000000330000003500000037000000320000002e0000002e0000002a",
            INIT_20 => X"000000fe000000c200000084000000a6000000830000003b0000001d0000001d",
            INIT_21 => X"00000032000000310000003300000032000000320000003d0000008d000000f1",
            INIT_22 => X"0000002a00000026000000270000002300000022000000270000002a0000002f",
            INIT_23 => X"000000330000002e00000032000000380000003b0000003e000000380000002d",
            INIT_24 => X"00000100000000d7000000800000008000000049000000220000001e00000030",
            INIT_25 => X"0000002d0000002e0000003400000034000000320000003600000042000000bb",
            INIT_26 => X"0000002e0000002b00000028000000280000002700000024000000290000002b",
            INIT_27 => X"000000530000004600000032000000360000003b000000400000003e0000003b",
            INIT_28 => X"000000f0000000e00000008000000042000000290000001f0000002300000034",
            INIT_29 => X"0000002f0000002c0000002c0000003600000038000000310000003a0000007c",
            INIT_2A => X"0000003a000000360000002d0000002c0000002c0000002b0000002b0000002e",
            INIT_2B => X"0000004c000000550000004900000033000000240000002b0000002e00000036",
            INIT_2C => X"000000d3000000ca0000004e0000002c000000230000001d0000002300000032",
            INIT_2D => X"0000002d00000028000000300000003a00000030000000360000004100000061",
            INIT_2E => X"000000300000002700000027000000330000002e0000002f000000300000002f",
            INIT_2F => X"000000330000002e0000004300000043000000280000001c000000270000002f",
            INIT_30 => X"000000aa000000680000002e0000002900000021000000200000002300000032",
            INIT_31 => X"0000002d000000360000003a0000003d00000035000000340000003600000040",
            INIT_32 => X"00000027000000280000002a0000002e000000310000002e000000290000002a",
            INIT_33 => X"000000330000000f0000001f0000002f0000003f0000002c0000002800000025",
            INIT_34 => X"000000470000002a0000002b00000025000000260000001f0000002a00000044",
            INIT_35 => X"000000350000003a0000003800000031000000260000001b0000001f00000031",
            INIT_36 => X"00000021000000270000002d0000003200000035000000390000003c00000038",
            INIT_37 => X"000000280000000d0000002600000038000000490000004f0000003e0000002a",
            INIT_38 => X"000000280000002c0000002a000000270000002b00000023000000310000003d",
            INIT_39 => X"0000002f000000240000001d0000001b0000001e000000170000001b0000002a",
            INIT_3A => X"0000002b0000002b00000031000000450000004b000000420000003e00000038",
            INIT_3B => X"000000140000001d0000001a0000003c0000005d0000006d000000550000003c",
            INIT_3C => X"000000260000002800000028000000280000002b0000002d0000003800000036",
            INIT_3D => X"00000012000000130000001d000000190000001d000000160000001a00000024",
            INIT_3E => X"0000002d0000003400000035000000420000004a0000003d0000002f00000020",
            INIT_3F => X"0000001500000022000000180000003000000059000000690000005900000043",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE1;


    MEM_IFMAP_LAYER0_INSTANCE2 : if BRAM_NAME = "ifmap_layer0_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000071000000730000006d0000007000000076000000740000006f00000070",
            INIT_01 => X"0000007700000075000000750000006f0000006f00000074000000710000006f",
            INIT_02 => X"0000006a0000006b0000006b0000006d000000700000006f0000007100000075",
            INIT_03 => X"000000550000005b0000005f000000610000006100000062000000650000006b",
            INIT_04 => X"0000007200000075000000710000007000000074000000720000006e00000070",
            INIT_05 => X"000000730000007500000077000000710000006e0000006f0000006e00000074",
            INIT_06 => X"0000006400000066000000680000006e00000073000000700000006f00000073",
            INIT_07 => X"000000580000005b0000005f0000006200000061000000660000006600000069",
            INIT_08 => X"0000007500000075000000730000006a0000006f0000006f0000006d0000006e",
            INIT_09 => X"0000007100000072000000730000006f0000006d000000720000007300000073",
            INIT_0A => X"000000550000004d0000004e0000005a000000600000006f0000007200000074",
            INIT_0B => X"000000590000005f000000620000006300000063000000670000006000000056",
            INIT_0C => X"0000007700000078000000750000006e000000700000006d0000006e0000006b",
            INIT_0D => X"00000072000000730000006f00000082000000920000007b0000007500000073",
            INIT_0E => X"0000003f0000004b0000005a0000005a00000057000000500000006f00000070",
            INIT_0F => X"0000005e00000063000000650000006600000062000000550000003e00000046",
            INIT_10 => X"000000740000007800000071000000720000007200000073000000720000006b",
            INIT_11 => X"0000006c0000006f000000720000009c000000d6000000800000007400000071",
            INIT_12 => X"0000005e00000066000000720000006e00000067000000450000003500000050",
            INIT_13 => X"0000005d0000005e000000650000006000000053000000490000004e00000048",
            INIT_14 => X"000000730000007400000071000000730000007000000064000000680000006d",
            INIT_15 => X"000000320000004b000000660000007a0000008a00000076000000740000006f",
            INIT_16 => X"00000060000000740000007a000000790000007100000053000000380000003a",
            INIT_17 => X"0000005f0000006200000069000000540000003a0000003a0000005b00000064",
            INIT_18 => X"000000760000007300000076000000750000004a000000250000005f00000064",
            INIT_19 => X"00000043000000570000006c000000620000006b000000780000007400000075",
            INIT_1A => X"0000006600000063000000760000008e00000082000000540000004b00000053",
            INIT_1B => X"0000005d00000063000000620000003d0000002f00000047000000530000006f",
            INIT_1C => X"0000007400000072000000750000006f000000400000002b0000006000000073",
            INIT_1D => X"000000570000006a000000830000006e0000005e0000006d0000007100000077",
            INIT_1E => X"000000620000005d0000007c00000099000000760000004d000000580000005f",
            INIT_1F => X"0000006100000067000000530000002f000000350000003c000000510000005d",
            INIT_20 => X"0000007a00000075000000710000007c000000790000003a00000069000000a1",
            INIT_21 => X"000000500000006f0000008f0000008d00000069000000590000008700000079",
            INIT_22 => X"0000004f00000067000000870000007d000000470000004e0000005500000051",
            INIT_23 => X"000000670000006a0000003b000000230000003900000049000000520000004d",
            INIT_24 => X"000000760000007400000074000000950000009a000000640000008b000000b0",
            INIT_25 => X"000000550000006e000000830000009900000083000000b4000000d6000000b4",
            INIT_26 => X"000000620000007c000000850000007d00000044000000390000004a00000054",
            INIT_27 => X"000000670000004b0000001e000000310000004c000000550000005500000051",
            INIT_28 => X"0000005900000076000000700000009c000000a90000009700000074000000b7",
            INIT_29 => X"0000006f0000006c000000890000009f00000087000000bf000000e0000000c5",
            INIT_2A => X"000000640000009300000093000000a5000000550000002c000000500000004c",
            INIT_2B => X"000000510000002e000000240000003b0000004f000000580000006600000053",
            INIT_2C => X"0000005d0000007b00000078000000a7000000af000000900000006c000000bf",
            INIT_2D => X"0000006b00000077000000ab000000a10000008e000000ab000000b60000005f",
            INIT_2E => X"000000590000008b00000098000000c900000079000000260000005400000062",
            INIT_2F => X"0000003800000037000000350000004b00000057000000680000005d00000050",
            INIT_30 => X"0000006d0000007b0000007b0000009c000000b40000008600000060000000c2",
            INIT_31 => X"0000007100000095000000ca000000a600000072000000900000009a00000044",
            INIT_32 => X"000000580000007600000095000000bb00000093000000320000007200000072",
            INIT_33 => X"000000370000004a0000004900000057000000570000005f0000005400000053",
            INIT_34 => X"000000740000007c0000006a0000006e000000bc0000009a0000005f000000c0",
            INIT_35 => X"00000083000000ac000000d8000000ae000000950000007d0000008400000048",
            INIT_36 => X"000000550000006e00000090000000b500000098000000470000007200000075",
            INIT_37 => X"0000004900000059000000580000006500000064000000500000004900000050",
            INIT_38 => X"0000007a00000077000000590000006d000000ba000000a70000006b000000c4",
            INIT_39 => X"0000008f0000008c000000a5000000b4000000b90000007b0000006a0000004a",
            INIT_3A => X"0000006d0000008000000085000000af00000098000000470000006400000088",
            INIT_3B => X"0000005f0000005500000060000000740000006e000000600000005d00000056",
            INIT_3C => X"0000007d000000780000005300000089000000b2000000a700000081000000c5",
            INIT_3D => X"00000079000000820000008a000000ec000000dd00000083000000780000005e",
            INIT_3E => X"000000550000006c000000930000009f00000086000000580000006800000070",
            INIT_3F => X"0000006800000060000000560000006e0000006d000000680000005800000048",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE2;


    MEM_IFMAP_LAYER0_INSTANCE3 : if BRAM_NAME = "ifmap_layer0_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000007e0000007d00000056000000aa000000b6000000a400000092000000cb",
            INIT_01 => X"0000006a0000006a0000008400000098000000a30000008f0000005000000079",
            INIT_02 => X"00000069000000820000008d0000008a0000008f0000005a0000006500000065",
            INIT_03 => X"000000680000006c00000058000000530000005b0000005d0000004f0000004c",
            INIT_04 => X"000000950000006000000066000000b6000000b8000000a7000000a6000000d7",
            INIT_05 => X"0000006e0000005b000000690000006600000069000000740000005d00000089",
            INIT_06 => X"000000450000007e00000078000000380000006000000080000000670000005b",
            INIT_07 => X"0000006e00000074000000700000005e0000005d000000460000003800000038",
            INIT_08 => X"0000008b0000005800000083000000b8000000b5000000af000000b8000000d3",
            INIT_09 => X"0000008f000000750000006f00000079000000400000005a0000008000000094",
            INIT_0A => X"0000003b00000044000000630000006d000000750000008b000000600000005c",
            INIT_0B => X"0000006f00000073000000780000007700000069000000450000003e00000029",
            INIT_0C => X"000000790000005a00000095000000b6000000b3000000b0000000bd000000c0",
            INIT_0D => X"000000b00000008600000061000000760000003b00000086000000880000007c",
            INIT_0E => X"000000330000003100000056000000810000007c000000770000004b00000076",
            INIT_0F => X"0000006b0000006f0000007100000079000000760000005b0000005a00000031",
            INIT_10 => X"00000087000000670000009d000000b5000000ad000000b2000000c10000009c",
            INIT_11 => X"000000b6000000ad000000760000005a0000004d0000005a00000069000000af",
            INIT_12 => X"000000210000002e000000340000003d0000004d0000004e0000006400000094",
            INIT_13 => X"00000069000000710000006d0000007b0000007d000000640000004700000039",
            INIT_14 => X"000000990000005700000090000000b3000000a9000000b2000000c800000078",
            INIT_15 => X"000000c0000000c4000000b60000009c0000008d0000008c000000de000000f7",
            INIT_16 => X"000000510000004600000036000000310000003e0000006d00000085000000ac",
            INIT_17 => X"0000005a0000005c000000600000006800000065000000630000005400000055",
            INIT_18 => X"000000d30000007000000092000000b1000000ac000000b7000000c500000069",
            INIT_19 => X"00000085000000850000008d000000840000008f000000e0000000fd000000fc",
            INIT_1A => X"0000005d00000055000000540000005400000052000000570000005d0000007c",
            INIT_1B => X"0000005f00000061000000610000006c00000068000000600000005b0000005e",
            INIT_1C => X"000000f5000000a6000000aa000000b6000000ae000000a80000008900000059",
            INIT_1D => X"000000480000004b0000004c000000500000005800000088000000e7000000fb",
            INIT_1E => X"00000057000000590000005a000000560000005200000051000000510000004f",
            INIT_1F => X"0000005a0000005f0000005e00000060000000600000005e0000005d00000059",
            INIT_20 => X"000000fa000000bd00000088000000b30000009900000066000000570000005b",
            INIT_21 => X"00000054000000530000005500000054000000540000005e0000009f000000f5",
            INIT_22 => X"000000590000005500000056000000530000004f000000520000005400000056",
            INIT_23 => X"000000670000005e00000063000000660000006500000067000000670000005c",
            INIT_24 => X"000000fd000000d500000088000000940000006a000000550000005e0000006f",
            INIT_25 => X"00000052000000530000005a0000005a000000580000005b0000005d000000c6",
            INIT_26 => X"0000005f0000005c000000590000005600000053000000500000005100000052",
            INIT_27 => X"000000890000007b000000690000006c0000006c0000006d0000006e0000006c",
            INIT_28 => X"000000f5000000e5000000910000005f00000053000000560000006300000072",
            INIT_29 => X"0000005300000052000000520000005c0000005e000000570000005c0000008f",
            INIT_2A => X"0000006e0000006a000000610000005a00000058000000560000005300000054",
            INIT_2B => X"0000007d0000008a000000820000006c0000005b0000005f0000006100000069",
            INIT_2C => X"000000e4000000db0000006a000000530000005600000059000000620000006e",
            INIT_2D => X"00000052000000500000005700000061000000570000005e000000680000007e",
            INIT_2E => X"000000660000005d0000005c0000006100000059000000590000005700000054",
            INIT_2F => X"00000060000000620000007e0000008100000065000000550000005d00000065",
            INIT_30 => X"000000c5000000850000005400000058000000580000005c000000610000006c",
            INIT_31 => X"000000530000006000000064000000670000005f0000005e0000006100000064",
            INIT_32 => X"0000005c0000005d0000005f0000005c0000005c00000058000000500000004f",
            INIT_33 => X"0000005d0000003c0000005a0000006e0000007d000000660000005d0000005a",
            INIT_34 => X"0000006b0000004f00000059000000570000005b00000058000000640000007c",
            INIT_35 => X"0000005c00000066000000640000005d00000052000000470000004d00000059",
            INIT_36 => X"00000053000000580000005e0000005f0000006100000063000000630000005e",
            INIT_37 => X"000000550000004000000061000000740000008300000084000000700000005b",
            INIT_38 => X"00000051000000580000005c0000005a0000005b000000550000006600000074",
            INIT_39 => X"000000560000005000000049000000470000004a000000430000004800000055",
            INIT_3A => X"00000058000000580000005f00000071000000770000006d000000650000005f",
            INIT_3B => X"00000040000000520000005200000073000000910000009c0000008200000069",
            INIT_3C => X"00000051000000570000005c000000590000005600000059000000690000006b",
            INIT_3D => X"0000003a0000003f00000049000000450000004900000042000000450000004f",
            INIT_3E => X"000000570000005f000000600000006f00000077000000680000005700000046",
            INIT_3F => X"00000043000000540000004d000000630000008700000092000000830000006d",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE3;


    MEM_IFMAP_LAYER0_INSTANCE4 : if BRAM_NAME = "ifmap_layer0_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002d0000002f000000290000002e00000035000000330000002f00000031",
            INIT_01 => X"0000002c0000002d00000029000000310000003400000029000000290000002c",
            INIT_02 => X"0000002b0000002d0000002d0000002c0000002b000000270000002600000028",
            INIT_03 => X"00000021000000240000002400000026000000290000002b000000270000002c",
            INIT_04 => X"0000002d0000002f0000002b00000031000000380000002d0000002800000033",
            INIT_05 => X"000000210000002800000029000000340000003600000029000000260000002e",
            INIT_06 => X"000000300000003400000037000000350000003200000029000000210000001e",
            INIT_07 => X"00000022000000200000001f00000022000000260000002d0000002e00000032",
            INIT_08 => X"0000002d0000002d0000002c0000002a0000003000000024000000210000002f",
            INIT_09 => X"0000002300000025000000260000003300000039000000300000002b0000002b",
            INIT_0A => X"000000320000002f000000320000003400000031000000360000002f00000027",
            INIT_0B => X"0000002100000022000000220000002300000027000000330000003700000030",
            INIT_0C => X"00000030000000300000002e0000002b0000002c0000001f0000002000000028",
            INIT_0D => X"000000360000002f000000290000004b0000005f000000390000002d0000002c",
            INIT_0E => X"0000003200000042000000540000004c000000410000002f000000430000003a",
            INIT_0F => X"0000002400000027000000270000002b0000002e0000002d0000002700000034",
            INIT_10 => X"0000002c0000002f000000280000002b0000002f000000310000003000000029",
            INIT_11 => X"000000470000003c000000380000006b000000a40000003b0000002a00000029",
            INIT_12 => X"0000005d00000069000000760000006f00000062000000380000001f00000032",
            INIT_13 => X"00000024000000240000002e000000300000002d0000002f0000004600000043",
            INIT_14 => X"0000002900000029000000270000002c00000035000000390000004000000036",
            INIT_15 => X"0000001f0000002b0000003a0000004e000000550000002a0000002700000025",
            INIT_16 => X"00000060000000740000007a000000780000006e0000004c0000002d0000002b",
            INIT_17 => X"000000280000002c0000003a00000031000000250000002f0000005600000061",
            INIT_18 => X"0000002b000000280000002b000000300000001c000000110000005000000039",
            INIT_19 => X"00000039000000460000004b0000003b0000003400000027000000250000002a",
            INIT_1A => X"0000005e0000005a0000006c00000084000000790000004a0000004000000048",
            INIT_1B => X"00000027000000300000003a0000002400000027000000450000004d00000067",
            INIT_1C => X"00000027000000240000002a0000003800000029000000260000005c0000005a",
            INIT_1D => X"0000004f0000005d0000006b0000004d00000031000000330000003300000031",
            INIT_1E => X"0000005800000051000000700000008c0000006b000000450000005200000058",
            INIT_1F => X"00000027000000330000003200000020000000310000003a0000004a00000054",
            INIT_20 => X"00000032000000290000002b00000052000000710000003b0000006900000090",
            INIT_21 => X"0000004a0000006500000080000000790000004e0000003b0000005f00000042",
            INIT_22 => X"000000460000005d0000007b000000700000003d00000049000000520000004d",
            INIT_23 => X"0000002d0000003b000000230000001b00000035000000430000004c00000045",
            INIT_24 => X"0000003c0000002f000000330000007000000095000000690000008f000000a3",
            INIT_25 => X"0000004f0000006b0000007d0000009100000077000000a6000000c600000092",
            INIT_26 => X"00000059000000720000007a000000700000003a00000035000000470000004f",
            INIT_27 => X"000000390000002c0000000f0000002b000000470000004e0000004e0000004a",
            INIT_28 => X"0000002f00000033000000320000007a000000a80000009e0000007a000000af",
            INIT_29 => X"0000006800000068000000840000009b00000083000000bc000000e2000000b3",
            INIT_2A => X"0000005c0000008a000000890000009a0000004d000000280000004d00000045",
            INIT_2B => X"0000002e0000001f000000210000003b000000490000004f000000600000004d",
            INIT_2C => X"0000002c000000370000003b00000088000000b20000009900000074000000bd",
            INIT_2D => X"0000005f0000006a0000009f0000009700000085000000a4000000bc00000050",
            INIT_2E => X"00000052000000820000008e000000c000000071000000220000004f00000059",
            INIT_2F => X"0000001a00000030000000370000004e000000510000005e000000580000004b",
            INIT_30 => X"0000002f000000350000004400000085000000b90000009000000069000000c2",
            INIT_31 => X"0000006200000081000000b7000000940000005e0000007e000000980000002c",
            INIT_32 => X"000000530000006f0000008c000000b20000008c0000002f0000006d00000069",
            INIT_33 => X"000000180000004000000049000000590000005100000055000000500000004f",
            INIT_34 => X"000000320000003a0000004200000062000000c0000000a300000067000000c1",
            INIT_35 => X"000000750000009d000000c80000009b0000007f000000670000007800000027",
            INIT_36 => X"000000500000006800000088000000ae00000093000000440000006d0000006b",
            INIT_37 => X"000000220000004500000051000000630000005e00000048000000460000004c",
            INIT_38 => X"000000370000003e000000430000006d000000bc000000ac00000070000000c4",
            INIT_39 => X"000000860000008c0000009f000000a9000000a9000000670000005800000022",
            INIT_3A => X"000000690000007a0000007f000000aa00000095000000460000005f0000007d",
            INIT_3B => X"0000002f00000035000000500000006f000000680000005a0000005b00000053",
            INIT_3C => X"0000004d000000580000004d0000008e000000b5000000ae00000088000000c5",
            INIT_3D => X"000000700000008200000089000000e6000000d3000000740000005d00000034",
            INIT_3E => X"00000050000000650000008a00000092000000760000004b0000005f00000065",
            INIT_3F => X"0000003000000030000000360000005d00000063000000630000005700000044",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE4;


    MEM_IFMAP_LAYER0_INSTANCE5 : if BRAM_NAME = "ifmap_layer0_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000710000007e0000005a000000ac000000bc000000b2000000a0000000cc",
            INIT_01 => X"0000005a00000058000000750000008d0000009b000000850000002500000052",
            INIT_02 => X"00000061000000760000007e0000006d000000680000003a000000570000005c",
            INIT_03 => X"0000002e000000370000002d00000037000000520000005e0000004d00000048",
            INIT_04 => X"000000910000006600000069000000ba000000c2000000b8000000b4000000d7",
            INIT_05 => X"000000620000004900000059000000590000005f000000690000003d0000006f",
            INIT_06 => X"0000003d00000073000000690000002000000040000000660000005f00000058",
            INIT_07 => X"000000360000004000000044000000400000004e000000410000003500000033",
            INIT_08 => X"0000008f0000006000000085000000bc000000c1000000bd000000c0000000cd",
            INIT_09 => X"0000008500000064000000600000006c00000037000000500000006f0000008d",
            INIT_0A => X"000000340000003a000000560000005c0000005d000000780000005d0000005d",
            INIT_0B => X"0000002e0000002d000000360000003e0000003b000000280000003c00000027",
            INIT_0C => X"000000840000006300000098000000b8000000b9000000b5000000bb000000b4",
            INIT_0D => X"000000a80000007b000000560000006c000000330000007e0000008700000082",
            INIT_0E => X"000000320000002c0000004e0000007600000069000000670000004900000076",
            INIT_0F => X"0000002e000000320000003400000040000000440000003c0000005d00000034",
            INIT_10 => X"000000920000006f000000a0000000b4000000ac000000af000000bb00000092",
            INIT_11 => X"000000b1000000ad000000740000005600000049000000570000006f000000b9",
            INIT_12 => X"000000290000003300000036000000390000003f000000420000006500000094",
            INIT_13 => X"0000003f000000450000003d0000004c000000520000004b0000005300000045",
            INIT_14 => X"0000009f0000005b00000093000000b3000000a8000000b0000000c80000007c",
            INIT_15 => X"000000c5000000d0000000c0000000a40000009300000090000000e1000000fa",
            INIT_16 => X"0000006600000057000000440000003a0000003e0000006d0000008f000000b5",
            INIT_17 => X"00000073000000700000007000000078000000770000007a0000006f0000006e",
            INIT_18 => X"000000d10000007100000096000000b6000000b1000000c0000000d500000085",
            INIT_19 => X"000000980000009c000000a2000000950000009d000000e8000000fc000000f7",
            INIT_1A => X"0000007d000000730000006e0000006f00000065000000680000007700000094",
            INIT_1B => X"0000008400000089000000840000008e0000008d000000870000008200000083",
            INIT_1C => X"000000ed000000a4000000ae000000c0000000bc000000bc000000a800000087",
            INIT_1D => X"000000650000006b00000069000000690000006f00000099000000e4000000f1",
            INIT_1E => X"000000800000007e0000007d0000007d00000074000000710000007800000073",
            INIT_1F => X"000000850000008b000000860000008700000089000000890000008b00000084",
            INIT_20 => X"000000f2000000b500000089000000bf000000b000000086000000820000008d",
            INIT_21 => X"00000074000000780000007900000077000000760000007f000000af000000f5",
            INIT_22 => X"000000820000007d0000007d0000007800000071000000730000007500000075",
            INIT_23 => X"000000950000008c00000090000000920000008e0000008e0000009100000086",
            INIT_24 => X"000000f9000000d10000008f000000a7000000880000007c0000008c000000a2",
            INIT_25 => X"00000073000000790000007f0000007f0000007d0000008000000076000000cd",
            INIT_26 => X"0000008a00000086000000830000007b00000075000000710000007000000071",
            INIT_27 => X"000000b6000000a7000000980000009a00000095000000930000009800000096",
            INIT_28 => X"000000f7000000ea000000a40000007e0000007a0000008200000093000000a5",
            INIT_29 => X"00000077000000770000007700000081000000830000007b0000007200000099",
            INIT_2A => X"0000009a000000960000008d000000830000007f0000007b0000007700000077",
            INIT_2B => X"000000a9000000b6000000b20000009e0000008a0000008c0000008d00000096",
            INIT_2C => X"000000ea000000e90000008a0000007e000000850000008a00000095000000a2",
            INIT_2D => X"00000077000000740000007b000000850000007c000000810000007e0000008c",
            INIT_2E => X"000000940000008b0000008a0000008c00000084000000820000007e0000007a",
            INIT_2F => X"0000008b0000008e000000b0000000b600000099000000850000008b00000093",
            INIT_30 => X"000000d30000009f0000007d0000008a0000008d0000008f00000093000000a1",
            INIT_31 => X"0000007800000083000000870000008b00000082000000800000007900000077",
            INIT_32 => X"000000880000008a0000008b0000008800000087000000820000007800000076",
            INIT_33 => X"00000088000000670000008c000000a4000000b2000000970000008a00000087",
            INIT_34 => X"0000008500000071000000840000008b000000920000008900000094000000b1",
            INIT_35 => X"0000008000000089000000870000008000000075000000690000006900000072",
            INIT_36 => X"0000007d0000008300000088000000890000008a0000008b0000008900000083",
            INIT_37 => X"0000007f0000006c00000092000000a8000000b5000000b30000009a00000085",
            INIT_38 => X"000000700000007d000000860000008b0000008f0000008400000094000000a8",
            INIT_39 => X"00000078000000730000006c0000006a0000006d000000660000006800000073",
            INIT_3A => X"0000007f0000007f00000086000000980000009c000000900000008700000080",
            INIT_3B => X"0000006b0000007e00000082000000a4000000be000000c5000000aa00000090",
            INIT_3C => X"000000730000007b0000008400000086000000860000008400000095000000a0",
            INIT_3D => X"00000059000000620000006c000000680000006c000000650000006900000072",
            INIT_3E => X"0000007b00000082000000830000009100000098000000890000007600000064",
            INIT_3F => X"0000006e000000810000007c00000091000000af000000b6000000a700000091",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE5;


    MEM_IFMAP_LAYER1_INSTANCE0 : if BRAM_NAME = "ifmap_layer1_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"00000021000000370000006c0000006000000000000000000000000000000000",
            INIT_07 => X"00000000000000170000000000000000000000000000004c0000000c00000038",
            INIT_08 => X"0000002b00000000000000070000001500000000000000000000002a0000000f",
            INIT_09 => X"000000290000000000000000000000000000001300000011000000610000005f",
            INIT_0A => X"0000005a000000b8000000460000004300000000000000730000005d00000000",
            INIT_0B => X"000000000000000000000023000000d600000017000000000000000000000000",
            INIT_0C => X"0000001f0000003a0000001c0000000000000000000000050000000000000000",
            INIT_0D => X"0000003800000024000000c20000001d000000000000000e0000013a00000027",
            INIT_0E => X"000000000000000000000022000001cf00000017000000000000006f00000080",
            INIT_0F => X"0000017a000000000000000000000000000000f2000000600000000000000016",
            INIT_10 => X"000000ce0000009d00000000000000000000000a000000000000000000000092",
            INIT_11 => X"0000000c0000007c000000000000007b00000000000000000000000d00000000",
            INIT_12 => X"00000000000000000000000f0000000000000000000000000000000300000000",
            INIT_13 => X"0000000000000011000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000360000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000380000000000000000",
            INIT_16 => X"0000009d000000000000007700000000000000000000004b0000000000000000",
            INIT_17 => X"000000000000000000000015000000000000002d000000000000000000000000",
            INIT_18 => X"0000000000000000000000060000000000000021000000000000001300000000",
            INIT_19 => X"000000000000000d000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000006a0000000000000000000000000000006e000000000000007900000000",
            INIT_1B => X"00000000000000cb000000000000000000000000000000060000000000000000",
            INIT_1C => X"0000000000000000000000370000001b000000390000003c0000000000000000",
            INIT_1D => X"000000b600000032000000000000000000000006000000000000000000000000",
            INIT_1E => X"000000000000006700000039000000000000000a000000000000000800000000",
            INIT_1F => X"00000015000000000000002a000000000000002e00000011000000200000000c",
            INIT_20 => X"0000000b00000009000000000000000000000000000000170000000900000036",
            INIT_21 => X"00000009000000290000000d0000000000000017000000000000000600000019",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_23 => X"000000090000000d000000000000001700000000000000000000000000000000",
            INIT_24 => X"000000000000000000000000000000130000001a000000260000001600000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000200000001000000000000000500000000000000000000000000000000",
            INIT_27 => X"0000000e000000000000001b0000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000011",
            INIT_29 => X"000000000000000000000000000000000000000f000000000000000000000000",
            INIT_2A => X"000000000000001500000018000000060000000100000000000000020000003b",
            INIT_2B => X"0000000000000005000000000000000b00000000000000000000000000000000",
            INIT_2C => X"0000001f0000000000000001000000400000001c000000060000001100000000",
            INIT_2D => X"000000080000001200000021000000080000002d00000017000000050000000c",
            INIT_2E => X"0000000000000031000000380000000000000000000000300000002200000013",
            INIT_2F => X"0000000000000000000000000000000000000008000000000000001a0000002e",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"00000000000000320000002a0000004a0000004a000000000000000000000022",
            INIT_32 => X"00000000000000000000003200000011000000000000000a0000000900000009",
            INIT_33 => X"000000000000001f00000019000000040000003e000000000000000500000000",
            INIT_34 => X"00000000000000160000000000000000000000000000004e000000000000005b",
            INIT_35 => X"000000000000005f00000083000000000000000d000000000000005b0000005d",
            INIT_36 => X"0000000000000000000000000000001c0000005b000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000190000000000000029000000000000000000000000",
            INIT_39 => X"00000000000000360000000000000017000000000000003c0000000000000000",
            INIT_3A => X"00000008000000000000001f0000000000000000000000000000001000000000",
            INIT_3B => X"0000003b000000aa000000000000000000000000000000000000000e00000017",
            INIT_3C => X"0000004d000000560000008700000027000000000000002f0000002700000056",
            INIT_3D => X"000000000000002d00000094000000510000006100000068000000720000004c",
            INIT_3E => X"0000000a0000000c00000018000000000000002500000038000000000000004d",
            INIT_3F => X"00000000000000000000001c0000000e000000000000002d0000009b00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE0;


    MEM_IFMAP_LAYER1_INSTANCE1 : if BRAM_NAME = "ifmap_layer1_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000001b0000003600000039000000390000007400000000",
            INIT_01 => X"00000092000000500000004d000000020000001d0000004b0000000000000013",
            INIT_02 => X"00000000000000000000009e0000002400000000000000000000000000000050",
            INIT_03 => X"00000000000000000000001c0000004b00000032000000150000001200000000",
            INIT_04 => X"000000000000004e000000000000000000000000000000000000000000000000",
            INIT_05 => X"000000000000000000000025000000000000002c000000370000000000000000",
            INIT_06 => X"0000001300000011000000000000003f00000000000000640000000000000000",
            INIT_07 => X"000000020000005f000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000400000053000000040000000b00000014000000000000000700000000",
            INIT_09 => X"00000000000000000000000000000000000000170000002e0000003200000018",
            INIT_0A => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"000000000000000000000000000000000000000000000000000000000000000d",
            INIT_0C => X"0000000e00000000000000160000000000000000000000000000000d00000000",
            INIT_0D => X"000000210000000100000000000000000000000600000000000000000000001e",
            INIT_0E => X"00000000000000000000001b0000001200000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000002e00000041000000380000003900000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000002200000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"000000000000001a00000000000000030000007c000000170000000000000023",
            INIT_14 => X"0000000000000017000000180000000600000015000000000000001a00000000",
            INIT_15 => X"00000092000000810000004000000035000000240000001e0000000c00000000",
            INIT_16 => X"0000000000000000000000000000003300000000000000190000006c00000027",
            INIT_17 => X"0000000000000000000000700000000000000000000000000000000000000000",
            INIT_18 => X"000000380000004f0000001c0000000000000000000000000000000500000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000360000000000000038",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000660000002600000065000000420000001c00000000",
            INIT_1E => X"0000004d00000000000000190000007700000056000000590000004e00000062",
            INIT_1F => X"00000025000000280000000c00000074000000b7000000470000003500000060",
            INIT_20 => X"000000840000006e000000500000003900000078000000850000003900000018",
            INIT_21 => X"000000bb000000ab0000009c00000092000000a90000008b0000009a0000008a",
            INIT_22 => X"0000005000000067000000a9000000b5000000a60000000a0000000000000000",
            INIT_23 => X"000000110000002d0000001c00000000000000000000004d0000009700000046",
            INIT_24 => X"0000001d000000680000001d000000000000002100000000000000000000001c",
            INIT_25 => X"0000002f0000002b000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000005600000067000000d100000024000000400000006a0000003400000037",
            INIT_27 => X"0000000000000000000000000000000000000061000000170000004200000073",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_2B => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000009b000000b3000000000000006800000000000000210000000000000000",
            INIT_2D => X"000000a900000098000000a00000007d000000c10000007c0000009c0000007d",
            INIT_2E => X"000000000000000000000000000000000000001c00000006000000b0000000c2",
            INIT_2F => X"0000000000000000000000000000000000000000000000110000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"00000050000000510000004b0000006100000062000000000000000000000000",
            INIT_35 => X"0000005a0000005e0000005b0000005300000088000000610000004100000049",
            INIT_36 => X"0000003c000000730000005f00000076000000600000005a000000680000002a",
            INIT_37 => X"0000005c0000005d00000041000000460000007b0000004e0000006d00000076",
            INIT_38 => X"0000002e0000002300000015000000100000004f0000003b0000004600000097",
            INIT_39 => X"000000000000000d00000000000000000000000000000000000000000000002f",
            INIT_3A => X"000000570000007b000000730000006300000000000000000000000000000000",
            INIT_3B => X"0000000500000040000000430000007000000045000000480000004b00000056",
            INIT_3C => X"00000024000000000000001e00000022000000320000002b0000004400000012",
            INIT_3D => X"00000021000000210000000000000009000000000000005d000000070000003c",
            INIT_3E => X"000000000000002b000000170000001900000015000000000000000600000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE1;


    MEM_IFMAP_LAYER1_INSTANCE2 : if BRAM_NAME = "ifmap_layer1_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004a0000005e0000005a0000000000000000000000000000000000000000",
            INIT_01 => X"0000002600000000000000360000003c0000004700000031000000260000002c",
            INIT_02 => X"0000003100000046000000020000000e000000500000003e0000003a00000026",
            INIT_03 => X"00000035000000440000005a00000026000000350000003f0000002d0000002e",
            INIT_04 => X"0000001d000000000000002c00000008000000000000001c0000004400000049",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000001100000032000000000000000a00000000000000170000000000000000",
            INIT_09 => X"000000000000002e00000000000000000000004c000000000000001100000000",
            INIT_0A => X"000000000000000000000011000000000000001c000000760000000000000002",
            INIT_0B => X"0000003e000000180000001a000000860000007b000000120000006e00000000",
            INIT_0C => X"000001160000004c0000004800000035000000330000003d000000af00000000",
            INIT_0D => X"000000f0000000be000000c10000006c00000074000000d1000000be0000010a",
            INIT_0E => X"0000007b0000003e000000550000002b00000003000000350000001500000096",
            INIT_0F => X"000000110000005700000064000000400000001000000000000000340000001c",
            INIT_10 => X"0000002f0000002700000030000000400000001f00000040000000000000000a",
            INIT_11 => X"0000000000000000000000000000000000000000000000370000007600000017",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"00000009000000000000006c000000000000002b000000000000000000000000",
            INIT_14 => X"000000000000006f000000840000006500000000000000970000000000000000",
            INIT_15 => X"0000000000000079000000c400000062000000b000000000000000ed00000000",
            INIT_16 => X"0000007600000025000000000000004600000000000000920000000000000053",
            INIT_17 => X"0000002400000000000000a20000000000000000000000000000001f00000053",
            INIT_18 => X"00000000000000000000000b0000000000000011000000060000000000000000",
            INIT_19 => X"00000024000000320000005c000000110000001e000000000000000600000000",
            INIT_1A => X"00000042000000260000002c00000046000000340000008a000000500000009e",
            INIT_1B => X"0000002a000000220000003600000022000000970000002e0000005900000036",
            INIT_1C => X"000000a6000000af000000170000001f00000000000000270000003500000031",
            INIT_1D => X"00000028000000bd0000009a0000001c0000002100000066000000370000002b",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000001f0000000b000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000001800000030000000000000000000000000000000000000000000000000",
            INIT_23 => X"000000860000007e000000470000000000000019000000200000002a00000005",
            INIT_24 => X"000000a3000000ae0000007d000000d0000000b0000000b3000000a70000008a",
            INIT_25 => X"0000000000000000000000000000000200000000000000e1000000bf000000ac",
            INIT_26 => X"0000004e000000000000002a0000002f00000004000000000000000000000000",
            INIT_27 => X"000000000000003a000000000000005300000000000000650000000000000000",
            INIT_28 => X"0000001c00000000000000250000000000000050000000000000000500000011",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000008b00000000",
            INIT_2A => X"0000001200000000000000000000000400000000000000220000000000000000",
            INIT_2B => X"000000000000000000000000000000000000000a000000240000000d00000018",
            INIT_2C => X"000000330000000000000000000000120000005000000004000000000000004d",
            INIT_2D => X"000000000000009100000000000000000000003f000000000000001e00000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000250000000000000000",
            INIT_2F => X"00000000000000000000007700000000000000000000000a0000004400000000",
            INIT_30 => X"00000000000000a6000000050000004200000067000000000000000000000000",
            INIT_31 => X"0000000000000003000000000000000b00000038000000410000003000000061",
            INIT_32 => X"000000230000004e000000290000000000000000000000000000000000000000",
            INIT_33 => X"000000000000006f0000002d0000000000000023000000000000002200000000",
            INIT_34 => X"00000000000000000000000000000000000000000000005c0000002e00000005",
            INIT_35 => X"0000000000000000000000000000002c0000002e000000030000002b00000000",
            INIT_36 => X"00000000000000530000005e0000005e00000000000000000000000000000000",
            INIT_37 => X"000000b000000090000000390000003000000036000000300000000000000000",
            INIT_38 => X"00000079000000b40000006a000000680000004a0000006700000067000000a2",
            INIT_39 => X"00000000000000420000006a0000003400000043000000140000003b00000025",
            INIT_3A => X"00000027000000000000002c0000002200000000000000240000000000000034",
            INIT_3B => X"0000000000000000000000080000001700000033000000000000003c00000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000046",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000001700000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000010000002d0000000a000000160000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE2;


    MEM_IFMAP_LAYER1_INSTANCE3 : if BRAM_NAME = "ifmap_layer1_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000008000000000000001e000000450000002f000000120000001700000003",
            INIT_01 => X"0000003a00000027000000390000004200000060000000000000000200000015",
            INIT_02 => X"000000880000007e0000007e000000480000000700000069000000260000003a",
            INIT_03 => X"000000ab000000a90000009e000000960000009200000066000000bb00000096",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE3;


    MEM_IFMAP_LAYER2_INSTANCE0 : if BRAM_NAME = "ifmap_layer2_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001d0000000f0000000d00000017000000140000000f0000001200000012",
            INIT_01 => X"00000016000000150000000c0000000600000001000000000000000a0000001d",
            INIT_02 => X"0000000000000003000000080000000400000013000000130000000f00000012",
            INIT_03 => X"0000000b000000000000000b0000000500000000000000000000000000000004",
            INIT_04 => X"00000000000000000000001e000000200000001b000000120000001b00000013",
            INIT_05 => X"0000000c00000000000000010000000100000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000110000000b00000019",
            INIT_07 => X"0000000300000003000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000001000000000000000000000000000000000000000000000000",
            INIT_0B => X"00000000000000000000001c0000000400000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000200000000000000000000000000000000",
            INIT_0E => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"000000000000000b000000000000000000000000000000000000000000000000",
            INIT_10 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"00000000000000000000000000000000000000000000000b0000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000020",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"000000000000000000000000000000000000000000000000000000000000000b",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"000000000000000d000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000070000000400000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000010000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000a0000003f0000000f0000001a0000000f000000000000000000000000",
            INIT_31 => X"0000002000000025000000380000003a00000032000000000000000000000000",
            INIT_32 => X"000000000000003a0000002c0000002000000027000000250000002900000022",
            INIT_33 => X"000000240000001f00000020000000200000001d0000001d0000001e00000000",
            INIT_34 => X"0000000e0000002f0000002f000000300000002100000028000000220000001e",
            INIT_35 => X"000000330000002f00000023000000220000001d00000019000000210000000f",
            INIT_36 => X"0000002a000000410000003100000033000000290000003a0000002800000034",
            INIT_37 => X"0000001a0000002d000000210000001c000000170000001f0000002a00000030",
            INIT_38 => X"000000000000000000000000000000000000000000000000000000290000001c",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"00000000000000000000000000000000000000060000000e0000001800000003",
            INIT_3E => X"000000000000000100000002000000000000000000000000000000000000000b",
            INIT_3F => X"0000001e0000000000000000000000000000000000000006000000000000001b",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER2_INSTANCE0;


    MEM_IFMAP_LAYER2_INSTANCE1 : if BRAM_NAME = "ifmap_layer2_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001d00000000000000030000000500000014000000110000000000000000",
            INIT_01 => X"00000000000000170000000f0000000300000000000000080000000000000010",
            INIT_02 => X"00000003000000440000000000000004000000060000000a0000001a00000000",
            INIT_03 => X"00000000000000000000000b0000001700000002000000000000000b00000000",
            INIT_04 => X"00000004000000000000003700000000000000000000000b0000001e0000000c",
            INIT_05 => X"000000060000000000000006000000140000002000000002000000110000000a",
            INIT_06 => X"000000110000000000000000000000200000000000000000000000000000002d",
            INIT_07 => X"00000000000000080000001100000004000000280000001d0000000000000008",
            INIT_08 => X"00000000000000060000000000000010000000000000000b0000000b00000000",
            INIT_09 => X"00000012000000090000000e0000002700000000000000240000001800000000",
            INIT_0A => X"00000000000000000000000c0000000000000000000000000000001500000012",
            INIT_0B => X"000000110000002d000000280000000d0000005800000000000000230000002b",
            INIT_0C => X"00000036000000000000000b0000001f000000220000001b0000000000000000",
            INIT_0D => X"0000001a000000210000001f0000000700000000000000450000001200000023",
            INIT_0E => X"000000380000002a0000002f0000002f0000002e00000028000000220000001e",
            INIT_0F => X"0000002a00000024000000240000002500000027000000000000002500000033",
            INIT_10 => X"000000520000002e0000002c0000003a0000002e0000002f000000360000002f",
            INIT_11 => X"0000002e0000002f0000002a0000002a000000260000002b0000001300000000",
            INIT_12 => X"000000190000002c000000330000002b00000028000000450000002a0000002f",
            INIT_13 => X"0000002e0000002d000000310000002e00000024000000230000002800000019",
            INIT_14 => X"00000000000000000000000000000000000000000000001f0000003a00000043",
            INIT_15 => X"00000000000000000000000a0000000200000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"00000000000000030000001c0000001f00000000000000170000000800000010",
            INIT_18 => X"0000002b00000000000000000000000000000000000000000000002a00000000",
            INIT_19 => X"00000000000000000000003f0000002d00000042000000000000000000000011",
            INIT_1A => X"0000002c00000028000000000000000e00000000000000000000000000000071",
            INIT_1B => X"0000006c000000000000002a0000003b000000260000005a0000000000000025",
            INIT_1C => X"0000003c000000480000005d0000002400000034000000000000002300000005",
            INIT_1D => X"0000003100000059000000000000003e0000001e000000520000002f00000000",
            INIT_1E => X"00000000000000600000003e000000610000002c000000000000000000000037",
            INIT_1F => X"0000001500000073000000480000002500000031000000120000005c00000073",
            INIT_20 => X"00000075000000000000006a0000004a0000005a000000000000000000000038",
            INIT_21 => X"0000003100000028000000650000004d000000370000000c0000001200000047",
            INIT_22 => X"000000500000004f0000000000000046000000380000008b0000000600000000",
            INIT_23 => X"0000002a0000000b000000840000004200000068000000130000002500000006",
            INIT_24 => X"000000040000005b0000001600000029000000000000002c0000002e00000013",
            INIT_25 => X"0000001800000064000000000000009f0000003a0000004a0000000000000000",
            INIT_26 => X"0000000000000000000000170000005a0000003b000000300000004d00000000",
            INIT_27 => X"000000200000004c0000009300000000000000940000003c0000000f0000000c",
            INIT_28 => X"0000003100000020000000230000001d0000001a000000410000008300000071",
            INIT_29 => X"0000003c0000003a00000073000000d8000000000000004e0000002b0000001d",
            INIT_2A => X"0000005f0000004f000000400000003e0000003c0000003d0000003800000047",
            INIT_2B => X"0000003e0000003f0000004900000042000000af000000820000000000000012",
            INIT_2C => X"000000450000006a0000003d0000004800000050000000400000003800000039",
            INIT_2D => X"000000410000003c000000420000004d000000390000005a000000cb00000000",
            INIT_2E => X"0000003e0000004b000000760000007b000000380000004e0000004d00000048",
            INIT_2F => X"0000005500000044000000380000004400000043000000350000004800000054",
            INIT_30 => X"00000008000000080000000000000000000000800000006f0000001a0000003a",
            INIT_31 => X"0000000000000000000000000000000400000000000000050000000300000006",
            INIT_32 => X"0000000a000000070000000c0000000a00000007000000050000000600000000",
            INIT_33 => X"0000000000000006000000240000000000000000000000000000001a00000049",
            INIT_34 => X"0000000000000007000000040000000400000000000000000000000400000000",
            INIT_35 => X"000000000000001700000007000000150000001a0000000d0000000000000000",
            INIT_36 => X"00000037000000000000000d0000000500000009000000250000002800000000",
            INIT_37 => X"000000000000000100000000000000000000000000000000000000050000001b",
            INIT_38 => X"0000000e0000000600000056000000800000000b000000130000005a00000026",
            INIT_39 => X"0000000000000000000000180000000f00000025000000250000000000000000",
            INIT_3A => X"0000001f0000001a0000002a0000000000000000000000000000000800000000",
            INIT_3B => X"000000070000000600000027000000090000000000000000000000000000003a",
            INIT_3C => X"00000011000000090000000a0000000000000021000000000000000400000000",
            INIT_3D => X"0000001c00000007000000150000001d00000017000000000000000b00000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000160000001900000010",
            INIT_3F => X"000000040000000b000000040000001000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER2_INSTANCE1;


    MEM_IFMAP_LAYER2_INSTANCE2 : if BRAM_NAME = "ifmap_layer2_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000000000000040000001a00000000000000000000001c",
            INIT_01 => X"00000011000000040000000900000000000000000000002f0000000300000000",
            INIT_02 => X"0000001b0000000000000000000000000000000c0000004a0000000000000000",
            INIT_03 => X"000000850000009c00000046000000000000000000000000000000000000001f",
            INIT_04 => X"000000000000001b000000410000002000000000000000000000000000000028",
            INIT_05 => X"000000000000000000000000000000460000000f000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000002",
            INIT_08 => X"0000000000000011000000000000000000000012000000070000000400000000",
            INIT_09 => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000001300000000000000000000000000000000",
            INIT_0B => X"0000001300000014000000000000000000000000000000000000000000000000",
            INIT_0C => X"000000a2000000a30000009d0000000000000022000000280000000000000004",
            INIT_0D => X"0000007c00000094000000ad000000b7000000ac0000009d000000a4000000a5",
            INIT_0E => X"000000ac000000a8000000ad000000a20000009200000092000000840000007c",
            INIT_0F => X"0000003e0000002e0000003a0000007a000000a0000000a90000008c000000a0",
            INIT_10 => X"000000af000000b0000000ac0000006a000000890000008b0000006e0000004e",
            INIT_11 => X"000000270000000a0000001e000000070000002d00000048000000730000008e",
            INIT_12 => X"00000059000000a2000000aa000000a40000002b0000004d000000670000003a",
            INIT_13 => X"000000250000001b0000002d000000330000000c00000015000000270000004d",
            INIT_14 => X"00000043000000470000004e00000060000000940000001f000000170000003a",
            INIT_15 => X"0000002f0000001c000000170000003900000031000000000000001f0000002f",
            INIT_16 => X"00000031000000450000003b00000025000000990000008e0000001200000016",
            INIT_17 => X"0000000e0000001700000012000000100000002a0000003e000000000000002d",
            INIT_18 => X"0000002f0000002d0000003e000000320000002f0000009f000000620000002a",
            INIT_19 => X"0000000a0000001c000000260000000e00000010000000280000003200000000",
            INIT_1A => X"0000001e00000029000000270000002e0000002600000037000000620000002c",
            INIT_1B => X"0000002b00000000000000140000004100000022000000090000002d0000002f",
            INIT_1C => X"00000042000000540000000d000000300000003600000022000000550000000e",
            INIT_1D => X"00000000000000240000000500000010000000790000002d0000000f00000026",
            INIT_1E => X"000000060000001d000000340000002d00000028000000080000002000000035",
            INIT_1F => X"00000017000000000000002300000015000000000000008a0000006200000009",
            INIT_20 => X"000000000000000000000000000000000000000600000000000000000000001a",
            INIT_21 => X"000000000000003a000000060000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000003400000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000002300000022000000000000000000000000000000000000000000000000",
            INIT_29 => X"000000170000001d0000002400000026000000270000001e0000002000000025",
            INIT_2A => X"0000002a0000002c00000023000000180000001e00000024000000260000001a",
            INIT_2B => X"000000000000001d0000000e0000001d0000000f00000020000000280000001f",
            INIT_2C => X"000000210000002800000039000000060000001c0000002b0000002000000009",
            INIT_2D => X"00000000000000000000002e0000002100000006000000000000001a00000027",
            INIT_2E => X"0000000f00000029000000210000004c000000000000002c0000002500000000",
            INIT_2F => X"0000000000000009000000000000004800000000000000000000000400000024",
            INIT_30 => X"0000000b00000009000000560000000200000026000000000000004a00000000",
            INIT_31 => X"0000000000000006000000000000000000000059000000000000000000000000",
            INIT_32 => X"00000000000000130000003e0000001a000000000000000a000000000000002b",
            INIT_33 => X"00000000000000000000001400000000000000000000008e0000000000000000",
            INIT_34 => X"0000000000000000000000360000003f00000000000000200000000000000000",
            INIT_35 => X"0000000000000000000000150000000a00000000000000000000006600000000",
            INIT_36 => X"0000000000000000000000000000004200000038000000000000000000000000",
            INIT_37 => X"0000000200000000000000080000000f0000001d000000000000000000000042",
            INIT_38 => X"0000000000000024000000000000000000000011000000040000002100000000",
            INIT_39 => X"00000000000000000000000000000023000000210000001e0000000000000025",
            INIT_3A => X"00000000000000050000000200000000000000270000000f000000000000002c",
            INIT_3B => X"0000007800000000000000040000002a0000001400000034000000300000000c",
            INIT_3C => X"0000000900000008000000000000000000000000000000220000000000000000",
            INIT_3D => X"0000000000000040000000000000001400000020000000000000000000000001",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000004300000021000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER2_INSTANCE2;


    MEM_IFMAP_LAYER2_INSTANCE3 : if BRAM_NAME = "ifmap_layer2_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"000000000000000000000000000000000000005d000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000002b00000000000000000000000400000000000000000000000000000000",
            INIT_05 => X"000000370000003a00000030000000290000002f0000002c0000002d00000030",
            INIT_06 => X"000000350000002c000000310000002a0000002700000026000000250000002a",
            INIT_07 => X"0000000c0000003b000000290000001f000000000000002d0000002e00000030",
            INIT_08 => X"0000002e000000290000001c000000250000001f0000000e0000000000000000",
            INIT_09 => X"000000000000000000000000000000230000002d0000003b0000003200000035",
            INIT_0A => X"000000320000002300000000000000000000001a000000040000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000001900000025",
            INIT_0C => X"0000000000000018000000120000000000000000000000110000000000000006",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000300000003000000380000000b00000000000000000000000500000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000070000003a00000007000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000200000000000000000000000000000000",
            INIT_13 => X"000000000000000d000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000050000001a00000000000000000000000000000000",
            INIT_15 => X"000000000000000000000008000000000000000400000018000000030000000f",
            INIT_16 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000001f00000000000000000000000a00000011",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000b0000000c0000000c000000040000000800000008000000110000000a",
            INIT_22 => X"00000000000000060000000800000011000000230000002d000000210000000b",
            INIT_23 => X"00000042000000230000000500000000000000080000000c0000000a0000000a",
            INIT_24 => X"00000033000000350000000a000000170000000a000000000000000000000000",
            INIT_25 => X"0000000000000000000000090000001600000037000000050000000800000005",
            INIT_26 => X"0000000500000000000000000000000c0000000e000000000000000000000000",
            INIT_27 => X"000000040000001a000000000000000200000000000000000000000800000008",
            INIT_28 => X"0000000e0000000200000000000000010000000e000000000000000600000010",
            INIT_29 => X"0000000000000000000000000000000700000000000000090000000000000000",
            INIT_2A => X"0000003e0000000300000006000000000000000f000000000000000000000000",
            INIT_2B => X"0000000700000015000000140000000000000000000000000000000000000028",
            INIT_2C => X"0000000000000012000000180000001c00000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000001100000000000000110000000000000031",
            INIT_2E => X"0000003500000035000000020000000000000000000000000000000000000000",
            INIT_2F => X"000000000000000e000000050000000000000009000000000000000e00000021",
            INIT_30 => X"0000000000000000000000260000000000000000000000000000000100000000",
            INIT_31 => X"0000000c00000000000000000000000000000030000000260000000000000000",
            INIT_32 => X"0000000000000000000000000000000900000023000000000000000400000000",
            INIT_33 => X"000000000000000300000018000000000000000000000011000000360000004e",
            INIT_34 => X"0000000000000037000000510000001e00000000000000000000000000000007",
            INIT_35 => X"0000000c00000021000000350000000a00000005000000000000000000000000",
            INIT_36 => X"0000000000000000000000030000000500000004000000280000005600000000",
            INIT_37 => X"0000001800000000000000160000000000000000000000000000000000000000",
            INIT_38 => X"000000000000000000000000000000000000000000000000000000000000003f",
            INIT_39 => X"0000000b0000004f000000180000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000300000000000000220000000000000000000000000000001400000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000012",
            INIT_3D => X"0000000800000015000000090000000e0000000a000000130000000d00000000",
            INIT_3E => X"0000000200000006000000130000001b000000220000001c0000000c00000006",
            INIT_3F => X"0000001a0000000f000000360000000f0000000d000000090000000b00000008",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER2_INSTANCE3;


    MEM_IFMAP_LAYER2_INSTANCE4 : if BRAM_NAME = "ifmap_layer2_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000260000000a0000001a000000210000002400000035000000340000001f",
            INIT_01 => X"00000020000000280000003300000051000000080000000a0000000b00000024",
            INIT_02 => X"00000014000000330000001a000000190000002b0000004b0000005e00000053",
            INIT_03 => X"0000005b000000360000002f000000450000002e00000019000000120000000e",
            INIT_04 => X"000000150000005e000000710000001b000000150000003b000000420000005d",
            INIT_05 => X"000000670000003b000000330000003b00000064000000440000007e00000035",
            INIT_06 => X"00000013000000280000009e0000007f00000001000000250000003900000038",
            INIT_07 => X"000000500000007f0000005b0000002e0000004b0000007d0000007e000000bd",
            INIT_08 => X"0000005a0000001700000043000000940000007a000000150000003c00000047",
            INIT_09 => X"0000003b0000004600000081000000780000004e00000065000000a800000075",
            INIT_0A => X"000000a5000000390000003900000040000000a50000008e000000330000004c",
            INIT_0B => X"0000004b000000480000004c000000780000005f000000500000006a00000085",
            INIT_0C => X"0000005900000066000000380000007300000066000000b8000000b000000026",
            INIT_0D => X"0000000e0000002b0000002c000000410000006500000033000000510000004e",
            INIT_0E => X"000000790000005f000000330000006f0000007500000086000000b3000000c0",
            INIT_0F => X"000000c700000027000000270000002f00000025000000400000005a00000042",
            INIT_10 => X"00000079000000b900000091000000650000009e000000a20000008b000000ab",
            INIT_11 => X"000000cb000000c100000068000000710000005a00000047000000400000003c",
            INIT_12 => X"0000006f0000007c000000850000008a000000a5000000e7000000c90000009d",
            INIT_13 => X"000000b1000000a10000008c0000008e0000008a000000880000008000000078",
            INIT_14 => X"00000084000000760000007100000070000000750000007a000000af000000e5",
            INIT_15 => X"000000ef000000a6000000850000009d000000a30000009a000000950000008c",
            INIT_16 => X"0000009b0000008c000000820000007700000073000000790000008000000088",
            INIT_17 => X"00000074000000a70000007f0000008f00000097000000ab000000a300000093",
            INIT_18 => X"0000009a0000008500000086000000880000007c0000007e000000890000007f",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000008d000000af",
            INIT_1A => X"00000000000000000000000b0000001c00000013000000000000000000000000",
            INIT_1B => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"00000000000000000000001e0000001400000000000000000000003300000014",
            INIT_1D => X"000000280000001c0000003e000000000000000000000000000000000000003f",
            INIT_1E => X"00000019000000000000001e0000000700000000000000000000000000000000",
            INIT_1F => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000e000000060000001a0000000000000000",
            INIT_21 => X"000000000000001d000000040000000f00000000000000000000000000000009",
            INIT_22 => X"00000002000000000000002f0000002500000000000000000000000800000000",
            INIT_23 => X"000000260000000000000006000000000000000000000000000000030000004f",
            INIT_24 => X"0000000d0000000d00000018000000000000000000000000000000000000001c",
            INIT_25 => X"0000000800000018000000000000000900000000000000050000000000000000",
            INIT_26 => X"0000000000000000000000070000000000000002000000000000000000000000",
            INIT_27 => X"000000000000001c0000000000000000000000000000001e0000003d00000000",
            INIT_28 => X"0000003200000022000000000000002e00000000000000000000000000000010",
            INIT_29 => X"000000000000000d0000003a0000002600000036000000000000000000000003",
            INIT_2A => X"000000000000001500000012000000000000000a000000000000000000000000",
            INIT_2B => X"00000008000000000000000000000001000000310000001f0000002e00000000",
            INIT_2C => X"0000001900000000000000000000000000000000000000220000000000000000",
            INIT_2D => X"0000004100000021000000160000000000000000000000000000000d0000000f",
            INIT_2E => X"0000000c000000370000003f00000052000000a2000000000000000000000000",
            INIT_2F => X"000000360000000d000000000000000000000000000000020000000000000006",
            INIT_30 => X"0000000000000000000000000000000200000000000000560000004100000000",
            INIT_31 => X"0000002500000000000000020000000000000000000000030000000000000000",
            INIT_32 => X"000000070000000000000000000000010000000000000000000000060000003e",
            INIT_33 => X"0000003600000018000000000000000c0000004200000000000000000000000a",
            INIT_34 => X"0000000000000005000000000000000000000000000000090000001300000024",
            INIT_35 => X"0000000000000000000000000000000000000000000000040000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"00000000000000000000000000000000000000000000001f0000000400000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_3C => X"0000000000000001000000020000000000000007000000000000002d00000005",
            INIT_3D => X"0000000200000000000000000000000000000000000000000000000000000002",
            INIT_3E => X"000000060000000100000010000000000000000300000000000000000000003b",
            INIT_3F => X"0000005d000000000000000000000000000000000000002c0000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER2_INSTANCE4;


    MEM_IFMAP_LAYER2_INSTANCE5 : if BRAM_NAME = "ifmap_layer2_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000000000000000000000000000000e0000000000000000",
            INIT_01 => X"00000000000000520000000000000000000000000000000f0000001c00000000",
            INIT_02 => X"0000000000000000000000000000000400000000000000130000001200000000",
            INIT_03 => X"00000000000000000000002d000000000000000500000000000000170000000c",
            INIT_04 => X"000000000000001100000000000000160000000000000000000000030000001d",
            INIT_05 => X"0000001b00000000000000110000000000000008000000000000000000000012",
            INIT_06 => X"00000003000000000000003b0000000000000019000000090000000000000000",
            INIT_07 => X"0000000000000012000000120000000000000000000000050000000000000010",
            INIT_08 => X"0000002d000000000000000000000058000000000000000d0000003300000000",
            INIT_09 => X"0000001d0000002c0000003e0000003300000028000000020000000000000004",
            INIT_0A => X"0000004e0000004e0000002e000000000000003b000000000000003600000070",
            INIT_0B => X"0000005a000000530000005a00000058000000560000004f0000004900000044",
            INIT_0C => X"0000004c0000004a00000048000000490000000000000008000000480000006f",
            INIT_0D => X"000000600000005a0000005e0000005d000000570000005b0000005b00000054",
            INIT_0E => X"00000057000000530000004d000000450000005000000031000000000000008a",
            INIT_0F => X"0000006700000067000000500000005e00000074000000610000006400000061",
            INIT_10 => X"00000052000000520000005200000049000000550000005f0000004900000041",
            INIT_11 => X"0000002e000000330000002e0000002f00000045000000530000006b0000005e",
            INIT_12 => X"000000270000001c000000230000002b0000002f000000310000002f0000002f",
            INIT_13 => X"000000340000002d000000350000003200000032000000240000002700000026",
            INIT_14 => X"0000002400000015000000130000002100000004000000250000001300000055",
            INIT_15 => X"0000002c000000380000002e000000340000003b0000001a000000280000002d",
            INIT_16 => X"00000027000000040000000b0000000a0000004f0000001a0000000000000000",
            INIT_17 => X"0000001a0000002300000025000000360000002c000000790000000000000039",
            INIT_18 => X"000000530000000e000000000000001200000000000000530000001800000008",
            INIT_19 => X"00000000000000000000001a0000002c000000490000000a0000006300000000",
            INIT_1A => X"0000000000000039000000000000001e000000000000000b0000005f00000008",
            INIT_1B => X"00000000000000000000000000000000000000490000002e0000000000000038",
            INIT_1C => X"00000015000000000000000d00000004000000230000000000000000000000bf",
            INIT_1D => X"000000a400000000000000000000000a0000005000000061000000000000000c",
            INIT_1E => X"0000000100000000000000000000000d000000270000001e0000000000000000",
            INIT_1F => X"000000000000007c000000000000000800000000000000680000004500000000",
            INIT_20 => X"0000003c00000000000000170000000000000012000000220000002a00000000",
            INIT_21 => X"000000000000002200000006000000310000001c000000000000000300000011",
            INIT_22 => X"000000000000004a00000000000000180000000a000000440000003a00000026",
            INIT_23 => X"0000004800000005000000000000000a000000170000000e0000002a00000019",
            INIT_24 => X"0000000b00000000000000a30000000000000011000000510000001c00000056",
            INIT_25 => X"0000001e0000002d000000280000001400000000000000000000000000000056",
            INIT_26 => X"0000000000000000000000000000009800000000000000280000004000000000",
            INIT_27 => X"00000000000000110000000e0000001000000010000000090000000000000000",
            INIT_28 => X"0000000a0000000500000009000000000000001f000000480000004100000003",
            INIT_29 => X"0000000000000017000000080000001000000017000000140000001000000008",
            INIT_2A => X"0000000d00000009000000000000001100000000000000000000007400000010",
            INIT_2B => X"0000000d00000000000000000000002600000000000000090000000d00000010",
            INIT_2C => X"0000001000000018000000090000000c00000016000000000000000000000019",
            INIT_2D => X"0000000000000000000000000000000000000003000000310000000b00000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000001000000000000000000000000000000000000000400000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000012000000040000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000005",
            INIT_35 => X"0000000000000008000000380000000000000000000000270000000100000000",
            INIT_36 => X"0000000000000004000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"000000000000000f000000000000000000000000000000000000001400000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000012000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER2_INSTANCE5;


    MEM_IFMAP_LAYER2_INSTANCE6 : if BRAM_NAME = "ifmap_layer2_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000300000001e000000000000000000000000000000000000000000000011",
            INIT_01 => X"00000001000000240000001c000000000000000000000000000000000000003e",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"000000360000002f000000000000000000000013000000000000000000000000",
            INIT_0A => X"0000002b000000360000003b0000003900000030000000350000003500000033",
            INIT_0B => X"0000003600000038000000300000002700000028000000250000002000000020",
            INIT_0C => X"000000020000000200000023000000390000003b000000420000003300000039",
            INIT_0D => X"0000003900000036000000130000003000000027000000110000000600000006",
            INIT_0E => X"00000000000000040000000000000000000000000000001e0000003d00000037",
            INIT_0F => X"0000004000000037000000320000000000000015000000170000000000000001",
            INIT_10 => X"0000000000000000000000170000000000000000000000000000001e00000012",
            INIT_11 => X"0000003300000044000000100000003400000012000000000000000000000000",
            INIT_12 => X"0000000000000000000000090000001000000000000000000000000600000025",
            INIT_13 => X"0000002b0000000d0000000b00000038000000310000000f0000000000000000",
            INIT_14 => X"000000000000000000000000000000000000002a000000000000000b00000008",
            INIT_15 => X"000000170000002e000000110000000e0000003d000000070000002c00000000",
            INIT_16 => X"0000000400000000000000000000000000000000000000130000000300000008",
            INIT_17 => X"000000000000000a0000002e0000002200000000000000250000000000000019",
            INIT_18 => X"0000001100000015000000000000000200000000000000000000000f00000013",
            INIT_19 => X"0000002c000000000000000c00000000000000000000001c0000000000000009",
            INIT_1A => X"000000140000000e000000160000002100000000000000000000000000000000",
            INIT_1B => X"0000000000000005000000060000001f00000000000000000000000300000000",
            INIT_1C => X"00000000000000150000001400000005000000280000001e0000000000000000",
            INIT_1D => X"000000000000000000000000000000000000001700000011000000060000002c",
            INIT_1E => X"0000003c00000032000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"00000000000000000000004f0000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000002800000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000002f0000002b00000028000000200000002c000000290000002300000022",
            INIT_27 => X"00000024000000280000002e000000290000001e0000001d0000002900000032",
            INIT_28 => X"000000050000002e00000030000000430000000e000000210000002c00000024",
            INIT_29 => X"00000028000000020000003f0000002c00000015000000190000002900000021",
            INIT_2A => X"0000001c00000000000000100000002400000028000000200000002a00000029",
            INIT_2B => X"000000240000002e000000000000005c0000000b0000001a000000320000000c",
            INIT_2C => X"0000001800000023000000000000001900000025000000270000000c00000038",
            INIT_2D => X"000000130000000000000041000000050000002c00000000000000260000001a",
            INIT_2E => X"0000001200000038000000140000000000000025000000240000002a00000027",
            INIT_2F => X"00000000000000000000002f0000003700000000000000240000001a0000002b",
            INIT_30 => X"0000001d000000070000002a0000003400000000000000430000002500000016",
            INIT_31 => X"000000150000000000000000000000460000000e000000240000001100000020",
            INIT_32 => X"00000025000000000000000d000000280000002b00000000000000390000001c",
            INIT_33 => X"0000000b0000003500000000000000020000003400000029000000060000000b",
            INIT_34 => X"0000000d0000000d00000011000000000000002c000000110000000000000018",
            INIT_35 => X"000000000000001b0000000e0000000000000034000000000000003f00000000",
            INIT_36 => X"00000000000000000000001a00000000000000000000002b000000050000003f",
            INIT_37 => X"0000000f0000002c0000001d00000000000000140000002a0000000000000039",
            INIT_38 => X"0000003800000000000000000000002f00000010000000000000000f0000002f",
            INIT_39 => X"0000000f0000002b000000270000000500000000000000320000002900000000",
            INIT_3A => X"0000000000000000000000000000000000000021000000110000000800000008",
            INIT_3B => X"0000000000000003000000070000000000000000000000000000000500000052",
            INIT_3C => X"0000002e00000022000000000000000000000014000000030000000000000000",
            INIT_3D => X"0000000200000000000000000000000100000005000000020000000600000000",
            INIT_3E => X"000000000000000d000000220000000000000000000000090000000000000000",
            INIT_3F => X"0000000000000000000000000000000100000000000000000000000600000009",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER2_INSTANCE6;


    MEM_IFMAP_LAYER2_INSTANCE7 : if BRAM_NAME = "ifmap_layer2_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000140000000400000000000000000000001300000015",
            INIT_01 => X"0000001a0000001200000000000000000000000c000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER2_INSTANCE7;


    MEM_GOLD_LAYER0_INSTANCE0 : if BRAM_NAME = "gold_layer0_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001d0000000f0000000d00000017000000140000000f0000001200000012",
            INIT_01 => X"00000016000000150000000c0000000600000001000000000000000a0000001d",
            INIT_02 => X"0000000000000003000000080000000400000013000000130000000f00000012",
            INIT_03 => X"0000000b000000000000000b0000000500000000000000000000000000000004",
            INIT_04 => X"00000000000000000000001e000000200000001b000000120000001b00000013",
            INIT_05 => X"0000000c00000000000000010000000100000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000110000000b00000019",
            INIT_07 => X"0000000300000003000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000001000000000000000000000000000000000000000000000000",
            INIT_0B => X"00000000000000000000001c0000000400000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000200000000000000000000000000000000",
            INIT_0E => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"000000000000000b000000000000000000000000000000000000000000000000",
            INIT_10 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"00000000000000000000000000000000000000000000000b0000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000020",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"000000000000000000000000000000000000000000000000000000000000000b",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"000000000000000d000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000070000000400000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000010000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000a0000003f0000000f0000001a0000000f000000000000000000000000",
            INIT_31 => X"0000002000000025000000380000003a00000032000000000000000000000000",
            INIT_32 => X"000000000000003a0000002c0000002000000027000000250000002900000022",
            INIT_33 => X"000000240000001f00000020000000200000001d0000001d0000001e00000000",
            INIT_34 => X"0000000e0000002f0000002f000000300000002100000028000000220000001e",
            INIT_35 => X"000000330000002f00000023000000220000001d00000019000000210000000f",
            INIT_36 => X"0000002a000000410000003100000033000000290000003a0000002800000034",
            INIT_37 => X"0000001a0000002d000000210000001c000000170000001f0000002a00000030",
            INIT_38 => X"000000000000000000000000000000000000000000000000000000290000001c",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"00000000000000000000000000000000000000060000000e0000001800000003",
            INIT_3E => X"000000000000000100000002000000000000000000000000000000000000000b",
            INIT_3F => X"0000001e0000000000000000000000000000000000000006000000000000001b",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE0;


    MEM_GOLD_LAYER0_INSTANCE1 : if BRAM_NAME = "gold_layer0_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001d00000000000000030000000500000014000000110000000000000000",
            INIT_01 => X"00000000000000170000000f0000000300000000000000080000000000000010",
            INIT_02 => X"00000003000000440000000000000004000000060000000a0000001a00000000",
            INIT_03 => X"00000000000000000000000b0000001700000002000000000000000b00000000",
            INIT_04 => X"00000004000000000000003700000000000000000000000b0000001e0000000c",
            INIT_05 => X"000000060000000000000006000000140000002000000002000000110000000a",
            INIT_06 => X"000000110000000000000000000000200000000000000000000000000000002d",
            INIT_07 => X"00000000000000080000001100000004000000280000001d0000000000000008",
            INIT_08 => X"00000000000000060000000000000010000000000000000b0000000b00000000",
            INIT_09 => X"00000012000000090000000e0000002700000000000000240000001800000000",
            INIT_0A => X"00000000000000000000000c0000000000000000000000000000001500000012",
            INIT_0B => X"000000110000002d000000280000000d0000005800000000000000230000002b",
            INIT_0C => X"00000036000000000000000b0000001f000000220000001b0000000000000000",
            INIT_0D => X"0000001a000000210000001f0000000700000000000000450000001200000023",
            INIT_0E => X"000000380000002a0000002f0000002f0000002e00000028000000220000001e",
            INIT_0F => X"0000002a00000024000000240000002500000027000000000000002500000033",
            INIT_10 => X"000000520000002e0000002c0000003a0000002e0000002f000000360000002f",
            INIT_11 => X"0000002e0000002f0000002a0000002a000000260000002b0000001300000000",
            INIT_12 => X"000000190000002c000000330000002b00000028000000450000002a0000002f",
            INIT_13 => X"0000002e0000002d000000310000002e00000024000000230000002800000019",
            INIT_14 => X"00000000000000000000000000000000000000000000001f0000003a00000043",
            INIT_15 => X"00000000000000000000000a0000000200000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"00000000000000030000001c0000001f00000000000000170000000800000010",
            INIT_18 => X"0000002b00000000000000000000000000000000000000000000002a00000000",
            INIT_19 => X"00000000000000000000003f0000002d00000042000000000000000000000011",
            INIT_1A => X"0000002c00000028000000000000000e00000000000000000000000000000071",
            INIT_1B => X"0000006c000000000000002a0000003b000000260000005a0000000000000025",
            INIT_1C => X"0000003c000000480000005d0000002400000034000000000000002300000005",
            INIT_1D => X"0000003100000059000000000000003e0000001e000000520000002f00000000",
            INIT_1E => X"00000000000000600000003e000000610000002c000000000000000000000037",
            INIT_1F => X"0000001500000073000000480000002500000031000000120000005c00000073",
            INIT_20 => X"00000075000000000000006a0000004a0000005a000000000000000000000038",
            INIT_21 => X"0000003100000028000000650000004d000000370000000c0000001200000047",
            INIT_22 => X"000000500000004f0000000000000046000000380000008b0000000600000000",
            INIT_23 => X"0000002a0000000b000000840000004200000068000000130000002500000006",
            INIT_24 => X"000000040000005b0000001600000029000000000000002c0000002e00000013",
            INIT_25 => X"0000001800000064000000000000009f0000003a0000004a0000000000000000",
            INIT_26 => X"0000000000000000000000170000005a0000003b000000300000004d00000000",
            INIT_27 => X"000000200000004c0000009300000000000000940000003c0000000f0000000c",
            INIT_28 => X"0000003100000020000000230000001d0000001a000000410000008300000071",
            INIT_29 => X"0000003c0000003a00000073000000d8000000000000004e0000002b0000001d",
            INIT_2A => X"0000005f0000004f000000400000003e0000003c0000003d0000003800000047",
            INIT_2B => X"0000003e0000003f0000004900000042000000af000000820000000000000012",
            INIT_2C => X"000000450000006a0000003d0000004800000050000000400000003800000039",
            INIT_2D => X"000000410000003c000000420000004d000000390000005a000000cb00000000",
            INIT_2E => X"0000003e0000004b000000760000007b000000380000004e0000004d00000048",
            INIT_2F => X"0000005500000044000000380000004400000043000000350000004800000054",
            INIT_30 => X"00000008000000080000000000000000000000800000006f0000001a0000003a",
            INIT_31 => X"0000000000000000000000000000000400000000000000050000000300000006",
            INIT_32 => X"0000000a000000070000000c0000000a00000007000000050000000600000000",
            INIT_33 => X"0000000000000006000000240000000000000000000000000000001a00000049",
            INIT_34 => X"0000000000000007000000040000000400000000000000000000000400000000",
            INIT_35 => X"000000000000001700000007000000150000001a0000000d0000000000000000",
            INIT_36 => X"00000037000000000000000d0000000500000009000000250000002800000000",
            INIT_37 => X"000000000000000100000000000000000000000000000000000000050000001b",
            INIT_38 => X"0000000e0000000600000056000000800000000b000000130000005a00000026",
            INIT_39 => X"0000000000000000000000180000000f00000025000000250000000000000000",
            INIT_3A => X"0000001f0000001a0000002a0000000000000000000000000000000800000000",
            INIT_3B => X"000000070000000600000027000000090000000000000000000000000000003a",
            INIT_3C => X"00000011000000090000000a0000000000000021000000000000000400000000",
            INIT_3D => X"0000001c00000007000000150000001d00000017000000000000000b00000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000160000001900000010",
            INIT_3F => X"000000040000000b000000040000001000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE1;


    MEM_GOLD_LAYER0_INSTANCE2 : if BRAM_NAME = "gold_layer0_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000000000000040000001a00000000000000000000001c",
            INIT_01 => X"00000011000000040000000900000000000000000000002f0000000300000000",
            INIT_02 => X"0000001b0000000000000000000000000000000c0000004a0000000000000000",
            INIT_03 => X"000000850000009c00000046000000000000000000000000000000000000001f",
            INIT_04 => X"000000000000001b000000410000002000000000000000000000000000000028",
            INIT_05 => X"000000000000000000000000000000460000000f000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000002",
            INIT_08 => X"0000000000000011000000000000000000000012000000070000000400000000",
            INIT_09 => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000001300000000000000000000000000000000",
            INIT_0B => X"0000001300000014000000000000000000000000000000000000000000000000",
            INIT_0C => X"000000a2000000a30000009d0000000000000022000000280000000000000004",
            INIT_0D => X"0000007c00000094000000ad000000b7000000ac0000009d000000a4000000a5",
            INIT_0E => X"000000ac000000a8000000ad000000a20000009200000092000000840000007c",
            INIT_0F => X"0000003e0000002e0000003a0000007a000000a0000000a90000008c000000a0",
            INIT_10 => X"000000af000000b0000000ac0000006a000000890000008b0000006e0000004e",
            INIT_11 => X"000000270000000a0000001e000000070000002d00000048000000730000008e",
            INIT_12 => X"00000059000000a2000000aa000000a40000002b0000004d000000670000003a",
            INIT_13 => X"000000250000001b0000002d000000330000000c00000015000000270000004d",
            INIT_14 => X"00000043000000470000004e00000060000000940000001f000000170000003a",
            INIT_15 => X"0000002f0000001c000000170000003900000031000000000000001f0000002f",
            INIT_16 => X"00000031000000450000003b00000025000000990000008e0000001200000016",
            INIT_17 => X"0000000e0000001700000012000000100000002a0000003e000000000000002d",
            INIT_18 => X"0000002f0000002d0000003e000000320000002f0000009f000000620000002a",
            INIT_19 => X"0000000a0000001c000000260000000e00000010000000280000003200000000",
            INIT_1A => X"0000001e00000029000000270000002e0000002600000037000000620000002c",
            INIT_1B => X"0000002b00000000000000140000004100000022000000090000002d0000002f",
            INIT_1C => X"00000042000000540000000d000000300000003600000022000000550000000e",
            INIT_1D => X"00000000000000240000000500000010000000790000002d0000000f00000026",
            INIT_1E => X"000000060000001d000000340000002d00000028000000080000002000000035",
            INIT_1F => X"00000017000000000000002300000015000000000000008a0000006200000009",
            INIT_20 => X"000000000000000000000000000000000000000600000000000000000000001a",
            INIT_21 => X"000000000000003a000000060000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000003400000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000002300000022000000000000000000000000000000000000000000000000",
            INIT_29 => X"000000170000001d0000002400000026000000270000001e0000002000000025",
            INIT_2A => X"0000002a0000002c00000023000000180000001e00000024000000260000001a",
            INIT_2B => X"000000000000001d0000000e0000001d0000000f00000020000000280000001f",
            INIT_2C => X"000000210000002800000039000000060000001c0000002b0000002000000009",
            INIT_2D => X"00000000000000000000002e0000002100000006000000000000001a00000027",
            INIT_2E => X"0000000f00000029000000210000004c000000000000002c0000002500000000",
            INIT_2F => X"0000000000000009000000000000004800000000000000000000000400000024",
            INIT_30 => X"0000000b00000009000000560000000200000026000000000000004a00000000",
            INIT_31 => X"0000000000000006000000000000000000000059000000000000000000000000",
            INIT_32 => X"00000000000000130000003e0000001a000000000000000a000000000000002b",
            INIT_33 => X"00000000000000000000001400000000000000000000008e0000000000000000",
            INIT_34 => X"0000000000000000000000360000003f00000000000000200000000000000000",
            INIT_35 => X"0000000000000000000000150000000a00000000000000000000006600000000",
            INIT_36 => X"0000000000000000000000000000004200000038000000000000000000000000",
            INIT_37 => X"0000000200000000000000080000000f0000001d000000000000000000000042",
            INIT_38 => X"0000000000000024000000000000000000000011000000040000002100000000",
            INIT_39 => X"00000000000000000000000000000023000000210000001e0000000000000025",
            INIT_3A => X"00000000000000050000000200000000000000270000000f000000000000002c",
            INIT_3B => X"0000007800000000000000040000002a0000001400000034000000300000000c",
            INIT_3C => X"0000000900000008000000000000000000000000000000220000000000000000",
            INIT_3D => X"0000000000000040000000000000001400000020000000000000000000000001",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000004300000021000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE2;


    MEM_GOLD_LAYER0_INSTANCE3 : if BRAM_NAME = "gold_layer0_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"000000000000000000000000000000000000005d000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000002b00000000000000000000000400000000000000000000000000000000",
            INIT_05 => X"000000370000003a00000030000000290000002f0000002c0000002d00000030",
            INIT_06 => X"000000350000002c000000310000002a0000002700000026000000250000002a",
            INIT_07 => X"0000000c0000003b000000290000001f000000000000002d0000002e00000030",
            INIT_08 => X"0000002e000000290000001c000000250000001f0000000e0000000000000000",
            INIT_09 => X"000000000000000000000000000000230000002d0000003b0000003200000035",
            INIT_0A => X"000000320000002300000000000000000000001a000000040000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000001900000025",
            INIT_0C => X"0000000000000018000000120000000000000000000000110000000000000006",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000300000003000000380000000b00000000000000000000000500000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000070000003a00000007000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000200000000000000000000000000000000",
            INIT_13 => X"000000000000000d000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000050000001a00000000000000000000000000000000",
            INIT_15 => X"000000000000000000000008000000000000000400000018000000030000000f",
            INIT_16 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000001f00000000000000000000000a00000011",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000b0000000c0000000c000000040000000800000008000000110000000a",
            INIT_22 => X"00000000000000060000000800000011000000230000002d000000210000000b",
            INIT_23 => X"00000042000000230000000500000000000000080000000c0000000a0000000a",
            INIT_24 => X"00000033000000350000000a000000170000000a000000000000000000000000",
            INIT_25 => X"0000000000000000000000090000001600000037000000050000000800000005",
            INIT_26 => X"0000000500000000000000000000000c0000000e000000000000000000000000",
            INIT_27 => X"000000040000001a000000000000000200000000000000000000000800000008",
            INIT_28 => X"0000000e0000000200000000000000010000000e000000000000000600000010",
            INIT_29 => X"0000000000000000000000000000000700000000000000090000000000000000",
            INIT_2A => X"0000003e0000000300000006000000000000000f000000000000000000000000",
            INIT_2B => X"0000000700000015000000140000000000000000000000000000000000000028",
            INIT_2C => X"0000000000000012000000180000001c00000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000001100000000000000110000000000000031",
            INIT_2E => X"0000003500000035000000020000000000000000000000000000000000000000",
            INIT_2F => X"000000000000000e000000050000000000000009000000000000000e00000021",
            INIT_30 => X"0000000000000000000000260000000000000000000000000000000100000000",
            INIT_31 => X"0000000c00000000000000000000000000000030000000260000000000000000",
            INIT_32 => X"0000000000000000000000000000000900000023000000000000000400000000",
            INIT_33 => X"000000000000000300000018000000000000000000000011000000360000004e",
            INIT_34 => X"0000000000000037000000510000001e00000000000000000000000000000007",
            INIT_35 => X"0000000c00000021000000350000000a00000005000000000000000000000000",
            INIT_36 => X"0000000000000000000000030000000500000004000000280000005600000000",
            INIT_37 => X"0000001800000000000000160000000000000000000000000000000000000000",
            INIT_38 => X"000000000000000000000000000000000000000000000000000000000000003f",
            INIT_39 => X"0000000b0000004f000000180000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000300000000000000220000000000000000000000000000001400000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000012",
            INIT_3D => X"0000000800000015000000090000000e0000000a000000130000000d00000000",
            INIT_3E => X"0000000200000006000000130000001b000000220000001c0000000c00000006",
            INIT_3F => X"0000001a0000000f000000360000000f0000000d000000090000000b00000008",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE3;


    MEM_GOLD_LAYER0_INSTANCE4 : if BRAM_NAME = "gold_layer0_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000260000000a0000001a000000210000002400000035000000340000001f",
            INIT_01 => X"00000020000000280000003300000051000000080000000a0000000b00000024",
            INIT_02 => X"00000014000000330000001a000000190000002b0000004b0000005e00000053",
            INIT_03 => X"0000005b000000360000002f000000450000002e00000019000000120000000e",
            INIT_04 => X"000000150000005e000000710000001b000000150000003b000000420000005d",
            INIT_05 => X"000000670000003b000000330000003b00000064000000440000007e00000035",
            INIT_06 => X"00000013000000280000009e0000007f00000001000000250000003900000038",
            INIT_07 => X"000000500000007f0000005b0000002e0000004b0000007d0000007e000000bd",
            INIT_08 => X"0000005a0000001700000043000000940000007a000000150000003c00000047",
            INIT_09 => X"0000003b0000004600000081000000780000004e00000065000000a800000075",
            INIT_0A => X"000000a5000000390000003900000040000000a50000008e000000330000004c",
            INIT_0B => X"0000004b000000480000004c000000780000005f000000500000006a00000085",
            INIT_0C => X"0000005900000066000000380000007300000066000000b8000000b000000026",
            INIT_0D => X"0000000e0000002b0000002c000000410000006500000033000000510000004e",
            INIT_0E => X"000000790000005f000000330000006f0000007500000086000000b3000000c0",
            INIT_0F => X"000000c700000027000000270000002f00000025000000400000005a00000042",
            INIT_10 => X"00000079000000b900000091000000650000009e000000a20000008b000000ab",
            INIT_11 => X"000000cb000000c100000068000000710000005a00000047000000400000003c",
            INIT_12 => X"0000006f0000007c000000850000008a000000a5000000e7000000c90000009d",
            INIT_13 => X"000000b1000000a10000008c0000008e0000008a000000880000008000000078",
            INIT_14 => X"00000084000000760000007100000070000000750000007a000000af000000e5",
            INIT_15 => X"000000ef000000a6000000850000009d000000a30000009a000000950000008c",
            INIT_16 => X"0000009b0000008c000000820000007700000073000000790000008000000088",
            INIT_17 => X"00000074000000a70000007f0000008f00000097000000ab000000a300000093",
            INIT_18 => X"0000009a0000008500000086000000880000007c0000007e000000890000007f",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000008d000000af",
            INIT_1A => X"00000000000000000000000b0000001c00000013000000000000000000000000",
            INIT_1B => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"00000000000000000000001e0000001400000000000000000000003300000014",
            INIT_1D => X"000000280000001c0000003e000000000000000000000000000000000000003f",
            INIT_1E => X"00000019000000000000001e0000000700000000000000000000000000000000",
            INIT_1F => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000e000000060000001a0000000000000000",
            INIT_21 => X"000000000000001d000000040000000f00000000000000000000000000000009",
            INIT_22 => X"00000002000000000000002f0000002500000000000000000000000800000000",
            INIT_23 => X"000000260000000000000006000000000000000000000000000000030000004f",
            INIT_24 => X"0000000d0000000d00000018000000000000000000000000000000000000001c",
            INIT_25 => X"0000000800000018000000000000000900000000000000050000000000000000",
            INIT_26 => X"0000000000000000000000070000000000000002000000000000000000000000",
            INIT_27 => X"000000000000001c0000000000000000000000000000001e0000003d00000000",
            INIT_28 => X"0000003200000022000000000000002e00000000000000000000000000000010",
            INIT_29 => X"000000000000000d0000003a0000002600000036000000000000000000000003",
            INIT_2A => X"000000000000001500000012000000000000000a000000000000000000000000",
            INIT_2B => X"00000008000000000000000000000001000000310000001f0000002e00000000",
            INIT_2C => X"0000001900000000000000000000000000000000000000220000000000000000",
            INIT_2D => X"0000004100000021000000160000000000000000000000000000000d0000000f",
            INIT_2E => X"0000000c000000370000003f00000052000000a2000000000000000000000000",
            INIT_2F => X"000000360000000d000000000000000000000000000000020000000000000006",
            INIT_30 => X"0000000000000000000000000000000200000000000000560000004100000000",
            INIT_31 => X"0000002500000000000000020000000000000000000000030000000000000000",
            INIT_32 => X"000000070000000000000000000000010000000000000000000000060000003e",
            INIT_33 => X"0000003600000018000000000000000c0000004200000000000000000000000a",
            INIT_34 => X"0000000000000005000000000000000000000000000000090000001300000024",
            INIT_35 => X"0000000000000000000000000000000000000000000000040000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"00000000000000000000000000000000000000000000001f0000000400000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_3C => X"0000000000000001000000020000000000000007000000000000002d00000005",
            INIT_3D => X"0000000200000000000000000000000000000000000000000000000000000002",
            INIT_3E => X"000000060000000100000010000000000000000300000000000000000000003b",
            INIT_3F => X"0000005d000000000000000000000000000000000000002c0000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE4;


    MEM_GOLD_LAYER0_INSTANCE5 : if BRAM_NAME = "gold_layer0_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000000000000000000000000000000e0000000000000000",
            INIT_01 => X"00000000000000520000000000000000000000000000000f0000001c00000000",
            INIT_02 => X"0000000000000000000000000000000400000000000000130000001200000000",
            INIT_03 => X"00000000000000000000002d000000000000000500000000000000170000000c",
            INIT_04 => X"000000000000001100000000000000160000000000000000000000030000001d",
            INIT_05 => X"0000001b00000000000000110000000000000008000000000000000000000012",
            INIT_06 => X"00000003000000000000003b0000000000000019000000090000000000000000",
            INIT_07 => X"0000000000000012000000120000000000000000000000050000000000000010",
            INIT_08 => X"0000002d000000000000000000000058000000000000000d0000003300000000",
            INIT_09 => X"0000001d0000002c0000003e0000003300000028000000020000000000000004",
            INIT_0A => X"0000004e0000004e0000002e000000000000003b000000000000003600000070",
            INIT_0B => X"0000005a000000530000005a00000058000000560000004f0000004900000044",
            INIT_0C => X"0000004c0000004a00000048000000490000000000000008000000480000006f",
            INIT_0D => X"000000600000005a0000005e0000005d000000570000005b0000005b00000054",
            INIT_0E => X"00000057000000530000004d000000450000005000000031000000000000008a",
            INIT_0F => X"0000006700000067000000500000005e00000074000000610000006400000061",
            INIT_10 => X"00000052000000520000005200000049000000550000005f0000004900000041",
            INIT_11 => X"0000002e000000330000002e0000002f00000045000000530000006b0000005e",
            INIT_12 => X"000000270000001c000000230000002b0000002f000000310000002f0000002f",
            INIT_13 => X"000000340000002d000000350000003200000032000000240000002700000026",
            INIT_14 => X"0000002400000015000000130000002100000004000000250000001300000055",
            INIT_15 => X"0000002c000000380000002e000000340000003b0000001a000000280000002d",
            INIT_16 => X"00000027000000040000000b0000000a0000004f0000001a0000000000000000",
            INIT_17 => X"0000001a0000002300000025000000360000002c000000790000000000000039",
            INIT_18 => X"000000530000000e000000000000001200000000000000530000001800000008",
            INIT_19 => X"00000000000000000000001a0000002c000000490000000a0000006300000000",
            INIT_1A => X"0000000000000039000000000000001e000000000000000b0000005f00000008",
            INIT_1B => X"00000000000000000000000000000000000000490000002e0000000000000038",
            INIT_1C => X"00000015000000000000000d00000004000000230000000000000000000000bf",
            INIT_1D => X"000000a400000000000000000000000a0000005000000061000000000000000c",
            INIT_1E => X"0000000100000000000000000000000d000000270000001e0000000000000000",
            INIT_1F => X"000000000000007c000000000000000800000000000000680000004500000000",
            INIT_20 => X"0000003c00000000000000170000000000000012000000220000002a00000000",
            INIT_21 => X"000000000000002200000006000000310000001c000000000000000300000011",
            INIT_22 => X"000000000000004a00000000000000180000000a000000440000003a00000026",
            INIT_23 => X"0000004800000005000000000000000a000000170000000e0000002a00000019",
            INIT_24 => X"0000000b00000000000000a30000000000000011000000510000001c00000056",
            INIT_25 => X"0000001e0000002d000000280000001400000000000000000000000000000056",
            INIT_26 => X"0000000000000000000000000000009800000000000000280000004000000000",
            INIT_27 => X"00000000000000110000000e0000001000000010000000090000000000000000",
            INIT_28 => X"0000000a0000000500000009000000000000001f000000480000004100000003",
            INIT_29 => X"0000000000000017000000080000001000000017000000140000001000000008",
            INIT_2A => X"0000000d00000009000000000000001100000000000000000000007400000010",
            INIT_2B => X"0000000d00000000000000000000002600000000000000090000000d00000010",
            INIT_2C => X"0000001000000018000000090000000c00000016000000000000000000000019",
            INIT_2D => X"0000000000000000000000000000000000000003000000310000000b00000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000001000000000000000000000000000000000000000400000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000012000000040000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000005",
            INIT_35 => X"0000000000000008000000380000000000000000000000270000000100000000",
            INIT_36 => X"0000000000000004000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"000000000000000f000000000000000000000000000000000000001400000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000012000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE5;


    MEM_GOLD_LAYER0_INSTANCE6 : if BRAM_NAME = "gold_layer0_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000300000001e000000000000000000000000000000000000000000000011",
            INIT_01 => X"00000001000000240000001c000000000000000000000000000000000000003e",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"000000360000002f000000000000000000000013000000000000000000000000",
            INIT_0A => X"0000002b000000360000003b0000003900000030000000350000003500000033",
            INIT_0B => X"0000003600000038000000300000002700000028000000250000002000000020",
            INIT_0C => X"000000020000000200000023000000390000003b000000420000003300000039",
            INIT_0D => X"0000003900000036000000130000003000000027000000110000000600000006",
            INIT_0E => X"00000000000000040000000000000000000000000000001e0000003d00000037",
            INIT_0F => X"0000004000000037000000320000000000000015000000170000000000000001",
            INIT_10 => X"0000000000000000000000170000000000000000000000000000001e00000012",
            INIT_11 => X"0000003300000044000000100000003400000012000000000000000000000000",
            INIT_12 => X"0000000000000000000000090000001000000000000000000000000600000025",
            INIT_13 => X"0000002b0000000d0000000b00000038000000310000000f0000000000000000",
            INIT_14 => X"000000000000000000000000000000000000002a000000000000000b00000008",
            INIT_15 => X"000000170000002e000000110000000e0000003d000000070000002c00000000",
            INIT_16 => X"0000000400000000000000000000000000000000000000130000000300000008",
            INIT_17 => X"000000000000000a0000002e0000002200000000000000250000000000000019",
            INIT_18 => X"0000001100000015000000000000000200000000000000000000000f00000013",
            INIT_19 => X"0000002c000000000000000c00000000000000000000001c0000000000000009",
            INIT_1A => X"000000140000000e000000160000002100000000000000000000000000000000",
            INIT_1B => X"0000000000000005000000060000001f00000000000000000000000300000000",
            INIT_1C => X"00000000000000150000001400000005000000280000001e0000000000000000",
            INIT_1D => X"000000000000000000000000000000000000001700000011000000060000002c",
            INIT_1E => X"0000003c00000032000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"00000000000000000000004f0000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000002800000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000002f0000002b00000028000000200000002c000000290000002300000022",
            INIT_27 => X"00000024000000280000002e000000290000001e0000001d0000002900000032",
            INIT_28 => X"000000050000002e00000030000000430000000e000000210000002c00000024",
            INIT_29 => X"00000028000000020000003f0000002c00000015000000190000002900000021",
            INIT_2A => X"0000001c00000000000000100000002400000028000000200000002a00000029",
            INIT_2B => X"000000240000002e000000000000005c0000000b0000001a000000320000000c",
            INIT_2C => X"0000001800000023000000000000001900000025000000270000000c00000038",
            INIT_2D => X"000000130000000000000041000000050000002c00000000000000260000001a",
            INIT_2E => X"0000001200000038000000140000000000000025000000240000002a00000027",
            INIT_2F => X"00000000000000000000002f0000003700000000000000240000001a0000002b",
            INIT_30 => X"0000001d000000070000002a0000003400000000000000430000002500000016",
            INIT_31 => X"000000150000000000000000000000460000000e000000240000001100000020",
            INIT_32 => X"00000025000000000000000d000000280000002b00000000000000390000001c",
            INIT_33 => X"0000000b0000003500000000000000020000003400000029000000060000000b",
            INIT_34 => X"0000000d0000000d00000011000000000000002c000000110000000000000018",
            INIT_35 => X"000000000000001b0000000e0000000000000034000000000000003f00000000",
            INIT_36 => X"00000000000000000000001a00000000000000000000002b000000050000003f",
            INIT_37 => X"0000000f0000002c0000001d00000000000000140000002a0000000000000039",
            INIT_38 => X"0000003800000000000000000000002f00000010000000000000000f0000002f",
            INIT_39 => X"0000000f0000002b000000270000000500000000000000320000002900000000",
            INIT_3A => X"0000000000000000000000000000000000000021000000110000000800000008",
            INIT_3B => X"0000000000000003000000070000000000000000000000000000000500000052",
            INIT_3C => X"0000002e00000022000000000000000000000014000000030000000000000000",
            INIT_3D => X"0000000200000000000000000000000100000005000000020000000600000000",
            INIT_3E => X"000000000000000d000000220000000000000000000000090000000000000000",
            INIT_3F => X"0000000000000000000000000000000100000000000000000000000600000009",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE6;


    MEM_GOLD_LAYER0_INSTANCE7 : if BRAM_NAME = "gold_layer0_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000140000000400000000000000000000001300000015",
            INIT_01 => X"0000001a0000001200000000000000000000000c000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE7;


    MEM_GOLD_LAYER1_INSTANCE0 : if BRAM_NAME = "gold_layer1_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000101000000bc00000051000001040000004000000012000000a0",
            INIT_01 => X"00000000000000ba00000000000000000000001c000000000000004700000000",
            INIT_02 => X"0000000000000092000000000000000000000031000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000200000000000000000000010400000000000000000000000000000000",
            INIT_05 => X"0000003800000000000000a80000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000037000000530000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"00000000000000000000000000000000000000000000000f0000000000000000",
            INIT_0A => X"000000b7000000820000011300000037000001340000017a000000a800000000",
            INIT_0B => X"000000620000014d00000000000000790000002d000000000000000000000035",
            INIT_0C => X"00000035000000100000007e0000000000000000000000000000000000000000",
            INIT_0D => X"00000000000000000000000000000000000000d1000000000000006a00000000",
            INIT_0E => X"00000081000000d20000007700000033000000a000000000000000b0000000b0",
            INIT_0F => X"000000650000000000000057000000a9000000080000000000000000000000c6",
            INIT_10 => X"000000000000007a00000058000000000000003c000000a100000000000000c8",
            INIT_11 => X"0000000000000000000000000000005c00000000000000060000000000000000",
            INIT_12 => X"000000ff00000000000000480000007700000000000000e60000002c00000000",
            INIT_13 => X"0000000000000000000000360000000000000019000000000000000000000024",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"00000000000000aa0000006c000000b50000004d0000005d0000000000000000",
            INIT_17 => X"000000300000001b000000000000003f00000000000000000000000000000000",
            INIT_18 => X"0000001200000000000000b30000011900000000000000000000000000000015",
            INIT_19 => X"000000000000000000000026000000b6000000bd00000000000000aa00000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000028",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000001700000068000000d00000014f0000014400000124000000c000000000",
            INIT_1D => X"0000000000000016000000570000000900000000000000000000004000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000005d000000cf",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"000000b800000001000000a80000000000000000000000000000000000000000",
            INIT_21 => X"000000000000000000000063000000150000009000000096000000280000001e",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000009e0000011b000000000000000000000000000000000000000000000000",
            INIT_24 => X"00000079000000000000000000000000000000000000006c0000000000000000",
            INIT_25 => X"00000000000000110000001200000067000000ff0000000400000043000000f8",
            INIT_26 => X"0000004e00000086000000000000004100000069000000000000001c00000000",
            INIT_27 => X"0000002600000017000000510000006c00000091000000000000000000000031",
            INIT_28 => X"000000000000007800000000000000e0000000fd000000b00000000000000046",
            INIT_29 => X"000000ab00000059000000000000000000000000000000000000000000000010",
            INIT_2A => X"000000530000003b000000db0000008f0000006a000000ef000000fb000000c1",
            INIT_2B => X"00000062000000ab000000460000007b00000000000000000000001000000014",
            INIT_2C => X"00000051000001230000007a0000008c0000006d000000a20000013c0000005a",
            INIT_2D => X"000000000000003c00000000000000000000000000000000000000a100000097",
            INIT_2E => X"0000010400000000000000000000000000000000000000000000000000000007",
            INIT_2F => X"0000012f000000a20000004f0000001e00000000000000000000000000000000",
            INIT_30 => X"000000a100000083000001610000013a0000015b00000000000000000000008c",
            INIT_31 => X"000000dc00000070000000880000000000000000000000120000013800000072",
            INIT_32 => X"000000000000000000000000000000ae000000cd0000013e000000ad000000e0",
            INIT_33 => X"0000001f000000c8000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000001e00000000000000260000001b0000004e0000004b00000046000000bf",
            INIT_35 => X"000000a5000000aa000000060000001e000000360000009f0000013b00000073",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000010100000076000000430000006a00000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000007c00000066",
            INIT_3C => X"0000005900000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000003d00000000000000000000000000000000000000310000000000000069",
            INIT_3E => X"0000000000000000000000ed0000007200000031000000100000000000000000",
            INIT_3F => X"0000012c00000070000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER1_INSTANCE0;


    MEM_GOLD_LAYER1_INSTANCE1 : if BRAM_NAME = "gold_layer1_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000003200000000000000000000000000000000000000d00000017f",
            INIT_01 => X"00000076000000440000006d000000de00000021000000390000000800000067",
            INIT_02 => X"0000000000000000000000000000000000000000000000eb0000014100000084",
            INIT_03 => X"0000003f0000006e00000078000000b200000000000000000000000000000000",
            INIT_04 => X"0000001c0000000000000000000000000000000000000000000000920000007f",
            INIT_05 => X"00000000000000000000014800000087000000340000001e0000000000000191",
            INIT_06 => X"0000004a00000058000000000000000000000000000000000000000000000000",
            INIT_07 => X"000000c5000000d7000000f30000000000000000000000000000000000000046",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER1_INSTANCE1;


    MEM_GOLD_LAYER2_INSTANCE0 : if BRAM_NAME = "gold_layer2_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"00000021000000370000006c0000006000000000000000000000000000000000",
            INIT_07 => X"00000000000000170000000000000000000000000000004c0000000c00000038",
            INIT_08 => X"0000002b00000000000000070000001500000000000000000000002a0000000f",
            INIT_09 => X"000000290000000000000000000000000000001300000011000000610000005f",
            INIT_0A => X"0000005a000000b8000000460000004300000000000000730000005d00000000",
            INIT_0B => X"000000000000000000000023000000d600000017000000000000000000000000",
            INIT_0C => X"0000001f0000003a0000001c0000000000000000000000050000000000000000",
            INIT_0D => X"0000003800000024000000c20000001d000000000000000e0000013a00000027",
            INIT_0E => X"000000000000000000000022000001cf00000017000000000000006f00000080",
            INIT_0F => X"0000017a000000000000000000000000000000f2000000600000000000000016",
            INIT_10 => X"000000ce0000009d00000000000000000000000a000000000000000000000092",
            INIT_11 => X"0000000c0000007c000000000000007b00000000000000000000000d00000000",
            INIT_12 => X"00000000000000000000000f0000000000000000000000000000000300000000",
            INIT_13 => X"0000000000000011000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000360000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000380000000000000000",
            INIT_16 => X"0000009d000000000000007700000000000000000000004b0000000000000000",
            INIT_17 => X"000000000000000000000015000000000000002d000000000000000000000000",
            INIT_18 => X"0000000000000000000000060000000000000021000000000000001300000000",
            INIT_19 => X"000000000000000d000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000006a0000000000000000000000000000006e000000000000007900000000",
            INIT_1B => X"00000000000000cb000000000000000000000000000000060000000000000000",
            INIT_1C => X"0000000000000000000000370000001b000000390000003c0000000000000000",
            INIT_1D => X"000000b600000032000000000000000000000006000000000000000000000000",
            INIT_1E => X"000000000000006700000039000000000000000a000000000000000800000000",
            INIT_1F => X"00000015000000000000002a000000000000002e00000011000000200000000c",
            INIT_20 => X"0000000b00000009000000000000000000000000000000170000000900000036",
            INIT_21 => X"00000009000000290000000d0000000000000017000000000000000600000019",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_23 => X"000000090000000d000000000000001700000000000000000000000000000000",
            INIT_24 => X"000000000000000000000000000000130000001a000000260000001600000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000200000001000000000000000500000000000000000000000000000000",
            INIT_27 => X"0000000e000000000000001b0000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000011",
            INIT_29 => X"000000000000000000000000000000000000000f000000000000000000000000",
            INIT_2A => X"000000000000001500000018000000060000000100000000000000020000003b",
            INIT_2B => X"0000000000000005000000000000000b00000000000000000000000000000000",
            INIT_2C => X"0000001f0000000000000001000000400000001c000000060000001100000000",
            INIT_2D => X"000000080000001200000021000000080000002d00000017000000050000000c",
            INIT_2E => X"0000000000000031000000380000000000000000000000300000002200000013",
            INIT_2F => X"0000000000000000000000000000000000000008000000000000001a0000002e",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"00000000000000320000002a0000004a0000004a000000000000000000000022",
            INIT_32 => X"00000000000000000000003200000011000000000000000a0000000900000009",
            INIT_33 => X"000000000000001f00000019000000040000003e000000000000000500000000",
            INIT_34 => X"00000000000000160000000000000000000000000000004e000000000000005b",
            INIT_35 => X"000000000000005f00000083000000000000000d000000000000005b0000005d",
            INIT_36 => X"0000000000000000000000000000001c0000005b000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000190000000000000029000000000000000000000000",
            INIT_39 => X"00000000000000360000000000000017000000000000003c0000000000000000",
            INIT_3A => X"00000008000000000000001f0000000000000000000000000000001000000000",
            INIT_3B => X"0000003b000000aa000000000000000000000000000000000000000e00000017",
            INIT_3C => X"0000004d000000560000008700000027000000000000002f0000002700000056",
            INIT_3D => X"000000000000002d00000094000000510000006100000068000000720000004c",
            INIT_3E => X"0000000a0000000c00000018000000000000002500000038000000000000004d",
            INIT_3F => X"00000000000000000000001c0000000e000000000000002d0000009b00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER2_INSTANCE0;


    MEM_GOLD_LAYER2_INSTANCE1 : if BRAM_NAME = "gold_layer2_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000001b0000003600000039000000390000007400000000",
            INIT_01 => X"00000092000000500000004d000000020000001d0000004b0000000000000013",
            INIT_02 => X"00000000000000000000009e0000002400000000000000000000000000000050",
            INIT_03 => X"00000000000000000000001c0000004b00000032000000150000001200000000",
            INIT_04 => X"000000000000004e000000000000000000000000000000000000000000000000",
            INIT_05 => X"000000000000000000000025000000000000002c000000370000000000000000",
            INIT_06 => X"0000001300000011000000000000003f00000000000000640000000000000000",
            INIT_07 => X"000000020000005f000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000400000053000000040000000b00000014000000000000000700000000",
            INIT_09 => X"00000000000000000000000000000000000000170000002e0000003200000018",
            INIT_0A => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"000000000000000000000000000000000000000000000000000000000000000d",
            INIT_0C => X"0000000e00000000000000160000000000000000000000000000000d00000000",
            INIT_0D => X"000000210000000100000000000000000000000600000000000000000000001e",
            INIT_0E => X"00000000000000000000001b0000001200000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000002e00000041000000380000003900000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000002200000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"000000000000001a00000000000000030000007c000000170000000000000023",
            INIT_14 => X"0000000000000017000000180000000600000015000000000000001a00000000",
            INIT_15 => X"00000092000000810000004000000035000000240000001e0000000c00000000",
            INIT_16 => X"0000000000000000000000000000003300000000000000190000006c00000027",
            INIT_17 => X"0000000000000000000000700000000000000000000000000000000000000000",
            INIT_18 => X"000000380000004f0000001c0000000000000000000000000000000500000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000360000000000000038",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000660000002600000065000000420000001c00000000",
            INIT_1E => X"0000004d00000000000000190000007700000056000000590000004e00000062",
            INIT_1F => X"00000025000000280000000c00000074000000b7000000470000003500000060",
            INIT_20 => X"000000840000006e000000500000003900000078000000850000003900000018",
            INIT_21 => X"000000bb000000ab0000009c00000092000000a90000008b0000009a0000008a",
            INIT_22 => X"0000005000000067000000a9000000b5000000a60000000a0000000000000000",
            INIT_23 => X"000000110000002d0000001c00000000000000000000004d0000009700000046",
            INIT_24 => X"0000001d000000680000001d000000000000002100000000000000000000001c",
            INIT_25 => X"0000002f0000002b000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000005600000067000000d100000024000000400000006a0000003400000037",
            INIT_27 => X"0000000000000000000000000000000000000061000000170000004200000073",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_2B => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000009b000000b3000000000000006800000000000000210000000000000000",
            INIT_2D => X"000000a900000098000000a00000007d000000c10000007c0000009c0000007d",
            INIT_2E => X"000000000000000000000000000000000000001c00000006000000b0000000c2",
            INIT_2F => X"0000000000000000000000000000000000000000000000110000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"00000050000000510000004b0000006100000062000000000000000000000000",
            INIT_35 => X"0000005a0000005e0000005b0000005300000088000000610000004100000049",
            INIT_36 => X"0000003c000000730000005f00000076000000600000005a000000680000002a",
            INIT_37 => X"0000005c0000005d00000041000000460000007b0000004e0000006d00000076",
            INIT_38 => X"0000002e0000002300000015000000100000004f0000003b0000004600000097",
            INIT_39 => X"000000000000000d00000000000000000000000000000000000000000000002f",
            INIT_3A => X"000000570000007b000000730000006300000000000000000000000000000000",
            INIT_3B => X"0000000500000040000000430000007000000045000000480000004b00000056",
            INIT_3C => X"00000024000000000000001e00000022000000320000002b0000004400000012",
            INIT_3D => X"00000021000000210000000000000009000000000000005d000000070000003c",
            INIT_3E => X"000000000000002b000000170000001900000015000000000000000600000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER2_INSTANCE1;


    MEM_GOLD_LAYER2_INSTANCE2 : if BRAM_NAME = "gold_layer2_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004a0000005e0000005a0000000000000000000000000000000000000000",
            INIT_01 => X"0000002600000000000000360000003c0000004700000031000000260000002c",
            INIT_02 => X"0000003100000046000000020000000e000000500000003e0000003a00000026",
            INIT_03 => X"00000035000000440000005a00000026000000350000003f0000002d0000002e",
            INIT_04 => X"0000001d000000000000002c00000008000000000000001c0000004400000049",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000001100000032000000000000000a00000000000000170000000000000000",
            INIT_09 => X"000000000000002e00000000000000000000004c000000000000001100000000",
            INIT_0A => X"000000000000000000000011000000000000001c000000760000000000000002",
            INIT_0B => X"0000003e000000180000001a000000860000007b000000120000006e00000000",
            INIT_0C => X"000001160000004c0000004800000035000000330000003d000000af00000000",
            INIT_0D => X"000000f0000000be000000c10000006c00000074000000d1000000be0000010a",
            INIT_0E => X"0000007b0000003e000000550000002b00000003000000350000001500000096",
            INIT_0F => X"000000110000005700000064000000400000001000000000000000340000001c",
            INIT_10 => X"0000002f0000002700000030000000400000001f00000040000000000000000a",
            INIT_11 => X"0000000000000000000000000000000000000000000000370000007600000017",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"00000009000000000000006c000000000000002b000000000000000000000000",
            INIT_14 => X"000000000000006f000000840000006500000000000000970000000000000000",
            INIT_15 => X"0000000000000079000000c400000062000000b000000000000000ed00000000",
            INIT_16 => X"0000007600000025000000000000004600000000000000920000000000000053",
            INIT_17 => X"0000002400000000000000a20000000000000000000000000000001f00000053",
            INIT_18 => X"00000000000000000000000b0000000000000011000000060000000000000000",
            INIT_19 => X"00000024000000320000005c000000110000001e000000000000000600000000",
            INIT_1A => X"00000042000000260000002c00000046000000340000008a000000500000009e",
            INIT_1B => X"0000002a000000220000003600000022000000970000002e0000005900000036",
            INIT_1C => X"000000a6000000af000000170000001f00000000000000270000003500000031",
            INIT_1D => X"00000028000000bd0000009a0000001c0000002100000066000000370000002b",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000001f0000000b000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000001800000030000000000000000000000000000000000000000000000000",
            INIT_23 => X"000000860000007e000000470000000000000019000000200000002a00000005",
            INIT_24 => X"000000a3000000ae0000007d000000d0000000b0000000b3000000a70000008a",
            INIT_25 => X"0000000000000000000000000000000200000000000000e1000000bf000000ac",
            INIT_26 => X"0000004e000000000000002a0000002f00000004000000000000000000000000",
            INIT_27 => X"000000000000003a000000000000005300000000000000650000000000000000",
            INIT_28 => X"0000001c00000000000000250000000000000050000000000000000500000011",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000008b00000000",
            INIT_2A => X"0000001200000000000000000000000400000000000000220000000000000000",
            INIT_2B => X"000000000000000000000000000000000000000a000000240000000d00000018",
            INIT_2C => X"000000330000000000000000000000120000005000000004000000000000004d",
            INIT_2D => X"000000000000009100000000000000000000003f000000000000001e00000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000250000000000000000",
            INIT_2F => X"00000000000000000000007700000000000000000000000a0000004400000000",
            INIT_30 => X"00000000000000a6000000050000004200000067000000000000000000000000",
            INIT_31 => X"0000000000000003000000000000000b00000038000000410000003000000061",
            INIT_32 => X"000000230000004e000000290000000000000000000000000000000000000000",
            INIT_33 => X"000000000000006f0000002d0000000000000023000000000000002200000000",
            INIT_34 => X"00000000000000000000000000000000000000000000005c0000002e00000005",
            INIT_35 => X"0000000000000000000000000000002c0000002e000000030000002b00000000",
            INIT_36 => X"00000000000000530000005e0000005e00000000000000000000000000000000",
            INIT_37 => X"000000b000000090000000390000003000000036000000300000000000000000",
            INIT_38 => X"00000079000000b40000006a000000680000004a0000006700000067000000a2",
            INIT_39 => X"00000000000000420000006a0000003400000043000000140000003b00000025",
            INIT_3A => X"00000027000000000000002c0000002200000000000000240000000000000034",
            INIT_3B => X"0000000000000000000000080000001700000033000000000000003c00000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000046",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000001700000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000010000002d0000000a000000160000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER2_INSTANCE2;


    MEM_GOLD_LAYER2_INSTANCE3 : if BRAM_NAME = "gold_layer2_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000008000000000000001e000000450000002f000000120000001700000003",
            INIT_01 => X"0000003a00000027000000390000004200000060000000000000000200000015",
            INIT_02 => X"000000880000007e0000007e000000480000000700000069000000260000003a",
            INIT_03 => X"000000ab000000a90000009e000000960000009200000066000000bb00000096",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER2_INSTANCE3;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE0 : if BRAM_NAME = "sampleifmap_layer0_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000009f000000a20000009c000000a0000000a6000000a50000009f0000009e",
            INIT_01 => X"000000aa000000a9000000a6000000a1000000a0000000a10000009f0000009e",
            INIT_02 => X"0000009400000096000000950000009c000000a0000000a0000000a2000000a7",
            INIT_03 => X"000000740000007e000000890000008f0000008d0000008c0000008f00000095",
            INIT_04 => X"000000a2000000a4000000a0000000a2000000a60000009f0000009700000098",
            INIT_05 => X"000000ab000000ab000000aa000000a30000009f0000009b0000009c000000a3",
            INIT_06 => X"0000008d0000008c0000008b00000091000000970000009a000000a0000000a9",
            INIT_07 => X"000000770000007d000000880000008f0000008e000000910000009300000095",
            INIT_08 => X"000000a5000000a5000000a3000000a0000000a70000009e0000009700000097",
            INIT_09 => X"000000a9000000a7000000a6000000a10000009d0000009e000000a2000000a3",
            INIT_0A => X"0000007200000065000000620000006e00000079000000910000009f000000aa",
            INIT_0B => X"00000078000000820000008b0000008e0000008c0000008f0000008600000078",
            INIT_0C => X"000000a9000000a9000000a7000000a7000000ae000000a00000009b0000009b",
            INIT_0D => X"000000a4000000a20000009d000000b1000000bf000000a7000000a5000000a5",
            INIT_0E => X"0000004a000000500000005c000000620000006700000068000000950000009e",
            INIT_0F => X"0000007f000000880000008c0000008c00000084000000710000005300000056",
            INIT_10 => X"000000a6000000a9000000a3000000a9000000aa000000a10000009c0000009b",
            INIT_11 => X"0000008e0000009200000097000000c3000000f6000000ad000000a4000000a4",
            INIT_12 => X"0000005d000000610000006a0000007000000071000000550000004e0000006f",
            INIT_13 => X"00000081000000850000008a000000800000006900000055000000540000004a",
            INIT_14 => X"000000a7000000a7000000a5000000a100000093000000820000008500000094",
            INIT_15 => X"0000004200000061000000800000009d000000b4000000a3000000a5000000a3",
            INIT_16 => X"0000005e00000072000000770000007a00000076000000590000004200000045",
            INIT_17 => X"000000860000008a0000008c0000006c000000430000003a0000005b00000063",
            INIT_18 => X"000000aa000000a8000000aa00000099000000580000002f0000006d0000007f",
            INIT_19 => X"00000044000000640000007f0000008100000093000000a4000000a6000000a9",
            INIT_1A => X"0000006b000000690000007c000000920000008400000053000000480000004e",
            INIT_1B => X"000000860000008d000000840000004f0000002e0000003f0000005500000073",
            INIT_1C => X"000000a8000000a5000000a70000008f000000460000002a0000006300000083",
            INIT_1D => X"00000058000000740000009000000082000000780000008c000000a1000000ab",
            INIT_1E => X"0000006a0000006600000088000000a30000007c0000004d000000550000005b",
            INIT_1F => X"000000880000008a0000006b0000003900000031000000360000005500000064",
            INIT_20 => X"000000a6000000a3000000a1000000990000007c0000003600000067000000aa",
            INIT_21 => X"00000056000000790000009c0000009d0000007d00000071000000ae000000a5",
            INIT_22 => X"0000005700000071000000920000008a00000051000000500000005400000052",
            INIT_23 => X"00000089000000850000004a0000002800000038000000470000005600000053",
            INIT_24 => X"000000990000009c0000009e000000ae0000009a0000005e00000086000000b4",
            INIT_25 => X"0000005d0000007d00000094000000ae0000009c000000cf000000ed000000cf",
            INIT_26 => X"0000006a000000850000008f000000890000004c0000003b0000004a00000056",
            INIT_27 => X"000000840000005f00000028000000320000004b000000540000005700000056",
            INIT_28 => X"0000007a0000009f0000009b000000b1000000a50000008e0000006c000000b7",
            INIT_29 => X"000000780000007d0000009c000000b7000000a4000000dc000000ed000000d5",
            INIT_2A => X"0000006b0000009b0000009d000000af0000005b0000002d000000500000004e",
            INIT_2B => X"000000680000003b000000290000003b0000004e000000580000006700000057",
            INIT_2C => X"00000086000000ad000000a6000000bb000000aa0000008700000064000000bc",
            INIT_2D => X"0000007500000086000000bd000000b9000000aa000000c7000000c200000075",
            INIT_2E => X"0000005d00000092000000a0000000d20000007d000000260000005400000066",
            INIT_2F => X"0000004c0000003e000000370000004900000055000000680000005e00000053",
            INIT_30 => X"0000009f000000b2000000a6000000ae000000af0000007f0000005a000000bd",
            INIT_31 => X"0000007b000000a0000000d8000000ba00000089000000a8000000a800000061",
            INIT_32 => X"0000005b0000007b0000009b000000c200000096000000320000007300000078",
            INIT_33 => X"000000490000004f0000004900000054000000560000005f0000005400000054",
            INIT_34 => X"000000a7000000ad0000008800000077000000b9000000980000005d000000bd",
            INIT_35 => X"0000008d000000b4000000e2000000bd000000a7000000910000009300000067",
            INIT_36 => X"000000570000007200000095000000ba0000009a00000047000000750000007e",
            INIT_37 => X"0000005e000000610000005a0000006400000063000000500000004800000050",
            INIT_38 => X"000000a70000009c0000006300000069000000ba000000a80000006c000000c2",
            INIT_39 => X"0000009a00000091000000ac000000be000000c60000008a0000007300000064",
            INIT_3A => X"0000006e0000008200000089000000b300000098000000470000006700000092",
            INIT_3B => X"000000750000006100000064000000730000006d0000005f0000005b00000055",
            INIT_3C => X"0000009b0000008c0000004e00000082000000b8000000ac00000084000000c5",
            INIT_3D => X"000000830000008700000091000000f2000000e60000008f0000008200000073",
            INIT_3E => X"000000570000007000000098000000a8000000900000005f0000006c00000079",
            INIT_3F => X"0000008800000079000000670000007800000070000000690000005700000047",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE0;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE1 : if BRAM_NAME = "sampleifmap_layer0_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000008a0000007e0000004e000000a8000000bf000000a800000092000000cb",
            INIT_01 => X"00000071000000710000008c000000a2000000ad0000009a000000600000008a",
            INIT_02 => X"0000006d00000087000000940000009c000000ab000000700000006900000065",
            INIT_03 => X"00000090000000970000007d0000006b000000650000005e0000004f0000004e",
            INIT_04 => X"0000009c000000600000005e000000b0000000b7000000a4000000a3000000d6",
            INIT_05 => X"0000007300000066000000740000007200000076000000810000006a00000094",
            INIT_06 => X"0000004b00000085000000800000004400000076000000900000006500000056",
            INIT_07 => X"0000008c000000960000008f0000007400000066000000470000003a0000003c",
            INIT_08 => X"0000008d000000560000007c000000b0000000ad000000a7000000b2000000d4",
            INIT_09 => X"00000093000000810000007c000000860000004d000000680000008700000099",
            INIT_0A => X"000000400000004b0000006b0000007500000084000000960000005c00000055",
            INIT_0B => X"000000970000009a000000a00000009b0000008500000056000000410000002c",
            INIT_0C => X"000000770000005600000090000000b1000000ae000000ab000000bb000000c7",
            INIT_0D => X"000000b8000000910000006c000000810000004600000090000000890000007a",
            INIT_0E => X"0000003400000033000000590000008600000089000000830000004900000074",
            INIT_0F => X"000000950000009e000000a4000000ab000000a3000000790000005a0000002f",
            INIT_10 => X"000000830000006300000098000000b5000000b1000000b3000000c3000000a5",
            INIT_11 => X"000000bf000000b20000007a0000005d000000500000005d00000067000000ab",
            INIT_12 => X"00000018000000260000002e0000003c00000057000000590000006400000096",
            INIT_13 => X"000000780000007f0000008000000090000000900000006c0000003c0000002e",
            INIT_14 => X"00000096000000530000008a000000b5000000b2000000b1000000c300000075",
            INIT_15 => X"000000c2000000be000000b0000000950000008600000085000000db000000f5",
            INIT_16 => X"0000003a0000003100000022000000230000003d0000006e0000007d000000a8",
            INIT_17 => X"000000370000003b000000450000004e00000048000000450000003a0000003d",
            INIT_18 => X"000000d30000006d0000008c000000b1000000b0000000ae000000af0000004f",
            INIT_19 => X"0000007a000000740000007c000000720000007c000000d0000000fc000000fd",
            INIT_1A => X"000000380000003300000032000000340000003c000000440000004400000068",
            INIT_1B => X"0000002a0000002b000000300000003b000000330000002b0000003300000038",
            INIT_1C => X"000000f6000000a5000000a5000000b2000000a8000000900000006000000029",
            INIT_1D => X"000000300000003100000031000000350000003c0000006e000000e3000000fd",
            INIT_1E => X"0000002b0000002e0000002e000000260000002a0000002e0000002a0000002d",
            INIT_1F => X"0000002d000000330000003500000037000000320000002e0000002e0000002a",
            INIT_20 => X"000000fe000000c200000084000000a6000000830000003b0000001d0000001d",
            INIT_21 => X"00000032000000310000003300000032000000320000003d0000008d000000f1",
            INIT_22 => X"0000002a00000026000000270000002300000022000000270000002a0000002f",
            INIT_23 => X"000000330000002e00000032000000380000003b0000003e000000380000002d",
            INIT_24 => X"00000100000000d7000000800000008000000049000000220000001e00000030",
            INIT_25 => X"0000002d0000002e0000003400000034000000320000003600000042000000bb",
            INIT_26 => X"0000002e0000002b00000028000000280000002700000024000000290000002b",
            INIT_27 => X"000000530000004600000032000000360000003b000000400000003e0000003b",
            INIT_28 => X"000000f0000000e00000008000000042000000290000001f0000002300000034",
            INIT_29 => X"0000002f0000002c0000002c0000003600000038000000310000003a0000007c",
            INIT_2A => X"0000003a000000360000002d0000002c0000002c0000002b0000002b0000002e",
            INIT_2B => X"0000004c000000550000004900000033000000240000002b0000002e00000036",
            INIT_2C => X"000000d3000000ca0000004e0000002c000000230000001d0000002300000032",
            INIT_2D => X"0000002d00000028000000300000003a00000030000000360000004100000061",
            INIT_2E => X"000000300000002700000027000000330000002e0000002f000000300000002f",
            INIT_2F => X"000000330000002e0000004300000043000000280000001c000000270000002f",
            INIT_30 => X"000000aa000000680000002e0000002900000021000000200000002300000032",
            INIT_31 => X"0000002d000000360000003a0000003d00000035000000340000003600000040",
            INIT_32 => X"00000027000000280000002a0000002e000000310000002e000000290000002a",
            INIT_33 => X"000000330000000f0000001f0000002f0000003f0000002c0000002800000025",
            INIT_34 => X"000000470000002a0000002b00000025000000260000001f0000002a00000044",
            INIT_35 => X"000000350000003a0000003800000031000000260000001b0000001f00000031",
            INIT_36 => X"00000021000000270000002d0000003200000035000000390000003c00000038",
            INIT_37 => X"000000280000000d0000002600000038000000490000004f0000003e0000002a",
            INIT_38 => X"000000280000002c0000002a000000270000002b00000023000000310000003d",
            INIT_39 => X"0000002f000000240000001d0000001b0000001e000000170000001b0000002a",
            INIT_3A => X"0000002b0000002b00000031000000450000004b000000420000003e00000038",
            INIT_3B => X"000000140000001d0000001a0000003c0000005d0000006d000000550000003c",
            INIT_3C => X"000000260000002800000028000000280000002b0000002d0000003800000036",
            INIT_3D => X"00000012000000130000001d000000190000001d000000160000001a00000024",
            INIT_3E => X"0000002d0000003400000035000000420000004a0000003d0000002f00000020",
            INIT_3F => X"0000001500000022000000180000003000000059000000690000005900000043",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE1;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE2 : if BRAM_NAME = "sampleifmap_layer0_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000071000000730000006d0000007000000076000000740000006f00000070",
            INIT_01 => X"0000007700000075000000750000006f0000006f00000074000000710000006f",
            INIT_02 => X"0000006a0000006b0000006b0000006d000000700000006f0000007100000075",
            INIT_03 => X"000000550000005b0000005f000000610000006100000062000000650000006b",
            INIT_04 => X"0000007200000075000000710000007000000074000000720000006e00000070",
            INIT_05 => X"000000730000007500000077000000710000006e0000006f0000006e00000074",
            INIT_06 => X"0000006400000066000000680000006e00000073000000700000006f00000073",
            INIT_07 => X"000000580000005b0000005f0000006200000061000000660000006600000069",
            INIT_08 => X"0000007500000075000000730000006a0000006f0000006f0000006d0000006e",
            INIT_09 => X"0000007100000072000000730000006f0000006d000000720000007300000073",
            INIT_0A => X"000000550000004d0000004e0000005a000000600000006f0000007200000074",
            INIT_0B => X"000000590000005f000000620000006300000063000000670000006000000056",
            INIT_0C => X"0000007700000078000000750000006e000000700000006d0000006e0000006b",
            INIT_0D => X"00000072000000730000006f00000082000000920000007b0000007500000073",
            INIT_0E => X"0000003f0000004b0000005a0000005a00000057000000500000006f00000070",
            INIT_0F => X"0000005e00000063000000650000006600000062000000550000003e00000046",
            INIT_10 => X"000000740000007800000071000000720000007200000073000000720000006b",
            INIT_11 => X"0000006c0000006f000000720000009c000000d6000000800000007400000071",
            INIT_12 => X"0000005e00000066000000720000006e00000067000000450000003500000050",
            INIT_13 => X"0000005d0000005e000000650000006000000053000000490000004e00000048",
            INIT_14 => X"000000730000007400000071000000730000007000000064000000680000006d",
            INIT_15 => X"000000320000004b000000660000007a0000008a00000076000000740000006f",
            INIT_16 => X"00000060000000740000007a000000790000007100000053000000380000003a",
            INIT_17 => X"0000005f0000006200000069000000540000003a0000003a0000005b00000064",
            INIT_18 => X"000000760000007300000076000000750000004a000000250000005f00000064",
            INIT_19 => X"00000043000000570000006c000000620000006b000000780000007400000075",
            INIT_1A => X"0000006600000063000000760000008e00000082000000540000004b00000053",
            INIT_1B => X"0000005d00000063000000620000003d0000002f00000047000000530000006f",
            INIT_1C => X"0000007400000072000000750000006f000000400000002b0000006000000073",
            INIT_1D => X"000000570000006a000000830000006e0000005e0000006d0000007100000077",
            INIT_1E => X"000000620000005d0000007c00000099000000760000004d000000580000005f",
            INIT_1F => X"0000006100000067000000530000002f000000350000003c000000510000005d",
            INIT_20 => X"0000007a00000075000000710000007c000000790000003a00000069000000a1",
            INIT_21 => X"000000500000006f0000008f0000008d00000069000000590000008700000079",
            INIT_22 => X"0000004f00000067000000870000007d000000470000004e0000005500000051",
            INIT_23 => X"000000670000006a0000003b000000230000003900000049000000520000004d",
            INIT_24 => X"000000760000007400000074000000950000009a000000640000008b000000b0",
            INIT_25 => X"000000550000006e000000830000009900000083000000b4000000d6000000b4",
            INIT_26 => X"000000620000007c000000850000007d00000044000000390000004a00000054",
            INIT_27 => X"000000670000004b0000001e000000310000004c000000550000005500000051",
            INIT_28 => X"0000005900000076000000700000009c000000a90000009700000074000000b7",
            INIT_29 => X"0000006f0000006c000000890000009f00000087000000bf000000e0000000c5",
            INIT_2A => X"000000640000009300000093000000a5000000550000002c000000500000004c",
            INIT_2B => X"000000510000002e000000240000003b0000004f000000580000006600000053",
            INIT_2C => X"0000005d0000007b00000078000000a7000000af000000900000006c000000bf",
            INIT_2D => X"0000006b00000077000000ab000000a10000008e000000ab000000b60000005f",
            INIT_2E => X"000000590000008b00000098000000c900000079000000260000005400000062",
            INIT_2F => X"0000003800000037000000350000004b00000057000000680000005d00000050",
            INIT_30 => X"0000006d0000007b0000007b0000009c000000b40000008600000060000000c2",
            INIT_31 => X"0000007100000095000000ca000000a600000072000000900000009a00000044",
            INIT_32 => X"000000580000007600000095000000bb00000093000000320000007200000072",
            INIT_33 => X"000000370000004a0000004900000057000000570000005f0000005400000053",
            INIT_34 => X"000000740000007c0000006a0000006e000000bc0000009a0000005f000000c0",
            INIT_35 => X"00000083000000ac000000d8000000ae000000950000007d0000008400000048",
            INIT_36 => X"000000550000006e00000090000000b500000098000000470000007200000075",
            INIT_37 => X"0000004900000059000000580000006500000064000000500000004900000050",
            INIT_38 => X"0000007a00000077000000590000006d000000ba000000a70000006b000000c4",
            INIT_39 => X"0000008f0000008c000000a5000000b4000000b90000007b0000006a0000004a",
            INIT_3A => X"0000006d0000008000000085000000af00000098000000470000006400000088",
            INIT_3B => X"0000005f0000005500000060000000740000006e000000600000005d00000056",
            INIT_3C => X"0000007d000000780000005300000089000000b2000000a700000081000000c5",
            INIT_3D => X"00000079000000820000008a000000ec000000dd00000083000000780000005e",
            INIT_3E => X"000000550000006c000000930000009f00000086000000580000006800000070",
            INIT_3F => X"0000006800000060000000560000006e0000006d000000680000005800000048",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE2;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE3 : if BRAM_NAME = "sampleifmap_layer0_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000007e0000007d00000056000000aa000000b6000000a400000092000000cb",
            INIT_01 => X"0000006a0000006a0000008400000098000000a30000008f0000005000000079",
            INIT_02 => X"00000069000000820000008d0000008a0000008f0000005a0000006500000065",
            INIT_03 => X"000000680000006c00000058000000530000005b0000005d0000004f0000004c",
            INIT_04 => X"000000950000006000000066000000b6000000b8000000a7000000a6000000d7",
            INIT_05 => X"0000006e0000005b000000690000006600000069000000740000005d00000089",
            INIT_06 => X"000000450000007e00000078000000380000006000000080000000670000005b",
            INIT_07 => X"0000006e00000074000000700000005e0000005d000000460000003800000038",
            INIT_08 => X"0000008b0000005800000083000000b8000000b5000000af000000b8000000d3",
            INIT_09 => X"0000008f000000750000006f00000079000000400000005a0000008000000094",
            INIT_0A => X"0000003b00000044000000630000006d000000750000008b000000600000005c",
            INIT_0B => X"0000006f00000073000000780000007700000069000000450000003e00000029",
            INIT_0C => X"000000790000005a00000095000000b6000000b3000000b0000000bd000000c0",
            INIT_0D => X"000000b00000008600000061000000760000003b00000086000000880000007c",
            INIT_0E => X"000000330000003100000056000000810000007c000000770000004b00000076",
            INIT_0F => X"0000006b0000006f0000007100000079000000760000005b0000005a00000031",
            INIT_10 => X"00000087000000670000009d000000b5000000ad000000b2000000c10000009c",
            INIT_11 => X"000000b6000000ad000000760000005a0000004d0000005a00000069000000af",
            INIT_12 => X"000000210000002e000000340000003d0000004d0000004e0000006400000094",
            INIT_13 => X"00000069000000710000006d0000007b0000007d000000640000004700000039",
            INIT_14 => X"000000990000005700000090000000b3000000a9000000b2000000c800000078",
            INIT_15 => X"000000c0000000c4000000b60000009c0000008d0000008c000000de000000f7",
            INIT_16 => X"000000510000004600000036000000310000003e0000006d00000085000000ac",
            INIT_17 => X"0000005a0000005c000000600000006800000065000000630000005400000055",
            INIT_18 => X"000000d30000007000000092000000b1000000ac000000b7000000c500000069",
            INIT_19 => X"00000085000000850000008d000000840000008f000000e0000000fd000000fc",
            INIT_1A => X"0000005d00000055000000540000005400000052000000570000005d0000007c",
            INIT_1B => X"0000005f00000061000000610000006c00000068000000600000005b0000005e",
            INIT_1C => X"000000f5000000a6000000aa000000b6000000ae000000a80000008900000059",
            INIT_1D => X"000000480000004b0000004c000000500000005800000088000000e7000000fb",
            INIT_1E => X"00000057000000590000005a000000560000005200000051000000510000004f",
            INIT_1F => X"0000005a0000005f0000005e00000060000000600000005e0000005d00000059",
            INIT_20 => X"000000fa000000bd00000088000000b30000009900000066000000570000005b",
            INIT_21 => X"00000054000000530000005500000054000000540000005e0000009f000000f5",
            INIT_22 => X"000000590000005500000056000000530000004f000000520000005400000056",
            INIT_23 => X"000000670000005e00000063000000660000006500000067000000670000005c",
            INIT_24 => X"000000fd000000d500000088000000940000006a000000550000005e0000006f",
            INIT_25 => X"00000052000000530000005a0000005a000000580000005b0000005d000000c6",
            INIT_26 => X"0000005f0000005c000000590000005600000053000000500000005100000052",
            INIT_27 => X"000000890000007b000000690000006c0000006c0000006d0000006e0000006c",
            INIT_28 => X"000000f5000000e5000000910000005f00000053000000560000006300000072",
            INIT_29 => X"0000005300000052000000520000005c0000005e000000570000005c0000008f",
            INIT_2A => X"0000006e0000006a000000610000005a00000058000000560000005300000054",
            INIT_2B => X"0000007d0000008a000000820000006c0000005b0000005f0000006100000069",
            INIT_2C => X"000000e4000000db0000006a000000530000005600000059000000620000006e",
            INIT_2D => X"00000052000000500000005700000061000000570000005e000000680000007e",
            INIT_2E => X"000000660000005d0000005c0000006100000059000000590000005700000054",
            INIT_2F => X"00000060000000620000007e0000008100000065000000550000005d00000065",
            INIT_30 => X"000000c5000000850000005400000058000000580000005c000000610000006c",
            INIT_31 => X"000000530000006000000064000000670000005f0000005e0000006100000064",
            INIT_32 => X"0000005c0000005d0000005f0000005c0000005c00000058000000500000004f",
            INIT_33 => X"0000005d0000003c0000005a0000006e0000007d000000660000005d0000005a",
            INIT_34 => X"0000006b0000004f00000059000000570000005b00000058000000640000007c",
            INIT_35 => X"0000005c00000066000000640000005d00000052000000470000004d00000059",
            INIT_36 => X"00000053000000580000005e0000005f0000006100000063000000630000005e",
            INIT_37 => X"000000550000004000000061000000740000008300000084000000700000005b",
            INIT_38 => X"00000051000000580000005c0000005a0000005b000000550000006600000074",
            INIT_39 => X"000000560000005000000049000000470000004a000000430000004800000055",
            INIT_3A => X"00000058000000580000005f00000071000000770000006d000000650000005f",
            INIT_3B => X"00000040000000520000005200000073000000910000009c0000008200000069",
            INIT_3C => X"00000051000000570000005c000000590000005600000059000000690000006b",
            INIT_3D => X"0000003a0000003f00000049000000450000004900000042000000450000004f",
            INIT_3E => X"000000570000005f000000600000006f00000077000000680000005700000046",
            INIT_3F => X"00000043000000540000004d000000630000008700000092000000830000006d",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE3;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE4 : if BRAM_NAME = "sampleifmap_layer0_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002d0000002f000000290000002e00000035000000330000002f00000031",
            INIT_01 => X"0000002c0000002d00000029000000310000003400000029000000290000002c",
            INIT_02 => X"0000002b0000002d0000002d0000002c0000002b000000270000002600000028",
            INIT_03 => X"00000021000000240000002400000026000000290000002b000000270000002c",
            INIT_04 => X"0000002d0000002f0000002b00000031000000380000002d0000002800000033",
            INIT_05 => X"000000210000002800000029000000340000003600000029000000260000002e",
            INIT_06 => X"000000300000003400000037000000350000003200000029000000210000001e",
            INIT_07 => X"00000022000000200000001f00000022000000260000002d0000002e00000032",
            INIT_08 => X"0000002d0000002d0000002c0000002a0000003000000024000000210000002f",
            INIT_09 => X"0000002300000025000000260000003300000039000000300000002b0000002b",
            INIT_0A => X"000000320000002f000000320000003400000031000000360000002f00000027",
            INIT_0B => X"0000002100000022000000220000002300000027000000330000003700000030",
            INIT_0C => X"00000030000000300000002e0000002b0000002c0000001f0000002000000028",
            INIT_0D => X"000000360000002f000000290000004b0000005f000000390000002d0000002c",
            INIT_0E => X"0000003200000042000000540000004c000000410000002f000000430000003a",
            INIT_0F => X"0000002400000027000000270000002b0000002e0000002d0000002700000034",
            INIT_10 => X"0000002c0000002f000000280000002b0000002f000000310000003000000029",
            INIT_11 => X"000000470000003c000000380000006b000000a40000003b0000002a00000029",
            INIT_12 => X"0000005d00000069000000760000006f00000062000000380000001f00000032",
            INIT_13 => X"00000024000000240000002e000000300000002d0000002f0000004600000043",
            INIT_14 => X"0000002900000029000000270000002c00000035000000390000004000000036",
            INIT_15 => X"0000001f0000002b0000003a0000004e000000550000002a0000002700000025",
            INIT_16 => X"00000060000000740000007a000000780000006e0000004c0000002d0000002b",
            INIT_17 => X"000000280000002c0000003a00000031000000250000002f0000005600000061",
            INIT_18 => X"0000002b000000280000002b000000300000001c000000110000005000000039",
            INIT_19 => X"00000039000000460000004b0000003b0000003400000027000000250000002a",
            INIT_1A => X"0000005e0000005a0000006c00000084000000790000004a0000004000000048",
            INIT_1B => X"00000027000000300000003a0000002400000027000000450000004d00000067",
            INIT_1C => X"00000027000000240000002a0000003800000029000000260000005c0000005a",
            INIT_1D => X"0000004f0000005d0000006b0000004d00000031000000330000003300000031",
            INIT_1E => X"0000005800000051000000700000008c0000006b000000450000005200000058",
            INIT_1F => X"00000027000000330000003200000020000000310000003a0000004a00000054",
            INIT_20 => X"00000032000000290000002b00000052000000710000003b0000006900000090",
            INIT_21 => X"0000004a0000006500000080000000790000004e0000003b0000005f00000042",
            INIT_22 => X"000000460000005d0000007b000000700000003d00000049000000520000004d",
            INIT_23 => X"0000002d0000003b000000230000001b00000035000000430000004c00000045",
            INIT_24 => X"0000003c0000002f000000330000007000000095000000690000008f000000a3",
            INIT_25 => X"0000004f0000006b0000007d0000009100000077000000a6000000c600000092",
            INIT_26 => X"00000059000000720000007a000000700000003a00000035000000470000004f",
            INIT_27 => X"000000390000002c0000000f0000002b000000470000004e0000004e0000004a",
            INIT_28 => X"0000002f00000033000000320000007a000000a80000009e0000007a000000af",
            INIT_29 => X"0000006800000068000000840000009b00000083000000bc000000e2000000b3",
            INIT_2A => X"0000005c0000008a000000890000009a0000004d000000280000004d00000045",
            INIT_2B => X"0000002e0000001f000000210000003b000000490000004f000000600000004d",
            INIT_2C => X"0000002c000000370000003b00000088000000b20000009900000074000000bd",
            INIT_2D => X"0000005f0000006a0000009f0000009700000085000000a4000000bc00000050",
            INIT_2E => X"00000052000000820000008e000000c000000071000000220000004f00000059",
            INIT_2F => X"0000001a00000030000000370000004e000000510000005e000000580000004b",
            INIT_30 => X"0000002f000000350000004400000085000000b90000009000000069000000c2",
            INIT_31 => X"0000006200000081000000b7000000940000005e0000007e000000980000002c",
            INIT_32 => X"000000530000006f0000008c000000b20000008c0000002f0000006d00000069",
            INIT_33 => X"000000180000004000000049000000590000005100000055000000500000004f",
            INIT_34 => X"000000320000003a0000004200000062000000c0000000a300000067000000c1",
            INIT_35 => X"000000750000009d000000c80000009b0000007f000000670000007800000027",
            INIT_36 => X"000000500000006800000088000000ae00000093000000440000006d0000006b",
            INIT_37 => X"000000220000004500000051000000630000005e00000048000000460000004c",
            INIT_38 => X"000000370000003e000000430000006d000000bc000000ac00000070000000c4",
            INIT_39 => X"000000860000008c0000009f000000a9000000a9000000670000005800000022",
            INIT_3A => X"000000690000007a0000007f000000aa00000095000000460000005f0000007d",
            INIT_3B => X"0000002f00000035000000500000006f000000680000005a0000005b00000053",
            INIT_3C => X"0000004d000000580000004d0000008e000000b5000000ae00000088000000c5",
            INIT_3D => X"000000700000008200000089000000e6000000d3000000740000005d00000034",
            INIT_3E => X"00000050000000650000008a00000092000000760000004b0000005f00000065",
            INIT_3F => X"0000003000000030000000360000005d00000063000000630000005700000044",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE4;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE5 : if BRAM_NAME = "sampleifmap_layer0_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000710000007e0000005a000000ac000000bc000000b2000000a0000000cc",
            INIT_01 => X"0000005a00000058000000750000008d0000009b000000850000002500000052",
            INIT_02 => X"00000061000000760000007e0000006d000000680000003a000000570000005c",
            INIT_03 => X"0000002e000000370000002d00000037000000520000005e0000004d00000048",
            INIT_04 => X"000000910000006600000069000000ba000000c2000000b8000000b4000000d7",
            INIT_05 => X"000000620000004900000059000000590000005f000000690000003d0000006f",
            INIT_06 => X"0000003d00000073000000690000002000000040000000660000005f00000058",
            INIT_07 => X"000000360000004000000044000000400000004e000000410000003500000033",
            INIT_08 => X"0000008f0000006000000085000000bc000000c1000000bd000000c0000000cd",
            INIT_09 => X"0000008500000064000000600000006c00000037000000500000006f0000008d",
            INIT_0A => X"000000340000003a000000560000005c0000005d000000780000005d0000005d",
            INIT_0B => X"0000002e0000002d000000360000003e0000003b000000280000003c00000027",
            INIT_0C => X"000000840000006300000098000000b8000000b9000000b5000000bb000000b4",
            INIT_0D => X"000000a80000007b000000560000006c000000330000007e0000008700000082",
            INIT_0E => X"000000320000002c0000004e0000007600000069000000670000004900000076",
            INIT_0F => X"0000002e000000320000003400000040000000440000003c0000005d00000034",
            INIT_10 => X"000000920000006f000000a0000000b4000000ac000000af000000bb00000092",
            INIT_11 => X"000000b1000000ad000000740000005600000049000000570000006f000000b9",
            INIT_12 => X"000000290000003300000036000000390000003f000000420000006500000094",
            INIT_13 => X"0000003f000000450000003d0000004c000000520000004b0000005300000045",
            INIT_14 => X"0000009f0000005b00000093000000b3000000a8000000b0000000c80000007c",
            INIT_15 => X"000000c5000000d0000000c0000000a40000009300000090000000e1000000fa",
            INIT_16 => X"0000006600000057000000440000003a0000003e0000006d0000008f000000b5",
            INIT_17 => X"00000073000000700000007000000078000000770000007a0000006f0000006e",
            INIT_18 => X"000000d10000007100000096000000b6000000b1000000c0000000d500000085",
            INIT_19 => X"000000980000009c000000a2000000950000009d000000e8000000fc000000f7",
            INIT_1A => X"0000007d000000730000006e0000006f00000065000000680000007700000094",
            INIT_1B => X"0000008400000089000000840000008e0000008d000000870000008200000083",
            INIT_1C => X"000000ed000000a4000000ae000000c0000000bc000000bc000000a800000087",
            INIT_1D => X"000000650000006b00000069000000690000006f00000099000000e4000000f1",
            INIT_1E => X"000000800000007e0000007d0000007d00000074000000710000007800000073",
            INIT_1F => X"000000850000008b000000860000008700000089000000890000008b00000084",
            INIT_20 => X"000000f2000000b500000089000000bf000000b000000086000000820000008d",
            INIT_21 => X"00000074000000780000007900000077000000760000007f000000af000000f5",
            INIT_22 => X"000000820000007d0000007d0000007800000071000000730000007500000075",
            INIT_23 => X"000000950000008c00000090000000920000008e0000008e0000009100000086",
            INIT_24 => X"000000f9000000d10000008f000000a7000000880000007c0000008c000000a2",
            INIT_25 => X"00000073000000790000007f0000007f0000007d0000008000000076000000cd",
            INIT_26 => X"0000008a00000086000000830000007b00000075000000710000007000000071",
            INIT_27 => X"000000b6000000a7000000980000009a00000095000000930000009800000096",
            INIT_28 => X"000000f7000000ea000000a40000007e0000007a0000008200000093000000a5",
            INIT_29 => X"00000077000000770000007700000081000000830000007b0000007200000099",
            INIT_2A => X"0000009a000000960000008d000000830000007f0000007b0000007700000077",
            INIT_2B => X"000000a9000000b6000000b20000009e0000008a0000008c0000008d00000096",
            INIT_2C => X"000000ea000000e90000008a0000007e000000850000008a00000095000000a2",
            INIT_2D => X"00000077000000740000007b000000850000007c000000810000007e0000008c",
            INIT_2E => X"000000940000008b0000008a0000008c00000084000000820000007e0000007a",
            INIT_2F => X"0000008b0000008e000000b0000000b600000099000000850000008b00000093",
            INIT_30 => X"000000d30000009f0000007d0000008a0000008d0000008f00000093000000a1",
            INIT_31 => X"0000007800000083000000870000008b00000082000000800000007900000077",
            INIT_32 => X"000000880000008a0000008b0000008800000087000000820000007800000076",
            INIT_33 => X"00000088000000670000008c000000a4000000b2000000970000008a00000087",
            INIT_34 => X"0000008500000071000000840000008b000000920000008900000094000000b1",
            INIT_35 => X"0000008000000089000000870000008000000075000000690000006900000072",
            INIT_36 => X"0000007d0000008300000088000000890000008a0000008b0000008900000083",
            INIT_37 => X"0000007f0000006c00000092000000a8000000b5000000b30000009a00000085",
            INIT_38 => X"000000700000007d000000860000008b0000008f0000008400000094000000a8",
            INIT_39 => X"00000078000000730000006c0000006a0000006d000000660000006800000073",
            INIT_3A => X"0000007f0000007f00000086000000980000009c000000900000008700000080",
            INIT_3B => X"0000006b0000007e00000082000000a4000000be000000c5000000aa00000090",
            INIT_3C => X"000000730000007b0000008400000086000000860000008400000095000000a0",
            INIT_3D => X"00000059000000620000006c000000680000006c000000650000006900000072",
            INIT_3E => X"0000007b00000082000000830000009100000098000000890000007600000064",
            INIT_3F => X"0000006e000000810000007c00000091000000af000000b6000000a700000091",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE5;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE6 : if BRAM_NAME = "sampleifmap_layer0_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000e8000000e8000000e8000000e8000000e8000000e8000000e7000000eb",
            INIT_01 => X"000000e9000000e9000000e9000000e9000000e9000000e9000000e8000000e8",
            INIT_02 => X"000000e9000000e8000000e8000000e8000000e6000000e7000000e8000000e9",
            INIT_03 => X"000000e8000000e9000000e9000000e8000000e8000000e8000000e9000000e8",
            INIT_04 => X"000000eb000000eb000000eb000000eb000000eb000000eb000000eb000000ee",
            INIT_05 => X"000000ec000000ec000000ec000000ec000000ec000000ec000000eb000000eb",
            INIT_06 => X"000000ec000000eb000000ea000000ea000000ea000000ec000000ec000000ed",
            INIT_07 => X"000000eb000000ec000000ec000000eb000000eb000000eb000000ec000000ec",
            INIT_08 => X"000000ea000000ea000000ea000000ea000000ea000000ea000000ea000000ed",
            INIT_09 => X"000000eb000000eb000000ea000000ea000000ea000000ea000000ea000000ea",
            INIT_0A => X"000000ea000000e7000000e7000000e3000000ea000000eb000000ec000000ec",
            INIT_0B => X"000000ea000000eb000000eb000000ea000000ea000000ea000000ea000000ea",
            INIT_0C => X"000000eb000000eb000000eb000000eb000000eb000000eb000000eb000000ee",
            INIT_0D => X"000000eb000000eb000000ea000000ea000000ea000000ea000000ea000000ea",
            INIT_0E => X"000000e4000000cf000000d1000000ba000000df000000e4000000e8000000e9",
            INIT_0F => X"000000eb000000eb000000eb000000ea000000ea000000ea000000ea000000ec",
            INIT_10 => X"000000eb000000eb000000eb000000eb000000eb000000eb000000ea000000ed",
            INIT_11 => X"000000eb000000eb000000ea000000ea000000eb000000eb000000ea000000ea",
            INIT_12 => X"000000e6000000d6000000c3000000a3000000cb000000db000000e9000000ec",
            INIT_13 => X"000000ec000000ec000000ec000000eb000000eb000000eb000000eb000000ed",
            INIT_14 => X"000000eb000000eb000000ec000000ec000000ec000000ec000000ec000000ef",
            INIT_15 => X"000000e5000000eb000000e8000000ea000000ed000000ed000000eb000000ea",
            INIT_16 => X"000000e2000000cf000000b8000000a5000000ae000000b9000000c2000000d0",
            INIT_17 => X"000000ed000000ed000000ed000000ec000000ec000000ec000000ec000000ec",
            INIT_18 => X"000000ec000000ed000000ed000000ea000000e7000000e8000000e4000000e4",
            INIT_19 => X"000000dd000000e9000000e0000000e1000000ef000000ef000000ed000000ed",
            INIT_1A => X"000000c60000009c0000008f000000900000009a0000009f000000a1000000b7",
            INIT_1B => X"000000ef000000ed000000ec000000eb000000eb000000eb000000ec000000e9",
            INIT_1C => X"000000ee000000ed000000ea000000e5000000e3000000e6000000e0000000d4",
            INIT_1D => X"000000d6000000e9000000db000000c9000000f0000000ef000000ef000000ef",
            INIT_1E => X"000000ba000000a20000009f000000a5000000ad000000b8000000b9000000c1",
            INIT_1F => X"000000ee000000ed000000ec000000ea000000e9000000e9000000ea000000e5",
            INIT_20 => X"000000ee000000ec000000e7000000e3000000e1000000e1000000dd000000d8",
            INIT_21 => X"000000e6000000e9000000dc000000c5000000ef000000ed000000ee000000ee",
            INIT_22 => X"000000da000000d9000000d2000000d1000000d0000000db000000d1000000d1",
            INIT_23 => X"000000ee000000ed000000eb000000e6000000e6000000e4000000e4000000e1",
            INIT_24 => X"000000ed000000eb000000e1000000ac000000880000007c0000007700000076",
            INIT_25 => X"000000ec000000e8000000e2000000d6000000e9000000eb000000eb000000ec",
            INIT_26 => X"000000b9000000c9000000d9000000e1000000e1000000e7000000e3000000e4",
            INIT_27 => X"000000ee000000ec000000eb000000df000000ba000000a7000000a7000000ac",
            INIT_28 => X"000000e5000000e3000000de000000920000006f0000006c000000670000006d",
            INIT_29 => X"000000e6000000e8000000e7000000e5000000e6000000e7000000ea000000ec",
            INIT_2A => X"0000008900000092000000a4000000bf000000df000000e5000000e7000000e7",
            INIT_2B => X"000000ed000000eb000000ea000000d800000095000000790000008000000086",
            INIT_2C => X"000000d3000000d5000000df000000d1000000c8000000c7000000bc000000c3",
            INIT_2D => X"000000dc000000d8000000d3000000d1000000d2000000db000000dc000000d8",
            INIT_2E => X"000000b2000000b5000000af000000b7000000da000000e1000000e2000000e1",
            INIT_2F => X"000000ec000000ea000000e7000000db000000b90000008e000000aa000000ba",
            INIT_30 => X"000000ab000000cb000000d6000000df000000d6000000ca000000bf000000c1",
            INIT_31 => X"0000007a0000006f000000650000005d00000062000000ae000000cf000000b1",
            INIT_32 => X"000000d9000000df000000dc000000da000000df000000ca0000009900000089",
            INIT_33 => X"000000eb000000e8000000dd000000db000000de000000c4000000d4000000dd",
            INIT_34 => X"000000be000000bf000000aa0000008a0000007d000000710000006f00000071",
            INIT_35 => X"0000004200000035000000310000002d000000360000009e000000d8000000d0",
            INIT_36 => X"000000cf000000df000000e3000000e9000000ea000000dd0000009f00000066",
            INIT_37 => X"000000dd000000d3000000bc000000b3000000c7000000d4000000d3000000ca",
            INIT_38 => X"000000c3000000970000008b0000007b000000440000003f000000450000003d",
            INIT_39 => X"000000b50000008a000000650000005f00000067000000a3000000ce000000d6",
            INIT_3A => X"00000083000000930000009e000000b7000000cd000000db000000dd000000cf",
            INIT_3B => X"000000c5000000b60000008a000000800000008500000088000000820000007d",
            INIT_3C => X"000000a30000007700000060000000840000007f000000550000003a00000028",
            INIT_3D => X"000000c8000000da000000c6000000b7000000b5000000b6000000b8000000ad",
            INIT_3E => X"000000630000005e000000620000007400000084000000910000009f000000ae",
            INIT_3F => X"000000b9000000bc0000009d000000960000008a0000007a0000006b00000069",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE6;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE7 : if BRAM_NAME = "sampleifmap_layer0_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ac0000008d000000760000008a000000ce000000860000001a0000000d",
            INIT_01 => X"000000b0000000e2000000e6000000e0000000e4000000dc000000cf000000b5",
            INIT_02 => X"0000009a00000095000000950000009a000000910000008e0000008a00000090",
            INIT_03 => X"0000009d000000a5000000b2000000be000000bb000000ad000000a00000009d",
            INIT_04 => X"000000e2000000d4000000c7000000c5000000e1000000c80000003a00000005",
            INIT_05 => X"000000d2000000dd000000df000000d1000000e6000000e8000000e9000000e5",
            INIT_06 => X"000000b8000000c0000000c2000000bd000000bc000000c1000000b4000000c6",
            INIT_07 => X"0000008a00000080000000830000008800000090000000a1000000ab000000ac",
            INIT_08 => X"000000c2000000c2000000c0000000b8000000ba000000be0000009100000027",
            INIT_09 => X"000000930000009a000000b4000000b1000000be000000c0000000bf000000c2",
            INIT_0A => X"0000006f0000007e000000840000007200000071000000920000009c00000091",
            INIT_0B => X"000000810000008100000079000000690000005e0000005d0000005b0000005c",
            INIT_0C => X"000000820000007f0000008000000083000000890000008f000000a20000007a",
            INIT_0D => X"00000064000000680000007c00000081000000810000007f0000008000000083",
            INIT_0E => X"00000053000000570000005e0000005e0000005e000000700000007600000066",
            INIT_0F => X"0000008200000079000000730000006c000000650000005d0000005300000050",
            INIT_10 => X"0000005a000000570000005700000054000000500000004d0000004c00000049",
            INIT_11 => X"00000078000000760000007600000073000000710000006b000000660000005e",
            INIT_12 => X"000000500000004f000000550000005f000000640000006a0000006e00000073",
            INIT_13 => X"000000880000007d000000710000005c00000052000000500000004d00000050",
            INIT_14 => X"000000160000001400000015000000120000001200000009000000030000000d",
            INIT_15 => X"00000046000000420000003c00000034000000300000002a000000220000001a",
            INIT_16 => X"000000390000003500000035000000370000003c000000430000004800000047",
            INIT_17 => X"0000008900000082000000780000006800000057000000480000003900000039",
            INIT_18 => X"0000000300000008000000160000002400000020000000080000000b00000024",
            INIT_19 => X"0000000300000001000000050000000600000000000000000000000000000001",
            INIT_1A => X"000000270000001e00000016000000150000001500000015000000180000000d",
            INIT_1B => X"00000099000000860000007a000000740000007b000000710000005500000039",
            INIT_1C => X"0000001b0000003100000046000000470000001b0000000d0000001a00000023",
            INIT_1D => X"0000000a0000001f00000039000000110000000000000002000000050000000f",
            INIT_1E => X"000000560000003e00000029000000190000000e000000070000000400000004",
            INIT_1F => X"000000ac0000009200000084000000750000007200000084000000900000007a",
            INIT_20 => X"0000002400000036000000410000002d00000003000000040000000d00000010",
            INIT_21 => X"00000083000000a1000000760000000700000000000000020000000400000012",
            INIT_22 => X"000000970000009a0000008a000000760000006d000000690000006900000070",
            INIT_23 => X"000000b8000000a40000008e00000081000000780000006a000000690000007f",
            INIT_24 => X"00000015000000200000001e0000000c00000000000000000000000c00000028",
            INIT_25 => X"000000cd000000b6000000440000000000000003000000020000000200000007",
            INIT_26 => X"000000670000007b00000096000000ac000000bb000000c3000000c2000000c4",
            INIT_27 => X"000000b9000000ab0000009800000084000000810000007a000000680000005f",
            INIT_28 => X"0000000c000000120000000c0000000400000001000000010000001a00000045",
            INIT_29 => X"000000cb00000099000000200000000100000004000000020000000200000004",
            INIT_2A => X"0000005e000000510000005b000000770000009b000000b3000000bf000000c3",
            INIT_2B => X"000000b8000000ad000000a200000090000000810000007d0000007d00000075",
            INIT_2C => X"0000000400000007000000050000000200000002000000010000002f00000053",
            INIT_2D => X"000000cd0000008e0000001b0000000100000003000000010000000100000001",
            INIT_2E => X"0000007900000066000000550000004a0000005500000079000000a9000000c6",
            INIT_2F => X"000000ba000000b0000000a50000009300000084000000790000007a00000080",
            INIT_30 => X"000000010000000100000001000000020000000300000006000000360000005c",
            INIT_31 => X"0000009d000000660000000f0000000000000001000000010000000100000001",
            INIT_32 => X"0000007c0000007a00000073000000630000004a000000380000004a00000075",
            INIT_33 => X"000000bc000000b1000000a20000009400000088000000800000007d0000007b",
            INIT_34 => X"000000020000000200000005000000080000000b000000130000002b00000057",
            INIT_35 => X"000000470000002a000000040000000000000002000000030000000300000003",
            INIT_36 => X"000000740000007b000000860000008400000071000000500000003900000035",
            INIT_37 => X"000000bc000000b6000000a90000009c0000008f0000008b0000008300000078",
            INIT_38 => X"0000001000000011000000160000001b0000001f000000240000002e00000052",
            INIT_39 => X"0000004000000025000000170000001300000013000000140000001300000012",
            INIT_3A => X"0000007300000075000000830000008b00000080000000740000006800000057",
            INIT_3B => X"000000bb000000b9000000ae0000009f000000940000008b000000830000007b",
            INIT_3C => X"000000300000002e0000002f00000033000000370000003a0000003e00000055",
            INIT_3D => X"0000006800000051000000440000003b00000037000000350000003300000031",
            INIT_3E => X"0000007a00000072000000760000007f0000007f000000850000007f00000074",
            INIT_3F => X"000000ba000000b4000000a80000009e000000950000008d0000008800000081",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE7;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE8 : if BRAM_NAME = "sampleifmap_layer0_instance8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000e8000000e8000000e8000000e8000000e8000000e8000000e7000000eb",
            INIT_01 => X"000000e8000000e9000000e9000000e9000000e9000000e9000000e8000000e8",
            INIT_02 => X"000000e9000000e8000000e7000000e8000000e9000000e9000000e7000000e7",
            INIT_03 => X"000000e8000000e9000000e9000000e8000000e8000000e8000000e9000000e9",
            INIT_04 => X"000000eb000000eb000000eb000000eb000000eb000000eb000000eb000000ee",
            INIT_05 => X"000000ec000000ec000000ec000000ec000000ec000000ec000000eb000000eb",
            INIT_06 => X"000000ec000000ec000000ea000000eb000000ec000000ec000000ea000000ea",
            INIT_07 => X"000000eb000000ec000000ec000000eb000000eb000000eb000000ec000000ec",
            INIT_08 => X"000000ea000000ea000000ea000000ea000000ea000000ea000000ea000000ed",
            INIT_09 => X"000000ea000000eb000000ea000000ea000000ea000000ea000000ea000000ea",
            INIT_0A => X"000000ea000000e9000000eb000000e6000000eb000000eb000000ea000000e9",
            INIT_0B => X"000000ea000000eb000000eb000000ea000000ea000000ea000000ea000000ea",
            INIT_0C => X"000000eb000000eb000000eb000000eb000000eb000000eb000000eb000000ee",
            INIT_0D => X"000000eb000000eb000000ea000000ea000000ea000000ea000000ea000000ea",
            INIT_0E => X"000000e4000000d2000000d8000000c0000000e2000000e6000000e8000000e9",
            INIT_0F => X"000000eb000000eb000000eb000000ea000000ea000000ea000000ea000000eb",
            INIT_10 => X"000000eb000000eb000000eb000000eb000000eb000000eb000000ea000000ed",
            INIT_11 => X"000000eb000000eb000000ea000000ea000000eb000000eb000000ea000000ea",
            INIT_12 => X"000000e5000000da000000cd000000ac000000d2000000e1000000ed000000ee",
            INIT_13 => X"000000ec000000ec000000ec000000ec000000eb000000eb000000eb000000eb",
            INIT_14 => X"000000eb000000ec000000eb000000eb000000eb000000eb000000eb000000ef",
            INIT_15 => X"000000e7000000ed000000e9000000eb000000ec000000ec000000eb000000ea",
            INIT_16 => X"000000e4000000d7000000c4000000b3000000bc000000c6000000cd000000d8",
            INIT_17 => X"000000ed000000ed000000ed000000ec000000ec000000ec000000ec000000eb",
            INIT_18 => X"000000ed000000ed000000ec000000e8000000e4000000e6000000e3000000e5",
            INIT_19 => X"000000e2000000ed000000e4000000e5000000ed000000ec000000eb000000eb",
            INIT_1A => X"000000ce000000a90000009f000000a3000000b0000000b4000000b4000000c5",
            INIT_1B => X"000000ed000000ed000000ee000000ec000000eb000000ec000000ed000000ee",
            INIT_1C => X"000000ed000000ee000000ed000000ea000000e8000000ea000000e6000000dc",
            INIT_1D => X"000000da000000ec000000de000000cc000000ee000000ec000000ed000000ed",
            INIT_1E => X"000000c7000000b0000000ae000000b6000000bf000000c9000000c9000000cc",
            INIT_1F => X"000000ee000000ef000000ef000000ef000000ee000000ee000000ef000000ef",
            INIT_20 => X"000000ec000000ed000000ee000000f0000000ef000000ee000000ec000000ea",
            INIT_21 => X"000000e7000000ea000000dd000000c6000000ef000000ed000000ec000000ec",
            INIT_22 => X"000000eb000000e9000000e0000000dd000000da000000e4000000d8000000d5",
            INIT_23 => X"000000ee000000f0000000f0000000f0000000f0000000ef000000ee000000f0",
            INIT_24 => X"000000ea000000ec000000ea000000bc0000009b0000008e0000008a0000008c",
            INIT_25 => X"000000ed000000ea000000e4000000d8000000ed000000ed000000eb000000e9",
            INIT_26 => X"000000cc000000db000000e9000000ed000000e8000000ec000000e6000000e6",
            INIT_27 => X"000000f0000000f0000000f1000000eb000000c7000000b4000000b3000000bd",
            INIT_28 => X"000000e2000000e4000000e50000009f0000007f0000007d0000007900000082",
            INIT_29 => X"000000eb000000ed000000eb000000ea000000ed000000ec000000ea000000e8",
            INIT_2A => X"0000009c000000a5000000b8000000ce000000e8000000ed000000ed000000ec",
            INIT_2B => X"000000f0000000f0000000f1000000e4000000a2000000850000008c00000095",
            INIT_2C => X"000000d1000000d5000000e3000000d9000000d3000000d3000000ca000000d4",
            INIT_2D => X"000000e5000000e1000000dd000000db000000dd000000e2000000de000000d5",
            INIT_2E => X"000000c2000000c8000000c6000000cc000000e7000000ed000000ec000000ea",
            INIT_2F => X"000000f0000000f1000000f0000000e6000000c300000097000000b2000000c5",
            INIT_30 => X"000000ae000000d0000000db000000e1000000d9000000d3000000ca000000cf",
            INIT_31 => X"0000008a00000081000000790000007200000070000000b8000000d5000000b4",
            INIT_32 => X"000000e2000000ea000000e9000000e8000000ec000000d8000000a700000098",
            INIT_33 => X"000000f1000000ef000000e6000000e3000000e6000000cb000000db000000e4",
            INIT_34 => X"000000c7000000c9000000b600000091000000830000007d0000007d00000082",
            INIT_35 => X"0000005400000049000000490000004600000047000000ac000000e6000000db",
            INIT_36 => X"000000d3000000e4000000e7000000ed000000ef000000e3000000a800000072",
            INIT_37 => X"000000e7000000dd000000c5000000ba000000ce000000db000000da000000d0",
            INIT_38 => X"000000c80000009d0000009b0000008d000000550000004f0000005600000051",
            INIT_39 => X"000000c000000097000000750000007000000079000000b4000000df000000e4",
            INIT_3A => X"0000008a0000009a000000a6000000ba000000cb000000db000000de000000d4",
            INIT_3B => X"000000d4000000c500000099000000890000008e000000920000008b00000085",
            INIT_3C => X"0000009e000000730000006b0000009700000090000000620000004600000035",
            INIT_3D => X"000000d2000000e4000000d1000000c2000000c1000000c2000000c2000000b4",
            INIT_3E => X"0000006f0000006a0000006f0000007d0000008800000096000000a5000000b5",
            INIT_3F => X"000000cb000000ce000000ae000000a400000097000000870000007900000076",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE8;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE9 : if BRAM_NAME = "sampleifmap_layer0_instance9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a2000000850000007b00000096000000d80000008c0000001d0000000f",
            INIT_01 => X"000000bd000000ee000000f1000000ea000000ea000000e0000000d1000000b5",
            INIT_02 => X"000000ab000000a5000000a5000000ab000000a30000009e0000009a0000009f",
            INIT_03 => X"000000af000000b7000000c4000000cf000000cc000000be000000b1000000ae",
            INIT_04 => X"000000e0000000d4000000cf000000cd000000e8000000cf0000003e00000005",
            INIT_05 => X"000000e4000000ee000000ee000000dd000000ee000000ee000000ec000000e6",
            INIT_06 => X"000000cc000000d4000000d6000000d4000000d5000000d8000000c8000000d9",
            INIT_07 => X"0000009a0000008f000000920000009c000000a5000000b5000000bf000000c1",
            INIT_08 => X"000000d0000000d3000000d3000000c5000000c4000000cc0000009b0000002d",
            INIT_09 => X"000000a9000000b0000000c6000000c1000000cf000000cf000000cb000000ce",
            INIT_0A => X"00000087000000960000009d0000008900000085000000a3000000ab000000a1",
            INIT_0B => X"0000008e0000008d000000850000007d00000074000000720000007000000073",
            INIT_0C => X"000000960000009600000098000000980000009a000000a0000000b300000087",
            INIT_0D => X"0000007a0000007e000000910000009500000095000000930000009300000096",
            INIT_0E => X"000000670000007000000075000000700000006d000000800000008600000078",
            INIT_0F => X"00000090000000850000007d00000079000000750000006f0000006700000061",
            INIT_10 => X"000000690000006600000066000000620000005d0000005a0000005a00000057",
            INIT_11 => X"00000085000000840000008800000089000000830000007c000000770000006f",
            INIT_12 => X"0000005c00000061000000650000006d000000770000007f0000008500000088",
            INIT_13 => X"000000950000008700000077000000680000006200000064000000640000005e",
            INIT_14 => X"0000001e00000019000000190000001a0000001a000000100000000b00000019",
            INIT_15 => X"0000004f0000004d0000004b000000450000003b000000330000002b00000024",
            INIT_16 => X"0000004500000045000000440000004300000048000000510000005800000057",
            INIT_17 => X"00000092000000880000007c0000007100000064000000590000004e00000047",
            INIT_18 => X"000000080000000b000000190000002d0000002c0000000d000000100000002e",
            INIT_19 => X"0000001700000013000000120000000d00000004000000020000000200000004",
            INIT_1A => X"0000003a000000320000002c000000260000001f00000021000000260000001d",
            INIT_1B => X"000000a00000008b0000007b000000730000007b000000730000005a00000046",
            INIT_1C => X"0000001f00000032000000460000005100000029000000130000001b00000029",
            INIT_1D => X"000000240000003200000040000000110000000000000002000000050000000f",
            INIT_1E => X"0000006100000047000000370000002b000000230000001e0000001e0000001e",
            INIT_1F => X"000000b300000098000000860000006f0000006900000078000000830000007c",
            INIT_20 => X"000000210000002b000000340000002c0000000c0000000a0000000a0000000f",
            INIT_21 => X"000000800000009e000000750000000800000001000000020000000400000012",
            INIT_22 => X"0000007e0000007e000000730000006b00000069000000670000006900000070",
            INIT_23 => X"000000c2000000ac0000009300000082000000740000005e000000560000006a",
            INIT_24 => X"0000000a0000000c0000000c0000000600000004000000030000000a00000028",
            INIT_25 => X"00000082000000800000003a0000000000000002000000010000000100000006",
            INIT_26 => X"000000420000004b000000600000006e00000071000000770000007b0000007f",
            INIT_27 => X"000000c5000000b6000000a20000008d00000084000000760000005d00000047",
            INIT_28 => X"0000000200000003000000020000000100000001000000010000001d0000004d",
            INIT_29 => X"0000002f0000002d0000000c0000000100000000000000000000000000000001",
            INIT_2A => X"0000004d00000030000000260000002a0000003100000032000000300000002e",
            INIT_2B => X"000000c6000000bb000000b00000009900000087000000800000007e0000006e",
            INIT_2C => X"000000000000000100000001000000000000000100000001000000340000005e",
            INIT_2D => X"0000002000000019000000030000000200000000000000000000000000000000",
            INIT_2E => X"000000710000005c00000042000000290000001d000000190000001900000019",
            INIT_2F => X"000000c9000000bf000000b30000009d0000008b0000007f0000007e0000007c",
            INIT_30 => X"0000000200000003000000030000000200000002000000070000003c00000066",
            INIT_31 => X"0000001f00000013000000010000000300000001000000000000000000000001",
            INIT_32 => X"0000007c0000007e000000730000005a0000003a0000001b0000000d00000011",
            INIT_33 => X"000000ca000000c0000000b00000009f0000009100000087000000820000007b",
            INIT_34 => X"000000070000000a0000000b0000000a0000000c000000170000003300000063",
            INIT_35 => X"000000150000000d000000050000000600000003000000040000000400000004",
            INIT_36 => X"0000007d0000007e0000007e00000071000000620000004d000000320000001b",
            INIT_37 => X"000000ca000000c5000000b8000000a80000009a000000940000008a00000080",
            INIT_38 => X"000000170000001a0000001c0000001e000000230000002c0000003900000060",
            INIT_39 => X"00000037000000280000001f0000001b00000017000000160000001500000015",
            INIT_3A => X"0000007f0000007a0000007a0000007900000070000000660000005800000046",
            INIT_3B => X"000000ca000000c8000000bd000000ac000000a0000000950000008b00000085",
            INIT_3C => X"000000370000003500000035000000380000003d000000430000004b00000065",
            INIT_3D => X"000000600000005400000047000000430000003e0000003a0000003800000037",
            INIT_3E => X"000000830000007d0000007c0000007f00000079000000740000006d00000067",
            INIT_3F => X"000000c8000000c3000000b7000000ab000000a2000000980000009100000088",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE9;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE10 : if BRAM_NAME = "sampleifmap_layer0_instance10" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000e8000000e8000000e8000000e8000000e8000000e8000000e7000000eb",
            INIT_01 => X"000000e9000000e9000000e9000000e9000000e9000000e9000000e8000000e8",
            INIT_02 => X"000000e6000000e8000000ea000000ea000000e8000000e9000000e9000000e9",
            INIT_03 => X"000000e8000000e9000000e9000000e8000000e8000000e8000000e9000000e7",
            INIT_04 => X"000000eb000000eb000000eb000000eb000000eb000000eb000000eb000000ee",
            INIT_05 => X"000000ec000000ec000000ec000000ec000000ec000000ec000000eb000000eb",
            INIT_06 => X"000000eb000000ed000000ee000000ed000000ea000000ea000000e9000000e9",
            INIT_07 => X"000000eb000000ec000000ec000000eb000000eb000000eb000000ec000000ea",
            INIT_08 => X"000000ea000000ea000000ea000000ea000000ea000000ea000000ea000000ed",
            INIT_09 => X"000000ea000000eb000000ea000000ea000000ea000000ea000000ea000000ea",
            INIT_0A => X"000000ea000000eb000000ee000000e9000000ec000000ea000000e7000000e7",
            INIT_0B => X"000000ea000000eb000000eb000000ea000000ea000000ea000000ea000000ea",
            INIT_0C => X"000000eb000000eb000000eb000000eb000000eb000000eb000000eb000000ee",
            INIT_0D => X"000000ea000000eb000000ea000000ea000000ea000000ea000000ea000000ea",
            INIT_0E => X"000000e6000000d5000000db000000c5000000e7000000e8000000e7000000e6",
            INIT_0F => X"000000eb000000eb000000eb000000ea000000ea000000ea000000ea000000eb",
            INIT_10 => X"000000eb000000eb000000eb000000eb000000eb000000eb000000ea000000ed",
            INIT_11 => X"000000eb000000eb000000ea000000ea000000eb000000eb000000ea000000ea",
            INIT_12 => X"000000e8000000dd000000d0000000b3000000db000000e6000000ed000000ec",
            INIT_13 => X"000000ec000000ec000000ec000000ec000000eb000000eb000000eb000000ed",
            INIT_14 => X"000000eb000000eb000000eb000000eb000000eb000000eb000000eb000000ee",
            INIT_15 => X"000000e8000000ed000000ea000000ec000000ec000000ec000000eb000000ea",
            INIT_16 => X"000000e8000000dc000000ca000000bd000000c8000000cf000000d2000000da",
            INIT_17 => X"000000ed000000ed000000ed000000ec000000eb000000eb000000eb000000ed",
            INIT_18 => X"000000eb000000eb000000ec000000e9000000e6000000e7000000e4000000e5",
            INIT_19 => X"000000e4000000ee000000e5000000e6000000ee000000ed000000ec000000ec",
            INIT_1A => X"000000d3000000b1000000ab000000b1000000be000000bf000000be000000cc",
            INIT_1B => X"000000ee000000ed000000ed000000ec000000eb000000e9000000ea000000ef",
            INIT_1C => X"000000ec000000eb000000ec000000ea000000ea000000ee000000e9000000de",
            INIT_1D => X"000000da000000eb000000dd000000cb000000ef000000ed000000ee000000ee",
            INIT_1E => X"000000cc000000b9000000bb000000c4000000cb000000d3000000d2000000d2",
            INIT_1F => X"000000ee000000ee000000ee000000ee000000ee000000ed000000ee000000f0",
            INIT_20 => X"000000eb000000eb000000ed000000f0000000f3000000f6000000f3000000f1",
            INIT_21 => X"000000e5000000e7000000da000000c4000000ef000000ed000000ed000000ed",
            INIT_22 => X"000000f1000000f0000000eb000000ea000000e3000000eb000000de000000d9",
            INIT_23 => X"000000ee000000ef000000ef000000ef000000f0000000f0000000f0000000f3",
            INIT_24 => X"000000e8000000e9000000e9000000bf000000a1000000990000009400000095",
            INIT_25 => X"000000ec000000e8000000e2000000d6000000eb000000ec000000eb000000ea",
            INIT_26 => X"000000d3000000e2000000f3000000f7000000ef000000f1000000eb000000e8",
            INIT_27 => X"000000ef000000ef000000ef000000eb000000c9000000b9000000ba000000c3",
            INIT_28 => X"000000e0000000e1000000e7000000a50000008900000089000000850000008d",
            INIT_29 => X"000000ec000000ee000000ec000000eb000000eb000000ea000000ea000000e9",
            INIT_2A => X"000000a3000000ac000000bf000000d5000000ee000000f1000000f0000000ee",
            INIT_2B => X"000000ef000000ee000000ef000000e5000000a60000008f000000990000009f",
            INIT_2C => X"000000ce000000d3000000e7000000e3000000df000000e0000000d7000000e0",
            INIT_2D => X"000000e9000000e6000000e1000000df000000db000000e1000000de000000d6",
            INIT_2E => X"000000ca000000cf000000cb000000d0000000ed000000f1000000ef000000ed",
            INIT_2F => X"000000ef000000ef000000ee000000e9000000ca000000a4000000c4000000d3",
            INIT_30 => X"000000ae000000d0000000e3000000f1000000ea000000e0000000d9000000de",
            INIT_31 => X"000000930000008b000000840000007e00000079000000bc000000d6000000b7",
            INIT_32 => X"000000e9000000f0000000ee000000eb000000ed000000dc000000ae000000a1",
            INIT_33 => X"000000f2000000f2000000e9000000ea000000ed000000d4000000e5000000ed",
            INIT_34 => X"000000cc000000cd000000c1000000a5000000970000008d0000009300000098",
            INIT_35 => X"000000620000005a0000005b0000005b0000005c000000b7000000ea000000e2",
            INIT_36 => X"000000d9000000e9000000ed000000f1000000f1000000e9000000b300000081",
            INIT_37 => X"000000ea000000e3000000cd000000c4000000d6000000df000000dc000000d4",
            INIT_38 => X"000000cf000000a4000000a40000009b0000006600000064000000720000006c",
            INIT_39 => X"000000cf000000a800000087000000830000008a000000be000000e4000000ea",
            INIT_3A => X"00000093000000a3000000ae000000c3000000d4000000e3000000e8000000df",
            INIT_3B => X"000000d8000000cb000000a0000000930000009700000098000000900000008c",
            INIT_3C => X"000000a1000000760000006e0000009c00000099000000740000005e0000004d",
            INIT_3D => X"000000d9000000ec000000d9000000ca000000c8000000c6000000c5000000b6",
            INIT_3E => X"0000007b000000760000007b0000008a000000950000009f000000ac000000ba",
            INIT_3F => X"000000d0000000d5000000b8000000ae000000a1000000910000008200000080",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE10;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE11 : if BRAM_NAME = "sampleifmap_layer0_instance11" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a2000000860000007b00000096000000dc000000970000002f00000023",
            INIT_01 => X"000000be000000ee000000f0000000e8000000e9000000e1000000d3000000b4",
            INIT_02 => X"000000bb000000b6000000b6000000bb000000b1000000aa000000a2000000a3",
            INIT_03 => X"000000b7000000c1000000d0000000da000000d9000000cc000000bf000000bd",
            INIT_04 => X"000000e5000000da000000d3000000d4000000ef000000d90000004f00000018",
            INIT_05 => X"000000ea000000f1000000ef000000dc000000ef000000f5000000f6000000ed",
            INIT_06 => X"000000e0000000e8000000ea000000e7000000e5000000e6000000d6000000e4",
            INIT_07 => X"000000a50000009e000000a1000000a9000000b3000000c5000000d1000000d4",
            INIT_08 => X"000000e3000000e6000000e5000000d9000000d8000000de000000b300000047",
            INIT_09 => X"000000bc000000c1000000d7000000cf000000dd000000e4000000e4000000e3",
            INIT_0A => X"0000009e000000ad000000b4000000a10000009c000000ba000000c3000000b8",
            INIT_0B => X"0000009c0000009e000000970000008c0000008300000085000000870000008a",
            INIT_0C => X"000000c1000000c0000000be000000bb000000bd000000c2000000cf000000a1",
            INIT_0D => X"0000009a000000a3000000ba000000bc000000bd000000bd000000be000000c0",
            INIT_0E => X"0000008800000090000000990000009400000091000000a3000000aa0000009a",
            INIT_0F => X"0000009c0000009400000092000000900000008d0000008b0000008600000082",
            INIT_10 => X"00000096000000930000008e000000860000007f0000007a000000710000006d",
            INIT_11 => X"000000af000000b4000000ba000000b5000000ac000000a5000000a000000098",
            INIT_12 => X"0000007f000000840000008b000000940000009b000000a3000000a8000000ac",
            INIT_13 => X"0000009c000000920000008a0000007e0000007a000000810000008500000081",
            INIT_14 => X"0000003d0000003a000000380000003400000030000000230000001900000029",
            INIT_15 => X"0000007e0000007e000000790000006a000000570000004d000000460000003e",
            INIT_16 => X"0000006600000067000000680000006a00000070000000780000007e0000007f",
            INIT_17 => X"000000950000008d000000880000008000000077000000730000006e00000069",
            INIT_18 => X"000000180000001e000000290000003a00000035000000130000001400000037",
            INIT_19 => X"0000003e0000003c000000380000002a000000140000000f0000000f00000011",
            INIT_1A => X"0000005a000000530000004f0000004e0000004c0000004d0000005100000047",
            INIT_1B => X"0000009e00000089000000800000007d0000008a0000008a0000007600000065",
            INIT_1C => X"00000025000000390000004c0000005400000029000000120000001a0000002d",
            INIT_1D => X"0000003e0000004e0000005b0000002300000007000000070000000b00000015",
            INIT_1E => X"0000007b00000063000000530000004a000000450000003f0000003e0000003c",
            INIT_1F => X"000000af00000092000000850000007400000072000000870000009500000092",
            INIT_20 => X"000000230000002f000000390000002e0000000b000000080000000900000011",
            INIT_21 => X"00000094000000b3000000860000000f00000003000000040000000700000014",
            INIT_22 => X"0000008d00000090000000850000007e0000007f0000007c0000007d00000083",
            INIT_23 => X"000000be000000a5000000900000008100000074000000610000005b00000074",
            INIT_24 => X"0000000c00000011000000110000000700000004000000030000000700000023",
            INIT_25 => X"0000009400000092000000400000000200000003000000020000000300000007",
            INIT_26 => X"00000045000000530000006a0000007a00000081000000890000008d00000090",
            INIT_27 => X"000000c2000000b00000009e000000870000007e000000710000005800000046",
            INIT_28 => X"0000000500000009000000050000000000000002000000010000001500000040",
            INIT_29 => X"000000440000003b0000000b0000000100000001000000000000000000000002",
            INIT_2A => X"000000470000002e0000002a000000310000003b000000430000004500000043",
            INIT_2B => X"000000c4000000b7000000ab0000009300000080000000780000007400000066",
            INIT_2C => X"0000000200000005000000020000000000000002000000010000002b00000052",
            INIT_2D => X"0000003600000026000000020000000000000000000000000000000000000000",
            INIT_2E => X"0000006900000052000000380000002700000022000000240000002b0000002e",
            INIT_2F => X"000000c7000000bb000000ae0000009600000083000000760000007300000073",
            INIT_30 => X"000000020000000300000001000000000000000100000003000000320000005d",
            INIT_31 => X"0000002f0000001c000000000000000200000001000000000000000000000001",
            INIT_32 => X"000000700000006f000000630000005100000037000000160000000c00000017",
            INIT_33 => X"000000c9000000bc000000ab00000097000000890000007e0000007700000071",
            INIT_34 => X"00000002000000040000000400000002000000040000000b0000002500000059",
            INIT_35 => X"000000180000000d000000020000000600000002000000010000000100000001",
            INIT_36 => X"0000006f000000700000007100000065000000520000003e0000002900000019",
            INIT_37 => X"000000c9000000c1000000b3000000a100000091000000890000007e00000073",
            INIT_38 => X"0000000c0000000d0000000f0000000f00000011000000160000002400000052",
            INIT_39 => X"0000002d0000001b00000015000000140000000f0000000e0000000d0000000c",
            INIT_3A => X"000000700000006b0000006e0000006900000058000000550000005100000043",
            INIT_3B => X"000000c8000000c4000000b7000000a4000000970000008a0000007f00000077",
            INIT_3C => X"0000002600000022000000210000002300000025000000260000003000000053",
            INIT_3D => X"0000004a0000003b000000300000002d0000002e0000002c0000002900000028",
            INIT_3E => X"000000750000006c0000006a0000006b00000061000000610000005c00000053",
            INIT_3F => X"000000c7000000bf000000b2000000a3000000990000008d000000850000007b",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE11;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE12 : if BRAM_NAME = "sampleifmap_layer0_instance12" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000c1000000bb000000b6000000a6000000840000008b0000009e0000009e",
            INIT_01 => X"000000e6000000e3000000df000000da000000ce000000d1000000cd000000c7",
            INIT_02 => X"000000ea000000ea000000e8000000ec000000eb000000e7000000e2000000d5",
            INIT_03 => X"000000ee000000ed000000e4000000e8000000ee000000e6000000e2000000ec",
            INIT_04 => X"000000c7000000c5000000c1000000ae0000008900000097000000ac000000aa",
            INIT_05 => X"000000ed000000e9000000e7000000e1000000d2000000d9000000d7000000ce",
            INIT_06 => X"000000f2000000ec000000ea000000f5000000f2000000e8000000e4000000db",
            INIT_07 => X"000000f6000000f6000000e8000000e9000000f3000000eb000000e4000000f1",
            INIT_08 => X"000000c7000000ce000000c9000000b50000008e0000009d000000b0000000ae",
            INIT_09 => X"000000ef000000e6000000e6000000e0000000d4000000da000000df000000d1",
            INIT_0A => X"000000f3000000ec000000d5000000e8000000ef000000e9000000e4000000dd",
            INIT_0B => X"000000f5000000fa000000e6000000ed000000f8000000ee000000e7000000f5",
            INIT_0C => X"000000cf000000d4000000cb000000ba00000093000000a0000000b2000000b4",
            INIT_0D => X"000000f0000000df000000e7000000dc000000d6000000dd000000e4000000d6",
            INIT_0E => X"000000f3000000e6000000ac000000b1000000e4000000e9000000e4000000e0",
            INIT_0F => X"000000f4000000f9000000e4000000ee000000fa000000ee000000e8000000f8",
            INIT_10 => X"000000cf000000d9000000cc000000bd00000093000000a5000000b9000000ba",
            INIT_11 => X"000000eb000000d3000000e7000000da000000d6000000de000000e7000000d3",
            INIT_12 => X"000000ed000000e0000000a80000009f000000d4000000e8000000e0000000e2",
            INIT_13 => X"000000f2000000f8000000ea000000e8000000f6000000eb000000e7000000f7",
            INIT_14 => X"000000d3000000db000000cb000000bf0000008e000000aa000000be000000c1",
            INIT_15 => X"000000cd000000c7000000e4000000d6000000d6000000dd000000ea000000d7",
            INIT_16 => X"000000e6000000de0000009e00000070000000c1000000eb000000ce000000cf",
            INIT_17 => X"000000eb000000f3000000e7000000e4000000f1000000e2000000e5000000f5",
            INIT_18 => X"000000d9000000de000000ca000000bf00000085000000ac000000bf000000c4",
            INIT_19 => X"000000b0000000bc000000e3000000d7000000d6000000da000000eb000000df",
            INIT_1A => X"000000b7000000ac0000008900000078000000bb000000cd000000ba000000bb",
            INIT_1B => X"000000eb000000f0000000e1000000e2000000eb000000d8000000df000000db",
            INIT_1C => X"000000e0000000e0000000da000000cb0000008c000000ae000000c5000000cc",
            INIT_1D => X"000000cd000000c9000000dd000000dc000000dc000000dc000000ed000000e8",
            INIT_1E => X"0000003c000000410000003e0000004700000053000000640000008a000000ac",
            INIT_1F => X"000000ec000000ef000000d4000000da000000e4000000d1000000b600000068",
            INIT_20 => X"000000c5000000af000000ba000000b0000000890000009d000000aa000000af",
            INIT_21 => X"000000c1000000c1000000c9000000d4000000d2000000ce000000d4000000d1",
            INIT_22 => X"000000450000005e00000053000000540000005b00000059000000690000008e",
            INIT_23 => X"000000c3000000cf000000a3000000ae000000b7000000a2000000790000004e",
            INIT_24 => X"000000800000006f0000006b0000006900000068000000710000007300000072",
            INIT_25 => X"0000009600000097000000930000009d0000009b00000097000000920000008b",
            INIT_26 => X"0000005300000056000000560000005500000063000000630000006400000076",
            INIT_27 => X"0000007b000000840000006d00000076000000990000009a000000800000008b",
            INIT_28 => X"0000005a000000540000005a00000053000000440000004b0000004c00000042",
            INIT_29 => X"0000006c000000720000006b0000006a00000067000000660000006a0000005d",
            INIT_2A => X"000000720000005f0000004200000048000000550000005b0000005a0000005a",
            INIT_2B => X"0000005e0000005c000000670000007d000000c7000000930000006e00000080",
            INIT_2C => X"00000046000000550000006a0000006f0000004d0000004b0000004100000035",
            INIT_2D => X"000000610000006b000000730000006c0000005d0000005f000000710000005d",
            INIT_2E => X"000000bb00000095000000550000005a00000061000000620000005f00000062",
            INIT_2F => X"00000055000000570000005f0000009a000000cc0000007000000092000000b3",
            INIT_30 => X"000000550000004d00000064000000640000004a0000005e000000560000003a",
            INIT_31 => X"00000057000000620000006e000000690000006c0000007f0000008500000078",
            INIT_32 => X"000000c3000000aa000000700000005f0000005f000000570000005100000051",
            INIT_33 => X"0000004f0000005500000050000000b2000000ad0000007f000000c1000000d0",
            INIT_34 => X"000000500000004700000044000000520000004b00000057000000590000004a",
            INIT_35 => X"00000062000000690000006a000000650000006f000000760000006700000059",
            INIT_36 => X"000000b8000000b40000008e000000720000006d000000620000006200000060",
            INIT_37 => X"000000430000003c00000050000000aa00000084000000a0000000c0000000bf",
            INIT_38 => X"0000005600000046000000480000004f0000004e000000520000004f0000004d",
            INIT_39 => X"000000830000008700000088000000890000008500000081000000790000006d",
            INIT_3A => X"000000b5000000b3000000a30000009400000096000000920000009400000092",
            INIT_3B => X"0000003b00000037000000490000005a00000065000000aa000000b0000000b9",
            INIT_3C => X"0000008a00000084000000830000006d000000680000006a0000005e00000060",
            INIT_3D => X"000000940000009e0000009b0000009b0000009a0000009b0000009800000090",
            INIT_3E => X"000000a9000000920000008200000077000000920000009c0000009d00000096",
            INIT_3F => X"0000004800000056000000620000004500000069000000a7000000a8000000b1",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE12;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE13 : if BRAM_NAME = "sampleifmap_layer0_instance13" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000008f0000009000000087000000810000008300000073000000650000006a",
            INIT_01 => X"0000009000000097000000990000009a0000009a0000009a0000009600000092",
            INIT_02 => X"0000009f00000092000000750000005e0000007f0000008b0000008600000082",
            INIT_03 => X"000000690000009a000000c00000009000000084000000a2000000a3000000a7",
            INIT_04 => X"00000091000000810000005d0000005f0000006d000000760000006c0000005f",
            INIT_05 => X"0000007b0000007a0000007e0000008600000090000000960000009700000095",
            INIT_06 => X"0000009c000000a20000009300000083000000940000009b000000850000007a",
            INIT_07 => X"000000940000009d000000a40000009f0000009500000099000000970000009d",
            INIT_08 => X"0000008c0000007b0000006f0000005600000046000000490000005900000066",
            INIT_09 => X"0000008d000000850000007e000000780000007500000078000000810000008f",
            INIT_0A => X"000000a1000000a50000009d000000970000009f000000990000008e00000096",
            INIT_0B => X"000000950000007d0000007900000083000000900000009a0000009800000099",
            INIT_0C => X"0000007b000000820000008a000000800000006e000000470000003d00000056",
            INIT_0D => X"000000990000009c000000980000008f00000084000000760000006c00000076",
            INIT_0E => X"000000a4000000a00000009a000000990000009a000000910000008900000095",
            INIT_0F => X"00000084000000560000004b0000005c000000690000007d0000009000000098",
            INIT_10 => X"000000760000007b0000007400000073000000720000006b0000006700000068",
            INIT_11 => X"00000075000000850000008d0000008f000000900000008d0000008600000074",
            INIT_12 => X"00000091000000980000009a0000009700000096000000820000005900000062",
            INIT_13 => X"00000041000000490000004700000041000000500000005a0000006000000075",
            INIT_14 => X"0000007e0000007d00000077000000720000006f0000006f0000006b00000063",
            INIT_15 => X"0000003d0000005b0000008200000083000000810000007d0000007d00000075",
            INIT_16 => X"0000005f00000072000000820000008b00000094000000730000003800000039",
            INIT_17 => X"0000001b000000330000004b0000003c0000003a000000490000005300000056",
            INIT_18 => X"0000005b0000006600000075000000740000007200000074000000680000003e",
            INIT_19 => X"0000004c000000600000008200000085000000700000004e0000005100000054",
            INIT_1A => X"000000510000005300000058000000600000006c0000006b0000005600000053",
            INIT_1B => X"000000180000001e0000002e000000340000002d000000330000003d00000046",
            INIT_1C => X"0000003500000041000000680000006b000000690000006a0000006000000039",
            INIT_1D => X"000000620000007300000085000000870000006e00000044000000400000003b",
            INIT_1E => X"00000037000000460000005000000051000000500000004e0000004f00000058",
            INIT_1F => X"000000180000001b0000001e00000022000000290000002d000000310000002c",
            INIT_20 => X"000000490000004f0000006d0000006d00000069000000680000005a00000041",
            INIT_21 => X"000000410000004400000053000000620000006a000000620000005800000055",
            INIT_22 => X"0000002c00000029000000330000004800000052000000510000004a00000046",
            INIT_23 => X"000000190000001b0000001e000000200000002300000027000000370000003d",
            INIT_24 => X"0000005100000058000000630000006600000067000000690000005700000043",
            INIT_25 => X"00000046000000420000003f0000003a000000390000003b000000450000004c",
            INIT_26 => X"0000002c000000310000002f0000002e000000360000003e0000004400000048",
            INIT_27 => X"0000001e00000018000000190000001d0000001c0000001e0000002e00000038",
            INIT_28 => X"0000002c0000002d00000032000000370000003a000000410000003a00000036",
            INIT_29 => X"0000003a0000003e000000400000003e0000003a00000037000000330000002e",
            INIT_2A => X"000000260000002a000000300000003100000030000000250000002600000033",
            INIT_2B => X"0000001f0000001c000000190000001b0000001c0000001b0000002000000029",
            INIT_2C => X"0000002700000021000000200000001f0000001b0000001a0000001d0000001e",
            INIT_2D => X"0000002800000026000000280000002e00000033000000350000003400000031",
            INIT_2E => X"0000002500000024000000250000002900000037000000420000002c00000026",
            INIT_2F => X"00000017000000210000001e0000001c0000001b0000001a0000001b0000001f",
            INIT_30 => X"000000200000001f0000001e0000001c0000001c0000001b0000001f00000021",
            INIT_31 => X"0000002d0000002900000027000000220000001e0000001e0000002100000023",
            INIT_32 => X"0000002000000026000000230000001e0000003100000049000000340000002a",
            INIT_33 => X"0000000d0000001a000000260000001e0000001d0000001b0000001a0000001b",
            INIT_34 => X"0000001b0000001a00000019000000190000001a0000001a0000001e0000001f",
            INIT_35 => X"0000002a00000028000000290000002a0000002800000025000000200000001d",
            INIT_36 => X"0000001d0000001e000000240000001c00000026000000400000002e00000027",
            INIT_37 => X"000000040000000900000025000000210000001c0000001b000000190000001a",
            INIT_38 => X"0000002500000022000000200000001e0000001c000000190000001b00000017",
            INIT_39 => X"000000210000001e000000230000002600000027000000280000002700000027",
            INIT_3A => X"0000001d0000001d0000001d0000001e0000002400000039000000240000001c",
            INIT_3B => X"000000050000000400000013000000240000001b000000170000001800000018",
            INIT_3C => X"0000002500000023000000220000002100000022000000200000001e0000001c",
            INIT_3D => X"0000000c0000000f000000180000001e00000022000000240000002600000026",
            INIT_3E => X"0000001c0000001b0000001b00000019000000200000002d0000001300000008",
            INIT_3F => X"0000000700000004000000050000001900000022000000140000001500000018",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE13;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE14 : if BRAM_NAME = "sampleifmap_layer0_instance14" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d8000000d3000000d0000000c10000009e000000a6000000bb000000be",
            INIT_01 => X"000000ed000000eb000000e8000000e5000000da000000de000000dd000000db",
            INIT_02 => X"000000f1000000f1000000ef000000f1000000ef000000ee000000e9000000dc",
            INIT_03 => X"000000f1000000ef000000e7000000ed000000f3000000eb000000e7000000f2",
            INIT_04 => X"000000da000000da000000d9000000c7000000a0000000b0000000c7000000c8",
            INIT_05 => X"000000f3000000ef000000ee000000e9000000db000000e5000000e5000000df",
            INIT_06 => X"000000f5000000ef000000ed000000f7000000f5000000ee000000ea000000e1",
            INIT_07 => X"000000f7000000f6000000e8000000ec000000f8000000ef000000e9000000f5",
            INIT_08 => X"000000d6000000df000000dc000000c9000000a2000000b3000000c8000000c9",
            INIT_09 => X"000000f4000000ea000000ea000000e5000000db000000e2000000e9000000dd",
            INIT_0A => X"000000f1000000ea000000d6000000eb000000f3000000ee000000e9000000e2",
            INIT_0B => X"000000f4000000f9000000e5000000ee000000fa000000f0000000e9000000f7",
            INIT_0C => X"000000d9000000e1000000d9000000c9000000a4000000b3000000c7000000cb",
            INIT_0D => X"000000f4000000e2000000e8000000dd000000d9000000e3000000eb000000df",
            INIT_0E => X"000000f1000000e4000000af000000b8000000eb000000ed000000e7000000e4",
            INIT_0F => X"000000f2000000f7000000e3000000ed000000fa000000ee000000e8000000f8",
            INIT_10 => X"000000d5000000e1000000d6000000c9000000a1000000b5000000cc000000cf",
            INIT_11 => X"000000ec000000d4000000e5000000d9000000d7000000e2000000ed000000d7",
            INIT_12 => X"000000ec000000e0000000ae000000aa000000e1000000ec000000e1000000e3",
            INIT_13 => X"000000ef000000f5000000e7000000e7000000f6000000eb000000e7000000f7",
            INIT_14 => X"000000d7000000e2000000d4000000c90000009a000000b7000000cd000000d0",
            INIT_15 => X"000000cd000000c7000000e5000000d7000000d7000000df000000ee000000da",
            INIT_16 => X"000000e9000000e3000000a70000007c000000cc000000ef000000d0000000d1",
            INIT_17 => X"000000e8000000f1000000e6000000e2000000ef000000e1000000e5000000f6",
            INIT_18 => X"000000d5000000dd000000cb000000c20000008b000000b3000000c7000000cc",
            INIT_19 => X"000000b0000000bc000000e6000000d8000000d4000000d8000000e9000000db",
            INIT_1A => X"000000be000000b70000009700000081000000c0000000d4000000c0000000be",
            INIT_1B => X"000000e0000000eb000000de000000db000000e5000000d6000000e0000000e0",
            INIT_1C => X"000000cc000000ce000000cb000000c00000008a000000af000000c6000000cd",
            INIT_1D => X"000000ce000000c7000000d8000000d5000000d2000000d0000000df000000d4",
            INIT_1E => X"000000450000005000000050000000550000005d0000007100000095000000b2",
            INIT_1F => X"000000d4000000dd000000c5000000d0000000de000000ce000000b70000006c",
            INIT_20 => X"000000b3000000a0000000ac000000a5000000850000009a000000a8000000ad",
            INIT_21 => X"000000c6000000c1000000bf000000c7000000c3000000bd000000c2000000be",
            INIT_22 => X"0000004f0000006e00000068000000680000006c0000006b0000007900000098",
            INIT_23 => X"000000af000000be00000095000000a3000000af0000009f0000007a00000052",
            INIT_24 => X"0000007f000000700000006e0000006d00000069000000720000007400000073",
            INIT_25 => X"000000a10000009e0000008f00000097000000930000008c0000008800000087",
            INIT_26 => X"0000005c000000660000006c0000006c00000078000000780000007700000086",
            INIT_27 => X"00000078000000820000006a0000006e0000009100000097000000800000008f",
            INIT_28 => X"000000640000006100000069000000630000005200000056000000570000004e",
            INIT_29 => X"0000007f0000008400000076000000720000006f0000006a0000006d00000065",
            INIT_2A => X"000000770000006c00000057000000600000006b0000006e0000006d0000006d",
            INIT_2B => X"00000068000000660000006f00000078000000bf000000900000006f00000084",
            INIT_2C => X"00000051000000620000007a00000080000000620000005f000000550000004a",
            INIT_2D => X"0000007b000000860000008b0000008400000073000000710000008100000068",
            INIT_2E => X"000000bd0000009e000000680000007100000077000000740000007300000078",
            INIT_2F => X"00000063000000630000006700000095000000c50000006d00000094000000b7",
            INIT_30 => X"000000660000005d00000073000000750000005d000000710000006b00000051",
            INIT_31 => X"000000710000007d000000880000008200000083000000950000009800000089",
            INIT_32 => X"000000c2000000af0000007f000000760000007b000000720000006c0000006c",
            INIT_33 => X"000000650000006200000050000000a7000000a200000076000000bd000000ce",
            INIT_34 => X"000000640000005900000054000000620000005d0000006a0000006e00000061",
            INIT_35 => X"0000007c00000082000000830000007e000000860000008a0000007b0000006e",
            INIT_36 => X"000000b4000000b50000009900000086000000870000007e0000007f0000007b",
            INIT_37 => X"00000059000000480000004d000000a00000007a00000097000000b7000000b8",
            INIT_38 => X"0000006b00000058000000580000005f00000061000000660000006500000066",
            INIT_39 => X"0000009d000000a1000000a4000000a30000009e000000970000008e00000082",
            INIT_3A => X"000000ae000000b1000000a9000000a2000000a9000000aa000000ad000000ab",
            INIT_3B => X"0000004b0000003f000000460000005700000062000000a4000000a8000000b0",
            INIT_3C => X"000000a000000098000000940000007e0000007c0000007f000000760000007b",
            INIT_3D => X"000000ae000000b9000000b8000000b7000000b4000000b3000000af000000a7",
            INIT_3E => X"000000a10000008e0000008500000080000000a0000000af000000b2000000ad",
            INIT_3F => X"00000052000000590000005f000000460000006c000000a6000000a2000000a9",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE14;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE15 : if BRAM_NAME = "sampleifmap_layer0_instance15" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a7000000a60000009a00000094000000980000008a0000007d00000085",
            INIT_01 => X"000000ab000000b5000000b9000000b9000000b6000000b3000000ae000000aa",
            INIT_02 => X"0000009b0000009000000078000000660000008b0000009a0000009800000098",
            INIT_03 => X"0000006c00000099000000bb0000009100000088000000a3000000a2000000a5",
            INIT_04 => X"000000aa000000980000007200000074000000830000008d000000850000007c",
            INIT_05 => X"000000970000009a000000a0000000a7000000ad000000b0000000af000000af",
            INIT_06 => X"0000009e000000a5000000980000008c000000a0000000a80000009600000090",
            INIT_07 => X"00000093000000980000009e0000009e000000970000009c0000009b000000a3",
            INIT_08 => X"000000a400000094000000870000006e0000005d000000600000007100000081",
            INIT_09 => X"000000a50000009f000000990000009400000092000000960000009f000000a9",
            INIT_0A => X"000000a4000000a8000000a4000000a1000000ac000000a8000000a0000000aa",
            INIT_0B => X"000000960000007d0000007900000084000000920000009e0000009e000000a0",
            INIT_0C => X"000000930000009c000000a50000009b00000087000000600000005500000070",
            INIT_0D => X"000000ab000000ae000000ad000000a7000000a0000000970000008d0000008e",
            INIT_0E => X"000000a6000000a3000000a1000000a3000000a8000000a20000009b000000a7",
            INIT_0F => X"0000008a0000005c00000052000000620000006f00000082000000970000009e",
            INIT_10 => X"0000008e000000960000008f0000008f0000008f000000870000008400000085",
            INIT_11 => X"0000008600000097000000a5000000a9000000ab000000a9000000a10000008a",
            INIT_12 => X"000000980000009f000000a3000000a3000000a4000000940000006b00000074",
            INIT_13 => X"00000048000000500000004e0000004b0000005b000000660000006c00000080",
            INIT_14 => X"000000960000009700000093000000900000008f000000900000008c00000084",
            INIT_15 => X"0000004e0000006e0000009c0000009f0000009a00000094000000920000008b",
            INIT_16 => X"0000006d0000007e0000008f00000099000000a3000000840000004a0000004b",
            INIT_17 => X"0000002100000039000000520000004b0000004c0000005a0000006400000067",
            INIT_18 => X"000000730000008100000091000000920000009200000094000000890000005e",
            INIT_19 => X"0000005d000000720000009a0000009d0000008700000063000000660000006a",
            INIT_1A => X"00000065000000660000006a000000710000007c0000007d0000006800000065",
            INIT_1B => X"0000001f0000002500000035000000430000003f000000450000004f00000058",
            INIT_1C => X"0000004d0000005c000000850000008900000086000000860000007d00000056",
            INIT_1D => X"00000073000000840000009600000099000000830000005c0000005900000052",
            INIT_1E => X"0000004f0000005f00000065000000630000006100000060000000610000006a",
            INIT_1F => X"0000001f00000022000000260000002f000000390000003c000000400000003c",
            INIT_20 => X"000000610000006a0000008a000000890000008300000081000000740000005a",
            INIT_21 => X"00000053000000540000005f000000710000007e0000007c000000740000006c",
            INIT_22 => X"00000045000000430000004a0000005c00000064000000620000005c00000059",
            INIT_23 => X"0000002000000023000000260000002b0000002e00000033000000420000004a",
            INIT_24 => X"000000660000006e000000780000007c0000007f00000082000000700000005c",
            INIT_25 => X"0000005b00000054000000500000004b0000004c000000500000005a00000061",
            INIT_26 => X"0000003d0000004300000041000000410000004900000051000000590000005f",
            INIT_27 => X"0000002500000023000000280000002a000000280000002a0000003a00000045",
            INIT_28 => X"0000003f00000040000000450000004a0000004e000000560000004f0000004c",
            INIT_29 => X"000000500000005100000052000000510000004d0000004a0000004600000041",
            INIT_2A => X"00000032000000360000003f0000004300000044000000370000003b00000049",
            INIT_2B => X"0000002500000027000000280000002900000028000000280000002d00000036",
            INIT_2C => X"0000003a0000003500000034000000310000002a000000280000002b0000002d",
            INIT_2D => X"0000003b0000003a0000003b0000004100000046000000480000004700000044",
            INIT_2E => X"0000002f0000002f000000330000003900000049000000550000003f00000038",
            INIT_2F => X"0000001d0000002a0000002a000000290000002800000027000000280000002c",
            INIT_30 => X"0000003200000031000000300000002c0000002600000024000000280000002b",
            INIT_31 => X"0000003d0000003e0000003b0000003500000031000000310000003400000035",
            INIT_32 => X"000000280000002f0000002e0000002c000000420000005e0000004500000037",
            INIT_33 => X"00000012000000200000002e000000290000002a000000280000002700000027",
            INIT_34 => X"0000002b00000029000000290000002700000024000000230000002700000028",
            INIT_35 => X"000000370000003c0000003d0000003d0000003a00000038000000330000002e",
            INIT_36 => X"00000024000000250000002e0000002800000036000000550000003c0000002e",
            INIT_37 => X"000000070000000d000000280000002b0000002a000000280000002600000026",
            INIT_38 => X"00000033000000310000002f0000002c00000028000000240000002600000022",
            INIT_39 => X"0000002b000000330000003700000039000000390000003b0000003900000036",
            INIT_3A => X"00000023000000230000002500000029000000320000004e000000300000001f",
            INIT_3B => X"0000000700000006000000140000002d00000029000000240000002500000025",
            INIT_3C => X"000000310000003000000030000000300000002f0000002d0000002b00000029",
            INIT_3D => X"000000110000001a00000022000000280000002d000000310000003300000032",
            INIT_3E => X"000000230000002200000022000000210000002c0000003f0000001b00000008",
            INIT_3F => X"0000000800000005000000060000001f0000002c000000220000002200000023",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE15;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE16 : if BRAM_NAME = "sampleifmap_layer0_instance16" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000f1000000ee000000ec000000de000000ba000000c2000000da000000de",
            INIT_01 => X"000000f5000000f2000000f1000000f0000000eb000000f4000000f5000000f3",
            INIT_02 => X"000000f3000000f3000000f3000000f9000000f8000000f5000000f0000000e3",
            INIT_03 => X"000000f6000000f3000000ea000000f1000000f7000000ef000000eb000000f5",
            INIT_04 => X"000000ee000000f0000000f0000000df000000b8000000c9000000e2000000e5",
            INIT_05 => X"000000f8000000f5000000f5000000f3000000e8000000f5000000f7000000f3",
            INIT_06 => X"000000f4000000ee000000ee000000fb000000fb000000f3000000ef000000e6",
            INIT_07 => X"000000fb000000fa000000ec000000f0000000fc000000f3000000ec000000f8",
            INIT_08 => X"000000e4000000ef000000ee000000db000000b5000000c7000000de000000e1",
            INIT_09 => X"000000f7000000ee000000ef000000eb000000e4000000ec000000f4000000eb",
            INIT_0A => X"000000ef000000e8000000d7000000ec000000f6000000f1000000ec000000e5",
            INIT_0B => X"000000f7000000fb000000e8000000f1000000fc000000f2000000eb000000f8",
            INIT_0C => X"000000e1000000eb000000e4000000d6000000b3000000c2000000d8000000de",
            INIT_0D => X"000000f7000000e6000000ec000000e1000000dd000000e6000000ef000000e5",
            INIT_0E => X"000000f1000000e5000000b0000000ba000000ee000000f0000000ea000000e6",
            INIT_0F => X"000000f3000000f8000000e4000000ee000000fb000000ef000000e9000000f8",
            INIT_10 => X"000000d9000000e7000000dd000000d2000000ac000000c1000000d9000000df",
            INIT_11 => X"000000ee000000d6000000e8000000db000000d7000000e1000000eb000000da",
            INIT_12 => X"000000ef000000e5000000b2000000b0000000e4000000ee000000e3000000e5",
            INIT_13 => X"000000f0000000f6000000e8000000e7000000f5000000ea000000e7000000f7",
            INIT_14 => X"000000d5000000e1000000d5000000ce000000a4000000bf000000d5000000dc",
            INIT_15 => X"000000ce000000c8000000e3000000d6000000d6000000da000000e6000000d6",
            INIT_16 => X"000000e9000000e6000000ad00000082000000cf000000ed000000ce000000d0",
            INIT_17 => X"000000e6000000f2000000e7000000dd000000e8000000db000000e1000000f4",
            INIT_18 => X"000000d0000000d9000000c9000000c400000096000000b9000000ca000000d4",
            INIT_19 => X"000000af000000b9000000dd000000d4000000d3000000d0000000db000000d3",
            INIT_1A => X"000000bb000000b80000009d00000089000000c5000000d2000000bd000000bb",
            INIT_1B => X"000000d8000000e7000000db000000d1000000da000000ce000000dc000000dd",
            INIT_1C => X"000000cb000000ce000000cc000000c500000093000000b3000000c9000000d3",
            INIT_1D => X"000000cb000000c0000000ce000000ce000000cd000000c6000000d2000000d0",
            INIT_1E => X"00000049000000580000005e000000640000006a0000007a0000009b000000b3",
            INIT_1F => X"000000c1000000ce000000b9000000c6000000d7000000ca000000b70000006f",
            INIT_20 => X"000000b3000000a1000000af000000aa0000008c000000a0000000ad000000b3",
            INIT_21 => X"000000c4000000ba000000b9000000c3000000bd000000b4000000b8000000bb",
            INIT_22 => X"0000005a000000800000007e0000007e0000008000000080000000890000009f",
            INIT_23 => X"0000009f000000b0000000890000009c000000ac0000009e0000007c00000058",
            INIT_24 => X"00000080000000720000007200000072000000700000007b0000007e0000007b",
            INIT_25 => X"000000a7000000a0000000920000009800000090000000890000008600000086",
            INIT_26 => X"000000680000007800000083000000820000008c000000900000008b00000093",
            INIT_27 => X"0000007500000080000000690000006a0000008d000000960000008300000095",
            INIT_28 => X"0000006a00000068000000730000006b00000058000000620000006600000059",
            INIT_29 => X"0000009200000097000000860000007b0000007300000071000000760000006b",
            INIT_2A => X"000000800000007a000000680000006f000000780000007f0000007f00000080",
            INIT_2B => X"000000700000006d0000007500000072000000b60000008b0000006e00000086",
            INIT_2C => X"0000005e00000071000000890000008e0000006a0000006e0000006800000058",
            INIT_2D => X"00000097000000a5000000a5000000940000007d0000007f0000009200000074",
            INIT_2E => X"000000bf000000a5000000720000007b0000007f0000007f000000820000008e",
            INIT_2F => X"0000006c0000006c0000006d0000008c000000b8000000640000008e000000b4",
            INIT_30 => X"000000760000006d000000820000008100000068000000840000008200000064",
            INIT_31 => X"0000008b0000009a000000a50000009b00000097000000a8000000ab0000009a",
            INIT_32 => X"000000c1000000b300000089000000860000008c000000810000007d00000082",
            INIT_33 => X"0000006d0000006900000054000000a00000009800000070000000b9000000cb",
            INIT_34 => X"000000790000006c00000065000000710000006a0000007e0000008600000078",
            INIT_35 => X"000000950000009e000000a1000000990000009f000000a10000009100000083",
            INIT_36 => X"000000b1000000b6000000a1000000960000009b000000910000009300000092",
            INIT_37 => X"000000600000004e000000500000009d0000007600000094000000b5000000b5",
            INIT_38 => X"00000086000000730000007100000074000000720000007d000000800000007f",
            INIT_39 => X"000000b9000000be000000bf000000be000000b8000000b0000000a80000009f",
            INIT_3A => X"000000a8000000af000000ad000000ac000000b8000000be000000c4000000c5",
            INIT_3B => X"0000005100000043000000470000005700000063000000a3000000a5000000ab",
            INIT_3C => X"000000c1000000b8000000b300000099000000910000009a0000009500000097",
            INIT_3D => X"000000c8000000d4000000d2000000d1000000d0000000cf000000cd000000c9",
            INIT_3E => X"0000009b0000008b0000008700000086000000ab000000c3000000c9000000c6",
            INIT_3F => X"000000560000005a0000005c0000004900000071000000a8000000a1000000a5",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE16;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE17 : if BRAM_NAME = "sampleifmap_layer0_instance17" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000c9000000c6000000b9000000af000000b0000000a70000009f000000a5",
            INIT_01 => X"000000be000000c9000000d0000000d2000000d2000000d2000000d0000000cd",
            INIT_02 => X"000000990000008e0000007a0000006c00000094000000a9000000aa000000aa",
            INIT_03 => X"0000006f00000098000000b5000000930000008e000000a7000000a5000000a7",
            INIT_04 => X"000000ca000000b60000008f0000008d0000009d000000ae000000aa0000009d",
            INIT_05 => X"000000a2000000a7000000b5000000bf000000ca000000d1000000d3000000d0",
            INIT_06 => X"000000a0000000a70000009d00000093000000a9000000b2000000a00000009b",
            INIT_07 => X"0000009400000096000000960000009e0000009c000000a1000000a2000000a9",
            INIT_08 => X"000000c2000000b1000000a40000008a000000790000008000000094000000a2",
            INIT_09 => X"000000b0000000ac000000ac000000aa000000ab000000b2000000bc000000c7",
            INIT_0A => X"000000ac000000af000000ad000000aa000000b5000000b0000000a8000000b4",
            INIT_0B => X"000000990000007d000000760000008500000096000000a3000000a5000000a8",
            INIT_0C => X"000000b0000000ba000000c5000000bc000000a60000007f000000750000008f",
            INIT_0D => X"000000ba000000bf000000be000000b9000000b2000000ab000000a3000000a9",
            INIT_0E => X"000000b2000000af000000ac000000ad000000b1000000ac000000a5000000b4",
            INIT_0F => X"0000009000000062000000570000006700000074000000880000009c000000a4",
            INIT_10 => X"000000aa000000b3000000ae000000b0000000b0000000a8000000a5000000a6",
            INIT_11 => X"00000096000000a8000000b5000000b9000000bd000000be000000b8000000a4",
            INIT_12 => X"000000a2000000ab000000ad000000ad000000ad0000009d0000007600000081",
            INIT_13 => X"0000004e0000005600000054000000500000005f0000006a0000007000000085",
            INIT_14 => X"000000b0000000b3000000b0000000ae000000af000000b1000000ac000000a5",
            INIT_15 => X"0000005e0000007e000000ab000000af000000ad000000ab000000ab000000a4",
            INIT_16 => X"000000750000008800000098000000a2000000ac0000008e0000005500000058",
            INIT_17 => X"000000270000003f000000580000004f000000500000005e000000680000006c",
            INIT_18 => X"0000008b0000009a000000ad000000af000000af000000b2000000a60000007c",
            INIT_19 => X"0000006c00000083000000a9000000ae0000009a0000007a0000007e00000082",
            INIT_1A => X"0000006c0000006d000000710000007900000085000000860000007200000072",
            INIT_1B => X"000000260000002b0000003b00000049000000450000004b000000560000005f",
            INIT_1C => X"00000064000000740000009e000000a30000009f000000a0000000960000006f",
            INIT_1D => X"0000008300000095000000a8000000ac00000097000000730000007000000068",
            INIT_1E => X"00000054000000640000006c0000006a0000006a0000006a0000006b00000077",
            INIT_1F => X"00000025000000280000002c0000003700000041000000440000004900000045",
            INIT_20 => X"0000007700000080000000a2000000a10000009a000000970000008a00000071",
            INIT_21 => X"0000006200000065000000720000008400000092000000900000008800000081",
            INIT_22 => X"0000004b0000004800000050000000630000006c0000006d0000006700000065",
            INIT_23 => X"00000027000000290000002d000000340000003a0000003d0000004d00000055",
            INIT_24 => X"0000007c000000840000008f00000094000000970000009a0000008800000074",
            INIT_25 => X"00000065000000630000005b00000056000000570000005b0000006700000076",
            INIT_26 => X"000000450000004a0000004800000048000000520000005e0000006300000065",
            INIT_27 => X"000000300000002f00000030000000330000003200000034000000440000004e",
            INIT_28 => X"0000005100000052000000560000005c000000630000006a0000006400000060",
            INIT_29 => X"000000580000005e0000005b0000005700000054000000510000004f00000052",
            INIT_2A => X"0000003b00000040000000480000004a0000004c00000044000000440000004d",
            INIT_2B => X"000000300000003400000030000000310000003200000031000000360000003f",
            INIT_2C => X"000000440000003e0000003d0000003c0000003700000036000000390000003b",
            INIT_2D => X"000000420000004500000044000000480000004d0000004f0000004f0000004e",
            INIT_2E => X"00000039000000380000003c000000410000005200000061000000470000003d",
            INIT_2F => X"0000002300000032000000320000003200000031000000300000003100000035",
            INIT_30 => X"000000370000003500000035000000310000002d0000002c0000003000000032",
            INIT_31 => X"0000004400000047000000420000003c00000038000000380000003b0000003a",
            INIT_32 => X"000000330000003a00000038000000350000004b000000680000004b0000003b",
            INIT_33 => X"0000001400000025000000350000003200000033000000310000003000000031",
            INIT_34 => X"000000300000002e0000002e0000002c00000029000000280000002c0000002d",
            INIT_35 => X"0000003d000000440000004400000044000000410000003f0000003900000033",
            INIT_36 => X"0000002f0000003000000038000000310000003f0000005d0000004200000032",
            INIT_37 => X"000000050000000e0000002e0000003400000033000000310000002f0000002f",
            INIT_38 => X"0000003b0000003800000036000000320000002d000000290000002b00000027",
            INIT_39 => X"000000310000003a0000003d000000400000004000000042000000400000003e",
            INIT_3A => X"0000002f0000002f00000030000000320000003b000000550000003500000024",
            INIT_3B => X"00000003000000030000001800000036000000320000002d0000002e0000002e",
            INIT_3C => X"0000003a0000003800000038000000380000003600000034000000320000002f",
            INIT_3D => X"000000140000001e000000270000002d0000003200000035000000370000003a",
            INIT_3E => X"0000002e0000002d0000002d0000002c0000003600000048000000210000000b",
            INIT_3F => X"00000007000000030000000800000025000000340000002b0000002c0000002c",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE17;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE18 : if BRAM_NAME = "sampleifmap_layer0_instance18" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a6000000a8000000a6000000b1000000be000000b0000000a70000009b",
            INIT_01 => X"000000b8000000b8000000bb000000bb000000bb000000bb000000b3000000aa",
            INIT_02 => X"000000bd000000bc000000bb000000bb000000ba000000b8000000b4000000b6",
            INIT_03 => X"000000c0000000ca000000c9000000c9000000c3000000bc000000bb000000bb",
            INIT_04 => X"0000009f0000009a0000009b000000b3000000bb000000ab000000a300000099",
            INIT_05 => X"000000a5000000a2000000ab000000a9000000af000000ab000000a50000009f",
            INIT_06 => X"000000a8000000a9000000ad000000a7000000a5000000a6000000a4000000aa",
            INIT_07 => X"000000bd000000cb000000ca000000cc000000ca000000be000000ad000000a9",
            INIT_08 => X"000000bc000000b0000000ae000000bb000000b8000000a8000000a00000009b",
            INIT_09 => X"000000b9000000bc000000c2000000c0000000be000000b1000000b3000000b6",
            INIT_0A => X"000000bf000000c1000000c5000000c3000000c2000000c1000000c2000000c1",
            INIT_0B => X"000000bd000000cc000000ce000000d0000000cf000000ce000000c5000000bf",
            INIT_0C => X"000000c5000000c7000000b9000000b4000000b1000000a60000009d00000097",
            INIT_0D => X"000000cb000000c4000000c5000000d2000000c6000000cd000000cc000000b6",
            INIT_0E => X"000000cc000000c5000000d2000000cf000000cb000000d2000000cf000000cd",
            INIT_0F => X"000000c0000000ce000000cf000000d1000000c9000000cc000000c6000000d0",
            INIT_10 => X"000000c4000000bf000000b5000000b1000000ae000000a80000009e00000097",
            INIT_11 => X"000000ca000000b9000000b9000000c4000000b9000000bd000000c2000000b7",
            INIT_12 => X"000000bc000000be000000c7000000c3000000c0000000c8000000c7000000c7",
            INIT_13 => X"000000c4000000cf000000cc000000ce000000c4000000c9000000c7000000c9",
            INIT_14 => X"000000c3000000c4000000ae000000ab000000ae000000a70000009c00000094",
            INIT_15 => X"000000bf000000bd000000bd000000bb000000b8000000bd000000be000000c0",
            INIT_16 => X"000000c1000000c0000000bc000000c0000000c6000000bb000000c3000000be",
            INIT_17 => X"000000c4000000d1000000d0000000d4000000d1000000cb000000ce000000cd",
            INIT_18 => X"000000c3000000cb000000b0000000a8000000ae000000a50000009900000094",
            INIT_19 => X"000000c3000000c5000000c2000000b6000000be000000bb000000bc000000bc",
            INIT_1A => X"000000c9000000c5000000c5000000c6000000cd000000c8000000c1000000c4",
            INIT_1B => X"000000c3000000cf000000cb000000c5000000c3000000c6000000c8000000c5",
            INIT_1C => X"000000d1000000c7000000bc000000ac000000ac000000a30000009b00000099",
            INIT_1D => X"000000c4000000bb000000bc000000c1000000bf000000bd000000be000000c4",
            INIT_1E => X"000000c8000000c4000000c9000000c2000000ce000000c4000000c2000000ca",
            INIT_1F => X"000000bd000000c7000000c4000000c8000000c9000000c8000000bb000000b5",
            INIT_20 => X"000000be000000b0000000b0000000ae000000ac000000a30000009f000000a0",
            INIT_21 => X"000000b6000000ac000000aa000000b5000000b0000000b0000000af000000b4",
            INIT_22 => X"000000bb000000b4000000bc000000b1000000bb000000b5000000b2000000bb",
            INIT_23 => X"000000b8000000c2000000c0000000c5000000bc000000bc000000c4000000c7",
            INIT_24 => X"000000b0000000b4000000ab000000aa000000ac000000a2000000a7000000ab",
            INIT_25 => X"0000009e0000009900000092000000960000009c000000960000009c0000009b",
            INIT_26 => X"000000a60000009c000000a20000009d0000009d000000a4000000a6000000a6",
            INIT_27 => X"000000b6000000c2000000c1000000c5000000bd000000bc000000c7000000c8",
            INIT_28 => X"000000ae000000b6000000b1000000ad000000b0000000a8000000b4000000af",
            INIT_29 => X"000000ad000000a8000000a30000009f0000009a0000009f000000a00000009c",
            INIT_2A => X"000000ac000000a7000000a8000000a0000000a2000000a0000000a4000000aa",
            INIT_2B => X"000000b7000000c1000000bf000000c5000000c4000000c4000000c3000000c2",
            INIT_2C => X"000000b6000000ae000000aa000000b7000000bb000000b2000000bb000000b5",
            INIT_2D => X"000000c1000000c1000000bb000000b8000000b5000000b4000000b3000000b3",
            INIT_2E => X"000000c0000000c0000000ba000000b8000000b9000000bc000000c0000000c1",
            INIT_2F => X"000000ba000000c4000000bf000000be000000bd000000c0000000bc000000bb",
            INIT_30 => X"000000c1000000950000008400000099000000ab000000ba000000be000000b9",
            INIT_31 => X"000000c4000000c3000000c1000000bf000000bc000000ba000000bf000000c6",
            INIT_32 => X"000000bf000000c0000000be000000bc000000bc000000be000000c0000000c3",
            INIT_33 => X"000000c1000000cc000000ca000000ca000000c5000000c3000000c1000000bf",
            INIT_34 => X"0000006d0000005e00000074000000840000009e000000bc000000c2000000ba",
            INIT_35 => X"000000c7000000c4000000c1000000bf000000c2000000c2000000b100000091",
            INIT_36 => X"000000c6000000c7000000c4000000c4000000c6000000c8000000c7000000c7",
            INIT_37 => X"000000b9000000c6000000c5000000c6000000c4000000c4000000c4000000c5",
            INIT_38 => X"0000005c0000008d000000b8000000c2000000c6000000c4000000c5000000ba",
            INIT_39 => X"000000cc000000cc000000c9000000c3000000b30000008e0000006800000054",
            INIT_3A => X"000000bf000000c2000000c2000000c2000000c7000000cc000000cc000000cc",
            INIT_3B => X"000000b5000000c0000000be000000bf000000be000000be000000be000000bd",
            INIT_3C => X"000000b1000000c9000000c8000000c5000000c8000000c6000000c7000000b8",
            INIT_3D => X"000000cd000000d0000000ca000000ad000000800000005d0000005400000075",
            INIT_3E => X"000000c3000000c5000000c4000000c3000000c7000000c7000000c8000000ca",
            INIT_3F => X"000000b2000000be000000bd000000bf000000bf000000c2000000c3000000c1",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE18;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE19 : if BRAM_NAME = "sampleifmap_layer0_instance19" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d6000000d0000000ce000000cd000000d0000000cb000000c9000000b9",
            INIT_01 => X"000000cb000000b50000008c000000690000005b0000004c0000005c000000af",
            INIT_02 => X"000000c2000000c2000000c2000000c1000000c2000000c5000000ca000000ce",
            INIT_03 => X"000000b4000000be000000be000000c1000000bf000000c1000000c3000000c2",
            INIT_04 => X"000000d0000000d3000000d4000000d4000000d6000000cf000000cc000000bb",
            INIT_05 => X"0000008400000063000000540000005400000057000000470000007c000000cb",
            INIT_06 => X"000000c4000000c5000000c0000000c3000000cb000000cb000000be000000a7",
            INIT_07 => X"000000b7000000c0000000bf000000c1000000bf000000c0000000c2000000c2",
            INIT_08 => X"000000d0000000d3000000d3000000d4000000d6000000cf000000cf000000be",
            INIT_09 => X"00000053000000560000005400000053000000570000004800000089000000d3",
            INIT_0A => X"000000cc000000cb000000b6000000a30000009b000000830000006b00000059",
            INIT_0B => X"000000b6000000bf000000c0000000c1000000bf000000c2000000c6000000ca",
            INIT_0C => X"000000d5000000d4000000d4000000d5000000d7000000d1000000d2000000bf",
            INIT_0D => X"0000005d000000570000004c0000003f0000003a0000002f00000071000000cc",
            INIT_0E => X"0000009f0000007a0000004d0000003a0000003e00000046000000500000005a",
            INIT_0F => X"000000b9000000c4000000c4000000c8000000c8000000c9000000c2000000b4",
            INIT_10 => X"000000d4000000d1000000d2000000d1000000d3000000cf000000d0000000bf",
            INIT_11 => X"000000580000004a00000044000000330000002500000041000000650000009d",
            INIT_12 => X"000000480000003e0000002e000000370000004900000055000000560000005b",
            INIT_13 => X"000000ba000000c4000000c3000000b80000009e000000850000006b0000004e",
            INIT_14 => X"000000c8000000d1000000ce000000cf000000d1000000cb000000ca000000ba",
            INIT_15 => X"0000006000000032000000350000002d00000064000000970000008c00000095",
            INIT_16 => X"000000420000005900000070000000620000004800000080000000a00000009c",
            INIT_17 => X"000000b2000000bc000000b7000000ad000000a3000000a60000008300000043",
            INIT_18 => X"000000d1000000d1000000d0000000d2000000d2000000ca000000c9000000b9",
            INIT_19 => X"000000a8000000940000009200000090000000bd000000d7000000d3000000d2",
            INIT_1A => X"0000009f000000b1000000b2000000a30000009a000000c0000000ce000000ca",
            INIT_1B => X"000000b0000000bc000000c1000000c4000000c2000000bf000000b20000009c",
            INIT_1C => X"000000b7000000b9000000bc000000c0000000c4000000c0000000bc000000b0",
            INIT_1D => X"000000ad000000ab000000aa000000aa000000ad000000b3000000b2000000b6",
            INIT_1E => X"000000aa000000a5000000a1000000a5000000a7000000a1000000a0000000a9",
            INIT_1F => X"0000009c000000a4000000a30000009d0000009600000098000000a0000000aa",
            INIT_20 => X"0000005d0000005e00000061000000660000006b0000006e0000006300000072",
            INIT_21 => X"00000065000000530000004e0000004d00000050000000580000005500000058",
            INIT_22 => X"000000710000006f0000006e0000006c0000006b0000006a0000006c00000071",
            INIT_23 => X"0000007c0000007a000000790000007800000077000000780000007700000075",
            INIT_24 => X"0000007100000072000000700000007300000075000000710000006d0000007a",
            INIT_25 => X"0000006c0000006e0000006d0000006e0000006d0000006f000000700000006f",
            INIT_26 => X"00000068000000650000006a0000006c0000006b000000690000007000000073",
            INIT_27 => X"000000650000005e00000066000000670000006d0000006d0000006b0000006a",
            INIT_28 => X"0000005e00000062000000680000006d000000700000006b0000006100000078",
            INIT_29 => X"0000004e000000500000004f0000005200000056000000580000005d0000005e",
            INIT_2A => X"0000004100000041000000420000004300000045000000480000004f00000050",
            INIT_2B => X"0000004d000000350000003f0000004300000040000000420000004100000040",
            INIT_2C => X"0000003d0000003f00000042000000420000004500000041000000370000005b",
            INIT_2D => X"0000003f0000003d0000003c00000039000000390000003c0000004000000042",
            INIT_2E => X"0000003c0000003b00000039000000380000003a00000040000000420000003f",
            INIT_2F => X"0000005c0000004b00000031000000340000003900000038000000390000003a",
            INIT_30 => X"0000004100000040000000430000004300000044000000420000003c0000005d",
            INIT_31 => X"0000003d0000003c0000003b0000003b0000003b0000003e0000004100000045",
            INIT_32 => X"00000038000000380000003700000037000000380000003a0000003f00000040",
            INIT_33 => X"00000051000000610000005d0000004100000035000000380000003a00000039",
            INIT_34 => X"0000003b000000390000003b00000039000000390000003d0000003900000059",
            INIT_35 => X"0000003d0000003b0000003d0000003c00000036000000380000003a0000003c",
            INIT_36 => X"0000003d0000003d0000003c0000003c000000390000003a0000003d00000041",
            INIT_37 => X"000000430000003b000000590000006100000046000000390000003e00000042",
            INIT_38 => X"0000003f0000003e0000003e0000003e0000003e0000003f0000003c00000059",
            INIT_39 => X"000000510000004e000000510000005400000052000000410000003d0000003e",
            INIT_3A => X"0000004000000042000000430000005000000053000000550000005400000058",
            INIT_3B => X"0000004b0000003d000000390000004c00000067000000560000003800000034",
            INIT_3C => X"0000004100000043000000420000003f0000003c0000003d0000003c0000005c",
            INIT_3D => X"0000004600000048000000490000004900000048000000410000004300000042",
            INIT_3E => X"0000003e00000040000000400000004b0000004b0000004b0000004a00000049",
            INIT_3F => X"00000049000000400000003c0000003900000040000000580000005600000041",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE19;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE20 : if BRAM_NAME = "sampleifmap_layer0_instance20" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ad000000ad000000ab000000b9000000c0000000b3000000b00000009c",
            INIT_01 => X"000000b5000000b6000000b8000000b9000000b8000000b6000000b3000000af",
            INIT_02 => X"000000bd000000bb000000ba000000ba000000b9000000b7000000b3000000b3",
            INIT_03 => X"000000b7000000ca000000c4000000c5000000c3000000bc000000bb000000bb",
            INIT_04 => X"000000a40000009f000000a2000000be000000c3000000b8000000b30000009b",
            INIT_05 => X"000000a7000000a4000000ae000000ab000000b0000000a9000000a5000000a3",
            INIT_06 => X"000000a9000000ab000000af000000a9000000a6000000a8000000a6000000ac",
            INIT_07 => X"000000be000000d7000000d0000000ce000000cc000000bf000000ae000000aa",
            INIT_08 => X"000000a8000000b2000000c1000000cb000000c4000000b9000000b20000009a",
            INIT_09 => X"000000bc000000be000000c5000000c3000000c4000000be000000af000000a0",
            INIT_0A => X"000000bf000000c1000000c6000000c4000000c3000000c2000000c3000000c4",
            INIT_0B => X"000000bf000000d7000000d0000000ce000000cd000000cd000000c4000000c0",
            INIT_0C => X"00000080000000bc000000c5000000ca000000c3000000bc000000b20000009a",
            INIT_0D => X"0000009400000095000000950000009e0000009b0000009a000000980000006c",
            INIT_0E => X"0000009f000000ae000000a3000000a8000000ad000000a3000000a1000000a7",
            INIT_0F => X"000000bc000000d4000000cd000000cc000000ce000000cc000000d0000000bc",
            INIT_10 => X"0000007e000000bd000000c4000000c6000000bf000000bb000000b10000009a",
            INIT_11 => X"000000710000007600000078000000730000006b0000006a0000008b00000080",
            INIT_12 => X"000000700000008800000070000000760000007e000000720000007200000077",
            INIT_13 => X"000000be000000d6000000cd000000ce000000ce000000c9000000cb000000a0",
            INIT_14 => X"00000093000000b7000000c8000000c5000000bd000000bb000000ae00000097",
            INIT_15 => X"0000009d0000009500000092000000aa000000a500000091000000a8000000a9",
            INIT_16 => X"000000b1000000bc000000b3000000b0000000bd000000b0000000b2000000b4",
            INIT_17 => X"000000be000000d8000000d1000000d0000000d0000000cf000000d0000000c4",
            INIT_18 => X"0000006000000093000000c6000000c2000000bd000000b9000000ac00000098",
            INIT_19 => X"0000008b00000080000000790000009800000098000000900000009700000095",
            INIT_1A => X"000000a400000096000000ad00000096000000a2000000aa000000970000009c",
            INIT_1B => X"000000bc000000d4000000cf000000d3000000d2000000cc000000a60000009c",
            INIT_1C => X"0000006500000077000000b5000000c2000000bb000000b6000000ac0000009b",
            INIT_1D => X"0000007f0000008700000087000000920000007800000083000000830000007b",
            INIT_1E => X"0000009f0000007b000000840000006d0000007b000000830000007b0000007b",
            INIT_1F => X"000000ba000000d0000000c9000000c9000000c7000000bf000000840000007b",
            INIT_20 => X"000000af000000ab000000ba000000c0000000b9000000b4000000af000000a1",
            INIT_21 => X"000000aa000000ad000000ac000000af000000a6000000ac000000a5000000a2",
            INIT_22 => X"000000be000000b2000000ac000000a3000000af000000b2000000b2000000ac",
            INIT_23 => X"000000b9000000d1000000c9000000c8000000cd000000c8000000b0000000ac",
            INIT_24 => X"000000b7000000c2000000c0000000be000000ba000000b4000000b7000000ac",
            INIT_25 => X"000000a2000000a40000009e0000009f000000a3000000a2000000a5000000a0",
            INIT_26 => X"000000b6000000a5000000a3000000a0000000a2000000ac000000ae000000a7",
            INIT_27 => X"000000b8000000d0000000ca000000ca000000cd000000ca000000c6000000c8",
            INIT_28 => X"000000b7000000c1000000c1000000c0000000be000000ba000000c4000000b1",
            INIT_29 => X"000000ac000000aa000000a6000000a40000009f000000a5000000a7000000a3",
            INIT_2A => X"000000b2000000ab000000ad000000a8000000ab000000a6000000a6000000a8",
            INIT_2B => X"000000b8000000d0000000c8000000c8000000c7000000c7000000c6000000c7",
            INIT_2C => X"000000c6000000be000000bb000000c9000000c8000000c3000000cc000000b7",
            INIT_2D => X"000000c6000000c6000000c2000000c1000000c1000000c1000000c1000000c2",
            INIT_2E => X"000000c5000000c4000000c4000000c5000000c6000000c3000000c3000000c6",
            INIT_2F => X"000000bb000000d1000000c8000000ca000000c9000000c9000000cb000000c9",
            INIT_30 => X"000000c40000009a0000008d000000a6000000b2000000c6000000cd000000b9",
            INIT_31 => X"000000ca000000c9000000c7000000c5000000c5000000c7000000ca000000ca",
            INIT_32 => X"000000c6000000c7000000c6000000c4000000c4000000c6000000c7000000c9",
            INIT_33 => X"000000bd000000d4000000ce000000cf000000ce000000cb000000ca000000c7",
            INIT_34 => X"0000006b0000005f0000007c00000090000000a5000000c8000000d0000000ba",
            INIT_35 => X"000000cc000000c9000000c6000000c5000000c7000000c7000000b30000008f",
            INIT_36 => X"000000cd000000cd000000c9000000c9000000cc000000ce000000cd000000cc",
            INIT_37 => X"000000b7000000cf000000ca000000ca000000cb000000cb000000cb000000cc",
            INIT_38 => X"0000005b0000008f000000c1000000ce000000cc000000d0000000d4000000ba",
            INIT_39 => X"000000cf000000cf000000cc000000c6000000b50000008e0000006500000051",
            INIT_3A => X"000000c5000000c6000000c5000000c5000000ca000000cf000000cf000000cf",
            INIT_3B => X"000000b5000000cc000000c5000000c4000000c5000000c5000000c5000000c5",
            INIT_3C => X"000000b3000000cf000000d4000000d1000000ce000000d2000000d6000000b8",
            INIT_3D => X"000000ce000000d2000000cb000000ae000000800000005d0000005300000074",
            INIT_3E => X"000000c9000000c9000000c7000000c6000000c9000000ca000000ca000000cc",
            INIT_3F => X"000000b4000000cb000000c6000000c6000000c7000000c9000000ca000000c8",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE20;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE21 : if BRAM_NAME = "sampleifmap_layer0_instance21" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d9000000d4000000d6000000d6000000d5000000d6000000d7000000ba",
            INIT_01 => X"000000cc000000b50000008a0000006500000056000000490000005b000000af",
            INIT_02 => X"000000c8000000c9000000c9000000c7000000c6000000c7000000cb000000d0",
            INIT_03 => X"000000b6000000cc000000c8000000ca000000c9000000c9000000ca000000c8",
            INIT_04 => X"000000d3000000d6000000d9000000db000000d9000000d8000000d8000000bb",
            INIT_05 => X"0000008200000061000000510000004f00000052000000440000007b000000cc",
            INIT_06 => X"000000c6000000c7000000c1000000c4000000ca000000c9000000bc000000a5",
            INIT_07 => X"000000b6000000cc000000c7000000c9000000c8000000c8000000c7000000c6",
            INIT_08 => X"000000d2000000d6000000d8000000d8000000d6000000d5000000d9000000bc",
            INIT_09 => X"0000004d00000050000000500000004e000000530000004600000088000000d4",
            INIT_0A => X"000000cc000000c9000000b20000009f000000970000007e0000006600000053",
            INIT_0B => X"000000b4000000c9000000c5000000c7000000c6000000c8000000c9000000cb",
            INIT_0C => X"000000d8000000d7000000d8000000d7000000d5000000d6000000da000000bb",
            INIT_0D => X"000000510000004d000000450000003a000000370000002d00000070000000cc",
            INIT_0E => X"000000a00000007c0000004f0000003b0000003e000000460000004d00000050",
            INIT_0F => X"000000b4000000ca000000c8000000cb000000cd000000cd000000c4000000b5",
            INIT_10 => X"000000d4000000d4000000d6000000d3000000d1000000d2000000d8000000bc",
            INIT_11 => X"0000004d000000410000003e00000030000000210000003a0000005f0000009a",
            INIT_12 => X"000000480000003f0000002f0000003800000048000000540000005400000052",
            INIT_13 => X"000000b6000000ca000000c1000000b50000009e000000840000006b0000004e",
            INIT_14 => X"000000c8000000d4000000d3000000d1000000cf000000ce000000d2000000b8",
            INIT_15 => X"0000005a0000002e000000320000002d000000610000008f0000008500000091",
            INIT_16 => X"00000041000000580000007000000061000000470000007f0000009e00000096",
            INIT_17 => X"000000b0000000c5000000b5000000a8000000a2000000a50000008200000043",
            INIT_18 => X"000000d2000000d5000000d4000000d3000000d0000000cd000000d2000000b7",
            INIT_19 => X"000000a6000000930000009300000094000000bf000000d4000000d1000000d1",
            INIT_1A => X"000000a2000000b4000000b5000000a60000009d000000c3000000d0000000c8",
            INIT_1B => X"000000b1000000c7000000c1000000c3000000c5000000c1000000b40000009f",
            INIT_1C => X"000000b9000000bb000000be000000c2000000c2000000c3000000c4000000ae",
            INIT_1D => X"000000ad000000ae000000b0000000b2000000b5000000b7000000b5000000b8",
            INIT_1E => X"000000b0000000aa000000a6000000aa000000ac000000a6000000a4000000aa",
            INIT_1F => X"0000009e000000af000000a30000009d0000009b0000009d000000a5000000af",
            INIT_20 => X"0000006000000061000000640000006700000069000000700000006c00000070",
            INIT_21 => X"00000067000000570000005300000054000000570000005e0000005a0000005c",
            INIT_22 => X"00000076000000740000007300000071000000700000006f0000007000000073",
            INIT_23 => X"0000007c000000840000007a000000790000007b0000007c0000007b0000007a",
            INIT_24 => X"00000071000000710000006f0000007100000070000000710000007300000075",
            INIT_25 => X"0000006b0000006e0000006d0000006e0000006e0000006f000000700000006f",
            INIT_26 => X"0000006b000000680000006d0000006f0000006e0000006c0000007300000073",
            INIT_27 => X"00000065000000620000005f0000006400000070000000700000006e0000006d",
            INIT_28 => X"0000005d00000061000000660000006a0000006a000000690000006600000071",
            INIT_29 => X"0000004e0000004f0000004e0000005200000055000000590000005e0000005f",
            INIT_2A => X"0000004100000041000000410000004300000044000000470000004f00000050",
            INIT_2B => X"0000006400000047000000370000003c00000041000000420000004200000041",
            INIT_2C => X"0000003c0000003e000000400000004000000040000000410000003c00000054",
            INIT_2D => X"0000003f0000003d0000003c00000039000000380000003d0000004000000042",
            INIT_2E => X"0000003c0000003b0000003a000000380000003b000000410000004300000040",
            INIT_2F => X"000000800000007500000048000000380000003800000038000000390000003a",
            INIT_30 => X"0000003f0000003d000000410000003f0000003e0000003f0000003b00000053",
            INIT_31 => X"0000003d0000003c0000003a0000003a000000390000003c0000003e00000043",
            INIT_32 => X"0000003d0000003e0000003c0000003d0000003e000000400000004400000041",
            INIT_33 => X"0000006300000089000000880000005b000000410000003d0000003a0000003a",
            INIT_34 => X"0000003c0000003a0000003b00000037000000390000003d000000350000004f",
            INIT_35 => X"0000003f0000003d0000003e0000003c00000037000000390000003c0000003d",
            INIT_36 => X"0000003f000000400000003e0000003e0000003b0000003c0000003f00000043",
            INIT_37 => X"0000004a0000004f000000770000008e0000006e000000470000003c0000003e",
            INIT_38 => X"0000003e0000003e0000003e0000003f00000041000000420000003a00000052",
            INIT_39 => X"0000004d0000004a0000004c0000004f0000004f000000410000003e0000003f",
            INIT_3A => X"000000410000003e0000003f0000004c0000004e000000500000005000000054",
            INIT_3B => X"000000450000004000000042000000660000008d0000007c0000005600000042",
            INIT_3C => X"000000390000003b0000003a0000003a0000003a0000003a000000340000004e",
            INIT_3D => X"00000045000000460000004700000047000000450000003a0000003b0000003a",
            INIT_3E => X"000000440000003f0000003f000000490000004a000000490000004800000048",
            INIT_3F => X"00000044000000410000003f000000420000005800000080000000800000005a",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE21;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE22 : if BRAM_NAME = "sampleifmap_layer0_instance22" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b4000000b5000000b7000000ca000000cd000000c1000000bb00000095",
            INIT_01 => X"000000bd000000bd000000c0000000c0000000c0000000c1000000bd000000b6",
            INIT_02 => X"000000be000000c0000000c1000000c1000000c0000000bd000000b9000000ba",
            INIT_03 => X"000000ab000000d4000000d1000000ca000000c3000000bc000000bb000000bb",
            INIT_04 => X"000000b3000000b3000000be000000e0000000e3000000d7000000cc0000009d",
            INIT_05 => X"000000b7000000b4000000be000000bb000000c3000000c3000000bb000000b3",
            INIT_06 => X"000000bc000000bc000000bf000000b9000000b7000000b8000000b7000000bc",
            INIT_07 => X"000000b7000000e3000000de000000df000000e0000000d3000000c2000000be",
            INIT_08 => X"000000b8000000c4000000d5000000df000000db000000d5000000c900000099",
            INIT_09 => X"000000ca000000cc000000d2000000d0000000d4000000d3000000c3000000b1",
            INIT_0A => X"000000d0000000d0000000d4000000d2000000d1000000d0000000d1000000d1",
            INIT_0B => X"000000b8000000e0000000d7000000da000000df000000de000000d5000000d0",
            INIT_0C => X"00000083000000c9000000dc000000e2000000de000000d3000000cf000000a6",
            INIT_0D => X"000000ab000000a6000000a7000000b2000000b1000000a60000009e00000077",
            INIT_0E => X"000000a5000000b4000000ba000000b9000000ba000000b2000000b2000000b7",
            INIT_0F => X"000000ba000000e6000000df000000e0000000dd000000dc000000e4000000cf",
            INIT_10 => X"0000008e000000d6000000e1000000e0000000da000000ca000000cb000000a7",
            INIT_11 => X"000000830000007c0000007e0000008100000081000000780000009800000099",
            INIT_12 => X"0000007b0000008d00000088000000880000008a000000820000008400000086",
            INIT_13 => X"000000b9000000e3000000dc000000de000000d9000000da000000e3000000ba",
            INIT_14 => X"000000a5000000d1000000da000000dc000000d9000000cb000000c9000000a4",
            INIT_15 => X"000000ac000000a3000000a0000000b3000000b40000009c000000b5000000c4",
            INIT_16 => X"000000be000000c6000000c0000000bf000000c9000000be000000c1000000bf",
            INIT_17 => X"000000bc000000e8000000e1000000df000000e1000000e1000000e1000000d4",
            INIT_18 => X"00000068000000ac000000d6000000d9000000d9000000c8000000c6000000a4",
            INIT_19 => X"000000a00000009700000090000000a5000000af000000a6000000a50000009e",
            INIT_1A => X"000000b9000000ad000000b7000000aa000000b6000000bd000000ad000000b2",
            INIT_1B => X"000000bc000000e7000000e0000000dd000000e2000000dc000000b2000000a6",
            INIT_1C => X"0000006f00000092000000cb000000da000000d8000000c7000000c9000000a9",
            INIT_1D => X"000000900000008f0000008f0000009b000000900000009d0000009500000086",
            INIT_1E => X"000000b00000008e0000008d0000007f0000008e000000940000008e00000093",
            INIT_1F => X"000000ba000000e4000000dc000000d9000000dc000000d10000009500000089",
            INIT_20 => X"000000c5000000c1000000cd000000db000000d9000000c7000000ce000000b1",
            INIT_21 => X"000000bd000000bb000000ba000000c0000000b8000000bb000000b7000000b8",
            INIT_22 => X"000000c8000000bc000000ba000000b2000000bf000000c2000000c2000000c0",
            INIT_23 => X"000000b9000000e4000000dd000000db000000db000000d6000000c6000000c1",
            INIT_24 => X"000000d2000000dc000000d6000000d7000000d6000000c5000000d4000000ba",
            INIT_25 => X"000000ba000000b9000000b4000000b6000000ba000000b6000000bb000000b9",
            INIT_26 => X"000000c6000000b6000000b6000000b5000000b8000000c3000000c6000000c1",
            INIT_27 => X"000000b7000000e3000000de000000df000000df000000dd000000de000000de",
            INIT_28 => X"000000cc000000d6000000d4000000d7000000d8000000c8000000de000000bc",
            INIT_29 => X"000000bf000000bc000000b8000000b5000000b0000000b6000000b8000000b5",
            INIT_2A => X"000000c9000000ba000000b8000000b6000000b9000000b8000000ba000000bd",
            INIT_2B => X"000000b8000000e3000000dc000000db000000db000000dc000000dd000000df",
            INIT_2C => X"000000de000000d7000000d1000000dc000000e0000000cf000000e2000000bf",
            INIT_2D => X"000000df000000df000000db000000d9000000d7000000d6000000d7000000d9",
            INIT_2E => X"000000db000000d9000000d6000000d8000000da000000db000000dd000000df",
            INIT_2F => X"000000ba000000e3000000db000000d7000000d6000000d9000000db000000db",
            INIT_30 => X"000000d9000000ac00000099000000b5000000ce000000d4000000dc000000bc",
            INIT_31 => X"000000e2000000e1000000df000000de000000dc000000dd000000e1000000e2",
            INIT_32 => X"000000da000000dc000000db000000d9000000da000000dc000000dd000000e1",
            INIT_33 => X"000000bb000000e6000000e0000000e0000000e0000000de000000dc000000d9",
            INIT_34 => X"00000073000000630000007e0000009d000000c1000000d6000000df000000bd",
            INIT_35 => X"000000e2000000df000000dc000000da000000dd000000dd000000c60000009d",
            INIT_36 => X"000000e0000000e0000000dd000000dc000000df000000e1000000e0000000e2",
            INIT_37 => X"000000b7000000e2000000dd000000dd000000de000000de000000de000000df",
            INIT_38 => X"0000005a00000092000000c4000000dc000000e9000000de000000e2000000bd",
            INIT_39 => X"000000e4000000e3000000e0000000da000000ca000000a10000007100000054",
            INIT_3A => X"000000d9000000d8000000d7000000d7000000dc000000e0000000e1000000e2",
            INIT_3B => X"000000b6000000e1000000da000000d7000000d8000000d8000000d8000000d8",
            INIT_3C => X"000000b3000000da000000e1000000e1000000ea000000e0000000e5000000bb",
            INIT_3D => X"000000e1000000e4000000dd000000c0000000910000006a0000005800000073",
            INIT_3E => X"000000db000000d9000000d6000000d6000000d9000000da000000db000000df",
            INIT_3F => X"000000b7000000e2000000dc000000d9000000da000000dc000000dd000000db",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE22;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE23 : if BRAM_NAME = "sampleifmap_layer0_instance23" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000e1000000e0000000e2000000e4000000e9000000de000000e9000000be",
            INIT_01 => X"000000d9000000c0000000920000006a0000005b0000005000000062000000b5",
            INIT_02 => X"000000d9000000da000000da000000d9000000da000000dd000000e1000000e0",
            INIT_03 => X"000000bc000000e3000000dc000000dd000000dd000000dd000000dd000000da",
            INIT_04 => X"000000dd000000e2000000e3000000e7000000e9000000dd000000ea000000bf",
            INIT_05 => X"0000008800000064000000500000004b0000004f0000004900000082000000d5",
            INIT_06 => X"000000de000000df000000d9000000d9000000dc000000d7000000c8000000ad",
            INIT_07 => X"000000bd000000e3000000db000000da000000db000000db000000dd000000dd",
            INIT_08 => X"000000dc000000e2000000e1000000e3000000e4000000d9000000e8000000bd",
            INIT_09 => X"0000004c0000004e0000004c0000004a000000500000004a00000090000000dd",
            INIT_0A => X"000000e2000000e1000000c9000000b0000000a1000000810000006400000053",
            INIT_0B => X"000000bb000000e1000000d9000000d7000000d7000000d9000000dc000000df",
            INIT_0C => X"000000e2000000e3000000e1000000e0000000e1000000d7000000e8000000bb",
            INIT_0D => X"000000520000004d000000450000003b000000380000003200000077000000d5",
            INIT_0E => X"000000a2000000850000005b000000410000003f000000420000004800000050",
            INIT_0F => X"000000bc000000e3000000dd000000dd000000df000000da000000cc000000b8",
            INIT_10 => X"000000e1000000e4000000e6000000df000000df000000de000000e7000000b7",
            INIT_11 => X"0000004e000000440000004300000035000000270000003c00000062000000a2",
            INIT_12 => X"000000430000003f000000310000003900000048000000530000005200000051",
            INIT_13 => X"000000c3000000df000000d7000000c6000000a80000008b0000006d0000004b",
            INIT_14 => X"000000d4000000e2000000e2000000de000000de000000e2000000e2000000b0",
            INIT_15 => X"0000005e0000003300000039000000350000006a000000960000008b0000009b",
            INIT_16 => X"000000430000005a00000072000000630000004900000082000000a10000009a",
            INIT_17 => X"000000be000000d0000000c5000000b7000000a9000000ab0000008600000045",
            INIT_18 => X"000000de000000de000000de000000df000000df000000e1000000e1000000af",
            INIT_19 => X"000000b3000000a00000009f0000009f000000cc000000e4000000e0000000de",
            INIT_1A => X"000000ad000000c0000000c1000000b2000000a9000000cf000000dc000000d6",
            INIT_1B => X"000000bd000000d2000000d1000000d8000000d6000000d2000000c3000000ab",
            INIT_1C => X"000000c7000000c9000000cc000000ce000000d1000000d7000000d4000000a6",
            INIT_1D => X"000000c4000000c2000000c1000000c0000000c2000000c5000000c3000000c7",
            INIT_1E => X"000000cd000000c8000000c4000000c8000000ca000000c4000000c2000000c4",
            INIT_1F => X"000000b5000000c9000000c5000000c5000000bf000000c0000000c5000000ce",
            INIT_20 => X"0000006a0000006b000000700000007600000078000000820000007800000065",
            INIT_21 => X"000000800000006c000000650000006200000063000000660000006200000065",
            INIT_22 => X"0000009e00000098000000960000009400000093000000920000009200000090",
            INIT_23 => X"00000092000000a7000000a5000000a8000000a8000000a8000000a6000000a4",
            INIT_24 => X"0000008800000089000000880000008a0000008600000086000000820000006f",
            INIT_25 => X"0000008300000083000000800000007f0000007e000000830000008600000084",
            INIT_26 => X"0000007e0000007c0000008000000081000000810000007f000000860000008a",
            INIT_27 => X"0000006000000073000000730000007700000084000000840000008200000081",
            INIT_28 => X"000000640000006c000000760000007a00000078000000780000007100000068",
            INIT_29 => X"0000005600000057000000550000005800000059000000550000005b00000060",
            INIT_2A => X"0000003c0000003f000000410000004200000043000000460000004f00000056",
            INIT_2B => X"0000004b0000003f00000032000000360000003b0000003c0000003c0000003b",
            INIT_2C => X"000000360000003b0000003f0000003a000000390000003d000000370000003d",
            INIT_2D => X"000000320000003100000032000000300000002f0000002f0000003300000038",
            INIT_2E => X"00000037000000320000002e0000002d0000002f000000350000003700000033",
            INIT_2F => X"00000068000000680000003a0000003000000034000000340000003400000036",
            INIT_30 => X"00000039000000370000003d0000003e0000003c000000410000003d00000044",
            INIT_31 => X"0000003600000038000000380000003b0000003a00000037000000380000003d",
            INIT_32 => X"0000003400000034000000330000003300000034000000370000003b00000039",
            INIT_33 => X"0000004b00000078000000710000004b00000039000000370000003500000033",
            INIT_34 => X"00000036000000340000003900000039000000350000003b000000340000003e",
            INIT_35 => X"0000003500000034000000380000003900000032000000300000003200000036",
            INIT_36 => X"0000003000000035000000370000003600000033000000340000003600000039",
            INIT_37 => X"000000320000003e000000650000007c0000005f0000003d0000003400000032",
            INIT_38 => X"0000003c0000003c0000003d0000003b000000370000003a000000350000003e",
            INIT_39 => X"0000004500000044000000480000004c0000004b0000003a0000003700000039",
            INIT_3A => X"00000035000000370000003a00000046000000490000004b0000004a0000004b",
            INIT_3B => X"00000033000000360000003a0000005b0000007f0000006b0000004500000033",
            INIT_3C => X"000000350000003900000038000000330000002e000000330000003300000040",
            INIT_3D => X"000000390000003c0000003e000000400000003e000000320000003300000034",
            INIT_3E => X"0000003700000034000000350000004000000040000000400000003e0000003c",
            INIT_3F => X"0000003200000034000000320000003500000048000000690000006700000046",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE23;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE24 : if BRAM_NAME = "sampleifmap_layer0_instance24" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002d0000002c00000028000000170000001e000000300000004600000041",
            INIT_01 => X"0000003000000033000000350000002c0000000f0000000a000000280000002d",
            INIT_02 => X"000000370000003c000000510000005f0000005b0000005d0000005a00000041",
            INIT_03 => X"0000004300000036000000330000004d00000044000000290000006f00000070",
            INIT_04 => X"000000310000003100000041000000290000001e0000003c0000004f00000045",
            INIT_05 => X"0000003100000037000000450000004100000019000000070000002300000031",
            INIT_06 => X"0000003b0000003700000051000000570000005000000053000000550000004d",
            INIT_07 => X"0000003d0000004100000036000000380000002f0000001f0000007900000083",
            INIT_08 => X"00000036000000320000004a0000004000000029000000480000005400000049",
            INIT_09 => X"000000270000002f000000430000003c000000240000000b0000002000000036",
            INIT_0A => X"0000003f0000003000000055000000530000003e0000003b0000004d0000004b",
            INIT_0B => X"00000030000000490000004e000000460000002900000017000000800000008b",
            INIT_0C => X"0000003f00000037000000440000005000000036000000500000004b00000058",
            INIT_0D => X"0000002700000028000000330000002b00000025000000110000001c0000003a",
            INIT_0E => X"00000044000000320000005400000056000000460000004b0000006200000055",
            INIT_0F => X"00000026000000410000005d000000640000004b0000002f000000890000008e",
            INIT_10 => X"000000440000003d0000003d00000051000000420000006f000000590000005f",
            INIT_11 => X"0000003f00000033000000230000001f000000160000000f000000160000003e",
            INIT_12 => X"0000004e00000033000000530000004d00000047000000480000004b00000048",
            INIT_13 => X"000000580000004b0000005f0000006300000057000000570000009c00000095",
            INIT_14 => X"00000039000000400000003a000000470000004d000000520000005300000052",
            INIT_15 => X"00000047000000470000003d000000320000001c00000011000000140000003b",
            INIT_16 => X"0000004e00000046000000530000002900000038000000440000004300000045",
            INIT_17 => X"00000063000000700000006f0000005e0000005900000062000000ac0000009c",
            INIT_18 => X"00000031000000490000004a000000480000003b000000200000004000000045",
            INIT_19 => X"0000003f0000005600000055000000520000003e0000001d0000001200000031",
            INIT_1A => X"0000004e000000550000005e000000190000002b0000005f0000003400000022",
            INIT_1B => X"0000002f00000056000000830000006c0000006b0000006d000000b4000000a6",
            INIT_1C => X"0000003d000000500000004e000000510000004600000019000000350000003b",
            INIT_1D => X"000000190000004b00000058000000570000005e000000350000000a00000028",
            INIT_1E => X"00000062000000590000006500000032000000390000005c0000002d0000000d",
            INIT_1F => X"0000001800000034000000800000007c0000007c00000078000000b300000090",
            INIT_20 => X"0000004f0000003f000000590000007700000066000000310000002f00000044",
            INIT_21 => X"0000000e000000290000005a0000005900000060000000510000002200000042",
            INIT_22 => X"000000730000006e000000710000006f00000047000000430000005c00000034",
            INIT_23 => X"000000160000001f000000730000007c0000007f000000790000009c00000088",
            INIT_24 => X"00000037000000410000007b000000800000007200000037000000350000004d",
            INIT_25 => X"0000002500000014000000450000006a0000006e0000006f000000520000004f",
            INIT_26 => X"0000005c0000007300000078000000760000006100000053000000690000005c",
            INIT_27 => X"000000170000000e0000005f000000770000007f0000007d0000009300000090",
            INIT_28 => X"0000003100000064000000840000008100000070000000360000003a00000055",
            INIT_29 => X"000000530000003f0000005d0000007d0000006d000000680000005400000027",
            INIT_2A => X"00000039000000550000007f0000006d0000006e000000680000005e00000061",
            INIT_2B => X"000000150000000c0000005d000000720000007c0000007b0000009600000098",
            INIT_2C => X"0000004b00000080000000830000007e0000006b00000032000000350000006c",
            INIT_2D => X"00000093000000810000006e0000008a0000006b000000550000005b00000033",
            INIT_2E => X"0000005d0000005a000000730000007500000077000000710000007800000084",
            INIT_2F => X"000000090000000e00000065000000790000007d000000710000008d000000a0",
            INIT_30 => X"0000007700000082000000800000006a0000005c0000002b0000002a00000060",
            INIT_31 => X"00000084000000690000006e0000009400000089000000720000007b00000078",
            INIT_32 => X"000000770000007e000000780000008c00000086000000800000008700000092",
            INIT_33 => X"000000280000001200000063000000820000006a000000630000009100000098",
            INIT_34 => X"00000088000000850000006f00000064000000590000003b0000004200000061",
            INIT_35 => X"0000007f00000083000000880000008e00000091000000960000008c00000093",
            INIT_36 => X"000000880000009c0000008e0000009700000093000000880000007b0000007d",
            INIT_37 => X"00000053000000320000005c00000082000000700000006d0000009000000092",
            INIT_38 => X"00000085000000850000005e000000680000005f0000004b0000004800000069",
            INIT_39 => X"00000098000000a000000096000000930000008500000080000000870000008f",
            INIT_3A => X"000000a5000000a20000008a0000008a00000087000000840000009000000091",
            INIT_3B => X"0000004d0000003b0000005f00000076000000770000007e0000007f000000a3",
            INIT_3C => X"000000830000007b00000062000000650000005b00000044000000440000005e",
            INIT_3D => X"000000a200000093000000930000007c0000004f0000008a000000c100000093",
            INIT_3E => X"000000b30000009400000079000000900000009000000098000000ab000000b4",
            INIT_3F => X"000000540000001a0000003f000000700000007b00000080000000a0000000b4",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE24;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE25 : if BRAM_NAME = "sampleifmap_layer0_instance25" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000008100000078000000780000006e000000590000004a0000004f00000058",
            INIT_01 => X"000000a6000000a40000009c0000007200000057000000c0000000b800000078",
            INIT_02 => X"0000008f00000094000000ad000000bb000000b6000000b7000000a10000009a",
            INIT_03 => X"00000076000000290000002c0000006b0000007c0000008e000000c3000000b5",
            INIT_04 => X"0000006a0000006f00000064000000740000006000000067000000590000005b",
            INIT_05 => X"000000ac000000ac000000990000008c000000a8000000bb0000008000000072",
            INIT_06 => X"0000009c000000ab000000a5000000a1000000a30000009d000000a4000000a7",
            INIT_07 => X"0000005e0000002a0000004a0000006a00000072000000a700000091000000a1",
            INIT_08 => X"0000005b0000005f0000004e000000720000007a000000780000006100000065",
            INIT_09 => X"00000099000000a000000089000000a7000000cc000000810000006e00000073",
            INIT_0A => X"000000a5000000a20000009c000000b3000000b2000000aa000000ba000000b3",
            INIT_0B => X"0000007200000046000000590000005400000048000000680000008c0000009c",
            INIT_0C => X"00000064000000480000004c0000005a000000600000007a0000006b0000006e",
            INIT_0D => X"000000b4000000a60000009f000000bd0000008c000000570000007f0000006d",
            INIT_0E => X"000000a1000000a200000099000000a2000000bc000000be000000ad000000ae",
            INIT_0F => X"0000008a000000700000003e000000420000004a0000004b0000009500000099",
            INIT_10 => X"000000670000003c00000047000000590000004e000000590000006a00000077",
            INIT_11 => X"000000be000000ae000000b50000007f00000042000000720000005f0000004b",
            INIT_12 => X"000000a5000000ab000000a0000000a4000000c1000000b8000000ab000000ba",
            INIT_13 => X"00000073000000700000005e0000004d0000005c000000680000008b00000092",
            INIT_14 => X"0000005f000000480000004c0000006a000000670000003a0000005e0000007e",
            INIT_15 => X"000000bc000000c4000000a10000005b0000006300000078000000410000005e",
            INIT_16 => X"000000a10000009a000000a0000000aa000000a7000000a7000000c1000000b6",
            INIT_17 => X"000000640000006d0000008800000069000000510000006e0000008a00000091",
            INIT_18 => X"00000054000000450000005e000000710000006800000046000000520000006f",
            INIT_19 => X"000000c8000000ba0000009b0000007f0000007d000000550000006d00000074",
            INIT_1A => X"000000a6000000a4000000a2000000940000009d000000b1000000bb000000bb",
            INIT_1B => X"00000061000000610000007300000078000000610000007900000095000000a2",
            INIT_1C => X"0000004c000000550000007b00000097000000b40000008c0000005c00000065",
            INIT_1D => X"000000c8000000ad000000af00000092000000540000005a0000007c00000067",
            INIT_1E => X"000000ad000000a3000000ac0000009f0000009f000000ad000000ad000000bc",
            INIT_1F => X"00000060000000640000005f0000007000000083000000830000008b000000a4",
            INIT_20 => X"0000006c0000007f0000009d000000c2000000d1000000c00000009000000077",
            INIT_21 => X"000000c5000000b0000000af0000007c0000006f0000006a0000005e0000006a",
            INIT_22 => X"000000a3000000af000000c50000009c000000a5000000b0000000aa000000b8",
            INIT_23 => X"000000660000006b0000006000000064000000650000007a0000008300000093",
            INIT_24 => X"00000088000000a0000000c4000000c5000000a90000008a000000740000006e",
            INIT_25 => X"000000a9000000b40000009f000000920000008a0000005c0000006300000081",
            INIT_26 => X"00000097000000b3000000bc000000a6000000b2000000af0000008d0000008e",
            INIT_27 => X"0000004900000066000000650000005b0000003a000000700000009a0000008f",
            INIT_28 => X"000000a3000000bf000000b9000000a50000006b0000004a000000570000005b",
            INIT_29 => X"00000074000000920000008400000076000000660000006a0000008000000086",
            INIT_2A => X"000000a7000000ad0000009f000000b7000000b6000000a1000000630000004d",
            INIT_2B => X"0000004d000000440000005c0000005b0000002b0000005e000000870000009c",
            INIT_2C => X"000000bb000000a6000000940000005f0000002c000000320000005f00000051",
            INIT_2D => X"0000006b000000770000007200000068000000720000007e00000090000000ae",
            INIT_2E => X"00000096000000a9000000b2000000a9000000b60000009d0000005200000051",
            INIT_2F => X"000000560000005000000045000000610000003f0000002c0000006c00000098",
            INIT_30 => X"000000b0000000920000006d0000001c00000015000000340000005f0000005a",
            INIT_31 => X"000000820000007200000077000000780000007f0000008e000000b5000000ca",
            INIT_32 => X"00000098000000b4000000ad0000009f000000a9000000900000007600000081",
            INIT_33 => X"0000006a000000a70000007200000033000000550000002c0000004400000077",
            INIT_34 => X"0000009c00000077000000310000001800000034000000390000005b0000005f",
            INIT_35 => X"0000007500000074000000850000008d0000009b000000ba000000cb000000bb",
            INIT_36 => X"0000007d0000009c000000a70000009f000000990000008b000000770000006d",
            INIT_37 => X"0000007a000000aa000000900000003700000040000000440000004100000065",
            INIT_38 => X"0000007300000036000000210000002e00000049000000200000004b0000005e",
            INIT_39 => X"00000092000000880000009b000000b1000000c2000000c3000000b000000096",
            INIT_3A => X"00000069000000600000005f00000065000000770000005e000000650000008b",
            INIT_3B => X"0000006a0000009a0000008f000000800000006d0000006b0000007600000083",
            INIT_3C => X"0000003b0000001b00000028000000410000004c00000018000000230000004e",
            INIT_3D => X"000000ba000000a5000000b7000000c0000000b0000000960000008800000078",
            INIT_3E => X"0000008c000000700000005500000042000000560000006b000000aa000000cf",
            INIT_3F => X"000000800000009a0000008f00000096000000890000008900000095000000a9",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE25;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE26 : if BRAM_NAME = "sampleifmap_layer0_instance26" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000500000004b00000039000000210000002e000000400000005100000044",
            INIT_01 => X"00000042000000460000004b0000004700000022000000140000004600000053",
            INIT_02 => X"00000052000000540000006c0000007e000000790000007c0000007800000057",
            INIT_03 => X"000000570000004c00000043000000600000005b0000003b0000008100000088",
            INIT_04 => X"00000054000000540000005c000000380000002f0000004a0000006600000050",
            INIT_05 => X"000000490000004d0000005c0000005d00000030000000120000003e00000058",
            INIT_06 => X"000000530000004d0000006c000000750000006a0000006f000000750000006b",
            INIT_07 => X"000000510000005a0000004200000047000000410000002d0000008b00000097",
            INIT_08 => X"0000005a00000056000000690000005400000038000000580000006d0000005f",
            INIT_09 => X"0000003c0000004200000058000000590000003c00000014000000350000005c",
            INIT_0A => X"00000056000000420000007200000072000000540000004e0000006600000067",
            INIT_0B => X"0000003b00000062000000620000005400000037000000230000008f0000009e",
            INIT_0C => X"0000006000000058000000660000006d00000049000000640000006400000074",
            INIT_0D => X"00000037000000360000004300000041000000380000001a0000002d0000005e",
            INIT_0E => X"0000005b0000004500000072000000760000006200000061000000750000006a",
            INIT_0F => X"000000320000005e0000007e000000780000005d0000004000000096000000a0",
            INIT_10 => X"0000005e0000005a0000005e000000720000005d000000800000006800000078",
            INIT_11 => X"0000005600000049000000370000002f000000240000001a000000270000005d",
            INIT_12 => X"000000670000004a0000006d00000067000000650000006b0000007100000069",
            INIT_13 => X"0000006c0000006700000084000000810000007400000070000000ac000000a2",
            INIT_14 => X"0000004e0000005b000000590000005f00000062000000620000006600000069",
            INIT_15 => X"0000006c0000006a0000005d0000004d0000002b0000001b0000002300000058",
            INIT_16 => X"00000066000000620000006e000000390000004e000000640000006500000067",
            INIT_17 => X"000000780000008400000090000000810000007f00000082000000ba000000a7",
            INIT_18 => X"0000003f0000005d000000640000005a0000004f00000030000000600000005e",
            INIT_19 => X"0000006300000082000000810000007e0000005a000000260000001d0000004a",
            INIT_1A => X"0000006a000000710000007b000000250000003900000073000000470000003a",
            INIT_1B => X"0000003b00000065000000a0000000890000008c0000008d000000c1000000b7",
            INIT_1C => X"000000470000005e0000006100000067000000690000002f0000005400000056",
            INIT_1D => X"00000029000000720000008c0000008a0000008b000000490000001400000038",
            INIT_1E => X"0000008c000000780000007d0000003b0000004f00000073000000410000001a",
            INIT_1F => X"000000180000003f0000009b000000900000009400000096000000c3000000b0",
            INIT_20 => X"0000005c0000005000000072000000950000008c0000004a0000004e00000062",
            INIT_21 => X"000000170000003f000000860000008800000090000000710000002c00000047",
            INIT_22 => X"000000a50000009b0000008b00000070000000560000005e0000007c00000045",
            INIT_23 => X"00000016000000290000008e000000920000009600000096000000b1000000aa",
            INIT_24 => X"00000045000000540000009b000000a3000000940000004e0000005100000074",
            INIT_25 => X"00000038000000210000005d0000008a0000008e000000890000005a00000051",
            INIT_26 => X"000000810000009c0000009c0000009700000080000000730000008f0000007c",
            INIT_27 => X"000000180000001600000079000000940000009a00000098000000ad000000a7",
            INIT_28 => X"000000410000007f000000a6000000a500000091000000490000004f00000078",
            INIT_29 => X"0000006c000000470000005d0000007e0000007f0000008e0000007200000036",
            INIT_2A => X"0000005700000075000000a50000009c000000a1000000920000008500000087",
            INIT_2B => X"000000170000001300000074000000910000009c00000097000000af000000a9",
            INIT_2C => X"0000005f000000a5000000a8000000a10000008a00000042000000450000007b",
            INIT_2D => X"000000a200000088000000660000006d000000700000008a0000008c0000004b",
            INIT_2E => X"0000008800000076000000850000007c00000087000000970000009a00000099",
            INIT_2F => X"0000000b0000001400000077000000940000009d00000092000000aa000000bd",
            INIT_30 => X"00000098000000ad000000a400000087000000790000003c000000390000006a",
            INIT_31 => X"0000008b000000660000005c00000073000000760000007f0000009300000090",
            INIT_32 => X"00000088000000770000006b0000007800000074000000850000008a0000008d",
            INIT_33 => X"0000002b0000001a00000072000000a10000009100000087000000ae000000b0",
            INIT_34 => X"000000ab000000ac0000008c0000007f000000740000004e0000005500000074",
            INIT_35 => X"0000006e00000071000000760000007700000078000000820000007c00000099",
            INIT_36 => X"00000075000000810000007a000000830000007d000000770000006c00000069",
            INIT_37 => X"0000005f0000004100000070000000a60000009a0000008d000000a200000090",
            INIT_38 => X"000000a8000000a5000000720000008200000078000000630000006000000084",
            INIT_39 => X"000000840000008e000000810000007c00000070000000680000006b0000008b",
            INIT_3A => X"000000900000008d00000076000000730000006f0000006b000000770000007a",
            INIT_3B => X"0000005e00000048000000700000009d0000009f000000920000007b0000008e",
            INIT_3C => X"000000a6000000970000007c0000007f000000760000005d0000005a00000079",
            INIT_3D => X"0000008b0000007b0000007c0000006b0000004500000079000000ab00000099",
            INIT_3E => X"000000a700000083000000670000007a0000007700000080000000900000009b",
            INIT_3F => X"00000068000000220000004b00000095000000a0000000800000008c0000009f",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE26;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE27 : if BRAM_NAME = "sampleifmap_layer0_instance27" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a300000095000000980000008d0000007e000000640000006400000070",
            INIT_01 => X"0000008d0000008b000000850000006400000047000000a6000000a30000008a",
            INIT_02 => X"0000007e0000007d00000097000000a30000009e000000a00000008800000081",
            INIT_03 => X"0000008b000000330000003d0000008f0000008f0000007a000000b1000000a9",
            INIT_04 => X"00000089000000900000007c0000009300000081000000830000007000000070",
            INIT_05 => X"00000093000000920000007f0000007a00000099000000a8000000790000008f",
            INIT_06 => X"00000086000000990000008f000000860000008a000000840000008b0000008d",
            INIT_07 => X"0000006f0000003a00000064000000860000007a000000920000008200000091",
            INIT_08 => X"000000760000007b000000610000008d0000008e000000950000007600000079",
            INIT_09 => X"00000082000000880000006e00000091000000bb000000790000007e0000008f",
            INIT_0A => X"000000910000009600000086000000970000009a00000094000000a10000009a",
            INIT_0B => X"0000008600000061000000770000006700000057000000610000007b00000086",
            INIT_0C => X"0000007d0000005d000000650000007a0000006f000000970000008700000088",
            INIT_0D => X"000000a00000009200000088000000a90000007d000000600000009900000086",
            INIT_0E => X"0000009100000090000000800000008d000000a7000000a60000009400000096",
            INIT_0F => X"000000a90000009500000057000000530000005e0000004b0000008200000084",
            INIT_10 => X"000000820000005400000068000000790000005e000000700000008c00000094",
            INIT_11 => X"000000aa0000009b000000a3000000760000004a0000008d0000007400000066",
            INIT_12 => X"00000091000000930000008900000092000000a70000009d00000095000000a5",
            INIT_13 => X"000000a10000009c0000007700000060000000710000006d0000007c0000007f",
            INIT_14 => X"000000790000006300000065000000810000007d000000480000007700000098",
            INIT_15 => X"000000a9000000b5000000960000005d0000007d0000009a0000005b00000078",
            INIT_16 => X"0000008b00000081000000870000008f0000008f00000091000000ad000000a2",
            INIT_17 => X"000000990000009a000000ab000000810000006600000075000000780000007d",
            INIT_18 => X"000000730000006200000076000000880000007b000000520000006800000088",
            INIT_19 => X"000000b3000000ad000000950000008100000094000000750000008d00000096",
            INIT_1A => X"0000008d0000008c0000008b0000007e0000008f0000009f000000a8000000a5",
            INIT_1B => X"0000009500000096000000a4000000980000006d0000007a0000008500000088",
            INIT_1C => X"0000006f000000790000009e000000ac000000bf000000960000006f0000007d",
            INIT_1D => X"000000ac0000009a000000a10000009400000069000000730000009900000091",
            INIT_1E => X"0000008f0000008800000093000000890000008d0000009c0000009b000000a1",
            INIT_1F => X"000000950000009e000000950000009c000000860000007b0000008c00000089",
            INIT_20 => X"00000093000000aa000000bd000000d1000000dc000000c8000000a200000095",
            INIT_21 => X"000000a4000000960000009f0000008b000000880000007d0000007a00000091",
            INIT_22 => X"0000008800000093000000a9000000850000008e0000009f0000009b0000009b",
            INIT_23 => X"0000009c000000a00000008f0000009a000000720000006b0000007e0000007f",
            INIT_24 => X"000000b0000000bf000000d7000000d5000000be0000009d000000890000008b",
            INIT_25 => X"0000008f0000009a00000097000000ad000000a30000007500000084000000a9",
            INIT_26 => X"0000007c00000095000000a3000000910000009800000099000000810000007c",
            INIT_27 => X"000000780000009700000095000000910000004a000000600000008300000077",
            INIT_28 => X"000000c1000000d3000000cf000000bf00000086000000610000006f00000073",
            INIT_29 => X"00000068000000860000008f000000900000007f00000091000000ad000000b1",
            INIT_2A => X"0000008e000000940000008a000000a10000009b0000008b0000005c00000049",
            INIT_2B => X"0000006d0000006f00000091000000920000003c000000550000007500000083",
            INIT_2C => X"000000d5000000c3000000b2000000780000004000000041000000720000006a",
            INIT_2D => X"0000007d0000008d000000960000008e00000099000000ad000000b9000000ca",
            INIT_2E => X"0000007f00000095000000a1000000900000009a0000008e000000600000006c",
            INIT_2F => X"00000075000000760000006c0000009300000061000000310000006200000083",
            INIT_30 => X"000000c7000000b40000008700000029000000260000003e0000007000000074",
            INIT_31 => X"000000a10000009e000000a4000000ab000000b2000000b7000000cc000000d4",
            INIT_32 => X"0000007e0000009c00000099000000870000008d000000870000008b0000009d",
            INIT_33 => X"00000083000000c500000088000000540000007c0000003b0000004200000067",
            INIT_34 => X"000000bf0000009500000042000000250000004e0000004f0000007b0000007f",
            INIT_35 => X"0000009f000000a5000000b4000000b8000000c2000000d6000000db000000d0",
            INIT_36 => X"0000007200000087000000930000008a000000830000007b0000007d00000087",
            INIT_37 => X"0000008f000000c9000000ac0000004e0000005b000000550000004f0000006c",
            INIT_38 => X"000000970000004e00000030000000430000006b00000034000000680000007d",
            INIT_39 => X"000000b6000000b4000000c3000000cd000000da000000d9000000cb000000bd",
            INIT_3A => X"0000006f0000005900000059000000610000007a0000005e00000074000000a5",
            INIT_3B => X"00000081000000bc000000b50000009f00000086000000820000008a00000096",
            INIT_3C => X"0000004e000000290000003a0000006000000073000000280000003300000066",
            INIT_3D => X"000000ce000000c4000000d2000000da000000cf000000b9000000b5000000a0",
            INIT_3E => X"000000a0000000840000006600000056000000710000007c000000b4000000d6",
            INIT_3F => X"0000009c000000b9000000b3000000b4000000a7000000a7000000a7000000ba",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE27;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE28 : if BRAM_NAME = "sampleifmap_layer0_instance28" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000390000003700000024000000160000001e0000002e0000004000000032",
            INIT_01 => X"00000032000000310000002c0000002b000000120000000c000000360000003b",
            INIT_02 => X"00000039000000380000004e000000530000004d000000510000004d0000003a",
            INIT_03 => X"000000420000003500000029000000410000003a0000001f0000005d00000061",
            INIT_04 => X"0000003c0000003b0000003d000000230000001d00000039000000510000003a",
            INIT_05 => X"0000002f0000003b0000003e000000380000001b000000070000002f00000040",
            INIT_06 => X"0000003c00000033000000510000004e000000440000004a0000004a00000044",
            INIT_07 => X"00000042000000450000002c0000002d0000002700000015000000600000006f",
            INIT_08 => X"000000410000003c000000480000003500000023000000460000005700000048",
            INIT_09 => X"0000002100000030000000410000003400000023000000070000002600000045",
            INIT_0A => X"0000003e0000002d000000520000004d00000037000000320000004200000043",
            INIT_0B => X"000000330000004d0000004b0000003f00000026000000100000006300000074",
            INIT_0C => X"0000004a0000004100000048000000470000002f000000500000004c0000005e",
            INIT_0D => X"0000001e000000230000003400000028000000220000000c0000001e00000048",
            INIT_0E => X"000000430000002e0000004d000000510000004500000044000000570000004b",
            INIT_0F => X"0000002200000044000000600000005f000000490000002a0000006b00000077",
            INIT_10 => X"0000004c00000048000000440000004b0000003c0000006a0000004f00000061",
            INIT_11 => X"0000003b00000033000000250000001c000000110000000c0000001800000049",
            INIT_12 => X"0000004d0000002d0000004900000047000000470000004b0000004f00000048",
            INIT_13 => X"0000005000000049000000610000005e00000055000000520000008100000080",
            INIT_14 => X"0000003d0000004d000000450000003d000000430000004b0000004d00000052",
            INIT_15 => X"00000049000000470000003b0000002c000000160000000d0000001300000043",
            INIT_16 => X"0000004d0000003e000000490000002200000035000000490000004800000048",
            INIT_17 => X"0000005c000000680000006e0000005c0000005b000000600000009300000088",
            INIT_18 => X"000000320000004f0000004f0000003e00000033000000190000004600000048",
            INIT_19 => X"0000003e0000004d0000004b0000004900000036000000180000000f00000038",
            INIT_1A => X"0000004a0000004800000058000000160000002a000000600000003300000022",
            INIT_1B => X"0000002b00000051000000830000006b0000006c00000068000000a100000095",
            INIT_1C => X"0000003a0000004b000000480000004d00000046000000150000003b0000003f",
            INIT_1D => X"000000120000003e0000004b0000004b000000510000002f0000000800000029",
            INIT_1E => X"00000053000000480000005e0000002a00000040000000590000002700000006",
            INIT_1F => X"000000150000003400000085000000760000007800000072000000a200000083",
            INIT_20 => X"0000004600000039000000580000007900000068000000310000003500000049",
            INIT_21 => X"00000007000000220000004f0000004e00000053000000470000001700000033",
            INIT_22 => X"0000005d0000005b00000063000000500000003e0000003c0000005100000028",
            INIT_23 => X"00000014000000210000007c0000007900000079000000780000008d00000073",
            INIT_24 => X"00000033000000400000007f0000008300000076000000380000003a00000056",
            INIT_25 => X"0000001c0000000d0000003a0000005e0000006300000061000000400000003b",
            INIT_26 => X"0000004a0000005f000000690000006200000050000000490000005d00000053",
            INIT_27 => X"000000170000000d000000650000007f0000007e000000770000008400000074",
            INIT_28 => X"0000003000000067000000870000008400000074000000350000003b0000005b",
            INIT_29 => X"00000049000000320000004a0000006600000061000000600000004b00000020",
            INIT_2A => X"00000031000000470000006c000000620000006100000059000000520000005a",
            INIT_2B => X"000000140000000a0000005b0000007b0000008a000000770000007c00000077",
            INIT_2C => X"000000480000008700000087000000810000006e0000002f0000003300000065",
            INIT_2D => X"0000008700000075000000560000005e0000004f00000052000000540000002e",
            INIT_2E => X"000000580000004a000000580000005c0000005e0000005d0000006600000078",
            INIT_2F => X"000000070000000b0000005b000000770000008d000000760000007300000084",
            INIT_30 => X"000000770000008b000000830000006b00000060000000280000002800000058",
            INIT_31 => X"0000006c000000510000004a0000005f0000005900000057000000660000006b",
            INIT_32 => X"0000005f0000005700000055000000660000005d000000640000006e00000076",
            INIT_33 => X"000000200000000f000000590000007b0000007100000065000000780000007c",
            INIT_34 => X"000000890000008b0000006e000000640000005c000000370000003f0000005f",
            INIT_35 => X"0000005600000056000000580000005a0000005c00000065000000610000007b",
            INIT_36 => X"0000005f0000006e0000006c000000720000006c000000640000005800000055",
            INIT_37 => X"0000004c000000310000005800000080000000730000006b000000750000006d",
            INIT_38 => X"000000870000008600000056000000680000006000000047000000450000006a",
            INIT_39 => X"0000006a0000006e000000600000006000000058000000510000005700000074",
            INIT_3A => X"000000800000007f0000006b000000610000005c000000570000005f00000062",
            INIT_3B => X"00000046000000350000005c0000007a00000077000000740000005e0000007a",
            INIT_3C => X"00000085000000790000005f000000670000005c000000400000004000000060",
            INIT_3D => X"0000007100000062000000650000005800000033000000640000009600000081",
            INIT_3E => X"000000980000007100000053000000600000005f000000650000007700000083",
            INIT_3F => X"000000480000000d00000039000000760000007c000000620000007800000094",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE28;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE29 : if BRAM_NAME = "sampleifmap_layer0_instance29" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000082000000780000007c000000730000005a000000470000004c00000057",
            INIT_01 => X"000000780000007700000074000000540000003a000000960000008e0000006e",
            INIT_02 => X"0000006e000000670000007e000000890000008600000085000000710000006c",
            INIT_03 => X"0000006b000000210000002a000000750000007200000063000000a30000009f",
            INIT_04 => X"000000690000007500000063000000750000005d000000640000005800000056",
            INIT_05 => X"00000081000000810000006f0000006b0000008b0000009b000000660000006e",
            INIT_06 => X"000000710000007c0000007600000071000000760000006d000000770000007c",
            INIT_07 => X"0000005700000027000000480000006900000063000000830000007500000083",
            INIT_08 => X"0000005600000063000000470000006d0000007300000078000000600000005f",
            INIT_09 => X"000000750000007b0000005e00000082000000b00000006a000000630000006c",
            INIT_0A => X"00000079000000780000006f0000008300000088000000810000008d00000089",
            INIT_0B => X"0000006e00000043000000510000004800000043000000500000006b00000075",
            INIT_0C => X"0000005e000000470000004800000058000000570000007d000000700000006d",
            INIT_0D => X"0000009400000087000000760000009800000073000000490000007900000064",
            INIT_0E => X"0000007a00000079000000710000007d00000095000000940000008200000085",
            INIT_0F => X"0000008a00000073000000380000003d0000004e0000003a0000007100000072",
            INIT_10 => X"000000660000003c000000480000005800000043000000590000007400000077",
            INIT_11 => X"0000009c0000008d0000009200000065000000370000006d0000005700000048",
            INIT_12 => X"0000007c0000007f0000007b00000086000000980000008c0000008800000098",
            INIT_13 => X"000000770000007a000000620000004d000000620000005d000000690000006d",
            INIT_14 => X"000000600000004b00000046000000600000005d00000032000000610000007e",
            INIT_15 => X"00000097000000a2000000830000004900000061000000760000003b0000005a",
            INIT_16 => X"000000750000006e000000760000007d0000007f00000084000000a300000096",
            INIT_17 => X"0000006a000000700000008e0000006b0000004f0000005e0000006600000069",
            INIT_18 => X"00000059000000450000004e0000005c00000059000000370000005100000070",
            INIT_19 => X"0000009c000000970000007d0000006b00000076000000530000006b00000077",
            INIT_1A => X"00000075000000780000007b0000006c0000007e000000940000009b00000094",
            INIT_1B => X"0000006900000063000000790000008100000056000000540000006600000072",
            INIT_1C => X"0000004e000000450000005f000000770000009a000000780000005600000062",
            INIT_1D => X"00000096000000840000008b0000007d0000004e000000570000007e00000073",
            INIT_1E => X"0000007b0000007600000084000000790000007e000000920000008e0000008d",
            INIT_1F => X"000000670000006a00000065000000790000006f000000520000005800000073",
            INIT_20 => X"0000005c00000060000000770000009f000000b6000000a70000008800000074",
            INIT_21 => X"0000008f0000008300000088000000700000006f000000660000005a00000066",
            INIT_22 => X"00000077000000840000009c0000007500000080000000960000008e00000086",
            INIT_23 => X"0000006c00000071000000600000006a000000530000004e0000005900000066",
            INIT_24 => X"000000690000007b0000009e000000a600000092000000710000006d0000006c",
            INIT_25 => X"0000007b000000860000007e000000910000008c000000550000005200000066",
            INIT_26 => X"0000006a0000008a0000009600000083000000890000008a0000007300000068",
            INIT_27 => X"0000004b0000006900000065000000600000002d0000004a0000006f00000061",
            INIT_28 => X"0000007e00000097000000970000008b00000056000000370000005500000058",
            INIT_29 => X"000000520000006e0000006e0000006f00000057000000570000006800000068",
            INIT_2A => X"0000007a0000008100000078000000910000008c000000790000004b00000035",
            INIT_2B => X"00000040000000410000006200000061000000200000003e0000006200000074",
            INIT_2C => X"0000009c00000086000000750000004b00000020000000220000005c00000052",
            INIT_2D => X"0000005f0000005b0000005a0000005200000057000000620000006d0000008d",
            INIT_2E => X"0000006b000000800000008f000000810000008b000000790000004600000052",
            INIT_2F => X"000000420000004700000047000000630000003f0000001d0000004e00000071",
            INIT_30 => X"00000094000000720000004e0000000f0000000d00000023000000560000005a",
            INIT_31 => X"00000071000000560000005b00000061000000620000006f0000008b000000a2",
            INIT_32 => X"0000006a0000008700000087000000760000007e000000730000006a00000078",
            INIT_33 => X"0000005300000099000000600000002c0000005b000000260000002a0000004f",
            INIT_34 => X"0000007a000000570000001f0000000d000000250000002d000000560000005c",
            INIT_35 => X"0000005c0000005d00000072000000750000007a0000009e000000ad00000096",
            INIT_36 => X"0000005b00000073000000850000007e0000007100000067000000550000004d",
            INIT_37 => X"00000062000000860000006c0000002a0000003c0000003b000000320000004e",
            INIT_38 => X"0000005400000023000000170000002400000038000000180000004700000052",
            INIT_39 => X"000000790000006f0000008200000096000000a5000000a50000009200000076",
            INIT_3A => X"0000005600000046000000450000004e000000620000003f000000420000006c",
            INIT_3B => X"000000590000007b000000740000007800000062000000600000006c00000075",
            INIT_3C => X"000000250000000f0000001d0000003400000040000000110000001b00000041",
            INIT_3D => X"0000009c0000008800000098000000aa00000096000000740000006400000059",
            INIT_3E => X"0000007f00000066000000470000002f0000004a0000004500000079000000a6",
            INIT_3F => X"0000007500000092000000880000009300000082000000830000008b0000009c",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE29;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE30 : if BRAM_NAME = "sampleifmap_layer0_instance30" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000970000009c0000009d0000008d000000580000004d0000008b000000b3",
            INIT_01 => X"0000007600000079000000880000009700000097000000900000009e0000009c",
            INIT_02 => X"000000530000005e000000620000006200000054000000540000006c0000007e",
            INIT_03 => X"0000004d0000004c00000057000000750000006000000054000000560000005a",
            INIT_04 => X"000000a70000009e0000009f0000009f000000920000008000000085000000b8",
            INIT_05 => X"0000007d0000008800000096000000960000009a00000099000000a2000000a5",
            INIT_06 => X"000000580000005e000000620000005d000000520000005a0000006d00000081",
            INIT_07 => X"0000005a0000005b00000062000000760000006a0000005b0000004c0000004e",
            INIT_08 => X"000000a40000009b00000098000000a4000000aa000000b000000098000000b4",
            INIT_09 => X"0000008c00000092000000970000009c0000009f000000a2000000aa000000a2",
            INIT_0A => X"0000006b00000067000000620000005500000047000000580000007c00000092",
            INIT_0B => X"0000005f0000005d000000650000006f0000006f0000006f0000006d00000065",
            INIT_0C => X"000000a3000000a400000098000000a8000000b5000000b8000000ae000000af",
            INIT_0D => X"000000a40000009f000000a2000000ae000000a8000000a7000000b3000000a6",
            INIT_0E => X"0000006b000000630000005a000000480000003a000000590000008900000097",
            INIT_0F => X"0000006f0000006d0000006100000069000000790000007d0000008000000075",
            INIT_10 => X"000000af000000b0000000a1000000a2000000ac000000a7000000ae000000af",
            INIT_11 => X"000000a4000000a0000000a8000000b0000000b4000000b3000000b2000000b2",
            INIT_12 => X"0000005e000000630000005a0000004200000045000000780000009c000000ad",
            INIT_13 => X"000000740000007100000068000000700000007b0000007f0000007c00000069",
            INIT_14 => X"000000b3000000b0000000a6000000a9000000aa00000090000000ae000000b5",
            INIT_15 => X"000000960000009f000000ae000000b0000000b5000000b4000000b4000000b4",
            INIT_16 => X"00000070000000830000007d00000060000000740000009b000000af000000b5",
            INIT_17 => X"0000007c000000760000007800000079000000790000007a0000007800000075",
            INIT_18 => X"000000af000000b0000000ae000000af000000b20000008a0000009c000000c0",
            INIT_19 => X"00000099000000ad000000bb000000bb000000b8000000ba000000b4000000b8",
            INIT_1A => X"00000079000000940000009500000096000000a7000000ad000000ad000000a6",
            INIT_1B => X"000000800000007b0000007a000000780000006f0000006d0000007500000073",
            INIT_1C => X"000000b8000000af000000af000000ad000000ab0000009c0000007d000000b9",
            INIT_1D => X"000000a6000000b8000000b9000000bd000000c2000000c1000000b7000000bc",
            INIT_1E => X"0000007a0000008f00000089000000aa000000b0000000b1000000ac000000a4",
            INIT_1F => X"0000007d0000007b000000760000007500000067000000600000006e0000006b",
            INIT_20 => X"000000b4000000b2000000ad000000ac000000a00000009f000000950000009b",
            INIT_21 => X"000000a0000000ac000000af000000bb000000bf000000ba000000ba000000bb",
            INIT_22 => X"00000085000000a60000009b000000b7000000b0000000a6000000970000009a",
            INIT_23 => X"0000007d0000007a0000007a0000007600000077000000700000006800000068",
            INIT_24 => X"000000aa000000b7000000b2000000b2000000a900000093000000980000009a",
            INIT_25 => X"000000a9000000a5000000a7000000ae000000c1000000c6000000bc000000b0",
            INIT_26 => X"0000008d000000ab000000a0000000b3000000a9000000920000008c0000009d",
            INIT_27 => X"0000007d000000760000007b000000740000007700000075000000680000005f",
            INIT_28 => X"000000ba000000b8000000b8000000ae000000b10000009f0000007000000086",
            INIT_29 => X"000000bb000000a70000009e0000009b000000b0000000bf000000c2000000ba",
            INIT_2A => X"0000007c0000009b0000009c000000a0000000970000008600000093000000ae",
            INIT_2B => X"0000007f0000007b000000750000006b0000006600000069000000660000004a",
            INIT_2C => X"000000be000000bf000000b1000000930000009d000000ae0000005b00000041",
            INIT_2D => X"000000a300000094000000ae000000b8000000b0000000ac000000b0000000bc",
            INIT_2E => X"0000005000000083000000950000009800000095000000850000009a000000b0",
            INIT_2F => X"0000007d00000078000000710000006700000066000000670000006100000042",
            INIT_30 => X"000000b6000000bd000000ca000000bc000000b1000000bf0000005c00000015",
            INIT_31 => X"0000007200000098000000ae000000c8000000bc000000a50000009c000000b3",
            INIT_32 => X"0000004e00000072000000880000009700000089000000780000007f0000005f",
            INIT_33 => X"0000007600000075000000710000006200000062000000590000004900000040",
            INIT_34 => X"000000bb000000bc000000c3000000c8000000ad000000a8000000630000002c",
            INIT_35 => X"0000009a000000a8000000a8000000b9000000c2000000b400000095000000a5",
            INIT_36 => X"00000048000000640000007f0000009c0000008a00000091000000920000006b",
            INIT_37 => X"0000006f0000006c0000006a0000006200000060000000530000004000000039",
            INIT_38 => X"000000bb000000b4000000be000000c40000009f000000750000007600000069",
            INIT_39 => X"000000bc000000b4000000a5000000ab000000c1000000c6000000ad000000ad",
            INIT_3A => X"000000480000006900000080000000a0000000b3000000ad000000bb000000ae",
            INIT_3B => X"000000660000006100000064000000630000006c000000570000004500000043",
            INIT_3C => X"000000a8000000b4000000c4000000c60000009d00000068000000710000008a",
            INIT_3D => X"000000c8000000c4000000bf000000d2000000cd000000cb000000bf000000b4",
            INIT_3E => X"000000500000007100000099000000a8000000be000000bc000000bb000000c0",
            INIT_3F => X"000000620000005a0000005a0000007800000087000000600000004000000046",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE30;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE31 : if BRAM_NAME = "sampleifmap_layer0_instance31" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000096000000b0000000bb000000be00000093000000730000008a00000096",
            INIT_01 => X"000000cb000000be000000c2000000d3000000c6000000d3000000c7000000ab",
            INIT_02 => X"0000004600000064000000a6000000be000000bd000000b8000000ba000000bf",
            INIT_03 => X"0000005e0000004a0000005c000000950000008f0000006a000000380000002f",
            INIT_04 => X"00000091000000bf000000c0000000bd000000a5000000920000009b0000009b",
            INIT_05 => X"000000a8000000b2000000c2000000c000000095000000a9000000d20000009c",
            INIT_06 => X"0000002b00000043000000750000009a000000a7000000aa000000b5000000a9",
            INIT_07 => X"000000500000003f0000006a0000009c0000008f000000680000003100000022",
            INIT_08 => X"00000089000000ba000000be000000c4000000a60000008a000000a2000000a5",
            INIT_09 => X"0000008f00000080000000b6000000d2000000a90000009d000000c900000074",
            INIT_0A => X"000000330000002f0000003800000052000000610000007f000000930000007c",
            INIT_0B => X"00000041000000390000007b0000009d0000009d00000069000000400000002b",
            INIT_0C => X"00000098000000be000000be000000be0000009e0000007800000096000000a9",
            INIT_0D => X"000000ce00000090000000a5000000c3000000b9000000bc000000990000003c",
            INIT_0E => X"000000500000004700000033000000370000003d0000006500000089000000b1",
            INIT_0F => X"00000032000000360000008e000000b0000000a00000006e0000004a00000037",
            INIT_10 => X"0000009a000000ba000000bc000000ba000000a600000096000000a0000000aa",
            INIT_11 => X"000000c00000008c0000008c0000009b000000920000007e0000003100000020",
            INIT_12 => X"000000570000005200000049000000490000003e000000610000009c000000cc",
            INIT_13 => X"0000003300000048000000a7000000bc000000a60000006b0000003e0000003a",
            INIT_14 => X"0000007c000000a3000000b2000000b50000009c00000097000000ab000000b2",
            INIT_15 => X"0000008200000065000000630000004e00000037000000280000001d00000024",
            INIT_16 => X"000000550000003c0000003300000034000000370000005f0000007b00000090",
            INIT_17 => X"0000003700000059000000b1000000bb00000099000000660000004d0000004e",
            INIT_18 => X"0000006900000095000000a7000000a90000009800000092000000ab000000b5",
            INIT_19 => X"000000780000005c000000470000002f0000002e000000420000005e0000004f",
            INIT_1A => X"000000370000001e00000022000000230000002900000038000000370000005a",
            INIT_1B => X"0000003c0000006a000000ae000000ad00000077000000610000005600000052",
            INIT_1C => X"0000008900000094000000a00000009c000000a30000009e0000009c000000b1",
            INIT_1D => X"000000670000007d0000006d0000006e0000006b00000066000000760000008f",
            INIT_1E => X"000000130000000e0000001c000000180000001300000010000000110000002f",
            INIT_1F => X"0000004300000085000000ad0000008c0000006300000060000000410000002b",
            INIT_20 => X"000000c0000000ab0000008c00000097000000b6000000a70000008b0000009e",
            INIT_21 => X"000000650000007f0000008d00000092000000880000008500000074000000ac",
            INIT_22 => X"0000000f0000000a000000110000001800000019000000200000002500000041",
            INIT_23 => X"000000690000009c00000094000000620000004e000000610000004200000014",
            INIT_24 => X"000000b100000094000000880000009e000000ab000000ae000000a4000000a0",
            INIT_25 => X"0000007d0000008e0000008b0000007f00000097000000a900000093000000b8",
            INIT_26 => X"0000001a0000001100000018000000210000002b0000003f0000004d00000067",
            INIT_27 => X"00000088000000780000005a0000004800000032000000480000003e0000001f",
            INIT_28 => X"000000780000008c000000a8000000b1000000a7000000a7000000a3000000a0",
            INIT_29 => X"00000091000000a60000009c0000007b00000082000000760000008f000000ab",
            INIT_2A => X"0000004300000038000000420000004c0000004e0000005b000000690000007c",
            INIT_2B => X"0000006a000000510000007b0000006400000049000000410000004100000046",
            INIT_2C => X"0000007b00000099000000aa000000b4000000930000008c0000009f0000009c",
            INIT_2D => X"000000a2000000a80000009e000000830000007e000000730000009c0000008b",
            INIT_2E => X"00000077000000690000006800000070000000780000007b000000770000007f",
            INIT_2F => X"000000680000005c000000860000007a0000006d000000680000006900000074",
            INIT_30 => X"0000008c0000008d0000009c000000ad0000008b0000007b0000009e000000a4",
            INIT_31 => X"000000a8000000a60000009d00000097000000a100000082000000790000008d",
            INIT_32 => X"000000940000008a0000008500000081000000840000008f0000008a00000090",
            INIT_33 => X"000000930000007300000064000000780000008400000086000000890000008f",
            INIT_34 => X"0000009e0000009e000000a1000000a7000000a800000090000000950000008e",
            INIT_35 => X"000000a20000009e000000a0000000a1000000a90000009700000090000000a5",
            INIT_36 => X"0000009e00000096000000950000008d0000007f000000890000009100000099",
            INIT_37 => X"0000009f0000008b000000770000007b0000008f00000094000000960000009f",
            INIT_38 => X"000000a8000000aa000000a7000000a7000000b9000000b3000000a600000098",
            INIT_39 => X"00000085000000890000009d000000a9000000b2000000ad000000a4000000a7",
            INIT_3A => X"0000009d00000098000000970000008c000000880000008c0000008f00000092",
            INIT_3B => X"0000009900000090000000830000008500000090000000990000009c000000a6",
            INIT_3C => X"0000009f000000910000007d0000008b000000ab000000b7000000b20000009f",
            INIT_3D => X"0000007300000083000000980000009e0000009c000000950000008b000000a2",
            INIT_3E => X"000000a10000009c0000009d000000900000008f000000940000008e00000084",
            INIT_3F => X"0000009800000099000000960000009c0000009c000000940000009f000000a7",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE31;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE32 : if BRAM_NAME = "sampleifmap_layer0_instance32" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000053000000540000005f000000600000003b000000310000006000000076",
            INIT_01 => X"0000004f0000004b000000520000005c0000005a00000053000000610000005f",
            INIT_02 => X"00000033000000380000003800000037000000320000003b000000500000005b",
            INIT_03 => X"0000002f0000002f000000350000004c0000003a00000033000000380000003c",
            INIT_04 => X"000000680000005d000000600000006c00000069000000590000005800000082",
            INIT_05 => X"000000480000004f00000057000000540000005b0000005a0000006200000065",
            INIT_06 => X"00000033000000370000003800000037000000320000003d0000004800000052",
            INIT_07 => X"000000390000003a0000003d0000004b0000004100000035000000280000002b",
            INIT_08 => X"0000006a0000005f000000590000006c0000007a000000810000006800000084",
            INIT_09 => X"0000004c0000004f00000050000000550000005e000000620000006900000062",
            INIT_0A => X"000000420000003f0000003a000000330000002a000000360000004c00000055",
            INIT_0B => X"00000039000000380000003e000000430000004200000043000000420000003c",
            INIT_0C => X"00000069000000680000005a0000007000000084000000880000007f00000081",
            INIT_0D => X"0000005d000000570000005a0000006700000066000000650000007100000065",
            INIT_0E => X"0000003e00000039000000330000002a0000001f000000330000004e0000004f",
            INIT_0F => X"0000004500000043000000370000003c0000004a0000004b0000004d00000046",
            INIT_10 => X"0000007200000072000000630000006d0000007f000000790000007f00000080",
            INIT_11 => X"0000005c00000059000000630000006c00000071000000700000006f0000006f",
            INIT_12 => X"0000002e0000003800000034000000270000002c0000004e000000590000005e",
            INIT_13 => X"00000047000000450000003b0000004200000049000000470000004300000035",
            INIT_14 => X"00000074000000710000006a000000760000007f000000680000008300000089",
            INIT_15 => X"000000540000005a000000690000006d00000071000000740000007500000073",
            INIT_16 => X"0000003d000000520000004d0000003a0000004f00000067000000680000006a",
            INIT_17 => X"0000004b00000046000000480000004900000046000000430000003f0000003e",
            INIT_18 => X"0000006f00000073000000750000007a00000087000000660000007700000098",
            INIT_19 => X"0000005c000000660000007100000073000000700000007c0000007b00000079",
            INIT_1A => X"000000430000005b000000570000005c0000006e0000006d0000006500000064",
            INIT_1B => X"0000004e0000004a00000048000000450000003b00000038000000400000003e",
            INIT_1C => X"000000790000007200000076000000780000007e000000780000005900000093",
            INIT_1D => X"000000640000006c0000006d00000073000000730000007c0000007a00000080",
            INIT_1E => X"00000048000000570000004b000000660000006a0000006d0000006800000065",
            INIT_1F => X"0000004b000000490000004400000042000000350000002e0000003c0000003b",
            INIT_20 => X"0000007700000075000000740000007700000072000000780000006f00000076",
            INIT_21 => X"0000005e0000006100000067000000730000006d0000006f0000007a00000080",
            INIT_22 => X"00000059000000720000005f0000006d0000006400000061000000590000005e",
            INIT_23 => X"0000004b00000048000000480000004600000047000000400000003a0000003e",
            INIT_24 => X"0000006f0000007b0000007a0000007c00000078000000690000007100000077",
            INIT_25 => X"0000006f000000650000006d00000076000000790000007d0000007b00000076",
            INIT_26 => X"000000670000007a000000640000006a00000060000000520000005500000069",
            INIT_27 => X"0000004b000000440000004b0000004700000049000000470000003e0000003d",
            INIT_28 => X"0000007e0000007c0000007f000000780000007e000000720000004800000064",
            INIT_29 => X"000000900000007800000077000000790000007b00000080000000810000007f",
            INIT_2A => X"0000005b0000006c000000610000005f000000580000004f0000006300000083",
            INIT_2B => X"0000004c0000004900000046000000400000003b0000003d0000003e0000002e",
            INIT_2C => X"00000083000000840000007a0000005d000000690000007f0000003400000022",
            INIT_2D => X"000000850000007400000097000000a60000008c000000780000007300000081",
            INIT_2E => X"00000031000000560000005c0000006000000061000000560000006e0000008d",
            INIT_2F => X"0000004a00000045000000420000003e0000003c0000003e0000003c0000002a",
            INIT_30 => X"000000840000008c0000009a0000008c0000007d0000008e0000004000000004",
            INIT_31 => X"000000530000007700000093000000b20000009c0000007b0000006b0000007f",
            INIT_32 => X"000000310000004d0000005c0000006f00000064000000530000005b00000040",
            INIT_33 => X"0000004400000042000000430000003b00000039000000370000002f00000029",
            INIT_34 => X"0000008d0000008f000000960000009c0000007b0000007a0000004800000018",
            INIT_35 => X"00000077000000800000008100000097000000a00000008f0000006a00000077",
            INIT_36 => X"0000002d000000440000005a0000007b0000006d00000073000000740000004d",
            INIT_37 => X"0000003e0000003a0000003e0000003b00000037000000330000002b00000023",
            INIT_38 => X"0000008f000000860000009100000096000000700000004a0000005200000045",
            INIT_39 => X"0000009700000085000000720000007d0000009c000000a10000008400000083",
            INIT_3A => X"0000002f0000004b0000005d000000810000009800000092000000a000000091",
            INIT_3B => X"00000039000000360000003c0000003c0000004400000038000000300000002f",
            INIT_3C => X"0000007d000000860000009600000098000000700000003b0000004100000057",
            INIT_3D => X"000000a00000008f000000840000009b000000a5000000a70000009b0000008f",
            INIT_3E => X"00000039000000540000007800000089000000a10000009f0000009e000000a2",
            INIT_3F => X"000000390000003600000037000000510000005f000000400000002b00000033",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE32;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE33 : if BRAM_NAME = "sampleifmap_layer0_instance33" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000006c000000810000008d0000009000000066000000400000004e00000058",
            INIT_01 => X"0000009f00000086000000860000009e0000009d000000af000000a50000008b",
            INIT_02 => X"0000003100000049000000870000009a0000009800000093000000940000009a",
            INIT_03 => X"000000390000002c0000003d0000006f000000670000004b000000230000001e",
            INIT_04 => X"0000006900000091000000930000008f00000074000000570000005700000056",
            INIT_05 => X"000000790000007a0000008b000000910000006c00000085000000b300000080",
            INIT_06 => X"000000180000002a0000005800000072000000790000007c000000870000007d",
            INIT_07 => X"0000002e00000027000000500000007500000066000000490000001d00000013",
            INIT_08 => X"0000006200000091000000990000009c000000760000004d0000005c0000005c",
            INIT_09 => X"000000620000004b00000083000000a50000007a00000074000000aa0000005c",
            INIT_0A => X"0000001b000000110000001b000000360000004000000055000000610000004c",
            INIT_0B => X"0000002800000024000000640000007f0000007500000045000000280000001a",
            INIT_0C => X"000000730000009b000000a30000009c0000006e0000003c000000540000005e",
            INIT_0D => X"0000009c00000057000000710000009500000089000000940000007c00000027",
            INIT_0E => X"0000002e000000220000001800000027000000270000003d0000005000000078",
            INIT_0F => X"00000020000000220000007b0000009900000078000000450000002d0000001f",
            INIT_10 => X"0000007500000098000000a20000009600000072000000590000005d00000061",
            INIT_11 => X"0000007c00000049000000560000007300000074000000640000001d0000000d",
            INIT_12 => X"000000320000003100000032000000310000001b0000002f0000005b00000086",
            INIT_13 => X"000000200000003800000096000000a20000007d000000420000001e00000019",
            INIT_14 => X"0000005700000081000000960000008d0000006300000057000000680000006a",
            INIT_15 => X"0000003e00000029000000390000003600000025000000160000000b0000000f",
            INIT_16 => X"000000330000002200000023000000200000001a000000360000004800000053",
            INIT_17 => X"0000001f0000004a0000009e0000009b000000700000003e0000002b00000028",
            INIT_18 => X"0000004200000073000000890000007b0000005a0000004f0000006800000070",
            INIT_19 => X"000000450000002c000000260000001b0000001700000028000000420000002f",
            INIT_1A => X"0000001f0000000f00000016000000190000001d000000260000001f00000036",
            INIT_1B => X"0000001f0000005700000094000000860000004e0000003a0000003300000031",
            INIT_1C => X"0000005e0000007300000081000000690000006000000059000000580000006d",
            INIT_1D => X"0000003c0000004b0000003e000000420000003c000000360000004700000061",
            INIT_1E => X"0000000c0000000b00000013000000110000000e000000090000000a0000001a",
            INIT_1F => X"0000002300000069000000880000005e0000003b0000003a0000001f00000017",
            INIT_20 => X"000000930000008900000068000000600000007000000060000000460000005b",
            INIT_21 => X"000000350000003f000000450000004a00000043000000450000003a00000075",
            INIT_22 => X"000000120000000d000000090000000c0000000d000000130000001900000029",
            INIT_23 => X"00000047000000790000006800000034000000270000003e000000240000000c",
            INIT_24 => X"0000008600000069000000560000006100000062000000620000005c0000005b",
            INIT_25 => X"000000490000004e0000004900000044000000610000007c0000006b0000008e",
            INIT_26 => X"000000140000000b0000000e000000160000001c000000260000002b0000003e",
            INIT_27 => X"0000006400000058000000380000002500000014000000300000002a00000014",
            INIT_28 => X"0000004c0000005b0000006f0000007100000062000000610000005e0000005b",
            INIT_29 => X"00000054000000630000005f0000004700000051000000500000006e00000084",
            INIT_2A => X"0000002b000000200000002b0000003500000033000000380000003d00000048",
            INIT_2B => X"00000042000000300000005a000000400000002800000025000000280000002e",
            INIT_2C => X"00000048000000620000006d0000007100000052000000500000006000000057",
            INIT_2D => X"00000058000000600000005e0000004a0000004600000045000000730000005c",
            INIT_2E => X"0000004b0000003d0000003c000000420000004a0000004c0000004700000045",
            INIT_2F => X"0000003a000000360000005e0000004c000000410000003f0000004000000049",
            INIT_30 => X"000000500000004e0000005a000000690000004c000000430000006100000060",
            INIT_31 => X"0000005a0000005d0000005c00000057000000620000004c0000004800000057",
            INIT_32 => X"000000570000004d00000048000000420000004600000055000000540000004f",
            INIT_33 => X"0000005e0000004600000035000000430000004f000000500000005200000053",
            INIT_34 => X"0000005b000000580000005b0000006100000065000000510000005400000049",
            INIT_35 => X"0000005a0000005d0000005d00000059000000630000005b0000005900000069",
            INIT_36 => X"0000005b0000005400000052000000490000003c000000490000005500000058",
            INIT_37 => X"000000640000005700000044000000430000005500000057000000560000005d",
            INIT_38 => X"0000005f000000600000005f00000060000000710000006a0000006000000053",
            INIT_39 => X"0000004a000000520000005a0000005b000000680000006d0000006900000066",
            INIT_3A => X"0000005c00000057000000550000004d0000004a0000004d0000004e00000052",
            INIT_3B => X"0000005a000000570000004d0000004e000000540000005a0000005900000064",
            INIT_3C => X"0000005c0000004d000000420000005200000068000000710000006b0000005c",
            INIT_3D => X"0000003d0000004d0000005b000000580000005a0000005b000000510000005f",
            INIT_3E => X"000000600000005b0000005c0000005300000052000000560000004d00000046",
            INIT_3F => X"000000570000005b0000005a0000005c0000005b000000570000005c00000065",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE33;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE34 : if BRAM_NAME = "sampleifmap_layer0_instance34" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000360000003a0000004300000041000000240000001a0000003d00000053",
            INIT_01 => X"000000340000002e000000350000003e0000003b00000034000000410000003f",
            INIT_02 => X"000000260000002d0000002f0000002f000000270000002b0000004100000047",
            INIT_03 => X"00000029000000290000002e00000045000000320000002a0000002d0000002f",
            INIT_04 => X"0000004d000000440000004300000046000000460000003a0000003500000061",
            INIT_05 => X"0000002e00000032000000390000003400000039000000380000004100000044",
            INIT_06 => X"000000280000002c0000002f0000002f000000260000002b000000340000003c",
            INIT_07 => X"00000031000000330000003500000043000000380000002b0000001e00000020",
            INIT_08 => X"0000004e000000440000003900000044000000510000005c0000004700000064",
            INIT_09 => X"000000300000003100000030000000340000003b0000003f0000004700000040",
            INIT_0A => X"0000003800000035000000300000002b0000001e00000021000000320000003b",
            INIT_0B => X"000000310000002f000000350000003900000038000000390000003800000033",
            INIT_0C => X"0000004800000049000000370000004900000059000000610000005f00000060",
            INIT_0D => X"0000003f00000036000000370000004300000042000000420000004e00000041",
            INIT_0E => X"000000350000002f0000002900000022000000120000001a0000002e0000002f",
            INIT_0F => X"0000003c0000003a0000002d000000300000003e00000040000000440000003d",
            INIT_10 => X"0000004b0000004c0000003f000000490000005700000054000000610000005c",
            INIT_11 => X"0000003b000000350000003b000000430000004b0000004b0000004a0000004a",
            INIT_12 => X"000000270000002e000000290000001f0000001e00000033000000340000003b",
            INIT_13 => X"0000003c0000003a00000030000000340000003d0000003d0000003b0000002e",
            INIT_14 => X"0000004c0000004c000000460000005100000059000000470000006600000065",
            INIT_15 => X"00000031000000350000004300000044000000470000004e000000510000004c",
            INIT_16 => X"00000032000000420000003e0000002b00000039000000480000004100000043",
            INIT_17 => X"000000410000003c0000003d0000003c0000003a000000380000003600000038",
            INIT_18 => X"0000004b00000051000000500000005300000063000000490000005900000078",
            INIT_19 => X"00000035000000430000004f0000004c00000042000000550000005700000051",
            INIT_1A => X"0000002f0000004100000040000000410000004d0000004a000000400000003c",
            INIT_1B => X"000000420000003f0000003d0000003a000000300000002d0000003600000035",
            INIT_1C => X"000000540000004f00000051000000510000005b0000005b0000003b00000075",
            INIT_1D => X"0000003f0000004a0000004c0000004d00000048000000560000005600000057",
            INIT_1E => X"0000002f000000380000002f00000047000000490000004c0000004900000042",
            INIT_1F => X"000000400000003e00000039000000370000002a00000023000000310000002c",
            INIT_20 => X"00000050000000500000004f00000053000000510000005b000000540000005c",
            INIT_21 => X"0000003d00000043000000480000005100000046000000490000005300000058",
            INIT_22 => X"0000003c0000004f000000400000004f00000046000000460000004100000043",
            INIT_23 => X"000000400000003d0000003d0000003a0000003b000000340000002d0000002c",
            INIT_24 => X"0000004700000053000000560000005b0000005a0000004c0000005800000061",
            INIT_25 => X"000000550000004d00000053000000580000005300000054000000520000004f",
            INIT_26 => X"0000004b00000059000000480000005000000046000000390000003e00000051",
            INIT_27 => X"00000040000000390000003f0000003a0000003c0000003a000000310000002b",
            INIT_28 => X"00000054000000520000005b0000005900000062000000560000003000000051",
            INIT_29 => X"0000007e00000067000000650000005e0000005000000050000000540000005b",
            INIT_2A => X"00000044000000510000004c0000004b0000004300000037000000490000006b",
            INIT_2B => X"000000410000003e0000003a000000330000002d0000002f0000003100000020",
            INIT_2C => X"0000005a0000005a00000056000000400000004d000000630000001f00000014",
            INIT_2D => X"0000007900000067000000880000008f0000005f00000045000000450000005f",
            INIT_2E => X"00000021000000420000004d00000052000000500000003f0000005200000076",
            INIT_2F => X"0000003f0000003b00000036000000300000002e000000300000003000000021",
            INIT_30 => X"00000062000000690000007a0000006e0000005c000000700000003200000000",
            INIT_31 => X"000000490000005f0000007d0000009d00000077000000540000004800000060",
            INIT_32 => X"0000002a000000410000004f0000006000000054000000410000004700000034",
            INIT_33 => X"0000003a00000039000000380000002d00000029000000290000002500000025",
            INIT_34 => X"0000006f00000070000000780000007d0000005c000000610000003c00000014",
            INIT_35 => X"0000006c00000062000000640000007f000000800000006e0000004c00000059",
            INIT_36 => X"000000290000003a0000004c0000006a0000005b000000620000006300000044",
            INIT_37 => X"0000003500000032000000340000002e00000026000000250000002300000021",
            INIT_38 => X"000000730000006a000000750000007b000000580000003a000000460000003b",
            INIT_39 => X"0000008900000066000000500000005f0000007d000000820000006700000066",
            INIT_3A => X"0000002a000000400000004e0000006f000000840000007e0000008c00000083",
            INIT_3B => X"000000310000002e000000320000002f000000320000002a000000280000002b",
            INIT_3C => X"000000620000006c0000007c0000007e0000005e000000320000003500000049",
            INIT_3D => X"0000008c00000071000000620000007b000000880000008a0000007d00000072",
            INIT_3E => X"000000330000004900000069000000750000008c0000008a000000890000008f",
            INIT_3F => X"000000320000002d0000002d000000430000004d00000032000000230000002f",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE34;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE35 : if BRAM_NAME = "sampleifmap_layer0_instance35" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000053000000690000007500000077000000560000003a0000004100000048",
            INIT_01 => X"000000870000006d0000006b000000820000008200000093000000890000006e",
            INIT_02 => X"0000002a0000003d0000007700000087000000830000007e0000007f00000084",
            INIT_03 => X"00000033000000240000003300000061000000550000003c0000001b0000001a",
            INIT_04 => X"000000500000007a0000007c0000007800000066000000510000004800000047",
            INIT_05 => X"0000005c00000065000000790000007c000000540000006a0000009700000063",
            INIT_06 => X"000000110000001f000000480000005e00000065000000680000007300000063",
            INIT_07 => X"000000290000001f0000004600000068000000550000003a000000150000000e",
            INIT_08 => X"0000004b0000007d000000880000008600000064000000440000004e0000004f",
            INIT_09 => X"0000004800000037000000710000008e000000610000005b0000009300000047",
            INIT_0A => X"000000160000000d000000140000002a00000032000000450000004f00000035",
            INIT_0B => X"000000230000001e0000005b0000006f00000060000000370000002300000014",
            INIT_0C => X"0000005d0000008a000000990000008700000058000000320000004800000051",
            INIT_0D => X"0000008d000000470000005c0000007c000000710000007f0000006f0000001f",
            INIT_0E => X"0000002c00000024000000190000002400000021000000330000004100000067",
            INIT_0F => X"0000001a0000001e000000730000008900000060000000360000002b0000001a",
            INIT_10 => X"000000620000008600000096000000820000005f0000004f0000005200000053",
            INIT_11 => X"00000074000000420000004c000000650000006300000056000000170000000a",
            INIT_12 => X"0000002e0000002f0000002f0000002e00000017000000270000004e0000007a",
            INIT_13 => X"000000190000002f000000890000009200000067000000340000001b00000014",
            INIT_14 => X"000000460000006e000000870000007b000000530000004e0000005c0000005c",
            INIT_15 => X"0000003800000025000000340000002f0000001d00000010000000080000000c",
            INIT_16 => X"0000002c0000001d0000001c00000019000000120000002b0000003900000046",
            INIT_17 => X"000000180000003d0000008d0000008c0000005e000000310000002600000021",
            INIT_18 => X"0000003000000060000000760000006b0000004e000000460000005d00000061",
            INIT_19 => X"0000003b000000260000001f0000001300000013000000220000003a00000025",
            INIT_1A => X"000000180000000a0000001100000011000000120000001b0000001300000027",
            INIT_1B => X"0000001800000046000000800000007800000040000000300000002c0000002a",
            INIT_1C => X"0000004b0000005f0000006b0000005b00000058000000520000004d0000005e",
            INIT_1D => X"0000003300000043000000350000003a0000003900000030000000370000004a",
            INIT_1E => X"0000000600000007000000130000000e00000008000000030000000400000010",
            INIT_1F => X"0000001b0000005700000073000000510000002f000000300000001700000011",
            INIT_20 => X"0000007e00000075000000520000005300000069000000570000003b0000004b",
            INIT_21 => X"0000002e000000390000003d000000420000003e000000390000002200000055",
            INIT_22 => X"0000000e0000000c0000000e0000000f0000000d000000120000001700000024",
            INIT_23 => X"0000003e0000006800000055000000280000001e000000360000001c00000007",
            INIT_24 => X"0000007000000057000000450000005500000056000000510000004d0000004d",
            INIT_25 => X"0000003a00000045000000430000003b0000004f000000640000004f0000006f",
            INIT_26 => X"0000000e000000060000000c0000001100000015000000200000002600000033",
            INIT_27 => X"0000005a0000004c0000002e0000001f0000000f00000029000000220000000f",
            INIT_28 => X"000000390000004a00000060000000650000005500000052000000510000004f",
            INIT_29 => X"000000440000005a000000580000003d0000003e0000003a000000570000006d",
            INIT_2A => X"0000002300000018000000230000002c0000002a0000002f000000350000003b",
            INIT_2B => X"000000380000002700000052000000390000001f0000001b0000001d00000026",
            INIT_2C => X"00000039000000530000005f000000660000004a0000004a000000570000004c",
            INIT_2D => X"0000004d00000057000000540000003f0000003a00000037000000630000004d",
            INIT_2E => X"0000003f00000031000000310000003b00000044000000430000003c00000039",
            INIT_2F => X"0000002f0000002d000000540000003f0000003300000030000000310000003c",
            INIT_30 => X"00000044000000410000004e0000005e00000045000000400000005a00000055",
            INIT_31 => X"00000051000000530000004e0000004a0000005a000000420000003c0000004c",
            INIT_32 => X"000000480000003e000000390000003b000000400000004c0000004700000043",
            INIT_33 => X"000000530000003d00000029000000320000003e000000400000004200000044",
            INIT_34 => X"000000500000004e00000051000000570000005c000000490000004b0000003d",
            INIT_35 => X"000000500000004e0000004c0000004a00000059000000500000004c0000005d",
            INIT_36 => X"0000004b000000440000004200000040000000350000003e000000450000004a",
            INIT_37 => X"000000590000004e00000038000000320000004400000048000000480000004d",
            INIT_38 => X"00000055000000570000005500000056000000640000005a0000005100000046",
            INIT_39 => X"0000003c0000003f000000460000004a0000005a0000005d0000005700000056",
            INIT_3A => X"0000004c0000004700000046000000410000003e0000003e0000003c00000042",
            INIT_3B => X"0000004f0000004d000000410000003e000000470000004e0000004d00000055",
            INIT_3C => X"00000051000000460000003900000046000000590000005f0000005d0000004f",
            INIT_3D => X"0000002f0000003d0000004c0000004a00000047000000470000004000000053",
            INIT_3E => X"000000500000004b0000004c0000004500000046000000480000003f00000038",
            INIT_3F => X"000000490000004f0000004c0000004f0000004e000000490000004f00000056",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE35;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE36 : if BRAM_NAME = "sampleifmap_layer0_instance36" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000f6000000f9000000f6000000e6000000d9000000d1000000b9000000a0",
            INIT_01 => X"000000c7000000d8000000dd000000da000000dd000000e6000000f3000000f8",
            INIT_02 => X"0000008b0000007900000090000000a6000000b4000000b8000000bb000000bc",
            INIT_03 => X"0000005e0000005b000000650000005e0000004f00000066000000660000006a",
            INIT_04 => X"000000eb000000f3000000f5000000e8000000e6000000f2000000ef000000e1",
            INIT_05 => X"000000ba000000c8000000cb000000c9000000cd000000d8000000e6000000ed",
            INIT_06 => X"000000870000007a0000008d0000008e0000007f000000a1000000ab000000af",
            INIT_07 => X"00000064000000610000006b0000005f00000034000000250000005200000076",
            INIT_08 => X"000000d6000000df000000e2000000d9000000dc000000f1000000f9000000fc",
            INIT_09 => X"000000a7000000b3000000b6000000b3000000b8000000c3000000cf000000d5",
            INIT_0A => X"00000072000000800000008c000000800000008100000094000000980000009f",
            INIT_0B => X"0000006900000069000000730000006300000026000000040000002800000057",
            INIT_0C => X"000000c0000000c8000000cb000000d3000000d3000000de000000e1000000e9",
            INIT_0D => X"00000099000000a0000000a5000000a0000000a4000000ae000000b7000000bb",
            INIT_0E => X"000000690000007f0000007d0000007d0000008a0000008c0000008d00000091",
            INIT_0F => X"0000006d000000700000007800000070000000370000001a000000250000003b",
            INIT_10 => X"000000ab000000b3000000b4000000be000000c9000000cf000000c3000000cf",
            INIT_11 => X"0000008d00000093000000970000009100000092000000990000009f000000a3",
            INIT_12 => X"0000005a000000840000007a0000008100000087000000830000008800000087",
            INIT_13 => X"0000006d00000072000000780000007500000056000000300000003d0000003a",
            INIT_14 => X"000000970000009f0000009c00000099000000a2000000aa000000ab000000b6",
            INIT_15 => X"0000008a0000008a0000008d0000008b0000008a0000008c0000008d00000090",
            INIT_16 => X"0000004500000066000000890000008c0000008a000000860000008c00000087",
            INIT_17 => X"0000006e00000070000000800000008100000074000000430000003e0000004b",
            INIT_18 => X"000000850000008c00000086000000880000008600000088000000880000008d",
            INIT_19 => X"000000910000008e000000920000008f0000008d0000008b0000008900000087",
            INIT_1A => X"000000210000002f0000006b0000008e0000008f0000008a0000009100000091",
            INIT_1B => X"000000700000006f00000084000000840000007f0000006c0000004b00000048",
            INIT_1C => X"000000840000008a000000830000008800000081000000800000007d00000076",
            INIT_1D => X"000000990000009a0000009e0000009600000093000000900000008c00000088",
            INIT_1E => X"000000110000000d000000420000008000000094000000930000009500000092",
            INIT_1F => X"0000007000000072000000800000007b0000007a000000800000007500000050",
            INIT_20 => X"000000890000008f000000870000008b00000085000000840000007e00000073",
            INIT_21 => X"000000aa000000a30000009a000000940000009800000095000000910000008b",
            INIT_22 => X"0000001e0000000e0000002c00000073000000940000009d000000a20000009e",
            INIT_23 => X"0000006f000000740000007a000000770000007e000000880000008b00000069",
            INIT_24 => X"0000008d00000091000000880000008d00000088000000880000008000000076",
            INIT_25 => X"000000a7000000a20000009a0000009d000000a50000009a000000930000008d",
            INIT_26 => X"000000370000002e00000038000000630000008a00000091000000930000009b",
            INIT_27 => X"0000006e0000007500000074000000730000007e0000007a0000007c0000006d",
            INIT_28 => X"0000008c00000090000000880000008e000000890000008b000000840000007d",
            INIT_29 => X"00000098000000900000008b000000830000009900000096000000900000008b",
            INIT_2A => X"0000002a000000450000005c00000080000000d6000000d3000000ba000000a6",
            INIT_2B => X"0000006b000000710000006f0000007000000073000000630000005f00000055",
            INIT_2C => X"0000008a0000008e000000880000008d0000008a0000008e0000008900000085",
            INIT_2D => X"000000cb000000c9000000b60000008e00000084000000880000008f00000089",
            INIT_2E => X"0000002a00000092000000bd000000a2000000c0000000cf000000ce000000d2",
            INIT_2F => X"000000680000006c0000006a0000006d0000007200000067000000280000001b",
            INIT_30 => X"000000890000008a0000008c0000008f0000008b0000008f0000008b0000008c",
            INIT_31 => X"0000007300000089000000a0000000ab000000a4000000900000008500000087",
            INIT_32 => X"0000005f000000c9000000dc0000006f0000003b0000004b0000005d0000006a",
            INIT_33 => X"00000064000000690000006500000063000000740000003e000000070000000d",
            INIT_34 => X"000000870000008200000092000000920000008c0000008f0000008a00000090",
            INIT_35 => X"00000013000000310000005c0000005e0000006e0000008c0000009100000082",
            INIT_36 => X"0000009d000000d2000000d1000000780000001200000019000000320000001d",
            INIT_37 => X"0000005f00000063000000520000004500000044000000130000000600000026",
            INIT_38 => X"00000080000000790000008e000000900000008e000000920000008b00000091",
            INIT_39 => X"000000160000002e000000520000005600000044000000540000007f00000085",
            INIT_3A => X"000000cb000000cd000000c9000000af000000410000001e0000003200000013",
            INIT_3B => X"000000580000004f000000380000002300000016000000120000001000000066",
            INIT_3C => X"000000830000008b000000840000008a00000090000000940000008b0000008f",
            INIT_3D => X"00000022000000280000004e0000006a00000056000000480000004200000075",
            INIT_3E => X"000000c3000000cd000000c5000000cb000000b6000000730000004600000024",
            INIT_3F => X"00000053000000640000004f0000001800000012000000250000003d0000006c",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE36;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE37 : if BRAM_NAME = "sampleifmap_layer0_instance37" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000007900000084000000720000008500000090000000930000008b0000008e",
            INIT_01 => X"0000009b000000530000004400000055000000450000003c0000005900000051",
            INIT_02 => X"00000072000000d3000000d7000000d7000000eb000000ed000000db000000c0",
            INIT_03 => X"000000540000008f0000008b0000004100000014000000350000005d00000030",
            INIT_04 => X"000000430000003a0000004500000074000000890000008e0000008d0000008f",
            INIT_05 => X"000000f20000008c00000019000000240000001c0000001d0000004b00000051",
            INIT_06 => X"0000003a00000095000000df000000db000000dc000000e3000000eb000000ec",
            INIT_07 => X"0000005b000000a7000000a1000000850000004e0000004e0000005400000039",
            INIT_08 => X"000000340000002d000000470000008d00000086000000880000008c0000008f",
            INIT_09 => X"000000d90000009b000000290000002f00000016000000170000002100000043",
            INIT_0A => X"00000067000000ad000000df000000dc000000d0000000bf000000be000000c7",
            INIT_0B => X"00000059000000a500000094000000980000009500000087000000730000005d",
            INIT_0C => X"0000002b000000210000004c000000bd000000b50000007e0000008c0000008f",
            INIT_0D => X"000000c20000009e000000420000003900000017000000100000001500000039",
            INIT_0E => X"000000b3000000de000000ce000000c2000000c9000000c4000000b3000000b6",
            INIT_0F => X"0000004200000088000000920000009600000097000000950000009c00000097",
            INIT_10 => X"0000002a000000260000005a000000b5000000ea0000009a000000850000008c",
            INIT_11 => X"000000ba000000a000000031000000140000000b0000000b0000000b00000034",
            INIT_12 => X"000000c4000000a10000005a0000004500000073000000b9000000b9000000b0",
            INIT_13 => X"000000260000004d000000880000009300000099000000a0000000aa000000b7",
            INIT_14 => X"0000002e0000002d0000006a0000008b000000a3000000a30000008000000082",
            INIT_15 => X"000000b4000000a2000000360000001e0000000f00000009000000030000001c",
            INIT_16 => X"000000950000003000000015000000140000001500000071000000be000000ac",
            INIT_17 => X"00000027000000150000004300000080000000850000008e000000ab000000bb",
            INIT_18 => X"00000030000000340000006c000000480000001a00000067000000840000007c",
            INIT_19 => X"000000b0000000a5000000630000005a0000003b0000000b0000000700000012",
            INIT_1A => X"000000460000000e000000260000002f0000001d0000002a000000a9000000b1",
            INIT_1B => X"00000030000000150000000e0000003c00000075000000750000008800000095",
            INIT_1C => X"0000001f00000044000000720000003b0000001e000000490000007c00000079",
            INIT_1D => X"000000bb000000bb0000006c0000004f00000048000000180000000e0000000d",
            INIT_1E => X"0000001b0000001c0000001b0000001e0000002b0000001b0000008b000000bf",
            INIT_1F => X"0000003b0000002a0000001500000016000000590000007b000000840000006c",
            INIT_20 => X"0000001c0000004d000000710000003c0000003f00000047000000660000006d",
            INIT_21 => X"000000b3000000bd000000880000004600000047000000300000001f00000010",
            INIT_22 => X"0000000e0000001b0000002900000035000000360000001f00000074000000b4",
            INIT_23 => X"0000003b0000003200000022000000120000003c0000007c0000008500000048",
            INIT_24 => X"000000150000004b000000690000003a0000003c0000003d0000005100000057",
            INIT_25 => X"000000a3000000a40000009100000061000000600000004c0000002e00000014",
            INIT_26 => X"00000011000000250000003100000047000000390000002000000071000000aa",
            INIT_27 => X"00000032000000280000001d0000000c00000021000000600000006c00000029",
            INIT_28 => X"0000002f000000570000005f000000390000003c000000400000004900000049",
            INIT_29 => X"000000b6000000b7000000b0000000a9000000a500000089000000620000003d",
            INIT_2A => X"0000001b000000330000005c0000006000000036000000220000007c000000b6",
            INIT_2B => X"000000280000001d00000012000000060000000c0000003b0000004600000011",
            INIT_2C => X"0000002f0000004500000059000000410000004e000000450000004900000049",
            INIT_2D => X"0000006000000062000000600000005b000000560000004a0000003c00000034",
            INIT_2E => X"000000140000001d0000003e0000003b0000003c000000200000005300000062",
            INIT_2F => X"00000021000000110000000a00000007000000030000000a0000001100000004",
            INIT_30 => X"000000040000000f000000270000002d0000003600000048000000530000004b",
            INIT_31 => X"0000000b0000000a000000080000000700000007000000050000000200000003",
            INIT_32 => X"0000000f000000380000002f0000004300000042000000080000000d0000000b",
            INIT_33 => X"000000200000000f0000000a0000000600000003000000010000000200000002",
            INIT_34 => X"00000019000000100000000a000000150000002f000000510000005900000050",
            INIT_35 => X"0000000c0000000e0000000e0000000e0000000e0000000e0000000a0000000e",
            INIT_36 => X"000000070000002a000000480000003e0000001700000006000000090000000a",
            INIT_37 => X"00000021000000150000000b0000000700000005000000050000000400000003",
            INIT_38 => X"0000003a0000003b0000002f0000002e00000037000000490000004f00000049",
            INIT_39 => X"0000001c0000001d000000200000001f0000001c00000019000000110000001a",
            INIT_3A => X"000000060000000800000016000000140000000c000000100000001500000018",
            INIT_3B => X"0000001f0000001b0000000f0000000b00000008000000080000000700000008",
            INIT_3C => X"000000380000004800000053000000580000004e0000004c0000004800000045",
            INIT_3D => X"0000003100000032000000330000002f0000002a0000002b0000002600000020",
            INIT_3E => X"0000000c0000001300000022000000220000001c0000001e000000260000002c",
            INIT_3F => X"0000001d0000001e0000001a000000120000000d0000000f000000100000000e",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE37;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE38 : if BRAM_NAME = "sampleifmap_layer0_instance38" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000051000000500000004e000000420000003a000000390000003100000025",
            INIT_01 => X"0000003800000043000000430000004100000042000000490000005200000056",
            INIT_02 => X"0000002700000032000000380000003400000073000000400000003200000032",
            INIT_03 => X"0000001300000015000000120000001d000000240000002e0000002200000016",
            INIT_04 => X"00000042000000480000004a00000043000000440000004d0000004800000043",
            INIT_05 => X"0000002e00000037000000360000003200000034000000390000004000000044",
            INIT_06 => X"000000210000001e000000230000002800000029000000270000002a00000029",
            INIT_07 => X"0000001200000016000000150000001c0000001b0000001e0000002e00000022",
            INIT_08 => X"00000031000000380000003d0000003a0000003e000000480000004400000048",
            INIT_09 => X"000000260000002b0000002a00000026000000280000002b0000002d00000030",
            INIT_0A => X"000000220000001f00000021000000230000001c0000001e0000002300000022",
            INIT_0B => X"000000110000001300000014000000150000000e0000000d0000002200000030",
            INIT_0C => X"000000240000002b000000300000003e0000003c0000003d0000003600000038",
            INIT_0D => X"0000002000000022000000210000001f00000020000000220000002300000023",
            INIT_0E => X"000000250000001d0000001c000000200000001d0000001b0000001e0000001d",
            INIT_0F => X"000000110000001000000013000000160000000f0000000b000000120000002a",
            INIT_10 => X"0000001b0000002000000024000000340000003b000000420000003900000039",
            INIT_11 => X"0000001e0000001c0000001a0000001a0000001a0000001c0000001d0000001c",
            INIT_12 => X"0000002a00000043000000300000001c0000001c0000001c0000001c0000001c",
            INIT_13 => X"00000011000000130000001f0000001b000000190000000d0000001200000019",
            INIT_14 => X"00000016000000190000001a0000001a000000210000002f0000003a0000003b",
            INIT_15 => X"0000001f0000001b0000001800000018000000190000001a0000001900000017",
            INIT_16 => X"0000003c0000005e0000005d000000210000001e000000210000001e0000001d",
            INIT_17 => X"00000013000000180000002d0000002b0000002c0000001e0000001b00000029",
            INIT_18 => X"0000001500000016000000170000001600000014000000170000001c00000022",
            INIT_19 => X"000000230000001d00000019000000180000001a000000190000001600000016",
            INIT_1A => X"000000250000003700000059000000330000001e000000230000001f00000020",
            INIT_1B => X"00000015000000170000001e000000240000002d0000002b0000002800000038",
            INIT_1C => X"0000001600000016000000170000001600000012000000100000001100000011",
            INIT_1D => X"000000270000001d0000001b000000190000001b0000001a0000001700000018",
            INIT_1E => X"0000000b00000012000000400000004100000030000000330000002d00000028",
            INIT_1F => X"00000015000000160000001600000019000000200000001f0000002500000022",
            INIT_20 => X"0000001700000017000000160000001500000012000000120000001200000011",
            INIT_21 => X"0000003b0000003300000038000000250000001e0000001c0000001800000019",
            INIT_22 => X"0000001000000011000000280000003d00000036000000370000003a0000003b",
            INIT_23 => X"0000001400000015000000170000001a0000001b00000018000000190000001a",
            INIT_24 => X"0000001800000016000000140000001500000012000000120000001200000013",
            INIT_25 => X"00000034000000390000004c0000003e00000031000000200000001900000018",
            INIT_26 => X"0000002c0000003000000031000000380000003a000000320000002e00000031",
            INIT_27 => X"0000001400000014000000180000001900000019000000190000002300000029",
            INIT_28 => X"0000001700000015000000150000001500000012000000130000001200000014",
            INIT_29 => X"0000004a0000003e000000420000003100000035000000240000001900000019",
            INIT_2A => X"000000210000004b000000680000007c000000b8000000a60000008900000068",
            INIT_2B => X"0000001300000012000000190000001800000019000000260000003d00000038",
            INIT_2C => X"0000001800000016000000180000001800000013000000140000001200000015",
            INIT_2D => X"000000be000000b20000009700000055000000300000001f0000001d00000019",
            INIT_2E => X"0000001600000098000000d0000000b2000000c5000000ca000000cd000000cd",
            INIT_2F => X"0000001100000011000000160000001500000028000000460000002500000018",
            INIT_30 => X"0000001a00000019000000180000001800000015000000160000001400000014",
            INIT_31 => X"000000750000008c0000009b0000009000000070000000420000002000000019",
            INIT_32 => X"0000004e000000d5000000e8000000750000003d000000470000005800000064",
            INIT_33 => X"0000001000000011000000150000001a00000046000000320000000a0000000f",
            INIT_34 => X"0000001a00000019000000170000001700000016000000190000001600000014",
            INIT_35 => X"000000120000003400000056000000500000005b00000067000000480000001a",
            INIT_36 => X"0000009b000000e0000000dd0000007c000000100000000f0000002200000011",
            INIT_37 => X"000000100000001200000013000000210000003b000000160000000700000024",
            INIT_38 => X"00000015000000130000001900000018000000160000001b0000001700000018",
            INIT_39 => X"00000018000000320000004e0000003d000000290000003a0000005500000037",
            INIT_3A => X"000000cd000000d1000000d8000000bf000000490000001e0000002b0000000b",
            INIT_3B => X"0000001200000014000000160000001b00000017000000100000000e00000067",
            INIT_3C => X"000000340000003c0000002500000019000000170000001a000000160000001a",
            INIT_3D => X"000000260000002e0000004d000000500000003b00000038000000340000004c",
            INIT_3E => X"000000d2000000d9000000d8000000df000000c40000007c0000004900000023",
            INIT_3F => X"000000110000003e000000470000001f0000000e000000150000003900000076",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE38;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE39 : if BRAM_NAME = "sampleifmap_layer0_instance39" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000005c00000060000000350000002100000017000000190000001400000019",
            INIT_01 => X"000000a20000005a0000004700000051000000420000003e0000005d00000049",
            INIT_02 => X"00000079000000de000000e4000000e3000000f5000000f5000000df000000c4",
            INIT_03 => X"00000013000000750000008c0000004800000009000000110000003b00000025",
            INIT_04 => X"00000045000000350000002c000000280000001a000000180000001500000019",
            INIT_05 => X"000000fb00000094000000200000003100000029000000250000005200000058",
            INIT_06 => X"0000001f0000008b000000e2000000e1000000e2000000e9000000f2000000f6",
            INIT_07 => X"0000002200000097000000a2000000850000004300000028000000190000000b",
            INIT_08 => X"000000360000002e000000460000005d00000026000000160000001300000016",
            INIT_09 => X"000000e3000000a300000031000000380000001b00000018000000260000004b",
            INIT_0A => X"0000004a000000a3000000e4000000e5000000da000000cb000000cd000000d6",
            INIT_0B => X"00000033000000a0000000960000009700000095000000800000005a00000039",
            INIT_0C => X"0000002a000000240000005a000000af0000007c000000260000000f00000013",
            INIT_0D => X"000000d0000000aa0000004f00000040000000150000000b000000170000003f",
            INIT_0E => X"000000b1000000e3000000d9000000ce000000d6000000d3000000c5000000c7",
            INIT_0F => X"0000002a00000088000000970000009a000000a2000000a7000000a800000098",
            INIT_10 => X"0000002e0000002f0000006f000000be000000dc000000650000000a00000012",
            INIT_11 => X"000000cc000000b1000000420000001f0000000e000000090000000a00000039",
            INIT_12 => X"000000d3000000ac000000660000004f0000007c000000c6000000ca000000c2",
            INIT_13 => X"000000110000004a0000008c0000009c000000a9000000b1000000b8000000c8",
            INIT_14 => X"00000034000000370000008000000096000000a500000084000000140000000e",
            INIT_15 => X"000000c6000000b4000000480000002d000000160000000a000000030000001e",
            INIT_16 => X"000000a3000000380000001e0000001a000000190000007b000000cd000000be",
            INIT_17 => X"000000110000000d0000004400000088000000930000009e000000b8000000ca",
            INIT_18 => X"000000350000003e00000082000000530000002100000053000000230000000a",
            INIT_19 => X"000000c2000000b7000000750000006c00000048000000100000000700000013",
            INIT_1A => X"0000004f000000140000002b000000310000001e0000002f000000b7000000c3",
            INIT_1B => X"00000018000000090000000a00000040000000810000008400000094000000a1",
            INIT_1C => X"000000240000004e00000088000000460000002300000037000000210000000a",
            INIT_1D => X"000000cd000000cd0000007e000000610000005800000022000000110000000f",
            INIT_1E => X"0000001f000000200000001f000000200000002b0000002000000098000000d0",
            INIT_1F => X"00000021000000190000000c00000017000000630000008a0000009100000075",
            INIT_20 => X"000000210000005700000088000000470000004100000036000000150000000a",
            INIT_21 => X"000000c5000000cf0000009a00000056000000570000003f0000002700000015",
            INIT_22 => X"0000000f0000001c0000002c00000037000000380000002500000081000000c6",
            INIT_23 => X"0000001f0000001c000000140000000e000000430000008b000000930000004d",
            INIT_24 => X"0000001c0000005600000080000000450000003e0000002f0000000e00000007",
            INIT_25 => X"000000b4000000b6000000a20000006f0000006f0000005e0000003c0000001e",
            INIT_26 => X"0000000f00000023000000350000004b0000003c000000290000007f000000bc",
            INIT_27 => X"00000016000000100000000d00000007000000260000006f0000007a0000002c",
            INIT_28 => X"0000003d0000006800000075000000460000003b00000027000000110000000b",
            INIT_29 => X"000000c7000000c9000000c3000000b9000000b70000009f0000007900000051",
            INIT_2A => X"0000001c0000003400000062000000660000003c0000002a00000088000000c6",
            INIT_2B => X"000000160000000c000000070000000300000010000000450000004f00000015",
            INIT_2C => X"0000003c000000550000006700000049000000430000001d0000001400000013",
            INIT_2D => X"0000006d000000710000007100000068000000640000005b0000005000000045",
            INIT_2E => X"000000170000001f00000042000000400000004100000025000000590000006d",
            INIT_2F => X"000000180000000b0000000600000006000000050000000e0000001400000008",
            INIT_30 => X"00000007000000160000002c0000002c000000250000001d0000001c00000017",
            INIT_31 => X"0000001000000011000000100000000d0000000c0000000c0000000a0000000a",
            INIT_32 => X"0000001000000038000000300000004400000043000000090000000f0000000f",
            INIT_33 => X"000000190000000e000000090000000600000004000000030000000300000004",
            INIT_34 => X"0000002000000019000000120000001700000020000000270000002500000021",
            INIT_35 => X"0000000f00000013000000150000001700000017000000170000001500000017",
            INIT_36 => X"0000000800000029000000470000003e00000018000000070000000a0000000b",
            INIT_37 => X"0000001d000000180000000e0000000900000006000000050000000500000004",
            INIT_38 => X"0000004d00000051000000430000003c00000032000000290000002500000023",
            INIT_39 => X"00000023000000270000002c00000031000000300000002d000000240000002c",
            INIT_3A => X"000000090000000a000000190000001700000010000000150000001b0000001d",
            INIT_3B => X"0000001e0000001f000000140000000e0000000b0000000a000000090000000b",
            INIT_3C => X"00000052000000660000006f0000006d000000570000003b0000002a0000002a",
            INIT_3D => X"0000004300000046000000480000004a00000047000000450000003e00000037",
            INIT_3E => X"00000012000000180000002c0000002f000000290000002b000000330000003b",
            INIT_3F => X"0000001e000000200000001c0000001600000013000000150000001600000014",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE39;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE40 : if BRAM_NAME = "sampleifmap_layer0_instance40" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000002000000050000000a000000090000000a0000000e0000000b0000000d",
            INIT_01 => X"0000000000000005000000060000000400000002000000010000000300000003",
            INIT_02 => X"000000080000001d000000170000001600000056000000230000000000000001",
            INIT_03 => X"000000050000000600000008000000130000001d000000270000001b0000000d",
            INIT_04 => X"00000000000000030000000800000007000000040000000a0000000c0000000d",
            INIT_05 => X"0000000100000004000000040000000200000001000000010000000200000004",
            INIT_06 => X"0000000700000006000000060000000700000013000000100000000100000001",
            INIT_07 => X"0000000600000004000000080000001300000016000000170000002e00000021",
            INIT_08 => X"0000000000000001000000040000000400000000000000030000000400000007",
            INIT_09 => X"0000000300000005000000060000000400000004000000040000000400000004",
            INIT_0A => X"0000000a000000060000000700000004000000090000000c0000000300000004",
            INIT_0B => X"0000000600000003000000060000000f0000000c0000000d0000002300000028",
            INIT_0C => X"000000030000000300000004000000120000000b000000080000000300000001",
            INIT_0D => X"0000000600000006000000090000000800000007000000080000000600000005",
            INIT_0E => X"00000017000000100000000a00000004000000090000000a0000000500000007",
            INIT_0F => X"0000000800000005000000060000000f0000000e00000011000000160000001e",
            INIT_10 => X"000000080000000700000006000000170000001a0000001d000000130000000c",
            INIT_11 => X"00000008000000070000000a0000000900000008000000090000000800000007",
            INIT_12 => X"0000002700000040000000250000000800000007000000080000000700000009",
            INIT_13 => X"000000090000000d0000000f0000000e000000150000000e0000001000000010",
            INIT_14 => X"000000080000000900000006000000090000000c000000160000001e00000018",
            INIT_15 => X"00000009000000070000000a0000000b0000000a000000090000000500000005",
            INIT_16 => X"0000003b0000005d0000005500000014000000070000000b0000000b0000000a",
            INIT_17 => X"00000009000000100000001b0000001700000020000000130000000e00000022",
            INIT_18 => X"000000070000000a0000000800000008000000070000000a0000000b0000000c",
            INIT_19 => X"0000000c0000000a0000000c0000000d0000000e0000000a0000000500000006",
            INIT_1A => X"000000280000003c0000005600000025000000070000000e0000000e00000009",
            INIT_1B => X"000000070000000600000010000000140000001c0000001c0000001c00000035",
            INIT_1C => X"000000090000000c0000000a0000000b00000007000000060000000600000003",
            INIT_1D => X"0000001300000010000000120000000e0000000e0000000c0000000800000009",
            INIT_1E => X"0000000a000000140000003e00000031000000160000001a0000001500000010",
            INIT_1F => X"000000070000000400000008000000090000000d000000100000001a0000001e",
            INIT_20 => X"0000000b0000000e0000000a0000000b00000008000000090000000a00000007",
            INIT_21 => X"000000280000002200000024000000130000000f0000000e0000000c0000000d",
            INIT_22 => X"000000090000000f0000002b0000003300000022000000220000002000000024",
            INIT_23 => X"000000080000000800000008000000080000000a000000090000000c00000014",
            INIT_24 => X"0000000d0000000e0000000a0000000c000000080000000b0000000c0000000c",
            INIT_25 => X"0000002600000028000000310000002700000022000000140000000e0000000e",
            INIT_26 => X"00000026000000340000003b0000003600000032000000270000001b00000020",
            INIT_27 => X"0000000a0000000b00000009000000060000000c0000000b0000001500000023",
            INIT_28 => X"0000000d0000000d0000000a0000000c000000090000000b0000000b0000000c",
            INIT_29 => X"0000003f000000320000003200000020000000280000001b000000100000000d",
            INIT_2A => X"00000022000000540000007100000079000000b4000000a10000007700000058",
            INIT_2B => X"0000000a0000000c0000000a00000009000000110000001d0000003100000032",
            INIT_2C => X"0000000c0000000d0000000c0000000e0000000b0000000e0000000a00000009",
            INIT_2D => X"000000ba000000af000000930000004d0000002700000018000000120000000c",
            INIT_2E => X"0000001c0000009e000000d5000000b1000000ca000000d2000000c8000000c8",
            INIT_2F => X"000000090000000b000000090000000a00000025000000460000002200000013",
            INIT_30 => X"0000000e0000000d0000000e000000100000000d0000000f0000000a00000008",
            INIT_31 => X"0000007d00000093000000a20000008e0000006c0000003e000000180000000c",
            INIT_32 => X"00000054000000d7000000f10000007e0000004a000000540000005e0000006e",
            INIT_33 => X"00000008000000090000000d000000190000004900000034000000090000000c",
            INIT_34 => X"0000000e0000000c00000010000000110000000e0000000f0000000b0000000b",
            INIT_35 => X"000000190000003d0000005f000000560000005d000000670000004400000014",
            INIT_36 => X"000000a7000000eb000000eb0000008900000017000000110000002300000016",
            INIT_37 => X"000000070000000900000011000000280000004200000017000000070000002a",
            INIT_38 => X"000000120000000b00000012000000100000000e000000120000000d0000000f",
            INIT_39 => X"0000001b0000003700000053000000440000002e0000003b0000005300000036",
            INIT_3A => X"000000e0000000e7000000e8000000c80000004c0000001c000000270000000c",
            INIT_3B => X"000000080000000d000000160000001f0000001a000000130000001600000073",
            INIT_3C => X"00000037000000390000001e0000000e0000000e000000130000000d00000010",
            INIT_3D => X"00000029000000320000004e000000520000003c00000039000000350000004f",
            INIT_3E => X"000000dd000000ec000000e6000000e7000000c80000007c0000004700000023",
            INIT_3F => X"000000090000003f00000049000000200000000e0000001a000000440000007e",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE40;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE41 : if BRAM_NAME = "sampleifmap_layer0_instance41" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000005c0000005d0000002f0000001800000011000000130000000e00000011",
            INIT_01 => X"000000a60000005e000000470000004c0000003d0000003c000000620000004f",
            INIT_02 => X"0000007c000000e7000000f0000000ed000000fc000000fa000000e2000000c6",
            INIT_03 => X"000000110000007e000000950000004c0000000c0000001c0000004a0000002a",
            INIT_04 => X"00000048000000380000002a0000002400000015000000120000001000000012",
            INIT_05 => X"000001000000009a000000220000002d00000024000000240000005800000060",
            INIT_06 => X"0000002700000096000000ee000000ed000000ed000000f4000000f9000000fa",
            INIT_07 => X"00000026000000a3000000ae0000008e0000004d0000003b0000002e00000015",
            INIT_08 => X"000000420000003c000000490000005c00000022000000100000001000000011",
            INIT_09 => X"000000f0000000ae000000370000003e000000210000001c0000002c00000054",
            INIT_0A => X"00000056000000b1000000ee000000ef000000e7000000d9000000d9000000e1",
            INIT_0B => X"00000037000000a9000000a1000000a4000000a4000000920000006a00000045",
            INIT_0C => X"000000380000003500000062000000b40000007d000000200000000a0000000d",
            INIT_0D => X"000000e0000000b900000059000000490000001b0000000e0000001c00000048",
            INIT_0E => X"000000c0000000f2000000e1000000d7000000e3000000e4000000d5000000d5",
            INIT_0F => X"0000002a0000008d0000009f000000a6000000b0000000b5000000b4000000a5",
            INIT_10 => X"000000390000003e0000007b000000c9000000e500000065000000070000000c",
            INIT_11 => X"000000da000000bf0000004f000000260000000f000000090000000f00000041",
            INIT_12 => X"000000e4000000b80000006d000000580000008a000000d8000000db000000d0",
            INIT_13 => X"0000000e0000004d00000093000000a6000000b5000000bf000000c9000000da",
            INIT_14 => X"0000003d000000450000008d000000a2000000b30000008b000000180000000d",
            INIT_15 => X"000000d4000000c200000056000000360000001b0000000b0000000400000023",
            INIT_16 => X"000000b10000004000000022000000200000002400000088000000db000000cc",
            INIT_17 => X"0000000d0000000f00000049000000900000009f000000ad000000cc000000dd",
            INIT_18 => X"0000003e0000004c0000008f00000060000000310000005b0000002700000009",
            INIT_19 => X"000000d0000000c5000000830000007900000051000000150000000700000015",
            INIT_1A => X"00000059000000190000002e000000370000002600000038000000c1000000d1",
            INIT_1B => X"00000014000000080000000e000000480000008d00000095000000a9000000b2",
            INIT_1C => X"0000002d0000005c0000009500000053000000300000003b0000002200000005",
            INIT_1D => X"000000db000000db0000008c0000006f000000640000002a000000130000000f",
            INIT_1E => X"000000270000002400000023000000250000003300000026000000a0000000de",
            INIT_1F => X"0000001e000000160000000c0000001d0000006e0000009b000000a400000082",
            INIT_20 => X"0000002a0000006500000094000000540000004d0000003a0000001700000007",
            INIT_21 => X"000000d3000000dd000000a800000064000000650000004a0000002b00000016",
            INIT_22 => X"0000001500000023000000340000003f000000400000002b00000089000000d4",
            INIT_23 => X"0000001c0000001800000012000000130000004e0000009a000000a200000056",
            INIT_24 => X"00000025000000650000008c000000520000004c000000370000001500000009",
            INIT_25 => X"000000c2000000c3000000b00000007e0000007f0000006c0000004300000021",
            INIT_26 => X"000000150000002e0000004100000056000000460000003000000087000000c9",
            INIT_27 => X"000000140000000b0000000a0000000b000000310000007b0000008300000032",
            INIT_28 => X"0000004b0000007800000084000000570000004900000031000000170000000b",
            INIT_29 => X"000000d5000000d4000000cf000000c8000000c8000000b1000000860000005d",
            INIT_2A => X"00000022000000400000006e00000071000000480000003500000094000000d6",
            INIT_2B => X"000000160000000d0000000900000007000000160000004c0000005500000018",
            INIT_2C => X"000000480000006000000073000000570000004e00000025000000160000000f",
            INIT_2D => X"0000007b0000007e0000007d0000007700000072000000690000005d00000052",
            INIT_2E => X"0000001b000000290000004e0000004b0000004c00000030000000660000007c",
            INIT_2F => X"000000190000000f0000000a0000000800000006000000100000001800000009",
            INIT_30 => X"0000000c0000001900000030000000320000002b000000230000001f00000015",
            INIT_31 => X"000000190000001a000000180000001400000011000000110000000e0000000e",
            INIT_32 => X"00000012000000410000003b0000004e0000004a0000000d0000001400000018",
            INIT_33 => X"0000001a0000000d000000090000000500000003000000040000000500000003",
            INIT_34 => X"000000250000001e000000170000001e000000250000002c0000002800000021",
            INIT_35 => X"0000001300000017000000180000001b0000001c0000001c000000190000001c",
            INIT_36 => X"000000080000002f00000053000000470000001c00000006000000090000000f",
            INIT_37 => X"0000001c000000150000000b0000000600000004000000050000000500000002",
            INIT_38 => X"000000590000005c0000004f000000490000003b000000300000002900000025",
            INIT_39 => X"000000280000002b00000030000000390000003b000000380000002f00000038",
            INIT_3A => X"0000000800000010000000250000002100000015000000150000001b00000023",
            INIT_3B => X"0000001c0000001d000000120000000d0000000a0000000a0000000900000008",
            INIT_3C => X"000000630000007600000080000000800000006500000046000000310000002c",
            INIT_3D => X"0000004f00000051000000530000005700000055000000540000004e00000047",
            INIT_3E => X"0000001300000020000000380000003a00000031000000310000003c00000047",
            INIT_3F => X"0000001c000000220000001f0000001900000015000000180000001800000013",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE41;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE42 : if BRAM_NAME = "sampleifmap_layer0_instance42" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000005c0000005b00000055000000510000004d000000510000005200000053",
            INIT_01 => X"0000004c0000005000000052000000570000005c000000650000005f0000005c",
            INIT_02 => X"0000002f00000034000000380000003c0000003e0000003f0000004100000044",
            INIT_03 => X"00000015000000190000001d000000240000002200000023000000250000002a",
            INIT_04 => X"0000005d0000005a00000054000000500000004d000000530000005300000054",
            INIT_05 => X"0000004c0000004e0000005200000058000000610000005f000000580000005a",
            INIT_06 => X"0000002e00000034000000360000003d00000042000000400000004400000047",
            INIT_07 => X"0000001f0000001d0000001e000000240000002300000024000000260000002a",
            INIT_08 => X"0000004c00000058000000540000004b0000004b000000500000005100000052",
            INIT_09 => X"0000004c0000004d000000580000006500000063000000570000005600000052",
            INIT_0A => X"0000002d00000034000000370000003a00000040000000400000004400000049",
            INIT_0B => X"000000350000003100000030000000310000002c00000029000000280000002b",
            INIT_0C => X"0000003200000050000000570000004a0000004e000000500000005100000053",
            INIT_0D => X"000000500000005800000066000000680000005b000000570000006100000055",
            INIT_0E => X"0000003a00000039000000380000003b0000003f0000003f0000004000000049",
            INIT_0F => X"0000004500000045000000470000004900000047000000440000003f0000003d",
            INIT_10 => X"000000370000004c000000530000004a0000004f0000004f0000004f0000004f",
            INIT_11 => X"000000570000005a000000590000004e0000004b0000004b0000005400000053",
            INIT_12 => X"0000005700000054000000500000004e00000046000000430000004200000053",
            INIT_13 => X"000000490000004f000000540000005800000059000000590000005600000057",
            INIT_14 => X"000000460000004600000049000000490000004d0000004b0000004a0000004c",
            INIT_15 => X"000000510000004e0000004e0000004b00000049000000470000004500000046",
            INIT_16 => X"000000680000006600000068000000640000006200000060000000590000005a",
            INIT_17 => X"000000420000004900000050000000570000005e000000610000005f00000063",
            INIT_18 => X"000000330000002b0000003e0000004a0000004900000047000000480000004a",
            INIT_19 => X"0000005e000000510000004a0000004b00000047000000440000004000000044",
            INIT_1A => X"0000006d000000680000006400000066000000720000006e0000006200000060",
            INIT_1B => X"0000004300000046000000490000004c00000050000000550000005b00000063",
            INIT_1C => X"000000290000002a0000003a0000004700000048000000470000004800000047",
            INIT_1D => X"000000600000005200000047000000410000003f0000003a0000003600000039",
            INIT_1E => X"000000610000006c0000006a00000067000000670000005d0000005e00000069",
            INIT_1F => X"0000004d0000004f000000500000005000000050000000540000005b0000005d",
            INIT_20 => X"0000002e000000570000006700000058000000520000004b0000004900000049",
            INIT_21 => X"000000570000005a000000570000005100000052000000450000003800000038",
            INIT_22 => X"000000660000006a00000066000000610000005b0000005e0000006300000062",
            INIT_23 => X"0000005f0000005b00000059000000590000005c00000061000000630000005e",
            INIT_24 => X"000000330000006800000099000000880000007b0000006d0000005f00000056",
            INIT_25 => X"0000005a000000660000006c0000006500000061000000490000003b0000003c",
            INIT_26 => X"0000006e00000069000000630000005d0000005d00000061000000610000005f",
            INIT_27 => X"0000006e0000006e0000006e0000006d0000006c0000006c0000006900000067",
            INIT_28 => X"0000003200000057000000a2000000a00000009d000000960000008b0000007f",
            INIT_29 => X"0000005a0000006b000000700000006500000058000000350000003800000043",
            INIT_2A => X"00000065000000600000005f00000060000000600000005e000000600000005e",
            INIT_2B => X"0000007000000074000000770000007b0000007e0000007d0000007100000068",
            INIT_2C => X"0000002c0000005a0000009f000000a0000000a20000009f0000009d00000098",
            INIT_2D => X"0000005c000000610000005a00000067000000560000003a0000004500000048",
            INIT_2E => X"0000005c0000005700000062000000630000005e0000005f000000600000005a",
            INIT_2F => X"0000006c00000074000000790000007f00000083000000830000007000000061",
            INIT_30 => X"000000300000007200000094000000980000009d000000a00000009e0000009b",
            INIT_31 => X"0000005d000000580000006000000073000000670000005e0000005800000044",
            INIT_32 => X"000000550000005400000065000000630000005e000000620000006500000059",
            INIT_33 => X"0000005f0000006b000000760000007f000000840000007d0000006e00000069",
            INIT_34 => X"00000050000000880000008e0000009000000092000000950000009400000094",
            INIT_35 => X"0000005e0000005c0000007100000072000000680000005e000000480000002f",
            INIT_36 => X"000000520000005500000061000000600000005d00000061000000670000005d",
            INIT_37 => X"0000004d000000570000006400000070000000790000006f0000006b0000006b",
            INIT_38 => X"0000008900000097000000930000008e0000008c0000008a0000008700000086",
            INIT_39 => X"000000620000005a0000005e000000590000003e00000032000000490000005d",
            INIT_3A => X"00000053000000560000005e0000005e00000061000000670000006900000066",
            INIT_3B => X"0000004b0000004a000000520000005f000000660000005c000000650000005f",
            INIT_3C => X"000000980000009a0000009f00000098000000900000008b0000008600000083",
            INIT_3D => X"000000660000005f00000064000000670000003900000035000000760000009e",
            INIT_3E => X"00000055000000570000005b000000610000006a0000006f000000740000006e",
            INIT_3F => X"0000005f0000005a000000550000005300000053000000550000006200000054",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE42;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE43 : if BRAM_NAME = "sampleifmap_layer0_instance43" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000007300000089000000a1000000a4000000a0000000980000009000000087",
            INIT_01 => X"00000067000000680000007a0000007b0000006e00000080000000910000009d",
            INIT_02 => X"00000057000000580000005a00000061000000680000006c0000006d00000069",
            INIT_03 => X"0000005e00000069000000690000006500000055000000570000005c0000004f",
            INIT_04 => X"0000007f000000b0000000b3000000aa000000a40000009f0000009a00000094",
            INIT_05 => X"00000067000000800000009100000071000000980000009d000000c5000000b0",
            INIT_06 => X"000000590000005b0000005f0000006100000066000000680000006500000067",
            INIT_07 => X"0000004600000056000000680000006d0000005b0000005b000000560000004f",
            INIT_08 => X"000000c4000000f8000000ee000000dd000000c5000000b2000000a40000009b",
            INIT_09 => X"0000006a000000890000008e0000006c000000b8000000b0000000c80000009c",
            INIT_0A => X"000000590000005f000000630000006500000065000000640000006300000064",
            INIT_0B => X"00000047000000490000005200000058000000530000005c0000005100000050",
            INIT_0C => X"000000f4000000fb000000f6000000fd000000f9000000eb000000d6000000bf",
            INIT_0D => X"0000006e0000008b0000007200000071000000c3000000ac0000009e000000a0",
            INIT_0E => X"0000005c00000066000000680000006700000063000000610000006200000062",
            INIT_0F => X"000000480000004a000000500000004b00000049000000550000004e00000053",
            INIT_10 => X"000000c9000000ba000000bb000000f3000000fe000000fd000000fc000000f5",
            INIT_11 => X"00000072000000800000006a000000740000009c000000970000008000000091",
            INIT_12 => X"0000005c000000690000006e0000006c00000067000000650000006700000068",
            INIT_13 => X"000000490000004d000000530000004e00000055000000540000004c00000052",
            INIT_14 => X"000000720000006b0000007e000000e900000100000000fc000000fc000000fb",
            INIT_15 => X"000000670000006800000063000000630000006e000000780000007300000069",
            INIT_16 => X"00000056000000600000006e000000700000006b0000006b0000006e0000006d",
            INIT_17 => X"0000004f00000052000000520000005b000000680000005a0000004c0000004e",
            INIT_18 => X"00000076000000720000007c000000c8000000eb000000f6000000f8000000f8",
            INIT_19 => X"000000440000004b00000056000000500000004f00000053000000570000005d",
            INIT_1A => X"000000610000006100000061000000620000006100000062000000640000005f",
            INIT_1B => X"0000005200000052000000550000006e0000006f0000005b000000570000005b",
            INIT_1C => X"0000008400000085000000880000008a00000096000000b5000000d6000000eb",
            INIT_1D => X"0000003a0000006000000059000000430000003c000000390000003d00000064",
            INIT_1E => X"0000006500000068000000650000005e00000050000000470000004500000033",
            INIT_1F => X"000000510000005100000062000000770000006d0000005e000000570000005d",
            INIT_20 => X"000000670000006f0000007a0000007c000000780000007a0000008200000099",
            INIT_21 => X"000000530000006a000000660000004500000034000000390000005a0000006a",
            INIT_22 => X"0000006d000000660000006700000064000000550000004d0000004700000040",
            INIT_23 => X"000000500000005c0000007300000071000000630000005d000000570000006a",
            INIT_24 => X"0000006d0000006600000061000000650000006d000000720000006f0000006d",
            INIT_25 => X"000000590000005f000000650000005d00000055000000670000007800000075",
            INIT_26 => X"000000660000006900000077000000720000005a000000520000004b0000004a",
            INIT_27 => X"0000004f0000006b0000007500000065000000620000005e0000006b0000006f",
            INIT_28 => X"000000710000006f0000006a000000630000005b0000005d0000006200000069",
            INIT_29 => X"0000005c000000540000004c000000500000005f000000610000006800000070",
            INIT_2A => X"0000005e000000690000007b00000075000000590000004f0000004800000051",
            INIT_2B => X"0000005a0000006f000000690000006000000065000000670000006700000060",
            INIT_2C => X"000000640000006b0000006e0000006c000000650000005e0000005700000057",
            INIT_2D => X"0000005c0000004c000000490000005d0000006800000056000000510000005b",
            INIT_2E => X"000000560000005d000000640000005b0000004f0000004f0000004d00000058",
            INIT_2F => X"0000006500000066000000600000006000000060000000610000005c00000057",
            INIT_30 => X"00000050000000560000005f000000650000006900000067000000600000005a",
            INIT_31 => X"0000005d0000006000000055000000620000006a000000600000005500000051",
            INIT_32 => X"0000005b000000540000004c000000470000004c0000004f0000005100000058",
            INIT_33 => X"000000600000005b00000060000000620000005a00000053000000560000005c",
            INIT_34 => X"0000004f0000004f0000004f00000050000000560000005f0000006300000064",
            INIT_35 => X"000000590000006100000060000000630000006c000000620000005300000052",
            INIT_36 => X"00000059000000520000004a0000004c000000510000004f000000540000005c",
            INIT_37 => X"00000053000000530000005c0000005d0000005600000052000000550000005a",
            INIT_38 => X"0000005300000059000000570000004d00000047000000490000004e00000057",
            INIT_39 => X"0000005c0000005900000067000000640000006a000000610000004f00000051",
            INIT_3A => X"00000053000000540000004f0000005200000059000000580000005700000060",
            INIT_3B => X"000000490000004f000000560000005600000053000000560000005a00000056",
            INIT_3C => X"0000005100000053000000560000005400000049000000460000003f0000003e",
            INIT_3D => X"000000580000005b000000680000005f0000006b0000005e0000004a0000004e",
            INIT_3E => X"000000530000005500000050000000550000005900000058000000580000005b",
            INIT_3F => X"000000480000004c0000004d0000004c00000050000000560000005900000054",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE43;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE44 : if BRAM_NAME = "sampleifmap_layer0_instance44" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000060000000600000005a0000005a000000590000005d0000005e0000005e",
            INIT_01 => X"0000005200000055000000580000005e000000650000006e0000006600000061",
            INIT_02 => X"000000380000003d000000410000004500000048000000490000004b0000004e",
            INIT_03 => X"000000190000001d000000220000002800000027000000290000002e00000033",
            INIT_04 => X"000000620000005f0000005900000059000000590000005f0000005f00000060",
            INIT_05 => X"000000520000005500000059000000600000006b0000006a0000006000000061",
            INIT_06 => X"000000350000003b0000003d0000004400000049000000470000004b0000004f",
            INIT_07 => X"0000001f0000001f000000200000002600000025000000270000002c00000031",
            INIT_08 => X"000000510000005d0000005a00000054000000570000005c0000005c0000005e",
            INIT_09 => X"000000540000005600000062000000700000006e000000630000006000000059",
            INIT_0A => X"00000030000000360000003a0000003f0000004600000044000000490000004f",
            INIT_0B => X"00000031000000300000002e0000002f0000002b000000290000002b0000002e",
            INIT_0C => X"00000039000000560000005d000000530000005a0000005c0000005d0000005f",
            INIT_0D => X"0000005a00000065000000720000007400000068000000630000006b0000005d",
            INIT_0E => X"0000003900000038000000380000003e0000004200000042000000430000004e",
            INIT_0F => X"0000003d0000003f000000410000004300000042000000410000003e0000003c",
            INIT_10 => X"0000003e0000005200000059000000530000005b0000005b0000005b0000005c",
            INIT_11 => X"0000006400000069000000680000005c00000058000000580000005f0000005c",
            INIT_12 => X"00000053000000500000004d000000500000004800000045000000460000005b",
            INIT_13 => X"0000003f000000460000004b0000004f00000050000000510000005100000053",
            INIT_14 => X"0000004d0000004c0000004f0000005200000059000000570000005600000058",
            INIT_15 => X"0000005f0000005e0000005e0000005a00000057000000550000005200000050",
            INIT_16 => X"0000006200000060000000640000006400000063000000620000005e00000063",
            INIT_17 => X"000000370000003e000000450000004c0000005300000058000000580000005d",
            INIT_18 => X"000000370000002a0000003d0000005100000054000000520000005400000055",
            INIT_19 => X"000000650000005d000000570000005b00000059000000580000005700000053",
            INIT_1A => X"0000006700000067000000670000006900000073000000700000006400000062",
            INIT_1B => X"00000036000000390000003f000000440000004a0000004e000000500000005b",
            INIT_1C => X"0000002c00000026000000370000004c00000054000000520000005300000052",
            INIT_1D => X"000000630000005b00000053000000500000005100000052000000550000004c",
            INIT_1E => X"0000005e00000071000000720000006d0000006c000000610000006000000067",
            INIT_1F => X"0000003b0000004000000044000000470000004b0000004d0000004d00000052",
            INIT_20 => X"0000003100000055000000680000005e0000005b000000540000005200000051",
            INIT_21 => X"0000005e000000650000006400000061000000630000005b0000005400000049",
            INIT_22 => X"00000067000000720000006f0000006a00000062000000650000006800000065",
            INIT_23 => X"0000004800000047000000460000004a0000004e000000520000005500000057",
            INIT_24 => X"00000036000000680000009d0000008e0000008000000073000000650000005c",
            INIT_25 => X"00000065000000750000007c00000075000000710000005d000000540000004b",
            INIT_26 => X"00000076000000740000006e00000068000000670000006b0000006a00000067",
            INIT_27 => X"0000005200000055000000550000005500000054000000550000005a00000064",
            INIT_28 => X"0000003500000059000000aa000000a6000000a0000000990000008e00000082",
            INIT_29 => X"0000006b0000007f000000820000007700000068000000460000004d00000050",
            INIT_2A => X"000000720000006e000000690000006a0000006a000000690000006c0000006a",
            INIT_2B => X"00000055000000590000005b0000005e00000060000000620000006200000069",
            INIT_2C => X"0000002e0000005d000000a9000000a7000000a4000000a20000009f0000009a",
            INIT_2D => X"000000720000007a000000700000007b000000670000004a0000005600000051",
            INIT_2E => X"0000006e00000067000000690000006b000000670000006a0000006d0000006a",
            INIT_2F => X"000000550000005a0000005e0000006000000063000000650000006100000066",
            INIT_30 => X"00000030000000750000009f0000009e0000009e000000a10000009f0000009d",
            INIT_31 => X"00000075000000740000007800000087000000780000006c0000006500000049",
            INIT_32 => X"00000069000000640000006a00000069000000660000006c000000730000006b",
            INIT_33 => X"0000004c000000550000005d0000006200000065000000600000006000000070",
            INIT_34 => X"0000004c00000087000000930000009300000093000000970000009800000099",
            INIT_35 => X"000000710000007300000085000000830000007500000067000000490000002c",
            INIT_36 => X"00000064000000650000006a0000006a0000006b00000071000000770000006c",
            INIT_37 => X"000000400000004a000000550000005d000000620000005d0000006900000075",
            INIT_38 => X"0000008300000095000000940000008f0000008e0000008e0000008e0000008f",
            INIT_39 => X"0000006d000000680000006b0000006300000046000000350000004100000054",
            INIT_3A => X"00000062000000650000006c0000006e000000750000007d0000007c00000072",
            INIT_3B => X"0000003f0000004100000048000000550000005a000000580000006f0000006c",
            INIT_3C => X"0000009300000099000000a000000099000000910000008e0000008d0000008c",
            INIT_3D => X"0000006e00000065000000680000006a0000003a000000340000006f00000097",
            INIT_3E => X"00000065000000680000006c000000730000008000000087000000890000007b",
            INIT_3F => X"0000004d0000004a000000480000004a0000004e000000590000006f00000063",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE44;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE45 : if BRAM_NAME = "sampleifmap_layer0_instance45" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000007200000088000000a0000000a40000009f0000009b000000950000008f",
            INIT_01 => X"0000006c000000660000007700000076000000680000007a0000008f0000009b",
            INIT_02 => X"0000006a0000006b0000006d0000007500000080000000850000008400000078",
            INIT_03 => X"000000440000004f000000540000005a00000056000000620000006c00000061",
            INIT_04 => X"00000081000000b0000000b1000000a7000000a10000009f0000009d0000009a",
            INIT_05 => X"0000006c0000007b00000089000000680000008e00000097000000c7000000b3",
            INIT_06 => X"0000006e00000070000000730000007700000080000000830000007e00000079",
            INIT_07 => X"00000027000000340000004a0000005c0000005e0000006a0000006900000063",
            INIT_08 => X"000000c7000000f7000000ec000000da000000c1000000b0000000a40000009d",
            INIT_09 => X"00000071000000860000008800000065000000b1000000ad000000ce000000a3",
            INIT_0A => X"00000071000000760000007a0000007d00000081000000820000007e00000077",
            INIT_0B => X"00000027000000250000002c0000003e000000500000006a0000006700000068",
            INIT_0C => X"000000f7000000fa000000f2000000fa000000f6000000e8000000d4000000c0",
            INIT_0D => X"000000780000008b000000700000006e000000c1000000ae000000aa000000a9",
            INIT_0E => X"000000740000007e0000007f0000008000000080000000800000007e00000076",
            INIT_0F => X"0000002b00000027000000250000002a0000003e00000060000000660000006c",
            INIT_10 => X"000000d2000000be000000ba000000f1000000fb000000fa000000fb000000f5",
            INIT_11 => X"0000007a00000087000000730000007d000000a00000009c00000092000000a1",
            INIT_12 => X"000000740000007d0000007f0000007f00000080000000810000007f00000078",
            INIT_13 => X"00000029000000290000002a0000002d0000004200000057000000620000006a",
            INIT_14 => X"000000820000007400000083000000ea000000fe000000fb000000fb000000fb",
            INIT_15 => X"0000006b00000072000000770000007a0000007c000000820000008a0000007f",
            INIT_16 => X"0000006c0000006f000000770000007d0000007f000000820000008000000076",
            INIT_17 => X"000000290000002c0000002f0000003d00000050000000520000005a00000063",
            INIT_18 => X"000000830000007b00000080000000cb000000ef000000f9000000fc000000fc",
            INIT_19 => X"0000004400000051000000690000006a00000067000000660000006c0000006f",
            INIT_1A => X"00000073000000700000006b0000006e00000074000000780000007500000066",
            INIT_1B => X"0000002d0000002d0000003400000051000000540000004b0000005900000068",
            INIT_1C => X"0000008a000000890000008900000090000000a0000000bf000000df000000f5",
            INIT_1D => X"0000003a00000063000000660000005a00000057000000510000004b0000006d",
            INIT_1E => X"000000740000007a000000740000006d000000650000005f000000560000003a",
            INIT_1F => X"0000002f0000002f000000420000005900000050000000460000004d00000061",
            INIT_20 => X"00000069000000700000007b0000008200000084000000860000008d000000a5",
            INIT_21 => X"000000560000006f0000006e00000053000000470000004a0000005e0000006b",
            INIT_22 => X"0000007c0000007b0000007b000000760000006c000000660000005a00000048",
            INIT_23 => X"000000300000003d00000054000000520000004400000042000000490000006c",
            INIT_24 => X"0000006a00000065000000610000006a000000750000007a0000007800000075",
            INIT_25 => X"0000006100000068000000680000005c000000570000006a0000007300000070",
            INIT_26 => X"0000007a000000820000008e00000086000000720000006c0000005f00000054",
            INIT_27 => X"000000320000004f000000570000004500000040000000450000006400000077",
            INIT_28 => X"0000006b0000006e0000006b000000650000005e00000060000000660000006c",
            INIT_29 => X"000000680000005d000000480000004200000051000000560000005d00000067",
            INIT_2A => X"0000007a000000850000009400000089000000710000006b0000005f0000005e",
            INIT_2B => X"0000003f000000550000004b0000004000000042000000510000006b00000072",
            INIT_2C => X"00000057000000650000006c0000006b000000630000005d0000005700000058",
            INIT_2D => X"0000005e0000004e0000003f0000004a00000053000000410000003c00000049",
            INIT_2E => X"000000720000007a0000007b000000690000005d0000005f0000005700000059",
            INIT_2F => X"0000004b0000004a0000003f0000003c0000003b0000004e000000680000006d",
            INIT_30 => X"0000003800000045000000540000005b0000005f000000610000005f0000005d",
            INIT_31 => X"0000004800000055000000490000005300000055000000420000003100000032",
            INIT_32 => X"0000006800000064000000580000004500000044000000430000003e0000003e",
            INIT_33 => X"000000450000003a000000360000003500000033000000400000005a00000065",
            INIT_34 => X"0000003000000034000000370000003b00000044000000510000005b00000060",
            INIT_35 => X"000000390000004d0000004f0000005200000052000000400000002e0000002f",
            INIT_36 => X"0000004a000000470000003f0000003a0000003a000000340000003200000035",
            INIT_37 => X"000000360000003000000031000000300000002e000000340000004100000048",
            INIT_38 => X"0000003000000034000000300000002c0000002b000000310000003c00000049",
            INIT_39 => X"000000350000003e0000004f0000004b000000490000003a0000002c00000030",
            INIT_3A => X"0000002f000000330000002f0000003400000039000000340000002e00000032",
            INIT_3B => X"0000002a0000002b0000002d0000002b0000002a0000002e000000310000002f",
            INIT_3C => X"0000002d00000029000000290000002a00000025000000270000002500000029",
            INIT_3D => X"0000002e0000003b0000004c0000004300000047000000360000002b0000002f",
            INIT_3E => X"0000002d000000310000002d0000002f000000300000002d0000002a0000002b",
            INIT_3F => X"00000026000000280000002800000025000000270000002a0000002d0000002b",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE45;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE46 : if BRAM_NAME = "sampleifmap_layer0_instance46" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000005f0000005d00000052000000500000004f000000530000005400000055",
            INIT_01 => X"0000004f000000540000004e0000004b000000480000004f000000550000005a",
            INIT_02 => X"00000033000000380000003b0000003c0000003d0000003c0000003e00000044",
            INIT_03 => X"00000015000000190000001e000000240000002300000025000000290000002e",
            INIT_04 => X"0000005d0000005a000000500000004e0000004f000000550000005500000056",
            INIT_05 => X"0000004800000047000000450000004400000047000000460000004900000054",
            INIT_06 => X"0000002e0000003400000035000000380000003e0000003e0000004300000046",
            INIT_07 => X"0000001b0000001a0000001b0000002100000020000000220000002500000029",
            INIT_08 => X"000000480000005600000050000000490000004e000000520000005300000054",
            INIT_09 => X"0000003c000000360000003f0000004800000043000000380000004100000046",
            INIT_0A => X"000000260000002d0000002f000000300000003a0000003d0000004100000042",
            INIT_0B => X"0000002c0000002a000000290000002a00000025000000220000002100000024",
            INIT_0C => X"0000002b0000004d000000520000004800000050000000520000005300000055",
            INIT_0D => X"0000002f000000320000003f0000004100000034000000320000004500000043",
            INIT_0E => X"0000002c0000002b0000002b0000002d00000036000000390000003400000032",
            INIT_0F => X"00000037000000380000003b0000003c0000003b00000038000000320000002f",
            INIT_10 => X"0000002c000000460000004c0000004800000051000000510000005100000052",
            INIT_11 => X"0000002300000026000000270000001f0000001d00000022000000330000003d",
            INIT_12 => X"00000044000000410000003d0000003d0000003b000000390000002b00000029",
            INIT_13 => X"000000380000003e000000430000004700000048000000470000004200000044",
            INIT_14 => X"000000380000003e00000042000000470000004f0000004c0000004c0000004d",
            INIT_15 => X"0000000e0000000f0000001400000016000000170000001a000000210000002c",
            INIT_16 => X"000000500000004e0000005200000053000000540000004f000000350000001f",
            INIT_17 => X"0000002e000000350000003c000000440000004b0000004d000000480000004c",
            INIT_18 => X"0000002000000020000000370000004700000048000000460000004700000049",
            INIT_19 => X"000000150000000e0000000b0000001200000013000000140000001800000026",
            INIT_1A => X"000000520000004f000000500000005600000059000000460000002900000018",
            INIT_1B => X"0000002a0000002d000000340000003b0000004300000048000000480000004b",
            INIT_1C => X"000000110000001c000000330000004300000045000000440000004500000044",
            INIT_1D => X"00000018000000110000000b000000090000000b0000000a0000000c00000017",
            INIT_1E => X"000000400000004d0000004f0000004d0000003f00000021000000160000001c",
            INIT_1F => X"0000002b0000002f000000360000003c00000042000000480000004900000041",
            INIT_20 => X"00000013000000460000005d000000520000004e000000470000004500000044",
            INIT_21 => X"0000001400000021000000210000002000000025000000190000000c00000012",
            INIT_22 => X"0000003b0000003c000000380000003100000021000000190000001800000016",
            INIT_23 => X"000000350000003400000034000000390000003f000000490000004b0000003b",
            INIT_24 => X"00000016000000550000008d0000008000000075000000670000005900000050",
            INIT_25 => X"0000001c000000350000003d0000003900000038000000210000000f00000015",
            INIT_26 => X"0000003a0000002d000000230000001800000014000000160000001600000015",
            INIT_27 => X"0000003d0000003f00000040000000410000004100000046000000480000003d",
            INIT_28 => X"00000018000000470000009800000098000000950000008e0000008300000077",
            INIT_29 => X"000000210000003f000000440000003c0000003100000015000000110000001e",
            INIT_2A => X"0000002b0000001c000000140000000f00000011000000150000001b00000019",
            INIT_2B => X"000000410000004400000047000000490000004a0000004d0000004600000037",
            INIT_2C => X"000000170000004f00000099000000990000009900000096000000940000008f",
            INIT_2D => X"0000002700000037000000300000003d0000002e000000190000002200000028",
            INIT_2E => X"0000001f000000120000001500000013000000150000001f000000240000001d",
            INIT_2F => X"000000450000004a0000004c0000004d0000004d0000004c0000003b0000002a",
            INIT_30 => X"000000200000006b000000920000009200000094000000970000009500000092",
            INIT_31 => X"000000290000002c00000034000000470000003b00000034000000370000002b",
            INIT_32 => X"00000019000000120000001c0000001a0000001e0000002c0000003200000022",
            INIT_33 => X"00000042000000490000004f000000510000005100000045000000320000002e",
            INIT_34 => X"000000400000007e000000890000008a0000008b0000008f0000008f00000090",
            INIT_35 => X"00000024000000280000004000000046000000410000003d0000002e0000001a",
            INIT_36 => X"00000013000000120000001d0000002100000028000000330000003600000024",
            INIT_37 => X"00000037000000400000004a0000004f0000004e0000003c000000330000002f",
            INIT_38 => X"0000007700000089000000880000008600000086000000860000008400000085",
            INIT_39 => X"00000022000000200000002a0000002e000000210000001b0000003100000047",
            INIT_3A => X"00000011000000110000001c00000027000000320000003d0000003900000028",
            INIT_3B => X"00000032000000360000003e0000004600000041000000300000003300000024",
            INIT_3C => X"0000008100000088000000910000008c00000085000000810000007f0000007d",
            INIT_3D => X"000000270000002700000033000000400000001e0000001e0000005a00000084",
            INIT_3E => X"00000013000000140000001c0000002c0000003d000000450000004500000031",
            INIT_3F => X"0000003d0000003c00000039000000350000002d000000290000003000000019",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE46;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE47 : if BRAM_NAME = "sampleifmap_layer0_instance47" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000005a000000750000009100000095000000910000008b000000840000007d",
            INIT_01 => X"00000028000000310000004d0000005700000050000000620000007200000080",
            INIT_02 => X"00000017000000190000001f0000002d0000003c000000440000003f0000002e",
            INIT_03 => X"000000320000003e00000042000000400000002d0000002b0000002a00000015",
            INIT_04 => X"000000680000009e000000a40000009a00000093000000900000008c00000088",
            INIT_05 => X"000000290000004b0000006700000050000000770000007a000000a600000095",
            INIT_06 => X"0000001b0000001f00000028000000300000003c00000041000000380000002d",
            INIT_07 => X"00000014000000230000003900000041000000320000002f0000002300000015",
            INIT_08 => X"000000b2000000eb000000e6000000d2000000b6000000a40000009700000090",
            INIT_09 => X"0000002d00000055000000670000004d000000950000008a000000ab00000085",
            INIT_0A => X"0000001d0000002700000030000000350000003c0000003f000000380000002b",
            INIT_0B => X"00000015000000160000001f00000027000000270000002f0000001d00000017",
            INIT_0C => X"000000e6000000f2000000f2000000f8000000f0000000e1000000cd000000b7",
            INIT_0D => X"00000031000000560000004d000000530000009f00000084000000840000008d",
            INIT_0E => X"000000210000002f00000037000000390000003a0000003c000000370000002a",
            INIT_0F => X"0000001b0000001c0000001d000000190000001c000000270000001a00000019",
            INIT_10 => X"000000b5000000ab000000b0000000ec000000f9000000f7000000f8000000f1",
            INIT_11 => X"00000034000000470000003c0000004d00000076000000720000006200000078",
            INIT_12 => X"0000002000000030000000390000003b0000003a00000039000000360000002e",
            INIT_13 => X"0000001a0000001f000000200000001c00000025000000250000001700000018",
            INIT_14 => X"00000055000000530000006a000000e0000000fd000000f9000000f9000000f8",
            INIT_15 => X"00000031000000340000002e0000003000000041000000510000004e00000047",
            INIT_16 => X"0000001b00000024000000330000003d00000039000000360000003700000033",
            INIT_17 => X"0000001c0000001f0000001f0000002800000036000000270000001600000015",
            INIT_18 => X"0000005e000000600000006d000000c2000000eb000000f5000000f8000000f7",
            INIT_19 => X"000000200000002d0000002b0000001c00000019000000230000003500000041",
            INIT_1A => X"000000290000002b0000002d000000300000002f0000002f000000330000002e",
            INIT_1B => X"0000001e0000001d00000021000000390000003a000000240000001e00000022",
            INIT_1C => X"000000740000007a000000810000008800000098000000b6000000d7000000ec",
            INIT_1D => X"00000022000000490000003400000014000000090000000d0000002300000051",
            INIT_1E => X"000000310000003b0000003b0000002f000000200000001a0000001c00000011",
            INIT_1F => X"0000001d0000001c0000002c0000003f00000034000000220000001a00000023",
            INIT_20 => X"0000005c00000068000000760000007b000000780000007a000000820000009a",
            INIT_21 => X"00000034000000450000003d0000001d000000120000001f000000460000005a",
            INIT_22 => X"0000003d00000041000000470000003a00000028000000240000002400000022",
            INIT_23 => X"0000001c000000270000003c00000038000000280000001f0000001700000030",
            INIT_24 => X"0000005d0000005b000000580000005f000000680000006d0000006b00000069",
            INIT_25 => X"000000310000002f00000038000000380000003e000000560000006200000060",
            INIT_26 => X"00000039000000480000005b0000004c000000300000002a0000002500000028",
            INIT_27 => X"0000001d000000370000003d0000002a000000230000001d0000002c00000036",
            INIT_28 => X"000000580000005b00000058000000560000005100000053000000590000005f",
            INIT_29 => X"000000340000002c00000023000000280000003e000000440000004900000053",
            INIT_2A => X"00000032000000470000005f0000005100000031000000270000001e00000028",
            INIT_2B => X"000000280000003a000000300000002200000023000000250000002a00000029",
            INIT_2C => X"000000400000004c0000005300000057000000550000004f000000490000004b",
            INIT_2D => X"000000310000002900000022000000320000003b0000002a0000002700000033",
            INIT_2E => X"0000002d0000003c000000450000003700000027000000240000001e00000026",
            INIT_2F => X"000000330000003000000024000000200000001d000000220000002600000026",
            INIT_30 => X"000000210000002c00000039000000440000004d0000004f0000004e0000004c",
            INIT_31 => X"000000260000003200000029000000370000003d0000002e0000001e0000001d",
            INIT_32 => X"000000300000002e000000250000001d0000001e0000001d0000001a0000001d",
            INIT_33 => X"0000002f00000024000000200000001e0000001800000019000000250000002e",
            INIT_34 => X"0000001b0000001e000000200000002600000032000000400000004a00000050",
            INIT_35 => X"0000001d0000002c0000002f000000350000003c0000002d0000001b0000001b",
            INIT_36 => X"000000250000002000000018000000190000001c00000017000000170000001c",
            INIT_37 => X"000000220000001c0000001e0000001a00000015000000150000001d00000023",
            INIT_38 => X"0000001c000000210000001d0000001a0000001a000000210000002d0000003a",
            INIT_39 => X"0000001c0000002100000032000000310000003300000027000000180000001b",
            INIT_3A => X"000000170000001900000015000000180000001d00000019000000150000001b",
            INIT_3B => X"00000017000000190000001a0000001500000012000000160000001a00000017",
            INIT_3C => X"0000001900000018000000190000001a0000001500000018000000170000001b",
            INIT_3D => X"0000001800000023000000330000002a0000003000000021000000160000001a",
            INIT_3E => X"000000190000001d000000170000001700000018000000150000001400000015",
            INIT_3F => X"0000001600000018000000160000001100000012000000160000001b00000018",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE47;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE48 : if BRAM_NAME = "sampleifmap_layer0_instance48" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b2000000b7000000bc000000a400000041000000150000001300000017",
            INIT_01 => X"000000b7000000b6000000b7000000b8000000ba000000ba000000ac000000aa",
            INIT_02 => X"000000c2000000990000006e0000006b0000005c0000007f000000a4000000b4",
            INIT_03 => X"000000c5000000c7000000c8000000c9000000c6000000c5000000c9000000c3",
            INIT_04 => X"000000b2000000bf000000ca000000990000002e000000150000001300000017",
            INIT_05 => X"000000b2000000b4000000b8000000ba000000b7000000a90000009e000000a4",
            INIT_06 => X"000000ce000000b40000006a0000004a000000560000008a000000ad000000b4",
            INIT_07 => X"000000ca000000cc000000cd000000cf000000ce000000d0000000d5000000cf",
            INIT_08 => X"000000a8000000b9000000c80000007f0000001f000000170000001400000017",
            INIT_09 => X"000000b2000000b3000000b2000000b2000000a20000009a0000009e0000009f",
            INIT_0A => X"000000d1000000c500000072000000470000007d000000b6000000be000000b5",
            INIT_0B => X"000000ce000000d0000000d3000000d4000000d3000000d5000000d8000000d5",
            INIT_0C => X"000000a0000000af000000bd0000006300000017000000180000001500000017",
            INIT_0D => X"000000c3000000bf000000ba000000aa00000095000000a6000000a8000000a8",
            INIT_0E => X"000000d6000000d200000092000000630000008d000000bc000000c8000000c3",
            INIT_0F => X"000000d6000000d7000000d9000000d9000000d5000000d4000000d4000000d5",
            INIT_10 => X"00000097000000a5000000aa0000004800000015000000170000001700000019",
            INIT_11 => X"000000bc000000a90000009d000000920000009b000000b9000000b7000000af",
            INIT_12 => X"000000db000000d3000000ac000000790000008d000000b2000000c4000000c5",
            INIT_13 => X"000000ce000000d1000000d4000000d6000000d9000000d9000000d9000000dd",
            INIT_14 => X"0000009a000000a40000008f00000031000000170000001a0000001b0000001a",
            INIT_15 => X"00000097000000800000007d00000082000000a6000000c8000000c2000000a9",
            INIT_16 => X"000000c9000000bc000000b6000000930000008f00000094000000a5000000a5",
            INIT_17 => X"000000d3000000d7000000d7000000dc000000db000000d5000000d9000000d4",
            INIT_18 => X"000000ab000000b40000007d00000025000000190000001b0000001a0000001e",
            INIT_19 => X"000000820000007a000000710000008b000000b3000000ca000000c5000000a9",
            INIT_1A => X"000000c9000000bf000000cb000000b90000008c0000007a0000008500000077",
            INIT_1B => X"000000e0000000dc000000da000000dc000000db000000d7000000da000000d7",
            INIT_1C => X"000000a8000000c1000000af00000064000000240000001f000000300000005e",
            INIT_1D => X"000000840000008e00000091000000ae000000c3000000c6000000c0000000a3",
            INIT_1E => X"000000d5000000bd000000d1000000c00000008b0000007a000000790000006a",
            INIT_1F => X"000000e5000000de000000d5000000d0000000e8000000ef000000ed000000f2",
            INIT_20 => X"000000a0000000be000000be000000b10000007a000000720000009e000000b4",
            INIT_21 => X"00000092000000a7000000b9000000c2000000c8000000c5000000ad00000085",
            INIT_22 => X"000000dc000000bd000000c9000000b10000008d000000850000008100000081",
            INIT_23 => X"000000ea000000e1000000c7000000bd000000d5000000e8000000eb000000f1",
            INIT_24 => X"0000009d000000c5000000c3000000c1000000ba000000b2000000c0000000c5",
            INIT_25 => X"00000097000000b2000000c3000000c1000000bf000000b9000000a300000080",
            INIT_26 => X"000000ea000000d0000000c2000000aa00000086000000830000008100000072",
            INIT_27 => X"000000eb000000d0000000bb000000b9000000c9000000eb000000f0000000ec",
            INIT_28 => X"00000097000000c5000000cd000000c8000000c0000000bb000000c4000000ca",
            INIT_29 => X"00000088000000a8000000bb000000c1000000bd000000b8000000af00000095",
            INIT_2A => X"000000f0000000cd000000b5000000a700000081000000800000008000000075",
            INIT_2B => X"000000dd000000c1000000bb000000ba000000ce000000ee000000f3000000f3",
            INIT_2C => X"000000a0000000c2000000d0000000cb000000c0000000c5000000cd000000cd",
            INIT_2D => X"0000007700000092000000ac000000c1000000bf000000c1000000bf000000a8",
            INIT_2E => X"000000ea000000bf000000b0000000a700000087000000850000008e0000007c",
            INIT_2F => X"000000c4000000b9000000b8000000ba000000d7000000ec000000f1000000f3",
            INIT_30 => X"000000b4000000bf000000c7000000c5000000c1000000c8000000cc000000ce",
            INIT_31 => X"0000008300000098000000ae000000ae000000ad000000b7000000b3000000ac",
            INIT_32 => X"000000e6000000bf000000ac000000a90000009a0000008e000000a60000008d",
            INIT_33 => X"000000c0000000b8000000ba000000c8000000e4000000ef000000f1000000f0",
            INIT_34 => X"000000ca000000b1000000b4000000c9000000bf000000c6000000ca000000d2",
            INIT_35 => X"0000009c00000093000000a8000000a80000008e0000008e0000009a000000ab",
            INIT_36 => X"000000e6000000c5000000a00000009e000000a400000096000000a9000000af",
            INIT_37 => X"000000d7000000c3000000bf000000e2000000f2000000f4000000f1000000f1",
            INIT_38 => X"000000d7000000a1000000aa000000cf000000c0000000c7000000c9000000d3",
            INIT_39 => X"0000007f00000089000000b1000000be000000ac000000ad000000ba000000bd",
            INIT_3A => X"000000ec000000c1000000b0000000af000000a000000096000000ae000000b4",
            INIT_3B => X"000000e1000000d4000000c9000000ef000000fb000000f3000000f2000000f5",
            INIT_3C => X"000000d90000009a000000b5000000d1000000c1000000c5000000c4000000d3",
            INIT_3D => X"00000098000000a6000000ad000000aa000000b9000000c3000000c5000000ce",
            INIT_3E => X"000000cc000000af000000b5000000c000000098000000a6000000b8000000a3",
            INIT_3F => X"000000e2000000e2000000d5000000df000000f7000000f4000000f3000000ee",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE48;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE49 : if BRAM_NAME = "sampleifmap_layer0_instance49" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000c60000009b000000c4000000c5000000b5000000b4000000c2000000d6",
            INIT_01 => X"000000b2000000ae000000a1000000ad000000b7000000ae000000c0000000d6",
            INIT_02 => X"000000760000009c000000b4000000a700000093000000bd000000a400000080",
            INIT_03 => X"000000e4000000ea000000d6000000ce000000eb000000ef000000d70000009d",
            INIT_04 => X"000000b9000000be000000ca000000b4000000a3000000a6000000c6000000d7",
            INIT_05 => X"000000ad000000b0000000ae000000c1000000d6000000cd000000d2000000cf",
            INIT_06 => X"00000087000000ab000000c8000000a300000099000000bf0000008900000081",
            INIT_07 => X"000000eb000000ef000000d2000000bb000000c1000000b80000009000000074",
            INIT_08 => X"000000c2000000d2000000cb000000b9000000a4000000ae000000cd000000d8",
            INIT_09 => X"000000b3000000be000000cb000000e1000000e2000000da000000d3000000bf",
            INIT_0A => X"000000ac000000aa000000c2000000a70000009e000000a80000007900000097",
            INIT_0B => X"000000ec000000de000000b8000000a2000000a900000099000000830000009a",
            INIT_0C => X"000000d2000000d1000000ca000000c5000000b4000000c0000000d0000000d8",
            INIT_0D => X"000000b5000000cf000000d5000000d1000000cc000000c5000000bd000000ba",
            INIT_0E => X"000000ab0000009c000000ae000000b7000000af0000009200000095000000b2",
            INIT_0F => X"000000cc000000ac000000a0000000a6000000b4000000a900000094000000a3",
            INIT_10 => X"000000ca000000c9000000cb000000bf000000b6000000ca000000d5000000da",
            INIT_11 => X"000000c7000000cf000000c6000000b2000000c0000000c1000000c3000000ca",
            INIT_12 => X"000000a6000000930000009b000000b1000000bb000000a6000000cb000000d3",
            INIT_13 => X"000000a70000009f0000009c0000009c000000af000000b6000000ab000000a7",
            INIT_14 => X"000000c8000000d0000000c8000000b3000000ba000000d1000000d7000000d9",
            INIT_15 => X"000000c2000000c4000000b6000000a1000000ba000000d2000000d7000000d1",
            INIT_16 => X"000000a60000009b0000008e0000009b000000b9000000be000000cf000000cb",
            INIT_17 => X"0000008f0000009e0000009e000000960000009f000000ad000000b3000000ac",
            INIT_18 => X"000000d9000000da000000c5000000a9000000c0000000d6000000d5000000d6",
            INIT_19 => X"000000bf000000c3000000b3000000aa000000c3000000d4000000d9000000d7",
            INIT_1A => X"000000aa000000a70000008e00000084000000aa000000c0000000c0000000be",
            INIT_1B => X"0000007d00000086000000930000009d0000009d000000ad000000b3000000aa",
            INIT_1C => X"000000de000000d8000000c1000000a8000000ca000000d3000000d1000000d5",
            INIT_1D => X"000000c6000000c9000000c2000000c2000000cd000000d3000000de000000df",
            INIT_1E => X"000000a7000000ab0000009b0000008600000099000000bc000000c4000000c6",
            INIT_1F => X"00000089000000850000008e000000a3000000a5000000b2000000bd000000a6",
            INIT_20 => X"000000d5000000d3000000bf000000af000000ca000000ce000000ce000000d3",
            INIT_21 => X"000000c9000000c9000000ce000000c2000000ab000000c6000000d8000000d6",
            INIT_22 => X"0000009d000000a70000009e0000009000000096000000b1000000c5000000c8",
            INIT_23 => X"00000090000000950000009600000098000000a8000000b0000000b50000009f",
            INIT_24 => X"000000d2000000d0000000bc000000b5000000c1000000c9000000cc000000d2",
            INIT_25 => X"000000c2000000c6000000d0000000b10000007a000000a0000000ce000000cd",
            INIT_26 => X"00000099000000a00000009c0000008b00000096000000a6000000b8000000c1",
            INIT_27 => X"000000830000008c00000098000000980000009b0000009f000000a00000009b",
            INIT_28 => X"000000d6000000cd000000b2000000ae000000bb000000c6000000ca000000d2",
            INIT_29 => X"000000b6000000bb000000ca000000b400000083000000a4000000cb000000d1",
            INIT_2A => X"000000900000009a00000099000000860000008b0000009d000000a9000000b6",
            INIT_2B => X"00000093000000960000009b0000009d0000008d000000830000008d00000097",
            INIT_2C => X"000000d7000000c4000000a8000000a8000000b5000000c2000000c8000000d2",
            INIT_2D => X"000000ac000000ad000000b9000000cb000000b8000000bd000000c7000000d4",
            INIT_2E => X"0000008d00000091000000940000008300000076000000930000009b000000a3",
            INIT_2F => X"0000009c000000a2000000a300000095000000850000007f0000008400000090",
            INIT_30 => X"000000d3000000bd0000009e000000a2000000b4000000bd000000c2000000d0",
            INIT_31 => X"000000a4000000a3000000ac000000bf000000c7000000c2000000c5000000d3",
            INIT_32 => X"000000910000009000000090000000890000006d00000082000000930000009e",
            INIT_33 => X"000000930000009f000000a200000097000000860000007c0000008400000090",
            INIT_34 => X"000000cd000000b30000008f0000009f000000b5000000b0000000b1000000c2",
            INIT_35 => X"000000a10000009c000000a5000000b5000000be000000c2000000c7000000d0",
            INIT_36 => X"000000920000008a000000850000008900000072000000700000008800000095",
            INIT_37 => X"0000008d00000094000000950000009600000090000000830000008300000092",
            INIT_38 => X"000000c70000009c00000085000000a7000000b2000000a50000009d000000ac",
            INIT_39 => X"0000008b0000008400000085000000a0000000c2000000c7000000c7000000ce",
            INIT_3A => X"000000950000008a00000081000000820000007e0000006b0000007e0000008c",
            INIT_3B => X"00000098000000950000008c000000880000008e000000910000008c0000008d",
            INIT_3C => X"000000b7000000820000007d0000009e0000009b000000900000008600000097",
            INIT_3D => X"000000690000005e0000006700000080000000a5000000b7000000bf000000c5",
            INIT_3E => X"0000008f0000008b0000007d000000790000007c000000750000007000000077",
            INIT_3F => X"000000960000009b00000095000000840000007d000000810000008c0000008b",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE49;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE50 : if BRAM_NAME = "sampleifmap_layer0_instance50" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000008e0000009300000093000000830000002f000000100000001500000013",
            INIT_01 => X"0000008f0000008c0000008c0000008d0000008e000000900000008900000087",
            INIT_02 => X"000000a4000000820000005d0000005f00000049000000600000007e0000008c",
            INIT_03 => X"00000097000000980000009b0000009e0000009d0000009b0000009c0000009b",
            INIT_04 => X"000000920000009b000000a10000007a0000001f000000110000001400000014",
            INIT_05 => X"00000097000000920000009600000098000000950000008b000000880000008a",
            INIT_06 => X"000000af0000009c00000058000000410000004900000075000000960000009f",
            INIT_07 => X"000000a3000000a4000000a8000000ac000000ad000000ab000000a9000000a8",
            INIT_08 => X"0000008c00000097000000a20000006600000015000000140000001400000014",
            INIT_09 => X"0000009f00000098000000990000009a0000008b00000088000000950000008d",
            INIT_0A => X"000000b7000000b1000000610000003a0000006d000000a1000000ab000000a6",
            INIT_0B => X"000000a6000000a9000000ad000000b1000000b2000000b1000000b2000000b3",
            INIT_0C => X"000000820000008c000000990000004f00000011000000150000001400000014",
            INIT_0D => X"000000b0000000a9000000a600000099000000870000009d000000a400000097",
            INIT_0E => X"000000c3000000c4000000850000005200000076000000a1000000af000000b0",
            INIT_0F => X"000000ab000000ad000000b1000000b3000000b3000000b4000000b7000000bd",
            INIT_10 => X"0000007700000082000000890000003800000013000000150000001400000015",
            INIT_11 => X"000000a7000000940000008b0000008400000092000000b3000000b20000009c",
            INIT_12 => X"000000d2000000ce000000a70000006d0000007800000098000000a9000000af",
            INIT_13 => X"000000ac000000b1000000b6000000ba000000bf000000c3000000c9000000d1",
            INIT_14 => X"0000007800000082000000730000002600000016000000170000001600000016",
            INIT_15 => X"000000840000006b0000006c000000760000009e000000c3000000b900000092",
            INIT_16 => X"000000c7000000be000000b70000008f00000084000000810000008f00000092",
            INIT_17 => X"000000c2000000c7000000ca000000d1000000d1000000cc000000d1000000cf",
            INIT_18 => X"00000094000000a1000000710000001e00000014000000150000001300000018",
            INIT_19 => X"00000071000000690000006200000080000000aa000000c2000000ba00000097",
            INIT_1A => X"000000c5000000c0000000ca000000b2000000800000006b0000007400000068",
            INIT_1B => X"000000da000000d7000000d6000000d8000000d7000000d1000000cf000000ce",
            INIT_1C => X"0000009c000000ba000000ae000000600000001d000000180000002900000058",
            INIT_1D => X"000000760000008100000084000000a4000000ba000000bd000000b500000095",
            INIT_1E => X"000000ce000000bb000000cc000000b40000007c0000006c0000006b0000005c",
            INIT_1F => X"000000e2000000dc000000d3000000cd000000e4000000e7000000e0000000e6",
            INIT_20 => X"00000093000000b7000000bd000000af000000750000006d00000099000000b1",
            INIT_21 => X"000000830000009a000000ad000000b8000000c0000000bc000000a100000078",
            INIT_22 => X"000000d8000000bc000000c5000000a60000007f000000770000007300000073",
            INIT_23 => X"000000e8000000e0000000c6000000bc000000d3000000e3000000e2000000e9",
            INIT_24 => X"00000090000000be000000c2000000bf000000b6000000af000000bc000000c2",
            INIT_25 => X"0000008a000000a4000000b6000000b7000000b6000000b10000009800000073",
            INIT_26 => X"000000e9000000d0000000bd000000a00000007b000000770000007600000066",
            INIT_27 => X"000000eb000000d1000000bd000000bb000000cb000000ea000000eb000000e8",
            INIT_28 => X"0000008a000000bf000000cd000000c6000000bb000000b7000000c0000000c7",
            INIT_29 => X"0000007c0000009a000000af000000b8000000b5000000b0000000a500000088",
            INIT_2A => X"000000f0000000cd000000b00000009e0000007800000077000000760000006b",
            INIT_2B => X"000000e0000000c6000000c0000000c0000000d4000000f2000000f4000000f3",
            INIT_2C => X"00000092000000bc000000d1000000c9000000bb000000c1000000c9000000c9",
            INIT_2D => X"0000006b000000840000009f000000b7000000b7000000b9000000b60000009b",
            INIT_2E => X"000000eb000000bd000000aa0000009e0000007e0000007c0000008500000073",
            INIT_2F => X"000000ca000000c0000000c0000000c2000000de000000f2000000f6000000f6",
            INIT_30 => X"000000a5000000b7000000c6000000c4000000bd000000c5000000c9000000cb",
            INIT_31 => X"000000780000008a000000a2000000a4000000a5000000b0000000aa0000009f",
            INIT_32 => X"000000e7000000bd000000a5000000a100000092000000870000009f00000085",
            INIT_33 => X"000000c7000000c1000000c3000000d0000000ea000000f7000000f8000000f4",
            INIT_34 => X"000000b90000009c000000a7000000c1000000b9000000c4000000ca000000d0",
            INIT_35 => X"0000008f000000890000009e000000a1000000870000008700000091000000a1",
            INIT_36 => X"000000e4000000c30000009d00000099000000a200000095000000a4000000a4",
            INIT_37 => X"000000de000000cc000000c7000000e8000000f5000000f9000000f7000000f2",
            INIT_38 => X"000000c10000007d0000008e000000bf000000b6000000c5000000cc000000d2",
            INIT_39 => X"0000007200000082000000aa000000b8000000a7000000a6000000b1000000b5",
            INIT_3A => X"000000e7000000bd000000ae000000ab0000009e00000098000000aa000000a5",
            INIT_3B => X"000000e9000000dd000000cf000000f2000000fb000000f5000000f4000000f2",
            INIT_3C => X"000000c00000007000000091000000bd000000b9000000c5000000c8000000d4",
            INIT_3D => X"00000089000000a0000000a7000000a4000000b4000000bd000000be000000c7",
            INIT_3E => X"000000c3000000a8000000b1000000b800000091000000a2000000b000000092",
            INIT_3F => X"000000eb000000ec000000dd000000e4000000f9000000f5000000f1000000e8",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE50;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE51 : if BRAM_NAME = "sampleifmap_layer0_instance51" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ad0000006e0000009b000000b0000000ae000000b6000000c7000000d8",
            INIT_01 => X"000000a4000000a70000009b000000a8000000b2000000a8000000ba000000d0",
            INIT_02 => X"0000006800000090000000ab0000009a00000086000000b1000000960000006e",
            INIT_03 => X"000000ed000000f3000000dd000000d2000000ed000000ee000000d100000091",
            INIT_04 => X"000000a200000095000000a7000000a30000009e000000a9000000ce000000db",
            INIT_05 => X"000000a1000000aa000000a8000000bc000000d1000000c8000000cd000000ca",
            INIT_06 => X"000000730000009b000000ba0000009300000087000000ad0000007800000070",
            INIT_07 => X"000000ef000000f3000000d4000000b9000000bc000000b20000008400000062",
            INIT_08 => X"000000b1000000b3000000b5000000af000000a1000000b3000000d6000000dd",
            INIT_09 => X"000000ab000000b8000000c5000000dc000000dd000000d4000000cf000000bd",
            INIT_0A => X"0000009300000094000000b1000000970000008c00000095000000670000008b",
            INIT_0B => X"000000ea000000d9000000b1000000970000009c0000008a0000007000000083",
            INIT_0C => X"000000c8000000be000000c2000000c2000000b2000000c6000000da000000df",
            INIT_0D => X"000000b1000000c8000000d0000000cb000000c7000000bf000000b8000000ba",
            INIT_0E => X"0000008f000000830000009b000000a80000009e0000007f00000087000000ab",
            INIT_0F => X"000000c50000009e00000090000000930000009f000000940000007e00000089",
            INIT_10 => X"000000c2000000be000000c7000000bf000000b7000000d0000000dd000000e1",
            INIT_11 => X"000000bf000000c6000000c1000000ab000000ba000000be000000bc000000c6",
            INIT_12 => X"0000008d0000007b00000087000000a0000000a900000094000000bf000000cf",
            INIT_13 => X"0000009a0000008c0000008800000087000000980000009f000000950000008e",
            INIT_14 => X"000000be000000c8000000c3000000b3000000be000000d6000000dd000000de",
            INIT_15 => X"000000b5000000b6000000b300000097000000b2000000d1000000cd000000c6",
            INIT_16 => X"00000093000000890000007c00000086000000a5000000ae000000c4000000c5",
            INIT_17 => X"0000007d0000008b0000008b000000830000008b00000099000000a100000099",
            INIT_18 => X"000000cf000000d2000000bf000000aa000000c6000000db000000da000000db",
            INIT_19 => X"000000b0000000b4000000ae0000009c000000b4000000cf000000ce000000cb",
            INIT_1A => X"00000098000000960000007d0000006f00000096000000b0000000b5000000b6",
            INIT_1B => X"0000006a00000073000000800000008a0000008a0000009a000000a100000098",
            INIT_1C => X"000000d5000000d2000000bc000000aa000000cf000000d9000000d6000000da",
            INIT_1D => X"000000b5000000ba000000ba000000ae000000b6000000c7000000d3000000d4",
            INIT_1E => X"000000950000009a000000890000007200000085000000ab000000b6000000ba",
            INIT_1F => X"00000076000000730000007b00000090000000920000009f000000ab00000094",
            INIT_20 => X"000000cd000000cf000000bd000000b3000000d1000000d4000000d4000000d8",
            INIT_21 => X"000000b6000000bb000000c3000000a70000008a000000b1000000cd000000cd",
            INIT_22 => X"0000008c000000960000008d0000007d000000820000009e000000b5000000b9",
            INIT_23 => X"0000007c000000820000008300000085000000950000009d000000a30000008d",
            INIT_24 => X"000000cc000000ce000000be000000bb000000c8000000d0000000d2000000d7",
            INIT_25 => X"000000ae000000b8000000c2000000910000005000000083000000c4000000c6",
            INIT_26 => X"000000880000008f0000008b000000780000008300000093000000a5000000ae",
            INIT_27 => X"00000070000000790000008500000085000000880000008c0000008e00000089",
            INIT_28 => X"000000d1000000cd000000b7000000b5000000c2000000cd000000d0000000d7",
            INIT_29 => X"000000a1000000ab000000ba0000008e0000005100000081000000c2000000cc",
            INIT_2A => X"0000007e000000890000008700000073000000780000008900000095000000a1",
            INIT_2B => X"0000008000000083000000880000008a0000007a000000700000007b00000085",
            INIT_2C => X"000000d4000000c6000000af000000b0000000bc000000c8000000cd000000d6",
            INIT_2D => X"000000950000009b000000a8000000aa0000008e000000a0000000c0000000d0",
            INIT_2E => X"0000007b000000800000008300000071000000640000007f000000850000008d",
            INIT_2F => X"00000089000000900000009000000082000000720000006c000000720000007e",
            INIT_30 => X"000000d2000000c0000000a6000000a9000000b7000000c0000000c4000000d2",
            INIT_31 => X"0000008c0000008d00000099000000ab000000b4000000b6000000c0000000d1",
            INIT_32 => X"0000007f0000007e0000007e000000780000005c0000006f0000007d00000086",
            INIT_33 => X"000000810000008d00000090000000850000007400000069000000720000007e",
            INIT_34 => X"000000cc000000b500000097000000a6000000b9000000b3000000b3000000c4",
            INIT_35 => X"000000880000008500000092000000a6000000b3000000ba000000c2000000cd",
            INIT_36 => X"00000080000000780000007300000078000000610000005d000000720000007e",
            INIT_37 => X"0000007b0000008200000083000000840000007e000000710000007100000080",
            INIT_38 => X"000000c30000009c0000008c000000ae000000b8000000aa000000a1000000b1",
            INIT_39 => X"000000730000006c0000007100000091000000b6000000bf000000c1000000c9",
            INIT_3A => X"000000830000007800000070000000720000006e000000590000006a00000076",
            INIT_3B => X"00000086000000820000007a000000750000007c0000007f0000007a0000007b",
            INIT_3C => X"000000b10000008000000082000000a6000000a1000000970000008c0000009d",
            INIT_3D => X"000000530000004700000053000000700000009a000000af000000b7000000bf",
            INIT_3E => X"0000007e000000790000006c0000006c0000006e000000650000005e00000063",
            INIT_3F => X"000000840000008900000084000000730000006b0000006f0000007a00000079",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE51;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE52 : if BRAM_NAME = "sampleifmap_layer0_instance52" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000740000006d000000730000007100000028000000130000001c00000017",
            INIT_01 => X"0000006b000000690000006900000069000000690000006a0000006700000071",
            INIT_02 => X"000000890000007200000056000000540000003a0000004c000000630000006a",
            INIT_03 => X"000000780000007a0000007d0000007f0000007d0000007c0000007d0000007c",
            INIT_04 => X"0000007c00000076000000820000006a0000001a000000140000001b00000018",
            INIT_05 => X"00000079000000720000007600000078000000750000006d000000720000007d",
            INIT_06 => X"000000960000008c000000510000003e000000440000006a0000008300000085",
            INIT_07 => X"0000008000000081000000850000008800000088000000890000008c0000008a",
            INIT_08 => X"0000007b00000074000000830000005800000012000000170000001a00000018",
            INIT_09 => X"000000840000007d0000007f0000008100000074000000740000008d0000008b",
            INIT_0A => X"0000009e0000009f000000590000003700000069000000980000009a0000008e",
            INIT_0B => X"00000084000000880000008b0000008e0000008e000000920000009700000097",
            INIT_0C => X"000000730000006a0000007c0000004500000012000000190000001900000018",
            INIT_0D => X"000000970000009500000094000000890000007800000092000000a60000009c",
            INIT_0E => X"000000a9000000b10000007a0000004a0000006d000000940000009c00000096",
            INIT_0F => X"0000008e00000091000000940000009600000095000000980000009d000000a1",
            INIT_10 => X"00000068000000600000006d0000003300000017000000190000001800000019",
            INIT_11 => X"0000009300000086000000800000007c0000008d000000b2000000b8000000a1",
            INIT_12 => X"000000b5000000b700000098000000600000006c000000890000009600000097",
            INIT_13 => X"00000093000000980000009c000000a0000000a4000000a8000000ae000000b3",
            INIT_14 => X"000000660000005f00000059000000230000001c0000001b0000001a0000001a",
            INIT_15 => X"000000760000006200000066000000740000009f000000c7000000c100000096",
            INIT_16 => X"000000aa000000a6000000a7000000840000007a000000770000008300000082",
            INIT_17 => X"000000a9000000af000000b1000000b7000000b7000000b3000000b7000000b2",
            INIT_18 => X"0000007b000000800000005c0000001d0000001a00000019000000160000001a",
            INIT_19 => X"0000006a000000630000005e0000007e000000ab000000c7000000c300000093",
            INIT_1A => X"000000b0000000aa000000c0000000ac0000007a000000650000006d00000060",
            INIT_1B => X"000000c2000000bf000000bf000000c5000000ca000000c5000000c4000000c3",
            INIT_1C => X"0000007e0000009b0000009a000000580000001900000011000000210000004d",
            INIT_1D => X"000000710000007b00000081000000a3000000b9000000c1000000be0000008c",
            INIT_1E => X"000000bd000000a5000000c6000000b100000079000000680000006700000058",
            INIT_1F => X"000000cd000000c4000000bb000000ba000000da000000e0000000db000000e4",
            INIT_20 => X"0000007700000099000000a70000009b00000060000000560000008000000095",
            INIT_21 => X"0000007f00000094000000aa000000b7000000bf000000bf000000a80000006f",
            INIT_22 => X"000000c1000000a2000000bb000000a30000007c000000740000007000000070",
            INIT_23 => X"000000d2000000c4000000a60000009d000000bb000000cf000000d5000000df",
            INIT_24 => X"000000750000009f000000a9000000a70000009b000000920000009e000000a1",
            INIT_25 => X"000000870000009f000000b4000000b6000000b5000000b30000009b00000068",
            INIT_26 => X"000000cc000000b2000000b20000009e00000079000000750000007400000064",
            INIT_27 => X"000000cf000000b00000009600000093000000a7000000cb000000d6000000d8",
            INIT_28 => X"00000070000000a0000000b0000000af000000a50000009e000000a5000000aa",
            INIT_29 => X"0000007900000095000000ac000000b6000000b4000000b1000000a40000007b",
            INIT_2A => X"000000d1000000af000000a60000009c0000007600000075000000740000006a",
            INIT_2B => X"000000ba0000009f0000009300000091000000a9000000cd000000d8000000de",
            INIT_2C => X"0000007a0000009d000000b0000000b0000000a6000000a9000000ae000000ac",
            INIT_2D => X"000000680000007f0000009d000000b6000000b6000000b9000000b10000008d",
            INIT_2E => X"000000ce000000a3000000a40000009f0000007d0000007b0000008400000073",
            INIT_2F => X"0000009c000000930000008e00000092000000b5000000cd000000d9000000e0",
            INIT_30 => X"0000008f00000099000000a4000000a5000000a0000000a5000000a7000000a7",
            INIT_31 => X"00000076000000850000009f000000a3000000a4000000ae000000a300000091",
            INIT_32 => X"000000cd000000a8000000a3000000a300000092000000870000009f00000086",
            INIT_33 => X"000000980000009000000090000000a3000000c7000000d6000000dc000000df",
            INIT_34 => X"000000a40000008300000088000000a30000009b000000a0000000a2000000a9",
            INIT_35 => X"00000092000000870000009e0000009f00000085000000840000008800000092",
            INIT_36 => X"000000cb000000b000000098000000980000009e00000090000000a2000000a7",
            INIT_37 => X"000000b6000000a20000009f000000c5000000da000000dd000000d8000000d7",
            INIT_38 => X"000000b20000006d00000078000000a80000009d000000a2000000a4000000ae",
            INIT_39 => X"0000007800000084000000ab000000b6000000a3000000a1000000a7000000a6",
            INIT_3A => X"000000cc000000aa000000a4000000a6000000950000008c000000a3000000a9",
            INIT_3B => X"000000c7000000bb000000b0000000d6000000e4000000da000000d5000000d3",
            INIT_3C => X"000000b70000006800000084000000aa0000009f000000a1000000a0000000af",
            INIT_3D => X"0000008d000000a3000000a8000000a2000000b0000000b8000000b6000000bc",
            INIT_3E => X"000000a900000096000000a5000000af0000008500000092000000a500000091",
            INIT_3F => X"000000c7000000c7000000ba000000c4000000dd000000d9000000d4000000ca",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE52;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE53 : if BRAM_NAME = "sampleifmap_layer0_instance53" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a80000006d00000097000000a100000094000000920000009f000000b3",
            INIT_01 => X"000000a6000000aa0000009c000000a5000000ae000000a4000000b5000000c7",
            INIT_02 => X"000000500000007e0000009e0000008f000000770000009f0000008800000069",
            INIT_03 => X"000000c5000000c9000000b7000000af000000cd000000d1000000b700000076",
            INIT_04 => X"0000009f00000097000000a5000000950000008300000085000000a4000000b5",
            INIT_05 => X"000000a2000000ac000000a8000000b9000000cd000000c4000000c7000000c2",
            INIT_06 => X"0000005c00000088000000ad00000086000000770000009b0000006900000068",
            INIT_07 => X"000000c8000000cb000000b0000000980000009e000000980000006f0000004b",
            INIT_08 => X"000000aa000000b1000000b00000009f000000850000008e000000ac000000b7",
            INIT_09 => X"000000aa000000bb000000c6000000d9000000d9000000cf000000c5000000b1",
            INIT_0A => X"0000007e00000082000000a20000008b0000007e000000850000005a00000083",
            INIT_0B => X"000000c7000000b8000000920000007c0000008400000076000000600000006f",
            INIT_0C => X"000000bc000000b6000000b7000000af00000095000000a1000000b0000000b9",
            INIT_0D => X"000000af000000ca000000d0000000c9000000c2000000b9000000aa000000aa",
            INIT_0E => X"0000007b000000710000008c0000009d00000091000000710000007b000000a4",
            INIT_0F => X"000000a600000084000000790000007f0000008e000000860000007000000077",
            INIT_10 => X"000000b2000000b1000000ba000000ab0000009b000000ad000000b7000000bd",
            INIT_11 => X"000000bd000000c3000000bc000000a4000000b1000000b2000000ac000000b4",
            INIT_12 => X"0000007c0000006a00000078000000930000009d00000088000000b6000000c9",
            INIT_13 => X"000000820000007a00000077000000780000008a000000940000008a00000080",
            INIT_14 => X"000000b0000000bb000000b70000009e000000a1000000b7000000bc000000bd",
            INIT_15 => X"000000b1000000ad000000a60000008b000000a4000000c0000000bf000000b8",
            INIT_16 => X"00000085000000790000006b0000007600000096000000a2000000bc000000c0",
            INIT_17 => X"0000006c0000007d0000007c000000750000007d0000008d000000960000008e",
            INIT_18 => X"000000c5000000c7000000b400000094000000a6000000bb000000ba000000ba",
            INIT_19 => X"000000aa000000a90000009f00000091000000a8000000c0000000c3000000c1",
            INIT_1A => X"0000008b000000860000006c0000005d00000086000000a3000000ac000000af",
            INIT_1B => X"0000005b00000065000000720000007c0000007c0000008e000000970000008d",
            INIT_1C => X"000000cf000000c9000000b00000008f000000ac000000b7000000b5000000ba",
            INIT_1D => X"000000ac000000ae000000ab000000a5000000af000000bd000000cb000000ce",
            INIT_1E => X"000000880000008a0000007800000061000000750000009e000000ab000000b2",
            INIT_1F => X"00000068000000640000006d000000820000008400000092000000a10000008a",
            INIT_20 => X"000000ca000000c6000000aa00000092000000a9000000af000000b2000000b8",
            INIT_21 => X"000000aa000000ab000000b4000000a100000088000000ab000000c5000000c8",
            INIT_22 => X"0000007e000000860000007c0000006c0000007300000090000000a8000000ad",
            INIT_23 => X"0000006f00000074000000750000007700000087000000910000009900000082",
            INIT_24 => X"000000c8000000c0000000a2000000930000009d000000a8000000b0000000b8",
            INIT_25 => X"0000009f000000a6000000b30000008d0000005200000081000000b9000000bf",
            INIT_26 => X"0000007a0000007f0000007a000000690000007400000084000000960000009f",
            INIT_27 => X"000000620000006b00000077000000770000007a00000080000000840000007f",
            INIT_28 => X"000000ca000000ba000000920000008600000094000000a3000000ac000000b8",
            INIT_29 => X"0000009000000098000000ac0000008c0000005800000082000000b2000000c0",
            INIT_2A => X"00000070000000790000007700000064000000690000007a0000008400000091",
            INIT_2B => X"00000072000000750000007a0000007c0000006c00000064000000710000007a",
            INIT_2C => X"000000cc000000b2000000840000007e0000008e0000009e000000a9000000b7",
            INIT_2D => X"000000830000008700000098000000a4000000900000009d000000af000000c3",
            INIT_2E => X"0000006d000000710000007300000061000000540000006f000000740000007c",
            INIT_2F => X"0000007b000000820000008200000074000000640000005f0000006600000072",
            INIT_30 => X"000000cc000000b20000007a000000770000008e00000099000000a1000000b1",
            INIT_31 => X"0000007b0000007a000000870000009d000000a8000000aa000000b4000000c5",
            INIT_32 => X"00000071000000700000006f000000680000004b0000005e0000006d00000077",
            INIT_33 => X"000000730000007e0000008200000077000000660000005c0000006400000070",
            INIT_34 => X"000000c8000000a90000006b00000074000000910000008d00000090000000a3",
            INIT_35 => X"00000079000000730000008100000096000000a3000000ac000000b7000000c2",
            INIT_36 => X"000000720000006a0000006500000068000000510000004e0000006400000070",
            INIT_37 => X"0000006e00000074000000750000007600000070000000630000006300000072",
            INIT_38 => X"000000c0000000910000005f0000007c0000008f000000830000007e0000008e",
            INIT_39 => X"000000650000005c0000006200000082000000a8000000b2000000b7000000be",
            INIT_3A => X"000000740000006a00000061000000630000005f0000004b0000005c00000068",
            INIT_3B => X"00000077000000740000006c000000670000006e000000710000006c0000006d",
            INIT_3C => X"000000ae0000007600000057000000740000007800000070000000680000007b",
            INIT_3D => X"000000460000003900000045000000630000008d000000a4000000ae000000b5",
            INIT_3E => X"000000700000006b0000005e0000005d00000060000000580000005100000057",
            INIT_3F => X"000000760000007b00000076000000650000005d000000610000006c0000006b",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE53;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE54 : if BRAM_NAME = "sampleifmap_layer0_instance54" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000bd000000cf000000d6000000da000000c7000000cd000000d2000000d9",
            INIT_01 => X"0000008f0000008c0000009a00000096000000a9000000a6000000ae000000bb",
            INIT_02 => X"000000e1000000e2000000d7000000db000000df000000db000000bf000000a7",
            INIT_03 => X"000000a2000000a1000000aa000000c8000000bb000000af000000be000000db",
            INIT_04 => X"000000b3000000d3000000e1000000d8000000d7000000dc000000dd000000de",
            INIT_05 => X"000000db000000d1000000ce000000c7000000bc000000be000000c0000000b4",
            INIT_06 => X"000000e5000000e1000000e2000000e9000000ec000000ec000000eb000000e5",
            INIT_07 => X"000000c8000000ba000000b7000000d8000000cd000000d0000000d4000000e7",
            INIT_08 => X"000000ad000000d9000000ef000000e9000000e8000000e7000000e9000000ea",
            INIT_09 => X"000000e0000000d4000000bc000000be000000b7000000ad000000b4000000a4",
            INIT_0A => X"000000e1000000d6000000df000000e5000000e1000000e3000000eb000000da",
            INIT_0B => X"000000d3000000d0000000ca000000d1000000d8000000e6000000e8000000ea",
            INIT_0C => X"0000009e000000e4000000f3000000f4000000f2000000f4000000f4000000f5",
            INIT_0D => X"0000009f000000a200000088000000910000009f000000830000009d00000092",
            INIT_0E => X"000000e2000000d0000000cb000000d1000000d3000000c3000000cb000000a9",
            INIT_0F => X"000000d4000000e0000000db000000c7000000d5000000e4000000e9000000e6",
            INIT_10 => X"00000075000000cf000000f1000000f5000000f4000000f4000000f3000000f5",
            INIT_11 => X"0000005c000000640000005b000000640000006b000000590000006c00000063",
            INIT_12 => X"000000e9000000ca000000b9000000b6000000950000007c0000007c00000066",
            INIT_13 => X"000000de000000e2000000d5000000c2000000cd000000e3000000e2000000e1",
            INIT_14 => X"0000007e000000d8000000ed000000f5000000f3000000f4000000f4000000f5",
            INIT_15 => X"000000630000006b0000006700000065000000660000005b0000005a00000048",
            INIT_16 => X"000000eb000000d8000000be0000007e0000005d0000005b0000005900000059",
            INIT_17 => X"000000ec000000d9000000bd000000ae000000c4000000d8000000df000000e7",
            INIT_18 => X"0000009e000000d9000000db000000f1000000f4000000f3000000f3000000f5",
            INIT_19 => X"0000008a0000008f000000840000008c00000097000000840000007200000050",
            INIT_1A => X"000000e9000000dd0000009b0000006e00000078000000720000007a00000082",
            INIT_1B => X"000000eb000000cc000000ab000000a7000000c0000000c6000000e0000000eb",
            INIT_1C => X"00000099000000d7000000c7000000e3000000f6000000f3000000f3000000f4",
            INIT_1D => X"00000083000000830000009e000000cf000000ca000000bb0000009200000051",
            INIT_1E => X"000000d70000009f000000840000009f00000084000000830000008d00000081",
            INIT_1F => X"000000dd000000b2000000ab000000c5000000d1000000d4000000d7000000e5",
            INIT_20 => X"00000082000000da000000ce000000e3000000f5000000f4000000f3000000f4",
            INIT_21 => X"0000007d0000007400000091000000b800000081000000800000008200000051",
            INIT_22 => X"000000c60000009000000093000000990000007d0000008e000000890000007c",
            INIT_23 => X"000000c9000000a9000000a4000000b8000000dc000000e9000000db000000d6",
            INIT_24 => X"0000006e000000a8000000be000000e4000000f2000000f4000000f3000000f3",
            INIT_25 => X"0000007800000073000000800000008f0000006e000000770000008600000053",
            INIT_26 => X"000000c40000008c0000009b000000950000007d00000092000000830000007d",
            INIT_27 => X"000000dc000000d7000000c8000000c8000000e9000000f0000000f0000000e9",
            INIT_28 => X"0000005f0000008200000085000000dc000000f5000000f4000000f1000000ef",
            INIT_29 => X"0000006c0000006d0000006b0000006d0000006c00000074000000740000004e",
            INIT_2A => X"000000a70000008f000000960000008800000073000000780000007800000073",
            INIT_2B => X"000000f4000000f5000000f5000000f4000000f3000000f5000000e4000000d0",
            INIT_2C => X"00000059000000a5000000a9000000d8000000f4000000f2000000e9000000de",
            INIT_2D => X"00000060000000620000005f0000005f000000640000005b000000430000003d",
            INIT_2E => X"0000007e000000810000007900000069000000610000005a0000005f00000060",
            INIT_2F => X"000000f4000000f4000000f4000000f4000000f3000000f8000000d80000009b",
            INIT_30 => X"00000064000000b5000000b7000000bf000000e3000000ec000000df000000d0",
            INIT_31 => X"0000005400000056000000630000006f00000065000000580000003800000037",
            INIT_32 => X"0000008100000070000000620000006d000000710000005d0000005400000052",
            INIT_33 => X"000000f4000000f4000000f4000000f4000000f4000000f5000000e2000000ae",
            INIT_34 => X"000000660000009c0000009a000000aa000000c3000000db000000cc000000c8",
            INIT_35 => X"000000550000005e0000007500000073000000660000006c0000006300000068",
            INIT_36 => X"0000007c0000006c00000068000000800000008c0000007a0000006a0000005a",
            INIT_37 => X"000000f4000000f4000000f5000000ef000000d4000000c3000000b300000096",
            INIT_38 => X"0000008a0000009300000094000000a4000000a9000000cf000000d2000000c8",
            INIT_39 => X"0000004d000000540000005d000000590000005d0000006a0000005c00000081",
            INIT_3A => X"000000520000004b0000004a0000004f0000005100000051000000510000004c",
            INIT_3B => X"000000f4000000f4000000f4000000bf0000008f0000008c0000007b00000065",
            INIT_3C => X"000000c0000000ba000000960000007000000077000000c4000000e2000000d2",
            INIT_3D => X"0000003f0000003c0000002f0000002d000000370000004d0000004d0000006c",
            INIT_3E => X"000000400000003d0000003200000031000000360000003b0000003f0000003b",
            INIT_3F => X"000000f4000000f6000000e100000087000000670000005b0000004b00000047",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE54;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE55 : if BRAM_NAME = "sampleifmap_layer0_instance55" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a1000000c0000000910000005d00000060000000b4000000c1000000c7",
            INIT_01 => X"000000470000004f0000004f00000068000000620000005c0000004900000056",
            INIT_02 => X"0000001c0000001600000032000000340000001b0000001e0000001c00000025",
            INIT_03 => X"000000f3000000f7000000ce00000080000000680000005b0000003500000018",
            INIT_04 => X"000000470000009f0000009d0000007800000071000000c2000000c7000000d3",
            INIT_05 => X"000000660000008000000079000000950000007c000000740000005a00000044",
            INIT_06 => X"000000630000005c00000093000000940000006400000070000000620000004e",
            INIT_07 => X"000000f5000000f2000000b70000009c0000008e000000870000006c0000005e",
            INIT_08 => X"0000001e00000084000000a50000006e00000066000000b7000000ca000000dc",
            INIT_09 => X"00000064000000810000006500000052000000530000006b0000006200000039",
            INIT_0A => X"000000a3000000a2000000a8000000ac0000009f0000009e000000ae00000099",
            INIT_0B => X"000000f7000000e40000008700000072000000770000009c000000af000000a0",
            INIT_0C => X"0000002a0000006f0000008d0000005300000062000000bc000000cf000000db",
            INIT_0D => X"0000005d0000004000000038000000350000003e0000004c000000480000003a",
            INIT_0E => X"00000067000000670000006b00000074000000650000005b0000007c000000a0",
            INIT_0F => X"000000f8000000d90000007600000051000000430000007e0000009b00000063",
            INIT_10 => X"0000003c0000005d000000580000003800000065000000c7000000d2000000d9",
            INIT_11 => X"0000004100000040000000360000003c000000460000003f0000002e00000038",
            INIT_12 => X"000000610000005d000000600000006400000067000000690000007200000063",
            INIT_13 => X"000000f9000000d4000000720000005200000049000000640000006f00000066",
            INIT_14 => X"0000004400000051000000460000005300000075000000ca000000cd000000d1",
            INIT_15 => X"0000003f000000570000004d00000044000000330000002b0000002300000032",
            INIT_16 => X"0000005d0000003e000000430000004000000048000000520000004700000034",
            INIT_17 => X"000000fa000000cc0000006c000000700000006c000000530000003c00000058",
            INIT_18 => X"00000049000000470000006f0000005d00000068000000c5000000ca000000cd",
            INIT_19 => X"0000004f0000008e000000630000004b0000002200000026000000290000003f",
            INIT_1A => X"000000990000006600000072000000630000007600000093000000560000001e",
            INIT_1B => X"000000f6000000c30000005a000000770000008d0000004a0000003f000000b2",
            INIT_1C => X"00000063000000610000006c0000003100000057000000b9000000c2000000c6",
            INIT_1D => X"000000370000005700000032000000280000002400000027000000330000005f",
            INIT_1E => X"0000009c00000074000000880000007a0000007f000000970000004f00000020",
            INIT_1F => X"000000f0000000c20000004e0000003e0000004a00000035000000370000009f",
            INIT_20 => X"000000900000006c0000003b000000250000004d000000a9000000b4000000b6",
            INIT_21 => X"000000210000001e0000001c0000001d000000200000002b0000003c0000006a",
            INIT_22 => X"000000750000007a000000790000006a000000580000003a0000002a00000027",
            INIT_23 => X"000000e1000000ba000000500000003300000032000000330000002f00000043",
            INIT_24 => X"0000008d0000006f000000600000005b0000007d000000a4000000a5000000a8",
            INIT_25 => X"0000001f0000001d0000001e0000001e00000024000000370000004a00000060",
            INIT_26 => X"000000b5000000b3000000cb000000cd000000ae000000400000001800000023",
            INIT_27 => X"000000d3000000ae0000005b00000042000000300000002b0000002600000057",
            INIT_28 => X"0000008d0000006c0000007600000098000000b4000000af000000a3000000a2",
            INIT_29 => X"0000001d000000190000001800000019000000300000004e000000530000005b",
            INIT_2A => X"000000a6000000a9000000b1000000b8000000a4000000470000002600000027",
            INIT_2B => X"000000ce000000a90000005f0000004e000000310000001e0000001e00000051",
            INIT_2C => X"00000092000000670000007500000092000000a6000000b3000000ac0000009a",
            INIT_2D => X"00000025000000210000001e0000002000000036000000520000005500000057",
            INIT_2E => X"000000890000008e000000790000006b00000065000000560000004d00000036",
            INIT_2F => X"000000c7000000a50000005b0000004e00000036000000210000001e0000003c",
            INIT_30 => X"0000007100000067000000850000008f000000940000009e000000a9000000a6",
            INIT_31 => X"0000002c0000002a000000270000002a0000003c0000004b000000510000004f",
            INIT_32 => X"0000008b000000830000006e0000005a0000004d000000410000003600000030",
            INIT_33 => X"000000c4000000a90000005b0000004600000036000000260000001d00000035",
            INIT_34 => X"0000004e0000006b00000085000000890000008d0000009300000097000000a2",
            INIT_35 => X"000000300000002e0000002a000000320000003c000000460000004e00000048",
            INIT_36 => X"0000007100000065000000590000004c000000420000003b0000003300000031",
            INIT_37 => X"000000ba000000ae000000620000003f00000034000000230000001d00000045",
            INIT_38 => X"0000003c0000006a0000008c0000008f0000008c0000008e0000008d00000094",
            INIT_39 => X"0000003a00000036000000340000003900000037000000420000004a00000042",
            INIT_3A => X"0000005d00000057000000500000004900000046000000410000003a0000003a",
            INIT_3B => X"000000b4000000b3000000830000004a0000003700000026000000250000004d",
            INIT_3C => X"0000003d0000007e000000920000009e000000a2000000a00000009500000090",
            INIT_3D => X"00000048000000490000004500000046000000430000003a0000003900000039",
            INIT_3E => X"0000006100000063000000610000005e00000062000000590000004900000044",
            INIT_3F => X"000000ba000000b6000000a40000007700000047000000400000004500000052",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE55;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE56 : if BRAM_NAME = "sampleifmap_layer0_instance56" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b9000000ca000000d1000000d7000000ca000000d0000000d0000000d7",
            INIT_01 => X"0000009d0000009a000000a70000009d000000a000000098000000a8000000b8",
            INIT_02 => X"000000e4000000e5000000db000000de000000e1000000e1000000cb000000b5",
            INIT_03 => X"000000a5000000b0000000b8000000d0000000c4000000b8000000c5000000dd",
            INIT_04 => X"000000ab000000cc000000dd000000d5000000d9000000e1000000e0000000e2",
            INIT_05 => X"000000e0000000d0000000cd000000c4000000b1000000b2000000bd000000b4",
            INIT_06 => X"000000e7000000e4000000e5000000ee000000f3000000f2000000f0000000ec",
            INIT_07 => X"000000c5000000bf000000be000000de000000d2000000d4000000d6000000e7",
            INIT_08 => X"000000a6000000d6000000ef000000ea000000eb000000ea000000ea000000eb",
            INIT_09 => X"000000df000000ce000000b7000000b8000000b1000000a8000000b1000000a6",
            INIT_0A => X"000000e0000000d9000000e4000000eb000000e8000000e3000000ec000000dc",
            INIT_0B => X"000000d2000000d1000000ce000000d9000000dd000000e6000000e9000000e9",
            INIT_0C => X"00000099000000e3000000f4000000f4000000f3000000f4000000f4000000f5",
            INIT_0D => X"000000a0000000a20000008a000000900000009f000000820000009b00000092",
            INIT_0E => X"000000e0000000d3000000d3000000de000000dc000000c2000000cd000000ac",
            INIT_0F => X"000000d4000000e2000000df000000cf000000db000000e5000000e9000000e6",
            INIT_10 => X"00000070000000cd000000f0000000f5000000f4000000f4000000f4000000f5",
            INIT_11 => X"0000005c000000640000005c000000650000006d0000005b0000006d00000062",
            INIT_12 => X"000000e3000000c9000000c2000000c20000009a0000007c0000007d00000068",
            INIT_13 => X"000000e1000000e8000000dc000000cb000000d3000000e3000000de000000dc",
            INIT_14 => X"0000007b000000d4000000eb000000f6000000f3000000f4000000f4000000f5",
            INIT_15 => X"000000660000006e0000006a00000067000000690000005f0000005d00000047",
            INIT_16 => X"000000e6000000d9000000c5000000810000005d0000005b000000590000005b",
            INIT_17 => X"000000ed000000e2000000c5000000b4000000c6000000d6000000da000000dd",
            INIT_18 => X"0000009c000000d5000000d6000000f0000000f4000000f3000000f3000000f5",
            INIT_19 => X"000000960000009b0000008b000000900000009a00000089000000770000004f",
            INIT_1A => X"000000e9000000e1000000a0000000720000007e00000079000000800000008e",
            INIT_1B => X"000000ec000000d4000000b0000000a5000000ba000000c0000000da000000e9",
            INIT_1C => X"00000096000000d3000000c1000000e2000000f7000000f3000000f3000000f4",
            INIT_1D => X"000000900000008d000000a5000000cd000000c8000000bc0000009800000051",
            INIT_1E => X"000000d6000000a30000008c000000a70000008f0000008d000000960000008e",
            INIT_1F => X"000000dc000000af000000ae000000c7000000d2000000d3000000d1000000e0",
            INIT_20 => X"0000007f000000d8000000ca000000e1000000f5000000f4000000f3000000f4",
            INIT_21 => X"000000870000007c00000097000000b900000087000000840000008600000051",
            INIT_22 => X"000000c00000008e0000009e000000a400000088000000960000009100000086",
            INIT_23 => X"000000c40000009c0000009e000000b1000000d7000000e7000000d8000000cf",
            INIT_24 => X"0000006e000000a8000000bd000000e3000000f2000000f4000000f2000000f2",
            INIT_25 => X"000000810000007c000000870000009300000076000000800000008c00000053",
            INIT_26 => X"000000c100000091000000a40000009e00000086000000970000008b00000085",
            INIT_27 => X"000000d7000000cc000000be000000c1000000e6000000ef000000ef000000e5",
            INIT_28 => X"0000005e0000008000000081000000da000000f4000000f3000000ef000000e8",
            INIT_29 => X"00000073000000730000007000000071000000700000007a0000007a0000004f",
            INIT_2A => X"000000aa000000990000009e000000900000007e0000007f000000800000007c",
            INIT_2B => X"000000f4000000f5000000f3000000f3000000f4000000f6000000e3000000ce",
            INIT_2C => X"000000580000009f000000a1000000d3000000f2000000f2000000e3000000cd",
            INIT_2D => X"00000066000000670000006100000062000000660000005e000000450000003c",
            INIT_2E => X"00000080000000890000007f00000071000000670000005f0000006400000068",
            INIT_2F => X"000000f4000000f4000000f4000000f4000000f3000000f8000000d700000099",
            INIT_30 => X"00000063000000ad000000aa000000b4000000dc000000e4000000d5000000bc",
            INIT_31 => X"00000055000000580000006700000072000000660000005a0000003900000037",
            INIT_32 => X"00000086000000760000006500000070000000730000005d0000005500000055",
            INIT_33 => X"000000f4000000f4000000f4000000f4000000f4000000f5000000e1000000b0",
            INIT_34 => X"000000630000008d0000008600000098000000b5000000ca000000bc000000b8",
            INIT_35 => X"00000056000000600000007800000076000000670000006f0000006600000067",
            INIT_36 => X"0000007f0000006e0000006a00000084000000920000007d0000006b0000005c",
            INIT_37 => X"000000f4000000f4000000f5000000ee000000d2000000c3000000b300000098",
            INIT_38 => X"0000007e0000007f0000007b0000009200000098000000bd000000c2000000b6",
            INIT_39 => X"0000004f000000550000005d0000005a0000005e000000690000005d0000007c",
            INIT_3A => X"000000530000004c0000004b000000510000005500000054000000530000004e",
            INIT_3B => X"000000f4000000f4000000f4000000bc0000008a0000008a0000007a00000065",
            INIT_3C => X"000000ae000000a90000007d0000006500000065000000a7000000cc000000bd",
            INIT_3D => X"0000003e0000003b0000002f0000002b000000360000004f0000004d00000067",
            INIT_3E => X"000000400000003d000000300000002f00000034000000390000003e0000003b",
            INIT_3F => X"000000f4000000f6000000df00000080000000610000005a0000004a00000046",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE56;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE57 : if BRAM_NAME = "sampleifmap_layer0_instance57" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000092000000ac0000007c000000520000005400000097000000a4000000ae",
            INIT_01 => X"000000440000004c0000004b000000640000005a000000570000004900000053",
            INIT_02 => X"00000019000000140000002f00000030000000170000001a0000001700000021",
            INIT_03 => X"000000f3000000f7000000ca0000007800000064000000560000003200000015",
            INIT_04 => X"000000400000008e000000870000006800000068000000b3000000b4000000c0",
            INIT_05 => X"000000620000007d0000007600000095000000780000006c0000005700000041",
            INIT_06 => X"00000060000000590000009000000090000000600000006a0000005900000046",
            INIT_07 => X"000000f4000000f1000000b2000000970000008b00000082000000670000005a",
            INIT_08 => X"0000001c0000007600000092000000620000005e000000ab000000bd000000d1",
            INIT_09 => X"0000005f0000008000000064000000530000004f000000670000005f00000036",
            INIT_0A => X"000000a1000000a0000000a8000000ab0000009e0000009b000000aa00000092",
            INIT_0B => X"000000f7000000e2000000800000006f000000770000009b000000ac0000009e",
            INIT_0C => X"00000028000000640000007f0000004c0000005b000000b0000000c1000000d0",
            INIT_0D => X"000000590000003d000000350000003200000039000000490000004400000035",
            INIT_0E => X"000000640000006300000068000000710000006200000057000000770000009c",
            INIT_0F => X"000000f8000000d6000000700000004d0000003f0000007a0000009800000060",
            INIT_10 => X"00000038000000530000004e000000330000005f000000be000000c3000000ca",
            INIT_11 => X"0000003d0000003b0000003300000039000000440000003c0000002700000033",
            INIT_12 => X"000000600000005c0000005f0000006300000065000000660000006e0000005f",
            INIT_13 => X"000000f9000000d00000006c0000004f00000046000000600000006c00000064",
            INIT_14 => X"0000003f000000490000003e0000004c0000006e000000c0000000c0000000c2",
            INIT_15 => X"0000003b00000053000000480000004100000030000000280000001d0000002e",
            INIT_16 => X"000000580000003b000000400000003c000000430000004d0000004300000030",
            INIT_17 => X"000000f9000000c9000000650000006b000000690000004e0000003600000052",
            INIT_18 => X"0000004300000041000000630000005500000061000000bb000000be000000c3",
            INIT_19 => X"0000004c0000008d00000060000000480000002000000023000000260000003a",
            INIT_1A => X"00000092000000610000006d0000005e000000710000008c0000004f00000019",
            INIT_1B => X"000000f4000000c000000053000000740000008a000000450000003a000000ab",
            INIT_1C => X"0000005e00000059000000630000002c00000052000000b0000000b7000000bd",
            INIT_1D => X"00000034000000550000002f000000260000002100000024000000300000005a",
            INIT_1E => X"000000970000007100000086000000770000007b000000910000004a0000001c",
            INIT_1F => X"000000ee000000c0000000470000003b0000004700000032000000330000009c",
            INIT_20 => X"0000008b00000065000000360000002200000048000000a3000000ad000000ae",
            INIT_21 => X"0000001e0000001a000000190000001a0000001e000000280000003a00000066",
            INIT_22 => X"0000007200000076000000750000006800000056000000350000002600000025",
            INIT_23 => X"000000df000000b80000004b0000002f0000002e000000300000002b0000003e",
            INIT_24 => X"00000088000000670000005900000057000000780000009e000000a0000000a2",
            INIT_25 => X"0000001d0000001b0000001b0000001c0000002200000034000000480000005c",
            INIT_26 => X"000000b4000000b1000000ca000000cf000000af0000003d0000001500000020",
            INIT_27 => X"000000d1000000ab000000570000003e0000002c000000280000002200000054",
            INIT_28 => X"00000088000000660000007000000093000000b0000000a80000009c0000009c",
            INIT_29 => X"0000001a0000001700000016000000160000002d0000004b0000005100000056",
            INIT_2A => X"000000a5000000a9000000b1000000b9000000a4000000450000002200000023",
            INIT_2B => X"000000cc000000a70000005c0000004b0000002d0000001a000000190000004e",
            INIT_2C => X"0000008e00000063000000710000008d000000a1000000ad000000a700000095",
            INIT_2D => X"000000220000001f0000001c0000001d000000330000004f0000005300000053",
            INIT_2E => X"000000850000008a000000740000006600000061000000510000004800000032",
            INIT_2F => X"000000c6000000a4000000590000004c000000320000001d0000001b00000037",
            INIT_30 => X"0000006c00000063000000820000008b000000900000009b000000a6000000a4",
            INIT_31 => X"000000290000002700000024000000260000003800000048000000500000004c",
            INIT_32 => X"000000830000007c0000006700000054000000480000003d000000330000002d",
            INIT_33 => X"000000c3000000a9000000590000004500000032000000210000001a00000031",
            INIT_34 => X"000000490000006600000082000000870000008d0000009200000094000000a0",
            INIT_35 => X"0000002d0000002b000000280000002f00000038000000420000004d00000045",
            INIT_36 => X"0000006a0000005e00000054000000460000003d00000036000000300000002e",
            INIT_37 => X"000000ba000000af000000620000003d000000300000001f0000001a00000040",
            INIT_38 => X"00000039000000680000008b0000008f0000008c0000008e0000008d00000093",
            INIT_39 => X"00000036000000330000003100000037000000340000003f0000004a00000040",
            INIT_3A => X"00000057000000510000004a00000044000000420000003d0000003600000036",
            INIT_3B => X"000000b5000000b6000000840000004800000034000000230000002100000048",
            INIT_3C => X"0000003a0000007c000000910000009d000000a3000000a10000009600000092",
            INIT_3D => X"0000004500000046000000420000004300000041000000390000003800000037",
            INIT_3E => X"0000005e000000600000005f0000005c0000005f000000570000004800000043",
            INIT_3F => X"000000b9000000b6000000a300000076000000460000003e0000004400000051",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE57;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE58 : if BRAM_NAME = "sampleifmap_layer0_instance58" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000af000000c6000000d1000000d1000000b6000000bf000000ca000000d1",
            INIT_01 => X"0000008f0000008d0000009a00000095000000a00000009d000000a5000000ab",
            INIT_02 => X"000000d6000000d9000000ca000000d1000000db000000d6000000bc000000a4",
            INIT_03 => X"00000095000000950000009d000000b7000000ad000000a1000000b1000000d0",
            INIT_04 => X"000000a3000000c8000000db000000cf000000cd000000d2000000d4000000d4",
            INIT_05 => X"000000d7000000cd000000c9000000c2000000b6000000b8000000b6000000a5",
            INIT_06 => X"000000d7000000d3000000d4000000dd000000e4000000e3000000e3000000df",
            INIT_07 => X"000000ba000000ad000000aa000000c6000000bb000000c3000000cd000000df",
            INIT_08 => X"000000a4000000d3000000ec000000e3000000e2000000e3000000e5000000e6",
            INIT_09 => X"000000e0000000cf000000bf000000bc000000b8000000b7000000ad0000009f",
            INIT_0A => X"000000d3000000c8000000d0000000d6000000d6000000e0000000e5000000db",
            INIT_0B => X"000000c6000000c5000000bc000000b9000000c5000000db000000e0000000de",
            INIT_0C => X"000000af000000e3000000f1000000f2000000f1000000f4000000f4000000f5",
            INIT_0D => X"000000b6000000b8000000a0000000ae000000bb000000a1000000b0000000a8",
            INIT_0E => X"000000d4000000c4000000ba000000b9000000ca000000d0000000d5000000b9",
            INIT_0F => X"000000c8000000d4000000c5000000a9000000bb000000d5000000dc000000d7",
            INIT_10 => X"00000084000000cd000000f1000000f5000000f4000000f4000000f3000000f5",
            INIT_11 => X"0000008d0000009b0000008b0000009f000000a70000008a000000a10000008b",
            INIT_12 => X"000000e0000000c4000000a9000000a9000000a400000099000000a60000008e",
            INIT_13 => X"000000d2000000cc000000b8000000a0000000b1000000d4000000d1000000d1",
            INIT_14 => X"00000081000000d7000000ee000000f6000000f3000000f4000000f4000000f5",
            INIT_15 => X"000000a7000000b1000000aa000000aa000000aa000000a00000009c00000071",
            INIT_16 => X"000000e4000000cd000000b3000000940000008f000000980000009d0000009d",
            INIT_17 => X"000000df000000c0000000a000000093000000aa000000c1000000ce000000da",
            INIT_18 => X"000000b4000000dd000000dd000000f1000000f4000000f3000000f3000000f5",
            INIT_19 => X"000000d3000000d9000000cb000000c8000000cf000000c4000000b400000083",
            INIT_1A => X"000000e1000000cd000000a6000000a3000000bf000000c0000000c3000000cc",
            INIT_1B => X"000000da000000b20000009200000091000000a9000000b1000000d5000000e3",
            INIT_1C => X"000000c0000000d9000000ca000000e6000000f7000000f2000000f2000000f4",
            INIT_1D => X"000000d1000000ce000000d7000000ea000000e8000000e0000000c200000086",
            INIT_1E => X"000000cc0000009a000000b4000000e0000000cf000000ca000000d0000000cf",
            INIT_1F => X"000000c70000009a00000092000000ab000000bc000000c4000000c9000000dc",
            INIT_20 => X"000000ae000000df000000d1000000e3000000f5000000f3000000f3000000f5",
            INIT_21 => X"000000c9000000c1000000cc000000dd000000c1000000c1000000ba00000087",
            INIT_22 => X"000000bc000000a3000000d0000000dc000000c6000000cd000000cd000000ca",
            INIT_23 => X"000000b2000000940000008b000000a1000000cb000000df000000d1000000cb",
            INIT_24 => X"000000a4000000c2000000cd000000e5000000f2000000f3000000f1000000f2",
            INIT_25 => X"000000c4000000c0000000c4000000ca000000b8000000bd000000c10000008c",
            INIT_26 => X"000000c8000000bc000000e0000000d7000000c6000000d0000000ca000000c7",
            INIT_27 => X"000000d3000000ca000000ba000000bc000000e3000000ed000000ee000000e6",
            INIT_28 => X"0000009c000000a9000000a0000000df000000f4000000f3000000ee000000ea",
            INIT_29 => X"000000b7000000b4000000ae000000ae000000ac000000b3000000b100000086",
            INIT_2A => X"000000c4000000d0000000dc000000cd000000be000000bc000000be000000bb",
            INIT_2B => X"000000f4000000f4000000f4000000f4000000f4000000f6000000e6000000d9",
            INIT_2C => X"00000097000000be000000b6000000d8000000f2000000f2000000e6000000d3",
            INIT_2D => X"000000aa000000a60000009f0000009e000000a0000000930000006e0000006a",
            INIT_2E => X"000000af000000c6000000bd000000ad000000a60000009e000000a3000000a9",
            INIT_2F => X"000000f4000000f4000000f4000000f4000000f3000000f8000000e0000000b7",
            INIT_30 => X"0000009f000000c3000000b4000000bd000000e1000000e9000000da000000c4",
            INIT_31 => X"0000008c0000008f000000a8000000ba000000a00000008d0000005c0000005d",
            INIT_32 => X"000000960000008f0000008300000098000000a700000092000000890000008b",
            INIT_33 => X"000000f4000000f4000000f4000000f4000000f4000000f3000000e3000000bc",
            INIT_34 => X"00000089000000a200000095000000a4000000c1000000d3000000c7000000c3",
            INIT_35 => X"00000092000000a6000000cd000000bd000000a6000000b2000000aa00000096",
            INIT_36 => X"0000008a0000008000000080000000af000000d3000000c0000000ac00000099",
            INIT_37 => X"000000f3000000f3000000f5000000ef000000d3000000bf000000b1000000a0",
            INIT_38 => X"000000890000008e000000880000009c000000a2000000c8000000cf000000c2",
            INIT_39 => X"0000008b00000095000000a3000000960000009f000000b1000000b2000000a2",
            INIT_3A => X"000000850000007f0000007c000000860000009300000092000000920000008d",
            INIT_3B => X"000000f4000000f3000000f5000000cc000000a6000000ad000000a300000095",
            INIT_3C => X"000000b9000000b40000008b000000710000006e000000ad000000d0000000c3",
            INIT_3D => X"0000005f000000590000004c00000049000000570000007f0000009a00000085",
            INIT_3E => X"00000067000000630000005600000056000000580000005e000000600000005c",
            INIT_3F => X"000000f5000000f5000000e8000000af0000009b0000008f000000740000006d",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE58;


    MEM_SAMPLEIFMAP_LAYER0_INSTANCE59 : if BRAM_NAME = "sampleifmap_layer0_instance59" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a1000000b5000000880000006000000065000000a1000000aa000000b7",
            INIT_01 => X"0000006a0000007d0000007d0000008c00000087000000810000008400000080",
            INIT_02 => X"0000002800000023000000470000004d000000270000002c0000002b00000035",
            INIT_03 => X"000000f3000000f6000000db000000a700000097000000910000005000000020",
            INIT_04 => X"000000490000009900000092000000780000007c000000c2000000c1000000ca",
            INIT_05 => X"00000083000000a90000009f000000b800000094000000830000008700000069",
            INIT_06 => X"000000730000006f000000aa000000af0000007a000000840000007600000066",
            INIT_07 => X"000000f4000000f2000000c5000000bb000000b5000000b2000000910000006f",
            INIT_08 => X"00000024000000820000009d0000007300000072000000b8000000c8000000d8",
            INIT_09 => X"000000840000009d000000810000006f0000006300000081000000950000004f",
            INIT_0A => X"000000bd000000ba000000c1000000c8000000b9000000b7000000c1000000b1",
            INIT_0B => X"000000f6000000e8000000a20000009400000097000000b6000000c7000000b5",
            INIT_0C => X"0000003d000000710000008b0000006000000071000000bb000000cc000000d9",
            INIT_0D => X"0000007d0000005e00000053000000550000005d00000073000000700000004e",
            INIT_0E => X"0000008f0000008c00000095000000a00000008a0000007f0000009f000000bf",
            INIT_0F => X"000000f7000000e20000009a00000073000000630000009f000000bd0000008a",
            INIT_10 => X"00000054000000630000005c0000004900000075000000c7000000d0000000d5",
            INIT_11 => X"0000005f00000067000000570000005f0000006900000061000000410000004b",
            INIT_12 => X"0000008f0000008900000090000000960000009700000099000000a200000086",
            INIT_13 => X"000000f7000000de00000092000000730000006f0000008f0000009900000093",
            INIT_14 => X"0000005a0000005c000000510000006500000083000000cc000000ce000000cc",
            INIT_15 => X"000000570000007d0000006f0000006200000045000000390000002d00000046",
            INIT_16 => X"0000007d0000005e00000065000000620000006700000070000000660000004a",
            INIT_17 => X"000000f8000000d4000000890000009a00000095000000710000005200000073",
            INIT_18 => X"0000005e000000560000007a0000006900000075000000ce000000d0000000d1",
            INIT_19 => X"00000063000000ad00000083000000660000002f000000330000003600000056",
            INIT_1A => X"000000ab0000007c0000008a00000079000000820000009e000000640000002d",
            INIT_1B => X"000000fa000000cf0000007500000098000000ab0000005f0000004b000000bb",
            INIT_1C => X"0000008000000072000000740000003b00000068000000cc000000d6000000dd",
            INIT_1D => X"0000004b0000006c00000046000000380000003000000034000000410000007c",
            INIT_1E => X"000000af0000008f000000a7000000910000008f000000a60000005f00000030",
            INIT_1F => X"000000fb000000d6000000680000005400000062000000480000004a000000af",
            INIT_20 => X"000000b000000080000000440000002f00000063000000c9000000d4000000d7",
            INIT_21 => X"0000002f0000002b00000027000000280000002d000000380000005000000087",
            INIT_22 => X"0000008b00000090000000930000007d0000006e000000500000003c00000037",
            INIT_23 => X"000000fb000000d90000006d000000450000004300000046000000430000005c",
            INIT_24 => X"000000aa0000008500000075000000730000009d000000cb000000cf000000cf",
            INIT_25 => X"0000002d0000002900000029000000280000003000000048000000650000007e",
            INIT_26 => X"000000c9000000c7000000dc000000da000000c0000000530000002700000032",
            INIT_27 => X"000000f7000000d20000007e0000005a0000003f00000038000000340000006b",
            INIT_28 => X"000000a1000000860000009a000000bf000000d8000000ce000000c0000000bc",
            INIT_29 => X"000000290000002300000022000000210000003e000000680000007300000079",
            INIT_2A => X"000000bb000000be000000c0000000c7000000b3000000550000003100000033",
            INIT_2B => X"000000f5000000d1000000850000006f00000042000000260000002700000060",
            INIT_2C => X"000000a0000000840000009e000000b5000000c6000000cd000000c6000000bf",
            INIT_2D => X"000000310000002c0000002600000027000000460000006f0000007600000072",
            INIT_2E => X"000000a6000000ad00000096000000870000007e000000690000005d00000044",
            INIT_2F => X"000000f2000000cf0000008200000071000000470000002a0000002800000048",
            INIT_30 => X"0000008500000082000000a3000000ab000000b8000000c6000000d1000000ce",
            INIT_31 => X"00000039000000350000002f000000320000004d000000680000006f0000006b",
            INIT_32 => X"000000b0000000a800000091000000780000006800000057000000480000003f",
            INIT_33 => X"000000ee000000d40000007e0000006600000047000000300000002800000045",
            INIT_34 => X"0000006500000086000000a6000000b2000000bd000000c2000000c2000000c7",
            INIT_35 => X"0000003e0000003b000000360000003e0000004f000000600000006900000063",
            INIT_36 => X"0000008f000000810000007400000064000000570000004e0000004500000041",
            INIT_37 => X"000000e8000000df0000008500000059000000470000002c0000002700000057",
            INIT_38 => X"0000005000000090000000bc000000bd000000bc000000be000000bc000000c1",
            INIT_39 => X"0000004e0000004a00000045000000490000004600000058000000630000005a",
            INIT_3A => X"000000720000006d00000066000000610000005d000000560000004e0000004e",
            INIT_3B => X"000000e7000000e8000000ad000000640000004a00000030000000300000005e",
            INIT_3C => X"00000055000000a5000000bb000000c8000000cd000000d0000000c7000000c4",
            INIT_3D => X"00000063000000620000005900000054000000540000004e0000004c0000004c",
            INIT_3E => X"0000007f00000080000000810000007d0000007c00000072000000630000005e",
            INIT_3F => X"000000df000000e1000000cc0000009400000060000000540000005b00000070",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYER0_INSTANCE59;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE0 : if BRAM_NAME = "samplegold_layer0_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001d0000000f0000000d00000017000000140000000f0000001200000012",
            INIT_01 => X"00000016000000150000000c0000000600000001000000000000000a0000001d",
            INIT_02 => X"0000000000000003000000080000000400000013000000130000000f00000012",
            INIT_03 => X"0000000b000000000000000b0000000500000000000000000000000000000004",
            INIT_04 => X"00000000000000000000001e000000200000001b000000120000001b00000013",
            INIT_05 => X"0000000c00000000000000010000000100000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000110000000b00000019",
            INIT_07 => X"0000000300000003000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000001000000000000000000000000000000000000000000000000",
            INIT_0B => X"00000000000000000000001c0000000400000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000200000000000000000000000000000000",
            INIT_0E => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"000000000000000b000000000000000000000000000000000000000000000000",
            INIT_10 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"00000000000000000000000000000000000000000000000b0000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000020",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"000000000000000000000000000000000000000000000000000000000000000b",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"000000000000000d000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000070000000400000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000010000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000a0000003f0000000f0000001a0000000f000000000000000000000000",
            INIT_31 => X"0000002000000025000000380000003a00000032000000000000000000000000",
            INIT_32 => X"000000000000003a0000002c0000002000000027000000250000002900000022",
            INIT_33 => X"000000240000001f00000020000000200000001d0000001d0000001e00000000",
            INIT_34 => X"0000000e0000002f0000002f000000300000002100000028000000220000001e",
            INIT_35 => X"000000330000002f00000023000000220000001d00000019000000210000000f",
            INIT_36 => X"0000002a000000410000003100000033000000290000003a0000002800000034",
            INIT_37 => X"0000001a0000002d000000210000001c000000170000001f0000002a00000030",
            INIT_38 => X"000000000000000000000000000000000000000000000000000000290000001c",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"00000000000000000000000000000000000000060000000e0000001800000003",
            INIT_3E => X"000000000000000100000002000000000000000000000000000000000000000b",
            INIT_3F => X"0000001e0000000000000000000000000000000000000006000000000000001b",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE0;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE1 : if BRAM_NAME = "samplegold_layer0_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001d00000000000000030000000500000014000000110000000000000000",
            INIT_01 => X"00000000000000170000000f0000000300000000000000080000000000000010",
            INIT_02 => X"00000003000000440000000000000004000000060000000a0000001a00000000",
            INIT_03 => X"00000000000000000000000b0000001700000002000000000000000b00000000",
            INIT_04 => X"00000004000000000000003700000000000000000000000b0000001e0000000c",
            INIT_05 => X"000000060000000000000006000000140000002000000002000000110000000a",
            INIT_06 => X"000000110000000000000000000000200000000000000000000000000000002d",
            INIT_07 => X"00000000000000080000001100000004000000280000001d0000000000000008",
            INIT_08 => X"00000000000000060000000000000010000000000000000b0000000b00000000",
            INIT_09 => X"00000012000000090000000e0000002700000000000000240000001800000000",
            INIT_0A => X"00000000000000000000000c0000000000000000000000000000001500000012",
            INIT_0B => X"000000110000002d000000280000000d0000005800000000000000230000002b",
            INIT_0C => X"00000036000000000000000b0000001f000000220000001b0000000000000000",
            INIT_0D => X"0000001a000000210000001f0000000700000000000000450000001200000023",
            INIT_0E => X"000000380000002a0000002f0000002f0000002e00000028000000220000001e",
            INIT_0F => X"0000002a00000024000000240000002500000027000000000000002500000033",
            INIT_10 => X"000000520000002e0000002c0000003a0000002e0000002f000000360000002f",
            INIT_11 => X"0000002e0000002f0000002a0000002a000000260000002b0000001300000000",
            INIT_12 => X"000000190000002c000000330000002b00000028000000450000002a0000002f",
            INIT_13 => X"0000002e0000002d000000310000002e00000024000000230000002800000019",
            INIT_14 => X"00000000000000000000000000000000000000000000001f0000003a00000043",
            INIT_15 => X"00000000000000000000000a0000000200000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"00000000000000030000001c0000001f00000000000000170000000800000010",
            INIT_18 => X"0000002b00000000000000000000000000000000000000000000002a00000000",
            INIT_19 => X"00000000000000000000003f0000002d00000042000000000000000000000011",
            INIT_1A => X"0000002c00000028000000000000000e00000000000000000000000000000071",
            INIT_1B => X"0000006c000000000000002a0000003b000000260000005a0000000000000025",
            INIT_1C => X"0000003c000000480000005d0000002400000034000000000000002300000005",
            INIT_1D => X"0000003100000059000000000000003e0000001e000000520000002f00000000",
            INIT_1E => X"00000000000000600000003e000000610000002c000000000000000000000037",
            INIT_1F => X"0000001500000073000000480000002500000031000000120000005c00000073",
            INIT_20 => X"00000075000000000000006a0000004a0000005a000000000000000000000038",
            INIT_21 => X"0000003100000028000000650000004d000000370000000c0000001200000047",
            INIT_22 => X"000000500000004f0000000000000046000000380000008b0000000600000000",
            INIT_23 => X"0000002a0000000b000000840000004200000068000000130000002500000006",
            INIT_24 => X"000000040000005b0000001600000029000000000000002c0000002e00000013",
            INIT_25 => X"0000001800000064000000000000009f0000003a0000004a0000000000000000",
            INIT_26 => X"0000000000000000000000170000005a0000003b000000300000004d00000000",
            INIT_27 => X"000000200000004c0000009300000000000000940000003c0000000f0000000c",
            INIT_28 => X"0000003100000020000000230000001d0000001a000000410000008300000071",
            INIT_29 => X"0000003c0000003a00000073000000d8000000000000004e0000002b0000001d",
            INIT_2A => X"0000005f0000004f000000400000003e0000003c0000003d0000003800000047",
            INIT_2B => X"0000003e0000003f0000004900000042000000af000000820000000000000012",
            INIT_2C => X"000000450000006a0000003d0000004800000050000000400000003800000039",
            INIT_2D => X"000000410000003c000000420000004d000000390000005a000000cb00000000",
            INIT_2E => X"0000003e0000004b000000760000007b000000380000004e0000004d00000048",
            INIT_2F => X"0000005500000044000000380000004400000043000000350000004800000054",
            INIT_30 => X"00000008000000080000000000000000000000800000006f0000001a0000003a",
            INIT_31 => X"0000000000000000000000000000000400000000000000050000000300000006",
            INIT_32 => X"0000000a000000070000000c0000000a00000007000000050000000600000000",
            INIT_33 => X"0000000000000006000000240000000000000000000000000000001a00000049",
            INIT_34 => X"0000000000000007000000040000000400000000000000000000000400000000",
            INIT_35 => X"000000000000001700000007000000150000001a0000000d0000000000000000",
            INIT_36 => X"00000037000000000000000d0000000500000009000000250000002800000000",
            INIT_37 => X"000000000000000100000000000000000000000000000000000000050000001b",
            INIT_38 => X"0000000e0000000600000056000000800000000b000000130000005a00000026",
            INIT_39 => X"0000000000000000000000180000000f00000025000000250000000000000000",
            INIT_3A => X"0000001f0000001a0000002a0000000000000000000000000000000800000000",
            INIT_3B => X"000000070000000600000027000000090000000000000000000000000000003a",
            INIT_3C => X"00000011000000090000000a0000000000000021000000000000000400000000",
            INIT_3D => X"0000001c00000007000000150000001d00000017000000000000000b00000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000160000001900000010",
            INIT_3F => X"000000040000000b000000040000001000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE1;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE2 : if BRAM_NAME = "samplegold_layer0_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000000000000040000001a00000000000000000000001c",
            INIT_01 => X"00000011000000040000000900000000000000000000002f0000000300000000",
            INIT_02 => X"0000001b0000000000000000000000000000000c0000004a0000000000000000",
            INIT_03 => X"000000850000009c00000046000000000000000000000000000000000000001f",
            INIT_04 => X"000000000000001b000000410000002000000000000000000000000000000028",
            INIT_05 => X"000000000000000000000000000000460000000f000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000002",
            INIT_08 => X"0000000000000011000000000000000000000012000000070000000400000000",
            INIT_09 => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000001300000000000000000000000000000000",
            INIT_0B => X"0000001300000014000000000000000000000000000000000000000000000000",
            INIT_0C => X"000000a2000000a30000009d0000000000000022000000280000000000000004",
            INIT_0D => X"0000007c00000094000000ad000000b7000000ac0000009d000000a4000000a5",
            INIT_0E => X"000000ac000000a8000000ad000000a20000009200000092000000840000007c",
            INIT_0F => X"0000003e0000002e0000003a0000007a000000a0000000a90000008c000000a0",
            INIT_10 => X"000000af000000b0000000ac0000006a000000890000008b0000006e0000004e",
            INIT_11 => X"000000270000000a0000001e000000070000002d00000048000000730000008e",
            INIT_12 => X"00000059000000a2000000aa000000a40000002b0000004d000000670000003a",
            INIT_13 => X"000000250000001b0000002d000000330000000c00000015000000270000004d",
            INIT_14 => X"00000043000000470000004e00000060000000940000001f000000170000003a",
            INIT_15 => X"0000002f0000001c000000170000003900000031000000000000001f0000002f",
            INIT_16 => X"00000031000000450000003b00000025000000990000008e0000001200000016",
            INIT_17 => X"0000000e0000001700000012000000100000002a0000003e000000000000002d",
            INIT_18 => X"0000002f0000002d0000003e000000320000002f0000009f000000620000002a",
            INIT_19 => X"0000000a0000001c000000260000000e00000010000000280000003200000000",
            INIT_1A => X"0000001e00000029000000270000002e0000002600000037000000620000002c",
            INIT_1B => X"0000002b00000000000000140000004100000022000000090000002d0000002f",
            INIT_1C => X"00000042000000540000000d000000300000003600000022000000550000000e",
            INIT_1D => X"00000000000000240000000500000010000000790000002d0000000f00000026",
            INIT_1E => X"000000060000001d000000340000002d00000028000000080000002000000035",
            INIT_1F => X"00000017000000000000002300000015000000000000008a0000006200000009",
            INIT_20 => X"000000000000000000000000000000000000000600000000000000000000001a",
            INIT_21 => X"000000000000003a000000060000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000003400000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000002300000022000000000000000000000000000000000000000000000000",
            INIT_29 => X"000000170000001d0000002400000026000000270000001e0000002000000025",
            INIT_2A => X"0000002a0000002c00000023000000180000001e00000024000000260000001a",
            INIT_2B => X"000000000000001d0000000e0000001d0000000f00000020000000280000001f",
            INIT_2C => X"000000210000002800000039000000060000001c0000002b0000002000000009",
            INIT_2D => X"00000000000000000000002e0000002100000006000000000000001a00000027",
            INIT_2E => X"0000000f00000029000000210000004c000000000000002c0000002500000000",
            INIT_2F => X"0000000000000009000000000000004800000000000000000000000400000024",
            INIT_30 => X"0000000b00000009000000560000000200000026000000000000004a00000000",
            INIT_31 => X"0000000000000006000000000000000000000059000000000000000000000000",
            INIT_32 => X"00000000000000130000003e0000001a000000000000000a000000000000002b",
            INIT_33 => X"00000000000000000000001400000000000000000000008e0000000000000000",
            INIT_34 => X"0000000000000000000000360000003f00000000000000200000000000000000",
            INIT_35 => X"0000000000000000000000150000000a00000000000000000000006600000000",
            INIT_36 => X"0000000000000000000000000000004200000038000000000000000000000000",
            INIT_37 => X"0000000200000000000000080000000f0000001d000000000000000000000042",
            INIT_38 => X"0000000000000024000000000000000000000011000000040000002100000000",
            INIT_39 => X"00000000000000000000000000000023000000210000001e0000000000000025",
            INIT_3A => X"00000000000000050000000200000000000000270000000f000000000000002c",
            INIT_3B => X"0000007800000000000000040000002a0000001400000034000000300000000c",
            INIT_3C => X"0000000900000008000000000000000000000000000000220000000000000000",
            INIT_3D => X"0000000000000040000000000000001400000020000000000000000000000001",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000004300000021000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE2;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE3 : if BRAM_NAME = "samplegold_layer0_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"000000000000000000000000000000000000005d000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000002b00000000000000000000000400000000000000000000000000000000",
            INIT_05 => X"000000370000003a00000030000000290000002f0000002c0000002d00000030",
            INIT_06 => X"000000350000002c000000310000002a0000002700000026000000250000002a",
            INIT_07 => X"0000000c0000003b000000290000001f000000000000002d0000002e00000030",
            INIT_08 => X"0000002e000000290000001c000000250000001f0000000e0000000000000000",
            INIT_09 => X"000000000000000000000000000000230000002d0000003b0000003200000035",
            INIT_0A => X"000000320000002300000000000000000000001a000000040000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000001900000025",
            INIT_0C => X"0000000000000018000000120000000000000000000000110000000000000006",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000300000003000000380000000b00000000000000000000000500000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000070000003a00000007000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000200000000000000000000000000000000",
            INIT_13 => X"000000000000000d000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000050000001a00000000000000000000000000000000",
            INIT_15 => X"000000000000000000000008000000000000000400000018000000030000000f",
            INIT_16 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000001f00000000000000000000000a00000011",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000b0000000c0000000c000000040000000800000008000000110000000a",
            INIT_22 => X"00000000000000060000000800000011000000230000002d000000210000000b",
            INIT_23 => X"00000042000000230000000500000000000000080000000c0000000a0000000a",
            INIT_24 => X"00000033000000350000000a000000170000000a000000000000000000000000",
            INIT_25 => X"0000000000000000000000090000001600000037000000050000000800000005",
            INIT_26 => X"0000000500000000000000000000000c0000000e000000000000000000000000",
            INIT_27 => X"000000040000001a000000000000000200000000000000000000000800000008",
            INIT_28 => X"0000000e0000000200000000000000010000000e000000000000000600000010",
            INIT_29 => X"0000000000000000000000000000000700000000000000090000000000000000",
            INIT_2A => X"0000003e0000000300000006000000000000000f000000000000000000000000",
            INIT_2B => X"0000000700000015000000140000000000000000000000000000000000000028",
            INIT_2C => X"0000000000000012000000180000001c00000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000001100000000000000110000000000000031",
            INIT_2E => X"0000003500000035000000020000000000000000000000000000000000000000",
            INIT_2F => X"000000000000000e000000050000000000000009000000000000000e00000021",
            INIT_30 => X"0000000000000000000000260000000000000000000000000000000100000000",
            INIT_31 => X"0000000c00000000000000000000000000000030000000260000000000000000",
            INIT_32 => X"0000000000000000000000000000000900000023000000000000000400000000",
            INIT_33 => X"000000000000000300000018000000000000000000000011000000360000004e",
            INIT_34 => X"0000000000000037000000510000001e00000000000000000000000000000007",
            INIT_35 => X"0000000c00000021000000350000000a00000005000000000000000000000000",
            INIT_36 => X"0000000000000000000000030000000500000004000000280000005600000000",
            INIT_37 => X"0000001800000000000000160000000000000000000000000000000000000000",
            INIT_38 => X"000000000000000000000000000000000000000000000000000000000000003f",
            INIT_39 => X"0000000b0000004f000000180000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000300000000000000220000000000000000000000000000001400000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000012",
            INIT_3D => X"0000000800000015000000090000000e0000000a000000130000000d00000000",
            INIT_3E => X"0000000200000006000000130000001b000000220000001c0000000c00000006",
            INIT_3F => X"0000001a0000000f000000360000000f0000000d000000090000000b00000008",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE3;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE4 : if BRAM_NAME = "samplegold_layer0_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000260000000a0000001a000000210000002400000035000000340000001f",
            INIT_01 => X"00000020000000280000003300000051000000080000000a0000000b00000024",
            INIT_02 => X"00000014000000330000001a000000190000002b0000004b0000005e00000053",
            INIT_03 => X"0000005b000000360000002f000000450000002e00000019000000120000000e",
            INIT_04 => X"000000150000005e000000710000001b000000150000003b000000420000005d",
            INIT_05 => X"000000670000003b000000330000003b00000064000000440000007e00000035",
            INIT_06 => X"00000013000000280000009e0000007f00000001000000250000003900000038",
            INIT_07 => X"000000500000007f0000005b0000002e0000004b0000007d0000007e000000bd",
            INIT_08 => X"0000005a0000001700000043000000940000007a000000150000003c00000047",
            INIT_09 => X"0000003b0000004600000081000000780000004e00000065000000a800000075",
            INIT_0A => X"000000a5000000390000003900000040000000a50000008e000000330000004c",
            INIT_0B => X"0000004b000000480000004c000000780000005f000000500000006a00000085",
            INIT_0C => X"0000005900000066000000380000007300000066000000b8000000b000000026",
            INIT_0D => X"0000000e0000002b0000002c000000410000006500000033000000510000004e",
            INIT_0E => X"000000790000005f000000330000006f0000007500000086000000b3000000c0",
            INIT_0F => X"000000c700000027000000270000002f00000025000000400000005a00000042",
            INIT_10 => X"00000079000000b900000091000000650000009e000000a20000008b000000ab",
            INIT_11 => X"000000cb000000c100000068000000710000005a00000047000000400000003c",
            INIT_12 => X"0000006f0000007c000000850000008a000000a5000000e7000000c90000009d",
            INIT_13 => X"000000b1000000a10000008c0000008e0000008a000000880000008000000078",
            INIT_14 => X"00000084000000760000007100000070000000750000007a000000af000000e5",
            INIT_15 => X"000000ef000000a6000000850000009d000000a30000009a000000950000008c",
            INIT_16 => X"0000009b0000008c000000820000007700000073000000790000008000000088",
            INIT_17 => X"00000074000000a70000007f0000008f00000097000000ab000000a300000093",
            INIT_18 => X"0000009a0000008500000086000000880000007c0000007e000000890000007f",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000008d000000af",
            INIT_1A => X"00000000000000000000000b0000001c00000013000000000000000000000000",
            INIT_1B => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"00000000000000000000001e0000001400000000000000000000003300000014",
            INIT_1D => X"000000280000001c0000003e000000000000000000000000000000000000003f",
            INIT_1E => X"00000019000000000000001e0000000700000000000000000000000000000000",
            INIT_1F => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000e000000060000001a0000000000000000",
            INIT_21 => X"000000000000001d000000040000000f00000000000000000000000000000009",
            INIT_22 => X"00000002000000000000002f0000002500000000000000000000000800000000",
            INIT_23 => X"000000260000000000000006000000000000000000000000000000030000004f",
            INIT_24 => X"0000000d0000000d00000018000000000000000000000000000000000000001c",
            INIT_25 => X"0000000800000018000000000000000900000000000000050000000000000000",
            INIT_26 => X"0000000000000000000000070000000000000002000000000000000000000000",
            INIT_27 => X"000000000000001c0000000000000000000000000000001e0000003d00000000",
            INIT_28 => X"0000003200000022000000000000002e00000000000000000000000000000010",
            INIT_29 => X"000000000000000d0000003a0000002600000036000000000000000000000003",
            INIT_2A => X"000000000000001500000012000000000000000a000000000000000000000000",
            INIT_2B => X"00000008000000000000000000000001000000310000001f0000002e00000000",
            INIT_2C => X"0000001900000000000000000000000000000000000000220000000000000000",
            INIT_2D => X"0000004100000021000000160000000000000000000000000000000d0000000f",
            INIT_2E => X"0000000c000000370000003f00000052000000a2000000000000000000000000",
            INIT_2F => X"000000360000000d000000000000000000000000000000020000000000000006",
            INIT_30 => X"0000000000000000000000000000000200000000000000560000004100000000",
            INIT_31 => X"0000002500000000000000020000000000000000000000030000000000000000",
            INIT_32 => X"000000070000000000000000000000010000000000000000000000060000003e",
            INIT_33 => X"0000003600000018000000000000000c0000004200000000000000000000000a",
            INIT_34 => X"0000000000000005000000000000000000000000000000090000001300000024",
            INIT_35 => X"0000000000000000000000000000000000000000000000040000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"00000000000000000000000000000000000000000000001f0000000400000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_3C => X"0000000000000001000000020000000000000007000000000000002d00000005",
            INIT_3D => X"0000000200000000000000000000000000000000000000000000000000000002",
            INIT_3E => X"000000060000000100000010000000000000000300000000000000000000003b",
            INIT_3F => X"0000005d000000000000000000000000000000000000002c0000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE4;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE5 : if BRAM_NAME = "samplegold_layer0_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000000000000000000000000000000e0000000000000000",
            INIT_01 => X"00000000000000520000000000000000000000000000000f0000001c00000000",
            INIT_02 => X"0000000000000000000000000000000400000000000000130000001200000000",
            INIT_03 => X"00000000000000000000002d000000000000000500000000000000170000000c",
            INIT_04 => X"000000000000001100000000000000160000000000000000000000030000001d",
            INIT_05 => X"0000001b00000000000000110000000000000008000000000000000000000012",
            INIT_06 => X"00000003000000000000003b0000000000000019000000090000000000000000",
            INIT_07 => X"0000000000000012000000120000000000000000000000050000000000000010",
            INIT_08 => X"0000002d000000000000000000000058000000000000000d0000003300000000",
            INIT_09 => X"0000001d0000002c0000003e0000003300000028000000020000000000000004",
            INIT_0A => X"0000004e0000004e0000002e000000000000003b000000000000003600000070",
            INIT_0B => X"0000005a000000530000005a00000058000000560000004f0000004900000044",
            INIT_0C => X"0000004c0000004a00000048000000490000000000000008000000480000006f",
            INIT_0D => X"000000600000005a0000005e0000005d000000570000005b0000005b00000054",
            INIT_0E => X"00000057000000530000004d000000450000005000000031000000000000008a",
            INIT_0F => X"0000006700000067000000500000005e00000074000000610000006400000061",
            INIT_10 => X"00000052000000520000005200000049000000550000005f0000004900000041",
            INIT_11 => X"0000002e000000330000002e0000002f00000045000000530000006b0000005e",
            INIT_12 => X"000000270000001c000000230000002b0000002f000000310000002f0000002f",
            INIT_13 => X"000000340000002d000000350000003200000032000000240000002700000026",
            INIT_14 => X"0000002400000015000000130000002100000004000000250000001300000055",
            INIT_15 => X"0000002c000000380000002e000000340000003b0000001a000000280000002d",
            INIT_16 => X"00000027000000040000000b0000000a0000004f0000001a0000000000000000",
            INIT_17 => X"0000001a0000002300000025000000360000002c000000790000000000000039",
            INIT_18 => X"000000530000000e000000000000001200000000000000530000001800000008",
            INIT_19 => X"00000000000000000000001a0000002c000000490000000a0000006300000000",
            INIT_1A => X"0000000000000039000000000000001e000000000000000b0000005f00000008",
            INIT_1B => X"00000000000000000000000000000000000000490000002e0000000000000038",
            INIT_1C => X"00000015000000000000000d00000004000000230000000000000000000000bf",
            INIT_1D => X"000000a400000000000000000000000a0000005000000061000000000000000c",
            INIT_1E => X"0000000100000000000000000000000d000000270000001e0000000000000000",
            INIT_1F => X"000000000000007c000000000000000800000000000000680000004500000000",
            INIT_20 => X"0000003c00000000000000170000000000000012000000220000002a00000000",
            INIT_21 => X"000000000000002200000006000000310000001c000000000000000300000011",
            INIT_22 => X"000000000000004a00000000000000180000000a000000440000003a00000026",
            INIT_23 => X"0000004800000005000000000000000a000000170000000e0000002a00000019",
            INIT_24 => X"0000000b00000000000000a30000000000000011000000510000001c00000056",
            INIT_25 => X"0000001e0000002d000000280000001400000000000000000000000000000056",
            INIT_26 => X"0000000000000000000000000000009800000000000000280000004000000000",
            INIT_27 => X"00000000000000110000000e0000001000000010000000090000000000000000",
            INIT_28 => X"0000000a0000000500000009000000000000001f000000480000004100000003",
            INIT_29 => X"0000000000000017000000080000001000000017000000140000001000000008",
            INIT_2A => X"0000000d00000009000000000000001100000000000000000000007400000010",
            INIT_2B => X"0000000d00000000000000000000002600000000000000090000000d00000010",
            INIT_2C => X"0000001000000018000000090000000c00000016000000000000000000000019",
            INIT_2D => X"0000000000000000000000000000000000000003000000310000000b00000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000001000000000000000000000000000000000000000400000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000012000000040000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000005",
            INIT_35 => X"0000000000000008000000380000000000000000000000270000000100000000",
            INIT_36 => X"0000000000000004000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"000000000000000f000000000000000000000000000000000000001400000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000012000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE5;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE6 : if BRAM_NAME = "samplegold_layer0_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000300000001e000000000000000000000000000000000000000000000011",
            INIT_01 => X"00000001000000240000001c000000000000000000000000000000000000003e",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"000000360000002f000000000000000000000013000000000000000000000000",
            INIT_0A => X"0000002b000000360000003b0000003900000030000000350000003500000033",
            INIT_0B => X"0000003600000038000000300000002700000028000000250000002000000020",
            INIT_0C => X"000000020000000200000023000000390000003b000000420000003300000039",
            INIT_0D => X"0000003900000036000000130000003000000027000000110000000600000006",
            INIT_0E => X"00000000000000040000000000000000000000000000001e0000003d00000037",
            INIT_0F => X"0000004000000037000000320000000000000015000000170000000000000001",
            INIT_10 => X"0000000000000000000000170000000000000000000000000000001e00000012",
            INIT_11 => X"0000003300000044000000100000003400000012000000000000000000000000",
            INIT_12 => X"0000000000000000000000090000001000000000000000000000000600000025",
            INIT_13 => X"0000002b0000000d0000000b00000038000000310000000f0000000000000000",
            INIT_14 => X"000000000000000000000000000000000000002a000000000000000b00000008",
            INIT_15 => X"000000170000002e000000110000000e0000003d000000070000002c00000000",
            INIT_16 => X"0000000400000000000000000000000000000000000000130000000300000008",
            INIT_17 => X"000000000000000a0000002e0000002200000000000000250000000000000019",
            INIT_18 => X"0000001100000015000000000000000200000000000000000000000f00000013",
            INIT_19 => X"0000002c000000000000000c00000000000000000000001c0000000000000009",
            INIT_1A => X"000000140000000e000000160000002100000000000000000000000000000000",
            INIT_1B => X"0000000000000005000000060000001f00000000000000000000000300000000",
            INIT_1C => X"00000000000000150000001400000005000000280000001e0000000000000000",
            INIT_1D => X"000000000000000000000000000000000000001700000011000000060000002c",
            INIT_1E => X"0000003c00000032000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"00000000000000000000004f0000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000002800000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000002f0000002b00000028000000200000002c000000290000002300000022",
            INIT_27 => X"00000024000000280000002e000000290000001e0000001d0000002900000032",
            INIT_28 => X"000000050000002e00000030000000430000000e000000210000002c00000024",
            INIT_29 => X"00000028000000020000003f0000002c00000015000000190000002900000021",
            INIT_2A => X"0000001c00000000000000100000002400000028000000200000002a00000029",
            INIT_2B => X"000000240000002e000000000000005c0000000b0000001a000000320000000c",
            INIT_2C => X"0000001800000023000000000000001900000025000000270000000c00000038",
            INIT_2D => X"000000130000000000000041000000050000002c00000000000000260000001a",
            INIT_2E => X"0000001200000038000000140000000000000025000000240000002a00000027",
            INIT_2F => X"00000000000000000000002f0000003700000000000000240000001a0000002b",
            INIT_30 => X"0000001d000000070000002a0000003400000000000000430000002500000016",
            INIT_31 => X"000000150000000000000000000000460000000e000000240000001100000020",
            INIT_32 => X"00000025000000000000000d000000280000002b00000000000000390000001c",
            INIT_33 => X"0000000b0000003500000000000000020000003400000029000000060000000b",
            INIT_34 => X"0000000d0000000d00000011000000000000002c000000110000000000000018",
            INIT_35 => X"000000000000001b0000000e0000000000000034000000000000003f00000000",
            INIT_36 => X"00000000000000000000001a00000000000000000000002b000000050000003f",
            INIT_37 => X"0000000f0000002c0000001d00000000000000140000002a0000000000000039",
            INIT_38 => X"0000003800000000000000000000002f00000010000000000000000f0000002f",
            INIT_39 => X"0000000f0000002b000000270000000500000000000000320000002900000000",
            INIT_3A => X"0000000000000000000000000000000000000021000000110000000800000008",
            INIT_3B => X"0000000000000003000000070000000000000000000000000000000500000052",
            INIT_3C => X"0000002e00000022000000000000000000000014000000030000000000000000",
            INIT_3D => X"0000000200000000000000000000000100000005000000020000000600000000",
            INIT_3E => X"000000000000000d000000220000000000000000000000090000000000000000",
            INIT_3F => X"0000000000000000000000000000000100000000000000000000000600000009",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE6;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE7 : if BRAM_NAME = "samplegold_layer0_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000140000000400000000000000000000001300000015",
            INIT_01 => X"0000001a0000001200000000000000000000000c000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000020000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000e00000000000000000000000000000000",
            INIT_1C => X"00000000000000000000000000000000000000000000001a0000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"000000000000002f0000003d0000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000120000001f00000013",
            INIT_28 => X"0000000000000000000000000000000000000009000000130000000000000000",
            INIT_29 => X"00000000000000000000000d0000004500000042000000000000000000000000",
            INIT_2A => X"00000000000000030000000000000000000000000000000a0000001f00000004",
            INIT_2B => X"000000000000000000000009000000090000000000000025000000100000000e",
            INIT_2C => X"0000000000000000000000000000000800000017000000190000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"00000020000000270000000e0000000000000000000000000000000000000000",
            INIT_2F => X"000000210000002a000000310000003a0000003e00000040000000370000001b",
            INIT_30 => X"000000370000000b0000000a000000120000002100000026000000140000001c",
            INIT_31 => X"000000420000004c0000005600000055000000500000004b0000003f00000041",
            INIT_32 => X"0000000a0000000200000000000000000000001e00000029000000320000003e",
            INIT_33 => X"000000020000000800000000000000010000000b000000030000000000000000",
            INIT_34 => X"0000001800000010000000000000000000000000000000000000000000000000",
            INIT_35 => X"000000000000000000000000000000000000002200000006000000060000000a",
            INIT_36 => X"000000040000000600000003000000000000000000000000000000000000000b",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000400000004",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_3A => X"0000002b0000002c0000002b0000002b0000002b0000002b0000000000000000",
            INIT_3B => X"0000002b0000002b0000002a0000002d0000002c0000002b0000002b0000002b",
            INIT_3C => X"0000002c0000002b0000002b0000002b0000002b0000002b0000002b0000002c",
            INIT_3D => X"0000002c0000002b0000002c00000031000000280000001c0000002b00000029",
            INIT_3E => X"000000230000002b0000002c0000002d0000002b0000002b0000002b00000029",
            INIT_3F => X"000000320000002c0000002b0000002b0000002b0000002c0000001a0000001c",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE7;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE8 : if BRAM_NAME = "samplegold_layer0_instance8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002c000000200000002f0000001f0000002c0000002b0000002c0000002d",
            INIT_01 => X"00000022000000190000002b0000002b0000002b00000046000000330000002d",
            INIT_02 => X"00000031000000330000002900000032000000200000002c000000290000002e",
            INIT_03 => X"0000002f00000038000000320000002b00000029000000170000001400000020",
            INIT_04 => X"0000002b0000001e0000001d0000001700000013000000120000002500000021",
            INIT_05 => X"00000027000000290000001f000000160000002e0000004b0000002600000032",
            INIT_06 => X"00000015000000200000002d000000550000003b00000021000000050000001b",
            INIT_07 => X"0000002700000034000000150000003b0000001e000000260000001400000019",
            INIT_08 => X"0000002f0000002a000000200000001c0000001900000021000000430000002e",
            INIT_09 => X"000000230000003200000037000000300000002a0000006b0000003b00000035",
            INIT_0A => X"00000014000000180000001e0000002500000023000000270000001700000028",
            INIT_0B => X"000000270000002b0000002900000027000000250000001d0000002e00000019",
            INIT_0C => X"0000002400000024000000290000001f0000002800000028000000300000002c",
            INIT_0D => X"00000022000000210000001900000014000000170000001a000000170000000c",
            INIT_0E => X"00000000000000250000002c00000029000000230000001f0000001c0000001d",
            INIT_0F => X"0000002d0000002f0000002b0000000d00000000000000000000000100000012",
            INIT_10 => X"00000000000000000000002400000018000000210000003c0000003600000031",
            INIT_11 => X"0000002000000026000000210000003f00000000000000000000000000000002",
            INIT_12 => X"00000000000000000000000000000026000000190000001f0000000e0000000e",
            INIT_13 => X"000000150000000700000012000000270000001b000000000000000000000000",
            INIT_14 => X"00000000000000000000000000000000000000230000001a0000000d00000017",
            INIT_15 => X"000000080000000d000000150000000a00000006000000030000000000000000",
            INIT_16 => X"0000004e0000004f0000004f0000004f00000052000000240000001a00000011",
            INIT_17 => X"0000004f0000004f00000051000000520000004d000000510000004f0000004f",
            INIT_18 => X"0000004f0000004e000000500000004f0000004f000000520000004e0000004f",
            INIT_19 => X"0000004e000000500000003a0000003100000080000000540000004f0000004d",
            INIT_1A => X"0000004a000000560000004c0000004f0000004e0000004e000000510000004e",
            INIT_1B => X"0000004f0000004e00000051000000270000003100000071000000640000006f",
            INIT_1C => X"0000006f0000002a00000079000000500000004e0000004c0000005100000045",
            INIT_1D => X"0000003f0000004e0000004f0000005200000011000000370000005000000043",
            INIT_1E => X"000000480000005700000035000000640000004f0000004b0000002100000022",
            INIT_1F => X"000000340000004900000048000000090000005b000000680000007a0000006a",
            INIT_20 => X"000000640000003e000000580000005e0000007f00000054000000540000004b",
            INIT_21 => X"0000003a0000001c00000051000000440000000000000060000000430000004b",
            INIT_22 => X"0000007400000062000000000000000000000003000000800000007c00000029",
            INIT_23 => X"0000000000000037000000140000000000000025000000660000005f00000074",
            INIT_24 => X"0000002700000040000000480000005000000076000000280000004c00000039",
            INIT_25 => X"0000004d00000040000000450000005d000000000000002a0000002300000016",
            INIT_26 => X"000000620000007c00000064000000690000005900000085000000610000006d",
            INIT_27 => X"00000054000000550000005a000000550000005e000000200000004900000055",
            INIT_28 => X"000000370000003c000000530000004d0000005b0000004c0000004d00000061",
            INIT_29 => X"0000004a0000002e0000003000000034000000380000000f0000002b00000028",
            INIT_2A => X"0000001c0000002b00000018000000330000004500000054000000540000004e",
            INIT_2B => X"0000002c00000000000000020000001d000000370000003a000000000000002e",
            INIT_2C => X"00000037000000060000002c0000003a0000001d000000000000000f00000017",
            INIT_2D => X"0000004400000046000000000000000800000012000000230000000a00000000",
            INIT_2E => X"0000000900000075000000060000000c0000000d0000001b0000004900000052",
            INIT_2F => X"000000060000003d000000220000000000000007000000090000000f00000006",
            INIT_30 => X"000000040000000a00000062000000100000000b0000001c0000000100000000",
            INIT_31 => X"0000001800000000000000000000000000000000000000000000000200000005",
            INIT_32 => X"000000000000000000000000000000000000001500000013000000130000001d",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000010000000000000000",
            INIT_39 => X"0000000000000000000000000000002d0000004a0000003a0000002800000000",
            INIT_3A => X"0000000500000019000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000007600000000000000000000000000000000000000000000000800000017",
            INIT_3C => X"000000000000000000000000000000000000000000000000000000170000007c",
            INIT_3D => X"00000000000000000000000000000056000000620000005f0000003200000000",
            INIT_3E => X"000000000000004e000000230000000000000000000000160000000000000000",
            INIT_3F => X"0000000000000072000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE8;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE9 : if BRAM_NAME = "samplegold_layer0_instance9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000000000000017000000a3000000790000000000000000",
            INIT_01 => X"0000004e00000066000000240000006f0000003d000000440000002800000013",
            INIT_02 => X"000000000000000000000000000000130000000000000000000000000000000b",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000004d00000000000000040000002000000019000000000000000000000009",
            INIT_08 => X"0000001c000000000000001d000000700000006300000055000000530000008e",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000020",
            INIT_0A => X"000000190000001e0000001c0000001900000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000003",
            INIT_0C => X"0000002200000000000000030000000a00000005000000440000004200000000",
            INIT_0D => X"0000005000000049000000000000000c0000001900000016000000140000001d",
            INIT_0E => X"0000001500000015000000170000000e000000100000000b000000000000001d",
            INIT_0F => X"0000001000000016000000170000001800000015000000150000001500000015",
            INIT_10 => X"0000001600000016000000160000001700000015000000150000001600000015",
            INIT_11 => X"0000000e00000000000000210000001a00000017000000150000001600000015",
            INIT_12 => X"0000001600000017000000150000001600000015000000160000001600000016",
            INIT_13 => X"00000016000000000000000000000000000000070000001f0000000f00000019",
            INIT_14 => X"000000270000001800000018000000120000000c000000070000001500000016",
            INIT_15 => X"0000000f0000000c000000000000000000000000000000000000001300000007",
            INIT_16 => X"0000001100000012000000160000001700000000000000000000000000000011",
            INIT_17 => X"00000009000000000000000200000000000000010000000a0000000800000011",
            INIT_18 => X"000000000000000000000019000000110000001f0000000b0000000000000000",
            INIT_19 => X"0000000000000004000000000000000000000000000000000000000000000000",
            INIT_1A => X"000000000000000000000000000000010000000d000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000080000000c00000010",
            INIT_1C => X"0000000000000002000000140000000000000000000000000000000200000001",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000001000000050000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000004000000070000000000000000000000060000000000000000",
            INIT_24 => X"0000000000000004000000000000000000000000000000000000000000000000",
            INIT_25 => X"00000000000000090000000a00000016000000150000000a0000002200000000",
            INIT_26 => X"00000000000000080000001d0000002000000044000000570000005900000052",
            INIT_27 => X"000000bc00000032000000090000000a0000000c0000000d0000000b00000030",
            INIT_28 => X"00000021000000000000000700000013000000220000002d0000004c000000a7",
            INIT_29 => X"00000032000000410000001b000000070000000b0000000a0000000d00000014",
            INIT_2A => X"000000000000000000000000000000030000000c000000140000002700000028",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000009",
            INIT_2F => X"0000001400000011000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"000000000000001d000000000000000000000000000000000000001000000000",
            INIT_32 => X"0000000000000000000000000000001900000014000000000000000000000000",
            INIT_33 => X"0000002500000000000000000000000000000000000000000000000000000006",
            INIT_34 => X"0000000000000000000000000000000000000000000000030000000000000000",
            INIT_35 => X"0000000000000031000000000000000000000000000000000000000400000000",
            INIT_36 => X"0000002000000008000000000000000000000009000000120000001b00000000",
            INIT_37 => X"000000360000001600000000000000000000000000000000000000000000003e",
            INIT_38 => X"00000000000000000000000b0000000000000000000000340000000000000015",
            INIT_39 => X"00000000000000a20000000d0000000600000008000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000010000000c00000000",
            INIT_3B => X"0000000000000000000000210000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000b0000000500000013000000000000000a000000030000000000000000",
            INIT_3E => X"0000000800000000000000000000000000000007000000060000001200000010",
            INIT_3F => X"0000000600000000000000000000003500000000000000120000000a00000013",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE9;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE10 : if BRAM_NAME = "samplegold_layer0_instance10" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000d0000001c0000001d0000000d0000000000000000000000380000001f",
            INIT_01 => X"000000130000000c00000009000000200000001b000000000000001e00000005",
            INIT_02 => X"00000016000000230000001b000000130000002100000032000000390000009d",
            INIT_03 => X"0000006c0000001200000012000000110000001600000010000000000000001a",
            INIT_04 => X"0000001100000014000000050000002600000037000000430000005700000081",
            INIT_05 => X"0000003f000000280000000f0000000f00000009000000090000000300000000",
            INIT_06 => X"000000000000000c0000000b0000000c000000000000000c000000350000003b",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000001b0000001a0000001e0000000000000000000000000000000000000000",
            INIT_1A => X"000000000000000000000000000000040000000f000000250000002600000023",
            INIT_1B => X"0000000100000000000000000000001300000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000001400000012",
            INIT_1D => X"0000001d0000002e000000300000001700000008000000000000000000000000",
            INIT_1E => X"0000000000000032000000400000003800000039000000430000000e0000001a",
            INIT_1F => X"000000190000001a0000001e0000001c00000017000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000059000000a5000000990000001f",
            INIT_21 => X"0000000b0000000c0000000e0000000a00000009000000070000000100000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000a00000045",
            INIT_23 => X"0000000200000002000000030000000200000001000000010000000100000002",
            INIT_24 => X"0000000200000001000000010000000200000002000000040000000300000001",
            INIT_25 => X"0000000200000000000000010000000000000001000000010000000100000001",
            INIT_26 => X"000000070000000a000000000000000000000000000000000000000e0000001c",
            INIT_27 => X"000000240000002a000000110000000600000004000000000000000000000001",
            INIT_28 => X"0000000000000000000000000000000100000001000000010000001600000025",
            INIT_29 => X"0000000000000000000000000000000000000002000000080000000200000002",
            INIT_2A => X"000000090000000c000000310000002a00000000000000000000000000000000",
            INIT_2B => X"00000040000000390000000c0000000000000002000000000000000100000004",
            INIT_2C => X"000000280000002d000000000000000000000000000000000000002a00000043",
            INIT_2D => X"0000000000000000000000000000000000000047000000780000008900000082",
            INIT_2E => X"00000000000000000000000200000034000000440000004d0000000100000000",
            INIT_2F => X"0000005200000069000000660000005500000025000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000800000039",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000001c00000004",
            INIT_32 => X"0000004b00000038000000240000001a00000000000000000000000e00000000",
            INIT_33 => X"0000003c0000001c0000003f000000560000004f000000410000004700000020",
            INIT_34 => X"0000000800000000000000120000002700000035000000480000004a0000005b",
            INIT_35 => X"000000000000000a000000000000000d00000005000000120000001100000005",
            INIT_36 => X"000000400000004c0000005e0000005f00000056000000470000003200000018",
            INIT_37 => X"000000080000001300000012000000000000000000000000000000110000002b",
            INIT_38 => X"0000000000000000000000000000000000000000000000010000000000000000",
            INIT_39 => X"000000170000001c000000000000000000000000000000010000001700000000",
            INIT_3A => X"0000001a00000057000000590000004d0000005d000000240000000000000003",
            INIT_3B => X"0000000000000001000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000001a00000078000000600000000500000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000030000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"000000f0000000f0000000ef000000ef000000ef000000ef000000ef00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE10;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE11 : if BRAM_NAME = "samplegold_layer0_instance11" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000f0000000ef000000f0000000ef000000f3000000f1000000ed000000ef",
            INIT_01 => X"000000ef000000f0000000f0000000f0000000f0000000f0000000f0000000f1",
            INIT_02 => X"000000f1000000f1000000f0000000ef000000f1000000ee000000e9000000ef",
            INIT_03 => X"000000ec000000ed000000f2000000f0000000f0000000f1000000f0000000f0",
            INIT_04 => X"000000f5000000f7000000f3000000f2000000f2000000f3000000cf000000de",
            INIT_05 => X"000000c4000000cd000000e5000000eb000000eb000000f2000000f2000000f6",
            INIT_06 => X"000000fd000000de000000d2000000f8000000f8000000fa000000d7000000b5",
            INIT_07 => X"000000f0000000f3000000ea000000f1000000e0000000f2000000f1000000f0",
            INIT_08 => X"000000dc000000d3000000ac000000aa000000fc000000f3000000e0000000e9",
            INIT_09 => X"000000b9000000d2000000f5000000fc000000f7000000f3000000e6000000ee",
            INIT_0A => X"000000d3000000d0000000df000000c9000000bd000000f7000000b7000000a2",
            INIT_0B => X"000000e7000000e4000000ee000000ec000000b6000000830000006b00000075",
            INIT_0C => X"000000b1000000de000000ad000000820000007500000056000000e9000000db",
            INIT_0D => X"000000a30000008e0000008f000000a0000000c2000000cf000000be000000a9",
            INIT_0E => X"000000ff000000f4000000e4000000c0000000b1000000d100000050000000ae",
            INIT_0F => X"000000c2000000c7000000c6000000c9000000d4000000c6000000c1000000e9",
            INIT_10 => X"000000ae000000c9000000d4000000d4000000d5000000d1000000cb00000092",
            INIT_11 => X"000000310000008a0000007f000000800000008f0000009a0000009b000000b4",
            INIT_12 => X"0000008a0000008b0000008b000000700000005c000000510000004c00000048",
            INIT_13 => X"000000170000000000000075000000680000006b000000680000006f0000007a",
            INIT_14 => X"00000029000000270000001a000000300000000000000000000000000000001a",
            INIT_15 => X"000000050000000000000000000000790000006b00000056000000420000002e",
            INIT_16 => X"0000003b0000002900000025000000450000003a000000000000000000000000",
            INIT_17 => X"00000000000000000000000000000009000000970000006a0000005300000051",
            INIT_18 => X"0000003f0000001f0000000e0000000000000000000000000000000000000000",
            INIT_19 => X"000000000000000000000000000000000000001e000000ad0000007f00000067",
            INIT_1A => X"000000760000006a0000004f0000002100000000000000010000000000000000",
            INIT_1B => X"000000000000000000000000000000000000000000000000000000b30000008c",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000350000000000000000",
            INIT_1F => X"0000001e00000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000160000001700000035",
            INIT_21 => X"0000000000000000000000000000001400000000000000000000000000000000",
            INIT_22 => X"0000004900000073000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000100000000000000000000000000000000000000610000004f00000032",
            INIT_25 => X"0000000000000000000000090000003b0000005400000075000000170000002f",
            INIT_26 => X"000000000000001f000000570000007b00000000000000000000000000000000",
            INIT_27 => X"000000510000003a000000120000000000000000000000000000003400000003",
            INIT_28 => X"00000000000000070000001f0000000000000000000000180000004c00000027",
            INIT_29 => X"00000000000000000000000f00000029000000460000002b0000000000000000",
            INIT_2A => X"0000001d00000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000004c0000003300000024000000000000000c000000000000000000000025",
            INIT_2C => X"0000002f00000031000000470000005300000059000000540000002f0000002a",
            INIT_2D => X"000000000000000200000001000000170000002e00000019000000200000001e",
            INIT_2E => X"0000005d000000640000006b0000006e000000660000005f000000300000005e",
            INIT_2F => X"00000006000000000000000000000000000000160000002f0000004900000050",
            INIT_30 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_31 => X"0000001800000017000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000700000000000000000000001400000003000000030000001a00000025",
            INIT_33 => X"000000030000000000000018000000000000000000000000000000110000003e",
            INIT_34 => X"0000000000000002000000460000001500000000000000000000000000000004",
            INIT_35 => X"0000000000000000000000000000000f00000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000b0000000a0000000a0000000a00000008000000000000000000000000",
            INIT_38 => X"0000000a000000090000000d0000000b0000000a000000080000000a0000000a",
            INIT_39 => X"0000000b0000000b0000000a0000000b0000000b000000090000000b0000000a",
            INIT_3A => X"0000000b0000000a0000001a0000002b000000060000000b0000000a0000000c",
            INIT_3B => X"00000010000000090000000b0000000a0000000b0000000b0000000a0000000c",
            INIT_3C => X"0000000c0000000c0000000a0000002a00000032000000100000001a00000009",
            INIT_3D => X"0000000000000022000000000000000a0000000a0000000e000000100000001a",
            INIT_3E => X"000000490000000e0000000f00000010000000360000001b0000001000000015",
            INIT_3F => X"000000140000000400000016000000000000000c0000000c000000310000004b",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE11;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE12 : if BRAM_NAME = "samplegold_layer0_instance12" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000100000000400000015000000430000002d000000270000001a0000000f",
            INIT_01 => X"0000000c0000002a000000280000002c00000015000000180000001200000012",
            INIT_02 => X"000000360000005c00000049000000180000004000000000000000090000000c",
            INIT_03 => X"000000130000001000000044000000460000004500000000000000000000001d",
            INIT_04 => X"000000470000001a00000032000000510000003e000000200000001d00000018",
            INIT_05 => X"0000002700000024000000290000002b0000000d000000150000000000000019",
            INIT_06 => X"000000190000000c00000002000000020000007f0000002d000000210000002b",
            INIT_07 => X"000000300000001d000000230000001e00000013000000000000002000000011",
            INIT_08 => X"000000470000004e0000004e0000005000000043000000590000003200000037",
            INIT_09 => X"000000350000003a000000340000004100000033000000420000003d00000039",
            INIT_0A => X"000000620000006100000057000000540000004b000000540000003c00000034",
            INIT_0B => X"0000002b0000002b000000450000004700000049000000480000004e0000005b",
            INIT_0C => X"0000001f0000004a0000002a000000130000000300000000000000340000000b",
            INIT_0D => X"0000000000000023000000160000001a0000001e0000002e0000003400000034",
            INIT_0E => X"00000000000000000000005f00000018000000110000000b0000001e00000027",
            INIT_0F => X"0000001200000000000000270000001a00000013000000120000000000000000",
            INIT_10 => X"0000000000000000000000000000002400000013000000120000001100000016",
            INIT_11 => X"0000000f000000050000000000000029000000200000000c0000000f00000003",
            INIT_12 => X"0000000400000009000000000000000300000022000000140000001000000010",
            INIT_13 => X"00000013000000130000001300000010000000250000001b000000140000000a",
            INIT_14 => X"0000001400000014000000130000001400000012000000130000001300000014",
            INIT_15 => X"000000130000001200000013000000130000000f000000150000001300000014",
            INIT_16 => X"000000120000001f000000210000000000000010000000120000001300000012",
            INIT_17 => X"0000001100000014000000120000001400000012000000100000001400000013",
            INIT_18 => X"0000001300000012000000330000003100000000000000000000000100000014",
            INIT_19 => X"0000002b00000000000000130000001400000017000000130000001a00000014",
            INIT_1A => X"0000001600000015000000130000004c0000001c000000090000001100000000",
            INIT_1B => X"0000000a0000002f0000000000000013000000120000003f0000000d00000000",
            INIT_1C => X"000000280000001d0000002c0000000000000000000000020000000c0000001f",
            INIT_1D => X"0000001a000000120000000e000000000000001900000003000000310000003f",
            INIT_1E => X"0000000a000000000000001f0000006b00000003000000190000000700000000",
            INIT_1F => X"000000140000005c000000350000001500000000000000010000002600000011",
            INIT_20 => X"00000001000000620000002c0000002100000005000000070000000000000002",
            INIT_21 => X"0000000000000000000000000000000e000000500000000e0000000a00000049",
            INIT_22 => X"000000390000002b0000001b000000c50000003b000000240000001e00000008",
            INIT_23 => X"000000080000001c000000120000001e0000000000000015000000080000002a",
            INIT_24 => X"000000000000000000000000000000000000006000000000000000020000000e",
            INIT_25 => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"000000000000000000000000000000000000000e000000000000002100000015",
            INIT_27 => X"0000001c00000017000000040000000000000000000000000000000000000000",
            INIT_28 => X"000000580000001d0000000b000000040000000b00000041000000000000002d",
            INIT_29 => X"0000003700000011000000250000003500000028000000160000000f00000005",
            INIT_2A => X"0000000000000088000000190000000c00000000000000100000002700000000",
            INIT_2B => X"0000000000000047000000350000002100000000000000000000000000000000",
            INIT_2C => X"00000000000000070000005500000019000000170000000f0000001c00000018",
            INIT_2D => X"0000001a000000000000003e0000003500000024000000440000002c00000000",
            INIT_2E => X"0000005300000026000000180000003e0000001e0000001d0000001c0000001f",
            INIT_2F => X"0000000000000000000000000000003d000000350000002e0000001f0000002e",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000100000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"000000000000000000000000000000000000000000000000000000220000002a",
            INIT_3A => X"0000000000000000000000000000001100000018000000000000000000000000",
            INIT_3B => X"0000000200000008000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000003f0000002d000000000000000000000000",
            INIT_3E => X"0000001a000000000000004d0000000000000010000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE12;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE13 : if BRAM_NAME = "samplegold_layer0_instance13" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000007000000120000000b00000000000000000000000000000000",
            INIT_05 => X"00000000000000000000003d0000004a0000003e0000003f0000006200000045",
            INIT_06 => X"0000000000000002000000000000000000000000000000000000001300000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000090000000900000001000000030000000b00000002",
            INIT_09 => X"000000000000000000000000000000000000000c000000200000000000000000",
            INIT_0A => X"0000002c000000000000000c0000001c0000001b000000190000001c00000020",
            INIT_0B => X"0000002c0000002c000000000000000000000000000000000000000000000024",
            INIT_0C => X"0000002d0000002c0000002d0000002c0000002c0000002c0000002c0000002c",
            INIT_0D => X"0000002c0000002c0000002c0000002c0000002c0000002c0000002c0000002a",
            INIT_0E => X"00000011000000300000002e0000002b0000002b0000002c0000002b0000002c",
            INIT_0F => X"0000002c0000002c0000002c0000002b0000002c0000002b0000002c00000020",
            INIT_10 => X"000000170000000d000000090000001700000031000000270000002f0000002c",
            INIT_11 => X"0000002e0000002d00000029000000260000001f0000002c0000002c0000002b",
            INIT_12 => X"00000027000000150000000a0000000f0000000e000000290000001900000039",
            INIT_13 => X"0000002a0000002b0000002b0000001000000000000000000000002a00000028",
            INIT_14 => X"0000000000000009000000110000001f0000002700000026000000280000002a",
            INIT_15 => X"0000000e000000190000002400000020000000360000001b0000001100000026",
            INIT_16 => X"00000024000000110000001a000000120000000b0000001f0000000f00000010",
            INIT_17 => X"0000000000000000000000000000003100000007000000000000000000000000",
            INIT_18 => X"00000000000000000000001e0000000c00000019000000220000002b00000000",
            INIT_19 => X"0000000c00000031000000170000000500000006000000040000000000000003",
            INIT_1A => X"00000026000000000000000c0000000000000000000000000000000000000000",
            INIT_1B => X"0000000c000000110000000c0000001d00000028000000290000002900000014",
            INIT_1C => X"00000000000000000000000e0000000000000000000000010000000e00000007",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000001c00000030000000380000002c00000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000002",
            INIT_25 => X"000000050000000000000004000000060000000000000001000000340000004a",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"00000000000000090000000300000000000000000000000d0000000400000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000700000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000010000000000000005000000000000000900000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_31 => X"0000001000000000000000000000000500000000000000000000000000000000",
            INIT_32 => X"0000000000000016000000000000000000000000000000000000000000000000",
            INIT_33 => X"00000000000000390000001e0000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000002a000000000000000000000000000000000000000e0000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000010000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000004",
            INIT_38 => X"0000000000000000000000000000000000000000000000090000000000000004",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000002b00000013000000000000001e00000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000700000024000000000000000c00000022",
            INIT_3E => X"0000001a00000016000000050000001600000049000000000000000000000000",
            INIT_3F => X"000000000000000000000000000000000000000000000000000000000000001a",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE13;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE14 : if BRAM_NAME = "samplegold_layer0_instance14" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001c0000001d0000001c000000190000001e0000005d0000000000000000",
            INIT_01 => X"000000000000000b0000000b0000000000000000000000000000000000000000",
            INIT_02 => X"0000000b0000001f0000001f00000024000000270000002c0000004b00000000",
            INIT_03 => X"0000000000000000000000030000000d00000012000000020000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000022000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000001000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000002e00000018000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000001e00000017000000200000000000000000000000160000003d0000002e",
            INIT_28 => X"0000000f00000004000000050000000b000000100000000f000000140000001a",
            INIT_29 => X"0000000800000000000000000000000a00000009000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000300000009000000000000000000000000",
            INIT_2B => X"0000000f0000001200000013000000070000000c000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000001000000002000000020000000000000000",
            INIT_2F => X"0000001900000015000000080000000a00000021000000250000000d00000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000007",
            INIT_31 => X"0000000000000000000000000000001000000013000000000000000000000012",
            INIT_32 => X"0000001b0000001600000011000000020000000000000000000000000000000c",
            INIT_33 => X"000000110000001e000000090000001c0000001b0000000b000000080000000d",
            INIT_34 => X"000000150000001e000000070000000d00000009000000180000001200000004",
            INIT_35 => X"0000000f0000000f0000000300000007000000070000000f0000001e00000015",
            INIT_36 => X"0000001f0000001b0000001a0000000d0000000f0000000a0000001b0000000a",
            INIT_37 => X"000000090000001d000000130000000500000010000000280000002400000019",
            INIT_38 => X"000000120000001900000025000000260000000a0000000e0000000e0000000e",
            INIT_39 => X"0000000b000000120000000000000005000000140000001b000000150000000f",
            INIT_3A => X"000000070000000b0000000b0000000900000008000000050000000a0000000d",
            INIT_3B => X"0000000b0000000b0000000b0000000a000000140000000c0000000a00000003",
            INIT_3C => X"000000350000003a0000003a0000003f0000003c0000002f000000080000000b",
            INIT_3D => X"0000002f0000002d0000002f0000002800000033000000330000002a00000032",
            INIT_3E => X"0000002d0000002b0000002f0000002f00000038000000340000002900000033",
            INIT_3F => X"000000320000002c0000002b000000320000002f000000190000002f00000029",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE14;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE15 : if BRAM_NAME = "samplegold_layer0_instance15" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000022000000200000002300000025000000240000002e0000002b00000021",
            INIT_01 => X"000000170000002d000000230000001f000000270000003c000000000000002a",
            INIT_02 => X"000000070000001900000017000000210000001a00000021000000270000002a",
            INIT_03 => X"0000000f0000000f0000001900000015000000250000001c0000001a0000000b",
            INIT_04 => X"00000019000000160000000e00000015000000120000000e0000001500000010",
            INIT_05 => X"000000110000002300000020000000150000000d0000001e0000002700000019",
            INIT_06 => X"000000300000001b0000001b0000001c0000002700000026000000240000001d",
            INIT_07 => X"0000002a000000180000001b0000002400000005000000160000000d0000002d",
            INIT_08 => X"00000022000000360000002d000000310000002f000000340000002a00000032",
            INIT_09 => X"0000003b0000003f000000380000002e0000002e00000000000000190000000b",
            INIT_0A => X"0000001b000000200000001900000011000000290000002e0000003500000037",
            INIT_0B => X"00000028000000350000003a000000390000001c000000310000002300000000",
            INIT_0C => X"0000001b0000001c000000210000002b000000190000002e0000002100000021",
            INIT_0D => X"0000002d000000320000002e0000002c00000031000000420000002d00000012",
            INIT_0E => X"00000009000000040000000c0000001c0000002600000021000000160000001f",
            INIT_0F => X"0000000f0000001500000023000000240000002100000031000000310000002e",
            INIT_10 => X"00000035000000030000000300000005000000080000000d0000001e0000002d",
            INIT_11 => X"000000140000000d0000001100000037000000260000001e0000001a0000002a",
            INIT_12 => X"000000180000002700000002000000050000000c000000010000000900000013",
            INIT_13 => X"000000060000000a0000001300000015000000110000000d0000001200000010",
            INIT_14 => X"0000000a0000000c0000000d0000000700000008000000010000000d0000000a",
            INIT_15 => X"0000000700000008000000150000000900000009000000050000000b0000000f",
            INIT_16 => X"0000000a000000080000000800000004000000090000000a0000000600000009",
            INIT_17 => X"000000090000000a0000000000000015000000030000000a0000000c0000000c",
            INIT_18 => X"0000005700000055000000440000002b00000078000000000000000a00000009",
            INIT_19 => X"0000005600000048000000560000005500000042000000670000005100000051",
            INIT_1A => X"0000005100000050000000570000003800000027000000720000004300000057",
            INIT_1B => X"0000005a0000005a0000003c000000110000008f000000430000005300000054",
            INIT_1C => X"000000670000004b0000004a0000004e0000002c000000220000006f0000003e",
            INIT_1D => X"000000370000004e000000610000003400000000000000ba0000003300000041",
            INIT_1E => X"000000640000005c0000003d000000500000003c00000044000000230000006c",
            INIT_1F => X"000000420000002b0000004e000000000000001a000000190000005a00000066",
            INIT_20 => X"000000500000006b00000039000000350000003a00000025000000390000002e",
            INIT_21 => X"000000180000001200000020000000560000000e0000001a000000300000004e",
            INIT_22 => X"0000003d0000003e0000005c0000003e0000002f000000270000000e00000050",
            INIT_23 => X"00000040000000380000002e0000005b0000001b000000730000001d00000000",
            INIT_24 => X"0000000a00000034000000330000003e00000041000000430000002600000009",
            INIT_25 => X"00000038000000310000003b0000003a00000071000000440000006b00000033",
            INIT_26 => X"00000021000000180000007c0000005300000063000000580000004f00000047",
            INIT_27 => X"0000006400000042000000200000005000000056000000150000006800000040",
            INIT_28 => X"00000040000000380000001a0000005d00000031000000460000005100000060",
            INIT_29 => X"000000420000003f00000054000000450000002600000049000000440000004c",
            INIT_2A => X"000000590000005b0000005f0000003f0000003e00000038000000610000004f",
            INIT_2B => X"00000073000000310000004a00000065000000540000004c000000330000002b",
            INIT_2C => X"0000003b000000360000004700000056000000560000003f000000000000004d",
            INIT_2D => X"0000004c000000730000001c00000027000000390000006f000000430000000e",
            INIT_2E => X"000000220000002d0000002a0000003400000033000000440000003800000029",
            INIT_2F => X"0000003800000033000000310000002f00000038000000440000006000000051",
            INIT_30 => X"00000022000000250000001f000000200000003e0000001f0000003000000031",
            INIT_31 => X"00000047000000040000002a0000002100000026000000290000001d00000024",
            INIT_32 => X"00000014000000110000001e000000210000001a000000230000002500000025",
            INIT_33 => X"0000001e000000510000000000000030000000230000001d0000001700000012",
            INIT_34 => X"000000000000000800000005000000080000003e000000160000001c00000021",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000002",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000008",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000a00000000000000000000000d00000021000000000000000000000000",
            INIT_3E => X"00000000000000000000000f0000002100000032000000000000000c0000001d",
            INIT_3F => X"0000000000000003000000060000000000000045000000690000002d00000008",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE15;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE16 : if BRAM_NAME = "samplegold_layer0_instance16" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000400000004f000000320000002000000010000000000000000000000000",
            INIT_01 => X"0000005e0000003a000000230000000000000000000000000000000000000034",
            INIT_02 => X"00000000000000000000000000000007000000160000001f0000002f00000059",
            INIT_03 => X"0000000000000000000000000000000000000072000000100000000000000000",
            INIT_04 => X"0000000c00000040000000200000000b00000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000170000004300000000000000000000000200000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000001100000019",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000002000000030000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"000000000000000000000001000000000000000000000000000000000000000b",
            INIT_0F => X"000000000000000000000000000000000000000b000000050000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000d0000000b000000020000000a00000001000000000000000000000000",
            INIT_12 => X"000000000000000000000000000000000000000b0000000e0000000f0000000d",
            INIT_13 => X"0000000f00000000000000250000000a00000009000000120000000d00000001",
            INIT_14 => X"0000001a00000013000000000000000000000000000000110000001600000019",
            INIT_15 => X"0000001d00000000000000000000002400000009000000110000002100000017",
            INIT_16 => X"00000024000000310000001f000000210000000700000010000000160000001e",
            INIT_17 => X"0000002300000000000000100000000000000000000000130000002400000023",
            INIT_18 => X"000000090000001c0000001f000000140000000d000000040000000100000024",
            INIT_19 => X"000000290000002e000000020000000000000000000000000000000000000001",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"000000000000001d000000140000003a00000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000190000003400000023000000190000000000000000",
            INIT_1E => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"00000000000000000000000000000012000000180000001a0000001800000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"000000000000000000000000000000000000001400000014000000080000000d",
            INIT_22 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000030000000c00000009",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"00000008000000000000000a0000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"000000040000000c000000000000000100000000000000000000000000000000",
            INIT_2F => X"0000002300000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"000000000000000b0000000f0000000000000005000000000000000000000009",
            INIT_31 => X"0000000e00000046000000000000000d00000001000000000000000000000000",
            INIT_32 => X"000000000000000f0000000e0000001900000000000000090000000000000000",
            INIT_33 => X"0000004100000015000000050000000000000000000000000000000000000004",
            INIT_34 => X"000000100000000d000000190000000300000009000000010000001700000000",
            INIT_35 => X"0000000000000019000000150000000000000000000000000000000000000006",
            INIT_36 => X"0000000000000000000000000000000c00000000000000110000000e00000012",
            INIT_37 => X"0000000000000018000000000000001200000025000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000a00000017000000000000000000000001",
            INIT_39 => X"0000000000000000000000040000000000000007000000210000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000030000000800000000",
            INIT_3B => X"0000000000000000000000080000000000000000000000170000001400000000",
            INIT_3C => X"0000000000000002000000000000000000000000000000000000000000000012",
            INIT_3D => X"0000000000000016000000000000000000000000000000000000000000000014",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000002000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE16;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE17 : if BRAM_NAME = "samplegold_layer0_instance17" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000002400000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000019000000000000000000000000",
            INIT_02 => X"000000000000000000000000000000000000000000000000000000000000001c",
            INIT_03 => X"0000000000000000000000000000000000000000000000110000000000000000",
            INIT_04 => X"0000000200000000000000020000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000600000000000000020000000000000000",
            INIT_06 => X"0000000300000005000000000000000100000000000000000000001100000000",
            INIT_07 => X"0000000000000000000000000000000200000004000000030000000800000002",
            INIT_08 => X"0000000000000000000000080000000400000004000000060000000000000022",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000400000000000000000000000000000001000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000010000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000003000000020000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000110000000500000000",
            INIT_27 => X"000000010000000a000000090000000200000000000000000000000000000000",
            INIT_28 => X"0000000000000004000000000000000800000005000000030000000e00000015",
            INIT_29 => X"0000001e0000001e000000230000000a00000004000000010000000000000000",
            INIT_2A => X"0000002d0000000f00000026000000090000000f000000110000002d00000012",
            INIT_2B => X"000000000000001a000000240000000f0000001d00000015000000250000002c",
            INIT_2C => X"0000003500000026000000270000003f0000003b0000003f0000004e00000012",
            INIT_2D => X"00000000000000030000000900000016000000390000003a0000004700000042",
            INIT_2E => X"0000000000000000000000000000000000000000000000170000000000000000",
            INIT_2F => X"00000000000000000000000000000000000000010000000d0000000000000000",
            INIT_30 => X"0000000000000000000000000000000400000000000000000000000c0000000d",
            INIT_31 => X"0000002f0000001b000000050000000000000000000000000000000000000000",
            INIT_32 => X"000000000000000000000000000000000000000000000000000000000000002c",
            INIT_33 => X"00000000000000000000000a0000000c000000100000001c0000001600000000",
            INIT_34 => X"00000000000000010000001a0000001300000001000000000000002300000016",
            INIT_35 => X"000000000000002f0000000e0000000100000000000000000000000000000000",
            INIT_36 => X"0000002b00000028000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000180000002e000000330000001c0000000000000004",
            INIT_38 => X"0000002600000000000000000000000000000013000000300000002300000000",
            INIT_39 => X"00000000000000000000000000000017000000120000001c0000002200000032",
            INIT_3A => X"0000001c00000004000000000000001e00000042000000000000000000000000",
            INIT_3B => X"0000002800000043000000370000001b00000004000000030000000000000005",
            INIT_3C => X"0000000500000002000000090000001b00000007000000040000000600000012",
            INIT_3D => X"0000000f00000005000000040000000a0000000400000000000000000000000e",
            INIT_3E => X"0000000000000001000000030000000000000000000000000000000000000010",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE17;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE18 : if BRAM_NAME = "samplegold_layer0_instance18" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000007000000020000000900000000",
            INIT_01 => X"000000f8000000f1000000fb000000f5000000f3000000c3000000df0000000d",
            INIT_02 => X"000000f4000000fd000000f5000000fb000000f600000100000000f4000000f9",
            INIT_03 => X"000000f9000000ef000000e5000000f4000000e9000000ec000000bf000000dd",
            INIT_04 => X"000000d4000000f1000000fe000000f3000000f8000000de000000ee000000f0",
            INIT_05 => X"000000e6000000da000000e0000000db000000e4000000da000000da000000b0",
            INIT_06 => X"0000009c000000c3000000ec000000ee000000ed000000f3000000bd000000d0",
            INIT_07 => X"000000a5000000a8000000b9000000ce000000cb000000cc000000cb000000c1",
            INIT_08 => X"000000930000007e00000097000000c8000000d2000000d30000008c0000007a",
            INIT_09 => X"00000074000000790000008d000000b8000000b2000000a9000000a400000097",
            INIT_0A => X"000000630000006c0000005e000000600000007d0000008d0000006800000064",
            INIT_0B => X"0000008e000000730000007c0000007d00000090000000910000007900000079",
            INIT_0C => X"000000a0000000740000006f0000006900000074000000580000009d0000006b",
            INIT_0D => X"000000ad000000b00000008f0000008b0000008600000092000000a2000000a0",
            INIT_0E => X"000000c6000000b8000000990000008a00000080000000860000005300000073",
            INIT_0F => X"00000065000000a2000000a200000098000000a5000000c4000000c2000000cf",
            INIT_10 => X"000000c8000000d0000000d2000000cf000000b00000009f000000a000000047",
            INIT_11 => X"0000009600000091000000a100000096000000810000009c000000a8000000ba",
            INIT_12 => X"000000af000000b5000000b5000000bb000000b5000000a9000000900000008b",
            INIT_13 => X"000000af000000640000007f00000096000000a7000000aa000000b4000000aa",
            INIT_14 => X"0000006f00000079000000ab000000bb000000a9000000a9000000b0000000b0",
            INIT_15 => X"000000a9000000940000003d00000050000000680000008b0000009e000000a4",
            INIT_16 => X"00000073000000660000006e0000009d0000009000000075000000790000009e",
            INIT_17 => X"0000008d0000008e0000007c0000002200000030000000410000005900000066",
            INIT_18 => X"00000044000000550000005800000057000000640000006f0000006a0000006d",
            INIT_19 => X"0000003c0000003c0000003d000000390000001b000000220000003500000038",
            INIT_1A => X"000000240000003100000037000000400000004000000045000000410000003f",
            INIT_1B => X"0000002b000000230000001f00000016000000180000001b0000001c00000021",
            INIT_1C => X"0000001b0000001a0000001f00000039000000370000002c000000320000002c",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000c0000001e",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"00000000000000000000000000000000000000000000003b0000000000000000",
            INIT_21 => X"0000001f00000008000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000001200000000000000000000000b00000003000000000000004500000007",
            INIT_23 => X"0000006e0000000b00000001000000000000000a000000000000001200000001",
            INIT_24 => X"00000040000000460000001f0000001d000000100000008b0000004600000046",
            INIT_25 => X"00000003000000040000003d0000003d0000004f00000050000000510000004a",
            INIT_26 => X"000000000000000000000000000000470000001b000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000800000000000000000000000000000000",
            INIT_28 => X"00000000000000110000000a0000000000000027000000000000000b00000000",
            INIT_29 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000380000005000000000",
            INIT_2B => X"0000000000000000000000110000003600000000000000020000000000000000",
            INIT_2C => X"0000001c00000011000000000000000500000027000000140000000000000000",
            INIT_2D => X"0000000000000002000000000000000000000000000000000000000000000015",
            INIT_2E => X"0000000000000000000000000000001a0000000000000000000000000000001f",
            INIT_2F => X"0000002c00000042000000360000001700000000000000000000000f00000022",
            INIT_30 => X"0000002c00000025000000000000002e00000017000000050000000000000000",
            INIT_31 => X"00000000000000230000001300000023000000360000003a0000001c00000002",
            INIT_32 => X"0000000f000000050000002000000003000000000000000e0000001c00000002",
            INIT_33 => X"0000002d0000000e0000000b0000001300000010000000160000002400000016",
            INIT_34 => X"0000001a000000230000000700000006000000290000002c0000001b00000028",
            INIT_35 => X"000000100000001f0000002c0000000000000003000000140000000b00000007",
            INIT_36 => X"0000000700000016000000000000001000000015000000150000000c00000005",
            INIT_37 => X"000000000000000000000000000000000000000000000000000000020000000b",
            INIT_38 => X"0000000200000005000000180000000000000012000000050000000000000000",
            INIT_39 => X"000000270000002e0000003b0000004500000024000000230000000000000000",
            INIT_3A => X"0000000c000000130000000e000000140000001d000000090000001900000020",
            INIT_3B => X"00000014000000190000001a00000030000000390000001a000000140000000e",
            INIT_3C => X"0000000a00000007000000160000003200000002000000170000001100000014",
            INIT_3D => X"000000030000000a0000000b00000009000000240000002d0000000d00000015",
            INIT_3E => X"000000170000000800000002000000250000005300000000000000210000001b",
            INIT_3F => X"0000000400000000000000060000000000000009000000110000002100000003",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE18;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE19 : if BRAM_NAME = "samplegold_layer0_instance19" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002a0000001000000007000000470000004b000000490000001e0000001f",
            INIT_01 => X"000000200000001200000026000000240000001f000000320000002800000033",
            INIT_02 => X"0000002c000000360000002800000000000000200000001c0000003500000028",
            INIT_03 => X"000000240000002c000000250000003400000026000000250000002d00000014",
            INIT_04 => X"000000260000002e0000003b000000000000000b000000000000001100000033",
            INIT_05 => X"00000033000000260000002b0000002d0000003600000031000000410000004d",
            INIT_06 => X"000000350000002b000000260000003200000000000000020000000000000014",
            INIT_07 => X"0000001a0000003000000011000000300000002e000000310000003300000034",
            INIT_08 => X"0000003e00000049000000550000003e00000040000000040000000000000007",
            INIT_09 => X"00000013000000120000001c000000000000002c0000002d0000003b0000003e",
            INIT_0A => X"000000350000003e0000003c0000003d00000047000000350000000800000009",
            INIT_0B => X"0000001300000017000000100000001f000000230000002f000000220000002a",
            INIT_0C => X"0000001f0000004400000042000000300000003d000000410000005000000023",
            INIT_0D => X"0000001b0000001a0000001c0000001c000000240000002f0000004b00000025",
            INIT_0E => X"00000020000000160000004b0000003d0000003a0000002c000000420000005f",
            INIT_0F => X"0000004b00000017000000230000002000000025000000230000002800000031",
            INIT_10 => X"0000002c0000002a0000002e000000390000003a000000350000002b00000038",
            INIT_11 => X"00000037000000380000002000000024000000190000002a000000210000002a",
            INIT_12 => X"000000160000003000000028000000300000002c0000002c0000003300000031",
            INIT_13 => X"00000026000000250000001d0000001f00000024000000210000002400000023",
            INIT_14 => X"000000250000000d000000410000001c00000027000000250000002600000028",
            INIT_15 => X"00000012000000280000001f000000000000000d000000250000002500000021",
            INIT_16 => X"0000001a00000007000000190000002300000009000000190000001100000019",
            INIT_17 => X"0000001e0000000c0000002a0000001e00000000000000160000001600000009",
            INIT_18 => X"00000005000000230000001f000000000000001b00000017000000170000000e",
            INIT_19 => X"0000000e000000210000000c0000002d00000016000000000000001b00000014",
            INIT_1A => X"00000017000000030000002800000059000000000000001e000000130000000c",
            INIT_1B => X"00000000000000170000000d0000001800000022000000180000000000000022",
            INIT_1C => X"000000190000001a00000037000000020000001200000000000000000000000e",
            INIT_1D => X"00000000000000000000000a0000000300000018000000000000000700000000",
            INIT_1E => X"0000002a000000130000000e0000003b00000022000000120000000800000000",
            INIT_1F => X"00000010000000000000001c00000015000000230000001c0000000a00000021",
            INIT_20 => X"0000000900000023000000000000003100000000000000460000003e0000000f",
            INIT_21 => X"0000001f0000001b000000060000000d000000030000001b0000003100000000",
            INIT_22 => X"000000270000001800000014000000000000000c00000000000000210000004c",
            INIT_23 => X"00000022000000000000000f0000000c00000013000000190000002200000032",
            INIT_24 => X"0000001a00000021000000000000000b00000025000000000000000900000020",
            INIT_25 => X"0000001b0000003d000000000000001c00000003000000040000000200000007",
            INIT_26 => X"0000000a000000070000002500000033000000000000000c000000070000000b",
            INIT_27 => X"000000000000000300000016000000170000000d0000000c0000001b0000001a",
            INIT_28 => X"0000001c00000015000000000000000f0000000f000000230000000400000000",
            INIT_29 => X"000000000000000000000000000000000000001f0000002f0000000000000000",
            INIT_2A => X"000000000000003e0000001100000000000000000000000c000000410000000b",
            INIT_2B => X"000000000000000b000000030000000000000003000000080000001800000004",
            INIT_2C => X"0000001700000004000000040000000a0000000b00000000000000080000002f",
            INIT_2D => X"0000000a0000000f0000000f000000000000001b00000005000000070000000d",
            INIT_2E => X"000000250000000a0000001000000014000000190000001a0000000d00000008",
            INIT_2F => X"0000001a0000001200000017000000170000000b0000000e0000000c00000005",
            INIT_30 => X"00000000000000390000000b0000001a0000001d0000001a0000001a0000001a",
            INIT_31 => X"000000000000000000000000000000000000001a000000150000000d00000014",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000d00000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000700000000000000000000000200000000",
            INIT_3C => X"0000000000000000000000000000000000000022000000180000000000000000",
            INIT_3D => X"0000001e0000000b000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000001200000003000000000000000000000000000000000000000000000013",
            INIT_3F => X"000000000000000000000000000000000000000000000000000000160000002c",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE19;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE20 : if BRAM_NAME = "samplegold_layer0_instance20" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000004500000000000000000000000000000000",
            INIT_01 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000006",
            INIT_0C => X"0000000000000000000000000000000100000001000000000000000000000000",
            INIT_0D => X"0000000000000005000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000002a000000240000002c0000002400000019000000190000000f00000008",
            INIT_0F => X"00000010000000000000000d000000240000002f000000280000002900000026",
            INIT_10 => X"000000000000003700000024000000290000002a000000210000002400000019",
            INIT_11 => X"0000002100000016000000000000001600000027000000320000002b0000002a",
            INIT_12 => X"0000001b0000000000000030000000150000001c00000031000000230000002e",
            INIT_13 => X"000000330000002400000026000000000000001c000000270000002e0000002d",
            INIT_14 => X"0000000000000000000000000000000000000010000000270000002900000026",
            INIT_15 => X"0000000700000006000000000000000000000000000000000000001c0000002a",
            INIT_16 => X"0000002700000008000000000000000000000000000000000000000400000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"000000000000000d0000002c0000000d00000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"00000000000000000000001d000000170000001d000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"000000000000000000000000000000000000001300000009000000000000000b",
            INIT_1D => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"00000000000000000000000000000014000000060000000a0000001400000008",
            INIT_1F => X"0000000800000001000000000000000400000000000000000000000000000000",
            INIT_20 => X"000000000000000000000000000000000000000000000000000000030000000d",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000003000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000038000000000000000000000002000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000300000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000010000001d00000010000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000100000000000000000000000c000000000000000c0000000000000000",
            INIT_33 => X"0000000b00000000000000000000001900000001000000000000000000000013",
            INIT_34 => X"0000000000000040000000000000000000000008000000040000000a00000000",
            INIT_35 => X"0000000000000000000000000000000000000007000000070000000000000038",
            INIT_36 => X"0000002600000026000000070000000000000000000000060000000600000000",
            INIT_37 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000006000000260000000000000000000000000000001b00000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"000000000000000000000007000000050000000000000004000000000000000a",
            INIT_3B => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_3C => X"00000000000000000000000000000002000000130000000e0000000800000000",
            INIT_3D => X"0000000700000000000000000000000f00000019000000000000000000000001",
            INIT_3E => X"000000000000001300000000000000000000001c00000012000000130000000c",
            INIT_3F => X"00000011000000180000000900000005000000080000000c0000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE20;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE21 : if BRAM_NAME = "samplegold_layer0_instance21" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000500000002000000020000000000000000000000170000001600000016",
            INIT_01 => X"0000001b0000000f000000120000000b000000140000000e0000000000000000",
            INIT_02 => X"0000001000000010000000070000000a000000020000000a0000001500000011",
            INIT_03 => X"0000001200000013000000140000000f0000003000000000000000120000000d",
            INIT_04 => X"0000001800000015000000120000001200000014000000120000001500000016",
            INIT_05 => X"0000002d0000000e00000014000000100000001200000029000000000000001b",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"000000000000000000000000000000000000001a000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000005000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000001c0000001d000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000002400000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"000000000000000000000000000000000000000000000000000000000000000d",
            INIT_31 => X"0000001e00000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000020000001400000029",
            INIT_33 => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000001300000026000000420000002d00000005",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"000000110000000f000000000000000000000000000000000000000000000000",
            INIT_37 => X"000000040000001f00000013000000010000000d000000200000001b00000016",
            INIT_38 => X"000000000000000000000000000000160000001f000000140000000100000011",
            INIT_39 => X"000000140000000f000000090000000600000000000000000000000000000000",
            INIT_3A => X"0000000b0000000f000000110000000a000000210000001a0000001b00000018",
            INIT_3B => X"0000000000000000000000000000000000000000000000010000000600000004",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000002e000000300000002a0000002900000035000000320000000d00000000",
            INIT_3F => X"00000032000000330000002c0000002e0000002e0000002d0000002e0000002b",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE21;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE22 : if BRAM_NAME = "samplegold_layer0_instance22" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000280000003200000042000000230000003100000039000000340000002e",
            INIT_01 => X"0000003400000034000000390000002e000000270000002d0000002a00000030",
            INIT_02 => X"0000002b0000001b0000002a0000001d00000026000000360000003600000034",
            INIT_03 => X"000000350000003600000033000000280000002c000000280000002100000020",
            INIT_04 => X"000000430000003c000000340000003b0000003d000000450000002700000038",
            INIT_05 => X"000000380000003200000037000000370000004c000000380000003d0000003a",
            INIT_06 => X"000000260000002b000000300000002a00000028000000280000002600000035",
            INIT_07 => X"00000026000000310000002e0000003500000033000000340000003600000029",
            INIT_08 => X"000000340000003300000035000000380000003900000035000000340000002e",
            INIT_09 => X"0000002d0000001f000000230000002f00000037000000330000003300000037",
            INIT_0A => X"000000340000003600000035000000380000003a0000003a0000002f0000002a",
            INIT_0B => X"0000001e0000000d0000002a0000003400000033000000350000003300000033",
            INIT_0C => X"0000003500000034000000340000003200000035000000300000002900000030",
            INIT_0D => X"0000001000000000000000290000003000000032000000320000003800000034",
            INIT_0E => X"00000033000000350000003700000032000000230000001e0000002200000018",
            INIT_0F => X"0000000c00000008000000000000002b00000032000000310000003000000037",
            INIT_10 => X"00000034000000240000001a00000019000000200000000c0000000b0000000c",
            INIT_11 => X"0000004500000026000000140000002d00000019000000320000003300000033",
            INIT_12 => X"0000001b0000003b000000390000004700000023000000260000002100000025",
            INIT_13 => X"0000002200000020000000140000000a0000001100000012000000130000001a",
            INIT_14 => X"00000020000000170000002e000000300000002a000000270000002600000023",
            INIT_15 => X"00000016000000150000001d000000170000001100000013000000150000001d",
            INIT_16 => X"000000090000000b000000030000001300000013000000170000001600000013",
            INIT_17 => X"0000000200000000000000030000000600000007000000040000000000000006",
            INIT_18 => X"0000000300000003000000040000000000000015000000000000000000000001",
            INIT_19 => X"0000000000000002000000050000000300000006000000070000000900000000",
            INIT_1A => X"0000003200000041000000640000004a0000001d000000000000001800000004",
            INIT_1B => X"0000003100000040000000410000003c0000003f000000390000004700000044",
            INIT_1C => X"0000004100000039000000700000006200000045000000260000004800000042",
            INIT_1D => X"00000050000000440000002d00000048000000490000004b000000380000004f",
            INIT_1E => X"000000430000003700000054000000540000006700000047000000270000004b",
            INIT_1F => X"0000004c00000054000000350000003b000000420000004b000000400000002a",
            INIT_20 => X"00000038000000490000003c0000003b00000042000000760000004400000031",
            INIT_21 => X"000000460000004c0000004e000000150000004200000037000000550000003e",
            INIT_22 => X"0000004e00000043000000400000004500000047000000700000005500000045",
            INIT_23 => X"0000006000000044000000500000005000000051000000290000003f00000052",
            INIT_24 => X"0000005200000059000000540000004b0000004e00000053000000470000005c",
            INIT_25 => X"00000063000000650000003a0000004a0000005000000052000000490000004c",
            INIT_26 => X"000000530000005d00000057000000560000004e00000043000000230000002f",
            INIT_27 => X"0000008400000064000000530000003300000050000000550000005500000059",
            INIT_28 => X"00000054000000510000005a000000590000004d000000230000000700000044",
            INIT_29 => X"000000cd00000062000000560000004d000000330000004f0000005500000053",
            INIT_2A => X"00000056000000550000003e0000004e000000390000001b0000000400000015",
            INIT_2B => X"00000016000000d20000007e000000530000004d000000310000005000000054",
            INIT_2C => X"000000410000003a00000038000000080000002800000016000000180000000f",
            INIT_2D => X"0000000000000064000000430000007800000050000000510000002b0000004c",
            INIT_2E => X"0000003d00000028000000000000001800000013000000340000003900000000",
            INIT_2F => X"0000003c000000590000007a0000005e0000006500000068000000690000003e",
            INIT_30 => X"000000290000005600000058000000550000005c000000560000006000000061",
            INIT_31 => X"0000004e00000034000000380000003a000000390000003e000000420000003b",
            INIT_32 => X"00000022000000250000003f0000004e00000044000000400000004600000043",
            INIT_33 => X"0000001c0000001f000000180000001a0000001a000000200000001900000028",
            INIT_34 => X"000000180000001900000022000000000000000a000000140000001700000014",
            INIT_35 => X"0000001700000011000000130000000800000016000000080000001600000013",
            INIT_36 => X"000000010000000900000007000000010000003b000000050000000000000016",
            INIT_37 => X"0000000200000008000000060000000c00000005000000060000000400000000",
            INIT_38 => X"00000000000000000000000000000000000000000000000d000000180000000d",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"000000310000000d000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000280000002f000000340000002e0000002400000012",
            INIT_3C => X"0000001200000005000000060000002000000000000000000000000600000000",
            INIT_3D => X"00000000000000000000000f0000000600000000000000000000000100000009",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000010",
            INIT_3F => X"0000000800000000000000000000001400000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE22;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE23 : if BRAM_NAME = "samplegold_layer0_instance23" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002b000000270000002c0000002e00000030000000000000000000000000",
            INIT_01 => X"0000000800000002000000030000000000000000000000180000002200000027",
            INIT_02 => X"000000050000000500000002000000000000000000000000000000000000001a",
            INIT_03 => X"0000002100000003000000010000000000000000000000000000000000000000",
            INIT_04 => X"000000000000000000000000000000000000000000000000000000140000007e",
            INIT_05 => X"0000000000000000000000000000000100000000000000000000000100000000",
            INIT_06 => X"0000000200000000000000000000000000000000000000000000000000000023",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"000000b70000007e000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000002f0000006d00000075000000a300000074000000a30000007d00000067",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000003",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000010000000b00000007000000090000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"00000000000000000000003b0000000000000000000000000000000000000000",
            INIT_11 => X"000000180000001300000014000000180000000c000000000000000000000000",
            INIT_12 => X"000000000000000000000000000000000000004e000000130000000400000010",
            INIT_13 => X"0000000700000005000000050000000200000007000000000000000000000007",
            INIT_14 => X"0000004800000000000000000000000000000000000000050000000000000005",
            INIT_15 => X"0000002000000030000000360000003c000000370000003b0000003300000046",
            INIT_16 => X"0000003900000039000000000000000000000000000000000000000000000000",
            INIT_17 => X"00000000000000310000003100000039000000320000003d0000004a0000003c",
            INIT_18 => X"0000002d000000370000005a0000000d00000000000000000000000000000000",
            INIT_19 => X"00000000000000220000003700000041000000490000003a0000003f0000003d",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"00000000000000000000000000000000000000000000001a0000001d00000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"00000000000000000000000000000000000000000000002b0000001a00000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000e00000015000000120000003f00000002",
            INIT_23 => X"0000001b00000002000000060000000000000000000000000000000000000000",
            INIT_24 => X"00000004000000060000001e0000001a000000150000000f000000130000002f",
            INIT_25 => X"0000000c00000007000000000000000100000000000000000000000000000000",
            INIT_26 => X"0000000000000012000000060000000f0000000f000000000000000c00000023",
            INIT_27 => X"0000000000000000000000020000000100000000000000000000000000000004",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000001300000013000000160000001b0000001200000012000000150000001f",
            INIT_2C => X"0000002000000000000000080000001100000012000000130000001500000015",
            INIT_2D => X"0000001600000013000000150000000d00000015000000140000001100000011",
            INIT_2E => X"0000000000000011000000020000000000000000000000180000001800000016",
            INIT_2F => X"0000000000000000000000030000000000000000000000060000000200000000",
            INIT_30 => X"00000000000000000000000f00000000000000050000000b0000000000000000",
            INIT_31 => X"0000001b0000001b0000001e0000002e00000015000000260000003f00000000",
            INIT_32 => X"0000001400000000000000000000000f00000000000000000000000600000025",
            INIT_33 => X"000000220000001c0000001c0000001d00000033000000260000002d0000000c",
            INIT_34 => X"0000002b00000039000000000000000000000008000000000000000000000010",
            INIT_35 => X"0000004000000021000000310000001e0000002b000000330000001800000029",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000002000000150000000300000000000000000000000300000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"000000000000000000000002000000290000001b000000000000000000000000",
            INIT_3B => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000220000003d00000000000000000000000000000000",
            INIT_3D => X"0000000000000008000000000000000000000000000000000000000000000000",
            INIT_3E => X"000000020000001c0000002e0000002300000016000000000000000000000000",
            INIT_3F => X"0000000000000000000000090000000000000000000000000000000000000007",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE23;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE24 : if BRAM_NAME = "samplegold_layer0_instance24" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000034000000050000000b000000150000001d000000140000000000000000",
            INIT_01 => X"0000000000000000000000000000000e00000000000000050000001600000021",
            INIT_02 => X"000000000000000600000000000000000000004f0000000f0000000000000000",
            INIT_03 => X"000000000000000000000000000000000000000f0000000c0000000e00000048",
            INIT_04 => X"0000000000000000000000010000000000000000000000120000000000000000",
            INIT_05 => X"0000000000000002000000010000000200000007000000060000000700000003",
            INIT_06 => X"0000000000000005000000070000000100000004000000000000000e00000007",
            INIT_07 => X"0000000d00000008000000030000000b000000080000000c0000000000000004",
            INIT_08 => X"000000170000000800000008000000090000000a00000003000000050000000c",
            INIT_09 => X"0000000f0000000800000010000000070000000d0000000a0000000800000000",
            INIT_0A => X"00000000000000000000000e0000000f00000003000000060000000700000004",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000a0000000f0000001000000012000000120000000b0000000400000000",
            INIT_0E => X"000000000000000000000000000000000000000000000000000000070000000a",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000010",
            INIT_10 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"000000000000000b0000000a0000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000001d0000000300000000000000030000000f000000060000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000b0000001f",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"000000100000000f0000000f0000001400000018000000140000000f00000002",
            INIT_24 => X"0000000000000001000000000000000400000005000000050000000b0000000c",
            INIT_25 => X"0000000000000000000000010000000000000000000000010000000600000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000003f000000380000003d00000042000000240000000d0000000000000000",
            INIT_2A => X"000000000000000000000003000000060000000a000000330000003f00000040",
            INIT_2B => X"00000010000000130000001d0000001a000000120000001a0000003a00000005",
            INIT_2C => X"00000001000000000000000000000004000000040000001a0000001300000011",
            INIT_2D => X"0000000100000004000000000000000000000001000000010000000600000000",
            INIT_2E => X"0000000500000000000000000000000000000005000000040000000000000000",
            INIT_2F => X"0000000100000000000000060000000b00000000000000000000000300000000",
            INIT_30 => X"0000000000000001000000300000001300000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"00000017000000610000002a0000000000000000000000000000000000000000",
            INIT_33 => X"0000000800000007000000080000000400000000000000000000000000000000",
            INIT_34 => X"0000004900000045000000000000000000000000000000000000000000000008",
            INIT_35 => X"000000000000000000000000000000010000000000000006000000020000000a",
            INIT_36 => X"0000005a00000009000000000000000300000004000000000000000100000000",
            INIT_37 => X"0000000000000001000000010000000000000000000000130000004500000075",
            INIT_38 => X"00000000000000050000000e00000013000000340000001a0000000300000005",
            INIT_39 => X"000000010000000100000009000000370000007400000082000000470000000c",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000001",
            INIT_3B => X"000000800000007a0000006e0000000000000000000000000000000000000000",
            INIT_3C => X"00000048000000510000005700000052000000700000008b0000008400000083",
            INIT_3D => X"00000018000000100000000c0000000c000000400000003a000000340000004a",
            INIT_3E => X"0000003e0000003c0000003a0000003400000027000000220000001f00000019",
            INIT_3F => X"00000004000000040000000c0000000b0000000a0000003f0000004300000043",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE24;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE25 : if BRAM_NAME = "samplegold_layer0_instance25" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000002000000000000000200000003",
            INIT_01 => X"0000000000000000000000000000000000000000000000020000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"000000bb000000c0000000b3000000a7000000bc000000d5000000c00000000d",
            INIT_04 => X"000000d4000000cb000000bf000000ba000000bc000000b9000000b5000000b8",
            INIT_05 => X"0000008d0000008e000000920000008a00000085000000e0000000e1000000c5",
            INIT_06 => X"000000c3000000db000000df000000d20000009e000000960000009800000091",
            INIT_07 => X"0000007e0000006c00000065000000730000008100000074000000e0000000de",
            INIT_08 => X"000000db000000be000000e4000000e2000000c0000000840000008100000083",
            INIT_09 => X"00000099000000970000008d0000008e000000940000009000000072000000cd",
            INIT_0A => X"000000d8000000d8000000c7000000e3000000e20000009e000000a200000095",
            INIT_0B => X"000000b0000000b8000000ba000000b5000000b4000000b2000000b1000000c0",
            INIT_0C => X"000000d6000000cf000000d6000000d6000000df000000dc000000cb000000cc",
            INIT_0D => X"000000cc000000c6000000c5000000c6000000ca000000c5000000c3000000c3",
            INIT_0E => X"000000d2000000980000008b000000c5000000db000000de000000dd000000df",
            INIT_0F => X"000000de000000dd000000da000000da000000de000000e1000000dd000000dd",
            INIT_10 => X"0000009f000000490000007d000000d7000000e7000000e1000000e3000000e0",
            INIT_11 => X"000000db000000db000000da000000d9000000dc000000df000000e2000000da",
            INIT_12 => X"0000005d0000003c00000064000000de000000e6000000e9000000e1000000de",
            INIT_13 => X"000000df000000dc000000da000000d8000000d8000000d4000000ce000000a9",
            INIT_14 => X"00000037000000350000002900000075000000dd000000e7000000e3000000e1",
            INIT_15 => X"000000e1000000da000000d8000000d3000000bf0000008b0000005f0000003e",
            INIT_16 => X"00000065000000530000002a0000002c0000007f000000d1000000e4000000de",
            INIT_17 => X"000000d0000000ce000000ca000000a300000073000000350000004000000043",
            INIT_18 => X"000000ba000000cb000000ae000000a3000000c6000000cc000000cd000000cf",
            INIT_19 => X"000000640000006b0000006b000000c8000000c9000000b8000000bc000000b9",
            INIT_1A => X"000000700000007000000071000000650000005800000058000000570000005d",
            INIT_1B => X"0000003d000000480000004900000046000000700000007b0000007b00000074",
            INIT_1C => X"0000002500000027000000280000003300000033000000330000003500000037",
            INIT_1D => X"0000002100000021000000240000002300000024000000400000002600000022",
            INIT_1E => X"0000002d0000001d0000001c0000001e00000022000000200000001e00000023",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000005300000050",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000002000000018000000170000002900000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000300000016000000140000001a00000013",
            INIT_23 => X"0000000000000000000000000000000000000000000000060000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000008",
            INIT_27 => X"0000000100000003000000000000000000000006000000000000000700000000",
            INIT_28 => X"0000001c0000000b000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000007400000015000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000015",
            INIT_2C => X"0000004c00000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000038",
            INIT_2E => X"000000070000002d000000000000000000000000000000000000000000000000",
            INIT_2F => X"00000000000000000000000000000000000000080000002a000000610000004d",
            INIT_30 => X"000000000000001e0000004f0000002000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000210000005f0000007c000000700000002400000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000003f00000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"000000480000002b0000001f0000003c000000630000005f0000005c00000052",
            INIT_35 => X"0000000000000000000000310000003b000000300000000d0000002a0000001a",
            INIT_36 => X"000000200000001e000000100000000000000000000000000000000000000000",
            INIT_37 => X"00000029000000320000003a00000039000000340000002f0000002d00000028",
            INIT_38 => X"000000050000000c0000000a00000012000000170000001e000000200000001c",
            INIT_39 => X"0000000000000000000000000000000a00000000000000000000000300000003",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000002700000017000000130000002b000000360000003e0000000000000000",
            INIT_3C => X"0000001d000000190000001b0000001c000000190000001c000000180000001d",
            INIT_3D => X"0000000500000007000000000000001a0000003b0000003b0000001700000016",
            INIT_3E => X"0000001c0000001f000000130000000200000000000000000000000800000000",
            INIT_3F => X"000000000000000000000000000000000000001b000000390000003c0000001d",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE25;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE26 : if BRAM_NAME = "samplegold_layer0_instance26" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000200000001e000000220000000000000000000000000000000000000000",
            INIT_01 => X"00000008000000000000000900000006000000000000000b0000003700000036",
            INIT_02 => X"0000002a0000002600000024000000260000000600000009000000000000000d",
            INIT_03 => X"0000002300000023000000260000002700000025000000120000002700000037",
            INIT_04 => X"000000240000002400000027000000220000001c0000002c000000220000001a",
            INIT_05 => X"0000001700000016000000170000001c0000001b00000019000000240000002a",
            INIT_06 => X"0000000b00000010000000250000002600000021000000240000002600000018",
            INIT_07 => X"000000210000001b0000001e00000022000000260000002e0000004a0000003e",
            INIT_08 => X"0000000000000000000000220000002b0000002700000023000000220000001f",
            INIT_09 => X"0000001f0000001e0000001a0000001c000000220000003f0000005200000012",
            INIT_0A => X"0000000000000002000000170000001d00000027000000290000002000000021",
            INIT_0B => X"000000200000001e0000002a0000002600000035000000460000003d0000001d",
            INIT_0C => X"0000001b00000000000000070000001800000018000000230000002800000022",
            INIT_0D => X"0000002900000035000000410000005b000000320000001e0000000f00000017",
            INIT_0E => X"000000150000000000000000000000000000001b000000190000002b00000025",
            INIT_0F => X"0000002800000020000000360000000300000003000000000000000000000026",
            INIT_10 => X"000000390000001d000000110000002e00000028000000250000002500000032",
            INIT_11 => X"0000001a000000350000003800000031000000240000002c000000270000002d",
            INIT_12 => X"000000230000002a0000001a000000120000001400000012000000140000001a",
            INIT_13 => X"0000002200000016000000390000002f00000034000000330000002c0000002b",
            INIT_14 => X"0000000e00000011000000180000001800000017000000110000001c0000001e",
            INIT_15 => X"0000000f00000011000000030000002500000016000000110000001100000012",
            INIT_16 => X"0000000600000007000000060000000c00000009000000100000000b0000000f",
            INIT_17 => X"0000000b00000000000000150000003400000010000000200000001e00000007",
            INIT_18 => X"000000090000000d0000000d0000000c0000000d000000080000000d00000018",
            INIT_19 => X"0000000e00000000000000010000001c00000031000000150000001b00000017",
            INIT_1A => X"0000001d00000004000000000000000000000000000000060000000000000000",
            INIT_1B => X"0000001b0000000000000000000000050000001a0000002f0000000e0000000c",
            INIT_1C => X"00000012000000210000001c00000017000000100000000f0000001900000000",
            INIT_1D => X"0000000000000002000000030000000000000000000000180000002900000011",
            INIT_1E => X"0000000f0000000f0000001f0000000500000005000000000000000000000006",
            INIT_1F => X"0000000e00000008000000080000000b000000000000000b0000001a0000001e",
            INIT_20 => X"0000001f0000000d000000100000000e00000023000000100000000100000007",
            INIT_21 => X"0000000d0000001100000019000000150000001300000015000000010000000e",
            INIT_22 => X"0000000000000025000000110000000d0000000d0000001d0000001700000013",
            INIT_23 => X"000000080000000a0000000b0000000f0000001a0000001f0000000d00000000",
            INIT_24 => X"00000000000000100000002f0000000c0000000c0000000d0000000b0000000f",
            INIT_25 => X"0000000d0000000300000005000000120000002d0000003c0000000000000000",
            INIT_26 => X"000000000000000d00000016000000340000000e0000000a0000000e0000000b",
            INIT_27 => X"000000090000001400000012000000190000001f0000002e0000002600000000",
            INIT_28 => X"00000000000000020000000d00000013000000320000000c0000000b00000009",
            INIT_29 => X"0000001d000000150000001b000000010000001b0000001c0000001f0000000c",
            INIT_2A => X"0000000000000000000000000000000f0000000d000000310000001000000019",
            INIT_2B => X"0000002b00000062000000110000002d0000000000000021000000530000001e",
            INIT_2C => X"0000001100000000000000000000000000000000000000000000002000000018",
            INIT_2D => X"0000000000000000000000080000000000000008000000000000000000000026",
            INIT_2E => X"0000001d000000170000001200000018000000100000000b0000000b00000014",
            INIT_2F => X"0000000000000004000000010000000a0000000d000000080000000c00000005",
            INIT_30 => X"0000001200000014000000100000000b000000080000000c0000000400000006",
            INIT_31 => X"0000001400000002000000450000001c00000018000000180000001800000011",
            INIT_32 => X"0000001a00000016000000210000001800000020000000140000001b00000015",
            INIT_33 => X"000000000000000000000000000000110000004d0000002d0000001d00000018",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE26;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE27 : if BRAM_NAME = "samplegold_layer0_instance27" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000002500000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000005100000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000003b0000004900000065000000510000005400000064000000480000005e",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000020000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000200000003000000030000000000000000000000000000000000000000",
            INIT_0F => X"0000000e00000007000000000000002400000005000000000000000000000007",
            INIT_10 => X"00000012000000130000000d00000014000000110000000e0000001100000010",
            INIT_11 => X"0000000c00000005000000010000001c0000001e000000110000001300000014",
            INIT_12 => X"000000270000002d0000002f000000260000002a000000280000002700000030",
            INIT_13 => X"000000250000001600000003000000000000001b0000001a0000001e0000001a",
            INIT_14 => X"00000038000000370000003a0000003300000034000000380000003000000035",
            INIT_15 => X"0000001e0000002a00000018000000020000000100000019000000190000001f",
            INIT_16 => X"000000160000002200000020000000240000001e000000260000002100000019",
            INIT_17 => X"000000070000000a0000001c00000007000000040000000a0000001400000012",
            INIT_18 => X"000000150000001d000000070000000f0000000d0000000d0000000e00000004",
            INIT_19 => X"0000001400000010000000130000000700000006000000100000000f00000012",
            INIT_1A => X"0000001200000014000000120000001600000015000000130000001500000018",
            INIT_1B => X"00000016000000130000000c00000000000000000000000d0000000d00000014",
            INIT_1C => X"0000001500000014000000150000001500000015000000150000001800000016",
            INIT_1D => X"0000001b0000001900000000000000000000000b000000250000001300000014",
            INIT_1E => X"0000001b00000018000000100000001300000014000000150000001600000016",
            INIT_1F => X"00000012000000000000000000000000000000000000001d0000001d0000001e",
            INIT_20 => X"0000001f0000001f0000001b000000110000001200000016000000180000000f",
            INIT_21 => X"000000000000000000000000000000000000000000000000000000100000002e",
            INIT_22 => X"0000001f0000001c0000001d0000001a000000160000000d0000000000000000",
            INIT_23 => X"0000000000000000000000000000001900000000000000000000001b00000000",
            INIT_24 => X"000000080000000b0000000e000000100000000c000000100000001a00000000",
            INIT_25 => X"0000000f000000010000000800000000000000070000000c0000000500000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000003",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000001000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000024000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"000000000000000000000000000000390000002f000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000300000063000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000d0000000e00000001000000000000000c0000004f0000000700000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000f0000002a0000001700000000000000100000004c0000000000000002",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE27;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE28 : if BRAM_NAME = "samplegold_layer0_instance28" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000025",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000500000003000000000000000000000002000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000004",
            INIT_04 => X"0000000f00000013000000050000000500000003000000140000000000000000",
            INIT_05 => X"0000000f0000001400000016000000140000001a000000130000000c0000000c",
            INIT_06 => X"000000170000000b000000160000001400000012000000140000001d00000006",
            INIT_07 => X"0000003e0000001c000000090000001d0000001e000000190000001b00000011",
            INIT_08 => X"0000000000000000000000000000000c00000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000001500000000000000070000000000000000",
            INIT_0A => X"000000000000000000000007000000000000000d000000000000000000000000",
            INIT_0B => X"000000000000000000000000000000000000002c000000000000000e00000000",
            INIT_0C => X"00000000000000000000000000000000000000000000000f0000000000000000",
            INIT_0D => X"000000000000000000000013000000000000000000000000000000000000000b",
            INIT_0E => X"0000000000000015000000000000003200000000000000000000000700000000",
            INIT_0F => X"0000000000000004000000000000000000000000000000000000000700000000",
            INIT_10 => X"0000000100000000000000000000000000000000000000240000000000000000",
            INIT_11 => X"000000000000000f0000000000000000000000000000001f0000000000000000",
            INIT_12 => X"0000000400000000000000080000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000002200000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000300000023",
            INIT_16 => X"0000002000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000016000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000005000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000004",
            INIT_1C => X"0000000700000000000000060000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000003000000020000000000000008000000000000000000000000",
            INIT_1F => X"000000000000000000000000000000000000000000000000000000000000000f",
            INIT_20 => X"00000007000000070000000a0000000000000000000000000000000000000000",
            INIT_21 => X"0000001200000000000000000000000000000000000000210000001100000008",
            INIT_22 => X"0000000000000003000000000000000000000009000000090000002b00000000",
            INIT_23 => X"0000000d0000000d000000170000000000000000000000000000001000000004",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"000000000000000b000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000009000000050000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000002000000040000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"000000000000000d0000001b0000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"00000000000000000000000d0000000000000000000000070000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE28;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE29 : if BRAM_NAME = "samplegold_layer0_instance29" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"000000000000000c000000000000001100000000000000000000000000000004",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_06 => X"0000001200000000000000000000000000000000000000000000000000000007",
            INIT_07 => X"0000000e00000000000000000000000000000000000000010000000000000000",
            INIT_08 => X"00000000000000000000000a0000000000000000000000010000000000000000",
            INIT_09 => X"000000000000000f000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_0B => X"0000000000000002000000080000000000000000000000000000000000000001",
            INIT_0C => X"0000000a00000006000000060000000500000006000000000000000000000000",
            INIT_0D => X"0000000000000000000000070000000200000000000000000000000000000000",
            INIT_0E => X"000000020000000f000000130000000b000000000000000d0000000500000002",
            INIT_0F => X"0000000000000012000000000000000000000001000000000000000000000000",
            INIT_10 => X"00000000000000050000000d000000050000000b0000000b0000000800000014",
            INIT_11 => X"0000000a00000015000000000000000000000000000000000000000200000000",
            INIT_12 => X"0000000500000000000000000000000400000009000000080000001400000014",
            INIT_13 => X"0000000f00000022000000000000000700000000000000000000000100000000",
            INIT_14 => X"0000000800000000000000000000000000000004000000080000000c0000000c",
            INIT_15 => X"000000100000000e0000000d0000000b00000000000000000000000000000008",
            INIT_16 => X"0000000000000000000000000000000000000000000000070000000f00000007",
            INIT_17 => X"0000000c00000006000000000000000100000001000000000000000000000000",
            INIT_18 => X"000000000000000000000000000000000000000000000000000000010000000f",
            INIT_19 => X"000000090000000c000000140000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000001000000000000000000000000000000030000000000000001",
            INIT_1B => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_1C => X"000000520000000800000000000000150000001b000000140000000000000000",
            INIT_1D => X"00000091000000000000003e000000000000000f000000000000001800000000",
            INIT_1E => X"000000000000004e0000000d0000001b00000010000000100000000000000000",
            INIT_1F => X"000000000000007c000000000000003f000000000000001d0000000000000008",
            INIT_20 => X"0000000000000000000000390000001e0000000e0000000c000000330000002b",
            INIT_21 => X"000000310000000c0000006000000000000000000000003d0000000000000022",
            INIT_22 => X"000000250000002c0000000000000000000000290000002f0000000000000033",
            INIT_23 => X"00000030000000840000001b0000004600000000000000000000002500000000",
            INIT_24 => X"00000008000000000000005600000006000000000000002d0000005d00000000",
            INIT_25 => X"0000000000000047000000ab0000002500000029000000000000001d00000000",
            INIT_26 => X"000000090000001a000000000000002b00000003000000000000004c00000020",
            INIT_27 => X"000000000000000000000038000000a90000001500000041000000000000001f",
            INIT_28 => X"0000001000000014000000190000000e00000011000000100000003000000033",
            INIT_29 => X"0000002a00000000000000000000002b00000084000000060000002a00000004",
            INIT_2A => X"00000003000000180000000e0000001f0000001a000000000000002200000020",
            INIT_2B => X"00000006000000170000001d0000000400000001000000730000001600000050",
            INIT_2C => X"000000520000001700000027000000170000001d000000200000000800000048",
            INIT_2D => X"0000000000000016000000040000002d00000027000000210000004a00000032",
            INIT_2E => X"0000001900000052000000320000001f0000003b000000250000001c00000022",
            INIT_2F => X"000000000000001e000000070000000000000032000000000000005c00000000",
            INIT_30 => X"0000001800000003000000360000002900000024000000400000003800000034",
            INIT_31 => X"0000002700000007000000000000002f00000000000000410000000500000000",
            INIT_32 => X"00000017000000170000000000000037000000310000001c000000460000002c",
            INIT_33 => X"0000000000000059000000220000000000000026000000280000002e00000000",
            INIT_34 => X"00000000000000450000001e00000000000000490000003c000000290000002a",
            INIT_35 => X"0000001f00000000000000200000000b00000010000000350000000800000000",
            INIT_36 => X"00000000000000190000005a0000000000000000000000670000004900000021",
            INIT_37 => X"000000320000002200000025000000080000001e000000230000001500000000",
            INIT_38 => X"0000000a00000039000000180000001c00000000000000000000002500000025",
            INIT_39 => X"00000005000000000000000000000000000000000000000d0000001b00000000",
            INIT_3A => X"000000000000000a00000003000000310000000a000000120000000000000005",
            INIT_3B => X"000000190000001100000000000000150000000c000000140000000000000000",
            INIT_3C => X"0000003400000000000000000000000000000000000000000000002100000058",
            INIT_3D => X"000000170000001f000000170000000000000000000000000000001300000052",
            INIT_3E => X"000000000000004c00000017000000010000001e000000390000000000000015",
            INIT_3F => X"000000000000000e000000000000002800000046000000070000001e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE29;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE30 : if BRAM_NAME = "samplegold_layer0_instance30" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004e000000000000000d0000002b00000000000000250000001200000007",
            INIT_01 => X"000000000000000000000000000000000000000000000011000000400000002a",
            INIT_02 => X"0000001e0000003b000000190000000000000048000000420000000000000000",
            INIT_03 => X"0000001400000025000000000000000000000000000000370000000000000000",
            INIT_04 => X"00000000000000000000000c0000002300000000000000000000000100000000",
            INIT_05 => X"0000001300000002000000000000000000000010000000000000001b00000010",
            INIT_06 => X"0000001f0000003a000000190000001000000000000000000000002a00000000",
            INIT_07 => X"0000000000000000000000230000001d00000000000000000000002e00000000",
            INIT_08 => X"0000000900000000000000000000001700000000000000110000003200000000",
            INIT_09 => X"00000000000000000000000000000000000000120000000a0000000000000000",
            INIT_0A => X"0000000000000000000000010000000a00000001000000250000000500000000",
            INIT_0B => X"0000000b00000015000000050000000d00000013000000000000000a00000016",
            INIT_0C => X"0000000b000000110000000000000000000000000000000e0000000300000002",
            INIT_0D => X"000000010000000000000000000000260000005700000095000000370000003d",
            INIT_0E => X"0000000000000011000000000000000600000014000000010000000000000000",
            INIT_0F => X"00000000000000000000000d000000140000003b000000130000000000000000",
            INIT_10 => X"0000000000000000000000000000000900000000000000000000000200000000",
            INIT_11 => X"0000002d00000019000000000000002100000036000000010000000000000000",
            INIT_12 => X"0000001900000000000000000000001800000000000000000000000100000000",
            INIT_13 => X"000000000000000000000004000000330000003b000000000000000000000000",
            INIT_14 => X"000000070000000c0000000f0000004f0000002e0000003e0000000000000000",
            INIT_15 => X"0000001e00000008000000180000000000000010000000000000001100000000",
            INIT_16 => X"000000000000000700000014000000020000000d000000020000004c00000000",
            INIT_17 => X"0000000000000019000000090000000d00000003000000030000000200000015",
            INIT_18 => X"000000100000000300000003000000070000001f000000110000000500000038",
            INIT_19 => X"0000003200000000000000000000002500000000000000190000000600000000",
            INIT_1A => X"00000009000000010000000f00000022000000000000000b000000160000000a",
            INIT_1B => X"0000000d0000001f000000150000000c000000060000000a0000000c00000027",
            INIT_1C => X"0000002e00000011000000000000002600000017000000000000000e00000030",
            INIT_1D => X"000000310000000a000000250000000700000024000000150000000b00000002",
            INIT_1E => X"00000009000000330000002e000000180000001100000000000000000000001b",
            INIT_1F => X"000000180000003c000000000000002f000000150000002b0000002700000023",
            INIT_20 => X"000000440000004600000046000000460000003e000000150000000000000000",
            INIT_21 => X"000000000000001100000026000000060000002d0000003c000000350000003f",
            INIT_22 => X"0000004c00000043000000520000003e00000053000000310000001500000009",
            INIT_23 => X"000000090000000b000000010000002a000000140000004c0000002d00000053",
            INIT_24 => X"0000005000000051000000520000004000000041000000380000002800000002",
            INIT_25 => X"0000000b0000001b0000000a00000012000000140000001b0000004400000047",
            INIT_26 => X"0000004f000000450000004c000000470000003f00000032000000250000000f",
            INIT_27 => X"000000130000000000000019000000090000001e000000000000001d00000043",
            INIT_28 => X"000000420000004c000000430000004e00000045000000400000002200000017",
            INIT_29 => X"0000000c0000000c0000000e0000003a00000025000000000000000600000005",
            INIT_2A => X"00000019000000510000005700000043000000450000003d0000004e00000030",
            INIT_2B => X"0000002c0000000b000000250000003c0000002d000000090000002000000000",
            INIT_2C => X"0000000c000000090000005900000050000000470000003b000000200000005c",
            INIT_2D => X"0000001e0000002c0000002a0000003d00000024000000050000002400000026",
            INIT_2E => X"00000027000000000000000d000000460000005b000000420000004400000026",
            INIT_2F => X"000000450000002c000000300000002f000000220000000f0000001500000015",
            INIT_30 => X"00000000000000000000001e0000000200000028000000260000003d00000037",
            INIT_31 => X"00000000000000000000000a000000000000002d000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000019000000000000003800000000",
            INIT_33 => X"0000000000000000000000000000001b000000000000001c0000000000000000",
            INIT_34 => X"00000000000000000000000000000000000000000000001d0000000000000048",
            INIT_35 => X"0000003e00000004000000000000000000000000000000000000001d00000000",
            INIT_36 => X"0000000800000000000000000000002000000000000000000000000000000000",
            INIT_37 => X"00000000000000150000000f000000000000002b000000000000000000000008",
            INIT_38 => X"000000000000002500000000000000000000002b000000000000000000000000",
            INIT_39 => X"0000000000000000000000050000000000000000000000000000002a00000000",
            INIT_3A => X"0000000100000002000000090000000000000000000000320000000000000000",
            INIT_3B => X"000000000000000000000000000000200000000000000000000000000000000b",
            INIT_3C => X"0000000d0000000f0000000e00000000000000000000000b0000001800000000",
            INIT_3D => X"000000000000000000000000000000000000001500000016000000160000000e",
            INIT_3E => X"000000090000001b00000027000000030000000500000000000000000000000c",
            INIT_3F => X"0000000000000000000000000000000000000000000000270000001200000012",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE30;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE31 : if BRAM_NAME = "samplegold_layer0_instance31" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000160000000f0000001400000026000000000000001b0000000000000000",
            INIT_01 => X"000000000000000000000000000000000000000000000000000000150000000e",
            INIT_02 => X"000000140000000000000017000000170000000d000000370000000000000005",
            INIT_03 => X"0000000100000000000000170000000000000011000000000000000000000000",
            INIT_04 => X"0000000a0000000e000000050000000300000002000000470000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_06 => X"000000000000000d000000140000000000000009000000130000001c0000000a",
            INIT_07 => X"0000000f0000000000000000000000000000001c000000000000000000000009",
            INIT_08 => X"0000000f0000000000000000000000140000000c000000340000000000000001",
            INIT_09 => X"00000000000000000000000000000000000000240000001d0000000000000000",
            INIT_0A => X"00000000000000210000000000000000000000130000001a0000002500000000",
            INIT_0B => X"000000000000000000000000000000000000001c0000003f0000000000000000",
            INIT_0C => X"00000000000000360000000000000000000000000000000e0000001300000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000070000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"00000000000000000000000000000000000000090000000f0000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000023000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000900000007000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000200000000000000000000000400000000",
            INIT_2B => X"0000000000000000000000020000000000000003000000000000000000000000",
            INIT_2C => X"0000000d00000015000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000800000000000000000000000000000000",
            INIT_30 => X"0000000200000000000000000000000000000010000000000000000a00000000",
            INIT_31 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"000000000000000000000000000000000000000c000000140000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000001800000000",
            INIT_34 => X"0000000b00000010000000000000000000000000000000000000000900000000",
            INIT_35 => X"000000000000000a000000000000000100000015000000010000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000009",
            INIT_37 => X"0000000f0000000000000000000000160000000000000000000000000000000c",
            INIT_38 => X"0000000e000000060000000000000018000000040000000b0000000000000000",
            INIT_39 => X"00000000000000000000002d0000003800000000000000120000000000000000",
            INIT_3A => X"0000000900000000000000000000003b0000000000000000000000000000000e",
            INIT_3B => X"0000000000000005000000000000000000000005000000090000000000000003",
            INIT_3C => X"0000001800000002000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000200000005",
            INIT_3E => X"00000000000000090000000d0000001000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000390000002000000000000000050000001100000010",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE31;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE32 : if BRAM_NAME = "samplegold_layer0_instance32" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000001500000003000000360000004a000000150000000800000000",
            INIT_01 => X"0000000000000000000000260000002000000000000000000000000400000014",
            INIT_02 => X"0000003000000019000000070000001200000000000000000000000000000000",
            INIT_03 => X"00000000000000030000001e00000003000000000000000f0000000000000000",
            INIT_04 => X"0000000000000000000000140000004f000000330000000c0000000000000000",
            INIT_05 => X"000000300000000a000000240000003c00000023000000120000003a00000000",
            INIT_06 => X"00000030000000240000004e00000041000000500000004f000000470000002a",
            INIT_07 => X"000000240000002f000000090000001a00000043000000450000002a0000004b",
            INIT_08 => X"000000520000004d0000002d00000062000000450000004b0000003e0000004e",
            INIT_09 => X"0000004c0000003e0000002e00000009000000110000003a0000004900000046",
            INIT_0A => X"0000003c00000037000000700000005f00000085000000520000004b00000032",
            INIT_0B => X"000000340000002f000000280000005b0000003a000000080000002c00000045",
            INIT_0C => X"0000006f0000006c000000370000007200000079000000a5000000650000003b",
            INIT_0D => X"0000006b000000540000004e00000018000000370000005e0000003100000030",
            INIT_0E => X"000000470000009800000069000000310000005f000000880000008d0000006d",
            INIT_0F => X"0000004e000000530000005a000000570000004f0000003e0000005700000041",
            INIT_10 => X"000000550000008f0000007e00000052000000340000004f0000008f00000086",
            INIT_11 => X"000000700000004d0000004e0000005100000051000000460000003e00000047",
            INIT_12 => X"0000002d0000006a000000930000006c000000600000004a0000005d0000007c",
            INIT_13 => X"000000750000005c000000780000004c00000047000000520000005f00000053",
            INIT_14 => X"0000005200000065000000830000007d000000720000005f0000005600000047",
            INIT_15 => X"000000420000005d0000007d000000600000006b0000006e0000005c00000067",
            INIT_16 => X"000000710000006a000000840000006d0000006300000055000000670000006e",
            INIT_17 => X"00000062000000540000003e0000005100000067000000630000007500000079",
            INIT_18 => X"0000008200000088000000800000005a000000570000005d0000004a00000051",
            INIT_19 => X"000000640000006800000070000000550000004d00000062000000660000007a",
            INIT_1A => X"0000006e0000008600000086000000780000006b000000760000005c00000057",
            INIT_1B => X"0000009c000000b60000007d0000008500000059000000510000005f00000067",
            INIT_1C => X"00000077000000760000007d0000006d000000820000007e0000006900000072",
            INIT_1D => X"000000a70000009b00000037000000480000007c0000003c000000470000005c",
            INIT_1E => X"0000005e00000075000000750000004b00000066000000770000006b00000076",
            INIT_1F => X"000000b30000009f0000002b000000140000004f000000670000003b0000003b",
            INIT_20 => X"00000034000000600000006f0000007000000068000000790000007600000083",
            INIT_21 => X"000000000000001d00000000000000000000000000000000000000680000003a",
            INIT_22 => X"0000000000000029000000000000001200000006000000140000000000000000",
            INIT_23 => X"00000003000000060000001c0000000000000002000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_25 => X"0000001800000000000000000000001200000017000000000000000000000038",
            INIT_26 => X"0000000300000000000000000000000000000000000000000000004500000000",
            INIT_27 => X"0000000000000028000000240000000000000000000000000000001000000000",
            INIT_28 => X"000000000000000a0000003c0000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000001e00000000000000000000002400000000",
            INIT_2A => X"0000000000000000000000260000004200000000000000000000000200000006",
            INIT_2B => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000027000000000000001500000000",
            INIT_2D => X"0000000000000000000000000000000300000003000000000000000000000007",
            INIT_2E => X"00000000000000000000000000000000000000080000000c0000000000000001",
            INIT_2F => X"0000000000000000000000040000000000000000000000000000000000000035",
            INIT_30 => X"0000000000000022000000060000002000000000000000000000004f00000000",
            INIT_31 => X"0000002c00000023000000090000000000000001000000000000000000000000",
            INIT_32 => X"0000000000000028000000000000000000000021000000230000000900000000",
            INIT_33 => X"0000000000000000000000070000000200000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000c00000000000000000000000000000033",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000001900000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"000000010000004d00000000000000000000000c000000020000000000000000",
            INIT_38 => X"0000000000000008000000570000000700000000000000000000000000000000",
            INIT_39 => X"000000000000006d000000180000001800000017000000110000000000000000",
            INIT_3A => X"0000000000000005000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000038000000000000001a00000000000000000000004500000023",
            INIT_3C => X"0000000000000035000000130000002400000000000000000000000000000000",
            INIT_3D => X"000000000000001b000000190000000000000003000000000000000000000000",
            INIT_3E => X"000000000000003400000000000000110000000a00000018000000060000002e",
            INIT_3F => X"0000002900000000000000180000000600000001000000070000000e00000025",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE32;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE33 : if BRAM_NAME = "samplegold_layer0_instance33" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001e00000000000000420000000000000013000000000000002500000012",
            INIT_01 => X"0000001400000020000000000000001100000011000000120000000f00000001",
            INIT_02 => X"000000000000000c000000000000003c00000012000000000000001d00000009",
            INIT_03 => X"00000000000000000000001c0000000e00000002000000000000002b00000000",
            INIT_04 => X"000000000000000000000006000000000000002c000000190000000000000035",
            INIT_05 => X"000000000000002000000000000000000000002100000000000000000000003d",
            INIT_06 => X"0000004400000000000000000000000d0000000000000010000000000000000e",
            INIT_07 => X"0000000000000000000000040000000000000000000000180000000000000009",
            INIT_08 => X"000000280000002d000000000000000000000017000000000000001d00000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"000000060000001e000000280000000000000000000000160000000000000000",
            INIT_0B => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"000000140000000e00000012000000110000000c000000000000000d00000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000001c0000000f000000200000000a00000008000000100000000000000000",
            INIT_0F => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000001f000000030000000f0000001a000000000000001f0000000000000018",
            INIT_11 => X"000000180000000a000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000008000000120000000100000022000000000000000000000000",
            INIT_13 => X"0000001f0000000f000000150000000000000000000000000000000000000000",
            INIT_14 => X"0000001600000000000000000000002100000000000000000000000000000023",
            INIT_15 => X"0000003100000000000000100000001a00000000000000000000000000000000",
            INIT_16 => X"000000000000001700000000000000050000000000000000000000000000002e",
            INIT_17 => X"0000003900000000000000000000000d0000002b000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000025",
            INIT_19 => X"000000310000004a0000000a0000002600000031000000060000000000000000",
            INIT_1A => X"0000006a0000000b000000300000003a000000390000002b0000006200000000",
            INIT_1B => X"00000000000000300000001e0000001c00000020000000270000004500000000",
            INIT_1C => X"00000000000000840000000a00000041000000270000004c0000001d0000004d",
            INIT_1D => X"00000058000000000000001500000022000000220000001d0000002700000060",
            INIT_1E => X"00000035000000050000007b0000004700000000000000320000002f00000052",
            INIT_1F => X"0000002d00000075000000190000000f0000001800000070000000000000002c",
            INIT_20 => X"000000000000002e00000014000000760000006b000000000000007000000000",
            INIT_21 => X"000000600000000000000038000000640000000a000000000000008800000008",
            INIT_22 => X"000000000000000000000029000000250000003f000000440000005e00000042",
            INIT_23 => X"0000002d0000005a000000030000002c00000067000000000000002d00000083",
            INIT_24 => X"0000006300000000000000000000003200000014000000730000000c00000029",
            INIT_25 => X"00000024000000150000002900000018000000260000000e0000002000000042",
            INIT_26 => X"000000410000004f00000008000000000000004700000005000000330000001e",
            INIT_27 => X"000000220000002300000019000000220000003500000000000000260000002d",
            INIT_28 => X"000000240000001b000000440000002f000000000000002f000000050000002e",
            INIT_29 => X"0000002c000000090000001a00000025000000140000002d0000000b0000003b",
            INIT_2A => X"000000280000004a0000000c0000000e00000034000000000000000a00000000",
            INIT_2B => X"00000000000000100000001100000017000000130000002d000000220000002f",
            INIT_2C => X"000000260000003f000000460000000d0000004f00000000000000430000001d",
            INIT_2D => X"00000020000000070000000d0000001800000002000000120000001c0000005d",
            INIT_2E => X"000000490000004200000011000000510000000e000000620000003000000051",
            INIT_2F => X"000000280000003f00000003000000120000002f000000000000000f0000001f",
            INIT_30 => X"00000000000000310000004f00000026000000290000001f0000004e0000003f",
            INIT_31 => X"0000000c000000380000002700000001000000000000001b000000130000002a",
            INIT_32 => X"00000054000000120000003e0000003b00000020000000360000006f00000048",
            INIT_33 => X"00000029000000000000003a0000006300000000000000000000001e00000029",
            INIT_34 => X"0000002a000000190000003a000000320000002b000000330000007a00000078",
            INIT_35 => X"0000001700000015000000080000009e0000003600000002000000000000001b",
            INIT_36 => X"0000000000000000000000000000000000000000000000120000000000000000",
            INIT_37 => X"00000000000000000000000f0000000200000001000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000003400000003",
            INIT_3A => X"000000000000000100000000000000000000000000000000000000310000002a",
            INIT_3B => X"0000001b00000018000000000000000000000029000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000001f00000002000000010000000000000000",
            INIT_3D => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000140000001300000035",
            INIT_3F => X"000000030000000000000000000000180000001e000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE33;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE34 : if BRAM_NAME = "samplegold_layer0_instance34" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"00000000000000000000000000000000000000000000000d0000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"00000000000000000000000000000018000000420000002f0000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000007",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000006",
            INIT_11 => X"00000000000000000000000f0000002a0000001e000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"00000000000000000000000000000000000000000000001e0000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000001600000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"000000000000000000000000000000000000000000000000000000000000001e",
            INIT_18 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000100000000000000000000001a00000000",
            INIT_1A => X"000000000000000d000000000000000500000000000000000000000000000004",
            INIT_1B => X"000000000000000200000000000000000000000000000000000000000000000e",
            INIT_1C => X"0000000d00000000000000170000000000000003000000070000000700000009",
            INIT_1D => X"0000001a0000000c000000170000001300000002000000000000000000000000",
            INIT_1E => X"00000000000000000000000000000005000000170000000d000000100000000b",
            INIT_1F => X"000000200000001a000000120000000f00000017000000000000000000000000",
            INIT_20 => X"000000000000000000000000000000000000002a0000000c0000001e0000001e",
            INIT_21 => X"0000001f0000002a0000001c00000019000000180000000c0000000000000000",
            INIT_22 => X"00000000000000000000000000000000000000030000001a0000002300000016",
            INIT_23 => X"000000160000003200000021000000210000001f000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000001600000023",
            INIT_25 => X"0000001c0000001d000000230000002500000030000000040000000000000000",
            INIT_26 => X"00000000000000000000000e0000001c00000000000000000000000000000013",
            INIT_27 => X"0000001b00000024000000280000001d000000220000002a0000001d00000000",
            INIT_28 => X"00000000000000000000000f0000001400000000000000000000000000000000",
            INIT_29 => X"000000000000001c00000023000000270000001c000000000000002b0000001a",
            INIT_2A => X"00000000000000000000001a0000000800000000000000000000000000000000",
            INIT_2B => X"00000000000000000000000c000000250000001a000000230000000000000000",
            INIT_2C => X"00000007000000090000001c0000000d00000000000000000000000000000000",
            INIT_2D => X"0000002b00000000000000000000000000000000000000160000001300000000",
            INIT_2E => X"0000003a000000180000003700000003000000540000002c0000002c00000034",
            INIT_2F => X"00000036000000260000001d0000000e0000007a00000000000000460000001f",
            INIT_30 => X"0000002c00000031000000130000001f0000001a000000510000002900000040",
            INIT_31 => X"00000024000000120000003400000040000000190000005d0000000000000046",
            INIT_32 => X"0000000700000051000000110000004d000000310000000a000000400000002e",
            INIT_33 => X"0000002c000000460000000300000041000000340000002f0000004600000000",
            INIT_34 => X"0000001b000000200000002500000009000000400000005e0000002e00000018",
            INIT_35 => X"00000000000000450000004800000000000000450000005e000000260000002c",
            INIT_36 => X"000000340000001d000000470000002a00000040000000020000006300000036",
            INIT_37 => X"00000017000000310000004f0000001700000000000000480000007300000023",
            INIT_38 => X"000000150000004b00000007000000300000002e000000370000001200000018",
            INIT_39 => X"0000000e0000000d0000002a000000290000000b000000100000003f00000078",
            INIT_3A => X"0000005f000000230000002b0000001500000000000000030000000f0000001e",
            INIT_3B => X"000000060000000000000037000000000000001e0000001a0000000d00000033",
            INIT_3C => X"00000018000000620000001d00000030000000000000001a000000110000000a",
            INIT_3D => X"0000000e0000000000000006000000010000000a0000001d0000002a0000002d",
            INIT_3E => X"000000280000002d0000003b00000028000000150000000f0000000900000001",
            INIT_3F => X"0000000f00000003000000000000000000000000000000150000001100000039",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE34;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE35 : if BRAM_NAME = "samplegold_layer0_instance35" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000044000000000000004c0000000a00000025000000290000001600000006",
            INIT_01 => X"00000000000000130000000200000009000000000000001e0000003600000012",
            INIT_02 => X"000000330000006500000029000000030000003100000014000000230000000a",
            INIT_03 => X"0000001100000000000000130000000000000000000000000000001400000030",
            INIT_04 => X"0000004d0000005c0000002f000000000000002000000035000000120000002a",
            INIT_05 => X"0000002e000000160000000700000000000000000000002b000000140000000c",
            INIT_06 => X"00000050000000610000001a0000000000000025000000450000004300000016",
            INIT_07 => X"0000000f00000043000000250000000000000000000000160000002a00000036",
            INIT_08 => X"0000005c000000510000001a000000000000001800000037000000550000000d",
            INIT_09 => X"0000000f000000310000003b000000070000000a000000010000003500000046",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000017",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000001",
            INIT_0C => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000100000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000100000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000018000000000000000000000002000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"000000000000000000000000000000000000000000000000000000000000000b",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_1A => X"00000000000000000000000000000000000000100000001f0000000000000000",
            INIT_1B => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000050000000000000000000000000000000000000009",
            INIT_1D => X"0000000000000018000000000000000d00000007000000000000003500000000",
            INIT_1E => X"0000000000000000000000000000001000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000500000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000001b00000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE35;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE36 : if BRAM_NAME = "samplegold_layer0_instance36" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_03 => X"0000000f00000008000000000000000200000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000500000001000000080000000600000006000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"00000000000000050000000300000009000000040000000e0000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000400000000000000080000000c00000000000000000000000000000000",
            INIT_0A => X"0000000500000000000000070000000000000000000000000000000000000000",
            INIT_0B => X"0000000b00000000000000150000000300000000000000020000000000000000",
            INIT_0C => X"00000000000000080000000000000003000000000000000a0000000000000000",
            INIT_0D => X"0000000000000000000000060000002700000007000000000000000400000000",
            INIT_0E => X"0000000000000000000000130000001b00000000000000000000000900000006",
            INIT_0F => X"0000000e00000001000000000000002000000002000000040000000300000005",
            INIT_10 => X"000000020000000000000000000000040000000b000000100000000600000003",
            INIT_11 => X"0000000800000003000000000000000c0000001c0000000b000000000000000a",
            INIT_12 => X"0000001600000011000000000000000000000000000000000000000000000000",
            INIT_13 => X"00000000000000090000000f000000000000000c000000250000000100000000",
            INIT_14 => X"00000000000000200000000c000000030000000200000000000000000000000f",
            INIT_15 => X"0000001100000000000000010000000c00000000000000030000001900000008",
            INIT_16 => X"0000000300000000000000210000000c00000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000120000000f00000000000000050000000300000014",
            INIT_18 => X"0000000e0000000f000000000000001100000007000000000000000000000000",
            INIT_19 => X"0000000100000001000000040000000f0000000000000000000000020000000f",
            INIT_1A => X"00000002000000130000000a00000015000000000000000b0000000300000000",
            INIT_1B => X"00000007000000080000000b00000001000000160000000c0000000000000007",
            INIT_1C => X"000000130000000a0000001a0000000d000000000000000f000000060000000f",
            INIT_1D => X"0000000c0000000c0000000b0000000300000003000000090000000f0000000a",
            INIT_1E => X"000000120000000a00000010000000000000002c0000000f0000000000000008",
            INIT_1F => X"00000001000000100000000b0000000900000033000000000000001100000009",
            INIT_20 => X"0000000a00000007000000090000000300000026000000140000002b00000000",
            INIT_21 => X"0000001f0000000b0000000d0000000000000012000000260000000200000014",
            INIT_22 => X"000000150000000c000000070000000600000006000000050000003a0000000c",
            INIT_23 => X"0000000f0000000f000000120000001c00000000000000260000000c00000000",
            INIT_24 => X"000000110000001a0000000b00000011000000000000000d0000000a00000028",
            INIT_25 => X"0000000f0000000c00000000000000110000002f0000000a0000000e00000002",
            INIT_26 => X"000000280000001000000018000000130000000b000000030000000e00000005",
            INIT_27 => X"00000013000000000000000e00000011000000010000005c0000000b00000000",
            INIT_28 => X"000000000000003f000000360000004b00000000000000160000001300000000",
            INIT_29 => X"0000002b0000000000000000000000040000000b00000000000000450000002a",
            INIT_2A => X"0000004f00000011000000000000002f0000002f000000190000000000000028",
            INIT_2B => X"000000130000003400000000000000240000000e000000030000000000000032",
            INIT_2C => X"000000410000006c0000002f0000002d00000015000000200000003100000000",
            INIT_2D => X"0000001800000039000000290000000000000027000000380000000000000000",
            INIT_2E => X"00000000000000220000006b0000003e00000027000000250000005c00000000",
            INIT_2F => X"0000001100000000000000a70000002d000000000000002c0000007900000000",
            INIT_30 => X"000000000000000000000020000000110000001e000000550000000000000062",
            INIT_31 => X"0000001600000001000000000000008f000000370000000000000037000000a5",
            INIT_32 => X"0000009000000000000000000000000700000014000000210000005100000000",
            INIT_33 => X"00000039000000070000000500000029000000340000000e0000001000000023",
            INIT_34 => X"0000000d00000018000000000000000000000000000000140000000900000018",
            INIT_35 => X"0000002400000032000000040000002e00000042000000030000001600000016",
            INIT_36 => X"000000000000002d000000000000000000000000000000000000001100000010",
            INIT_37 => X"0000001e0000001000000037000000000000000700000036000000030000003e",
            INIT_38 => X"00000023000000090000000f0000002400000003000000120000000100000011",
            INIT_39 => X"0000000a000000150000001b000000200000001c0000001b000000180000000e",
            INIT_3A => X"00000019000000050000005f0000001800000000000000270000001b00000008",
            INIT_3B => X"0000000e0000000000000000000000030000000b000000090000000c0000000b",
            INIT_3C => X"000000140000001000000008000000000000001100000006000000140000000b",
            INIT_3D => X"000000080000000000000000000000090000001c00000018000000190000001c",
            INIT_3E => X"0000000a0000001000000006000000110000000000000005000000030000000b",
            INIT_3F => X"0000000000000000000000220000004800000049000000180000000800000013",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE36;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE37 : if BRAM_NAME = "samplegold_layer0_instance37" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000001000000030000000e00000000000000000000000000000010",
            INIT_01 => X"000000010000000b000000000000001400000011000000000000000000000007",
            INIT_02 => X"0000002e000000030000000f0000000a000000040000000b0000000c00000000",
            INIT_03 => X"000000000000000000000000000000000000000000000002000000000000000d",
            INIT_04 => X"00000000000000000000002a0000001f000000000000000d0000002000000009",
            INIT_05 => X"000000000000002e000000000000000000000000000000000000000000000006",
            INIT_06 => X"0000003a00000066000000400000000000000010000000190000000400000000",
            INIT_07 => X"0000000000000005000000090000000000000006000000030000000000000001",
            INIT_08 => X"0000002700000008000000010000000f00000025000000120000001b00000000",
            INIT_09 => X"00000000000000110000001e00000019000000160000002f0000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000030000001200000003000000160000000b00000000",
            INIT_0C => X"000000030000002a0000000f00000000000000180000003c0000000000000000",
            INIT_0D => X"0000000000000014000000000000000000000000000000100000002800000015",
            INIT_0E => X"000000000000001a000000000000000000000000000000000000000000000000",
            INIT_0F => X"000000450000004f0000002d00000048000000000000001a0000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"000000370000000f0000000000000027000000000000000b0000000000000015",
            INIT_12 => X"00000001000000000000000000000015000000270000002f000000360000003a",
            INIT_13 => X"000000210000000c0000000b0000000f00000000000000000000000000000000",
            INIT_14 => X"0000003300000003000000000000003b000000440000004f0000003400000032",
            INIT_15 => X"000000000000000000000000000000050000001a000000250000002300000007",
            INIT_16 => X"0000008900000078000000740000002000000011000000170000001100000016",
            INIT_17 => X"0000004b0000004a00000069000000740000008c000000930000008f0000008b",
            INIT_18 => X"0000008d0000008a00000089000000800000004f000000520000004b00000051",
            INIT_19 => X"0000005400000045000000590000008a00000095000000a10000009a00000096",
            INIT_1A => X"00000096000000950000008f0000007500000085000000530000006200000056",
            INIT_1B => X"000000660000006c000000610000006e000000910000009d000000a6000000a0",
            INIT_1C => X"000000a60000009a000000900000008d00000074000000640000005d0000005e",
            INIT_1D => X"000000600000006000000087000000870000008e0000009000000099000000a5",
            INIT_1E => X"000000800000009d0000009d000000920000008b000000770000005e00000060",
            INIT_1F => X"0000005c0000005b000000510000007f00000083000000880000008e0000007d",
            INIT_20 => X"0000006600000066000000610000009300000091000000890000007b00000029",
            INIT_21 => X"0000004a0000005900000055000000430000005a00000078000000620000005e",
            INIT_22 => X"0000004e000000540000006300000076000000680000007b0000007a0000005a",
            INIT_23 => X"0000004b00000066000000590000005100000036000000460000006400000056",
            INIT_24 => X"00000052000000540000005f00000086000000730000005b0000006700000077",
            INIT_25 => X"0000006d0000004d0000007d000000640000004700000024000000450000006e",
            INIT_26 => X"000000560000006a0000006600000071000000990000005b0000005c00000076",
            INIT_27 => X"0000008a00000056000000560000008200000067000000420000002600000033",
            INIT_28 => X"000000410000003600000045000000890000005c000000770000005c00000022",
            INIT_29 => X"0000003c000000640000005c0000005e0000008900000063000000330000002f",
            INIT_2A => X"000000430000002f0000003200000041000000680000006e0000005100000045",
            INIT_2B => X"0000004f00000065000000670000005000000077000000780000005700000039",
            INIT_2C => X"000000570000002c000000210000001a00000023000000390000005d0000005c",
            INIT_2D => X"000000670000006d0000007f000000580000007500000076000000840000003f",
            INIT_2E => X"000000550000003c000000370000001a000000260000002d000000450000006e",
            INIT_2F => X"00000082000000710000006600000068000000690000007e0000006700000083",
            INIT_30 => X"000000700000004f0000005d0000005600000052000000500000005a00000060",
            INIT_31 => X"0000007900000079000000870000007f0000006d000000760000007d0000007e",
            INIT_32 => X"000000330000000400000062000000770000007a000000760000007600000073",
            INIT_33 => X"0000002300000003000000330000002c0000003200000029000000390000002a",
            INIT_34 => X"00000031000000140000002600000013000000390000002c000000200000002b",
            INIT_35 => X"00000038000000170000000e0000003b0000002d00000033000000340000002e",
            INIT_36 => X"000000340000002e0000002d000000030000002c000000200000003500000034",
            INIT_37 => X"0000002100000039000000050000003100000041000000280000003000000033",
            INIT_38 => X"0000002f000000390000002b00000027000000080000002d0000003300000035",
            INIT_39 => X"0000002a000000100000002700000033000000400000002f0000003200000035",
            INIT_3A => X"00000029000000330000002d0000002b0000003300000023000000330000003d",
            INIT_3B => X"0000002c0000003600000000000000370000004e0000001d0000002f00000029",
            INIT_3C => X"000000000000003d000000220000002a0000003a000000180000007f0000002f",
            INIT_3D => X"000000360000002b0000003600000000000000200000003d000000040000001c",
            INIT_3E => X"000000000000000800000021000000340000001200000015000000480000006b",
            INIT_3F => X"000000150000002c0000002d0000002c00000003000000000000001e0000002c",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE37;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE38 : if BRAM_NAME = "samplegold_layer0_instance38" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001000000026000000220000001100000034000000230000001200000071",
            INIT_01 => X"0000005c0000002d000000080000003400000033000000000000000000000008",
            INIT_02 => X"0000001500000022000000240000000700000034000000230000000a0000001c",
            INIT_03 => X"000000150000006b000000200000000000000047000000500000000900000000",
            INIT_04 => X"0000001d0000000e000000000000004900000000000000310000006800000000",
            INIT_05 => X"000000000000000b000000560000002500000000000000600000004a00000019",
            INIT_06 => X"0000002d0000001d0000001300000008000000510000002c0000002d0000002d",
            INIT_07 => X"0000000e0000000c000000250000003d0000002f00000000000000730000003d",
            INIT_08 => X"00000049000000260000000d0000001800000009000000000000003100000033",
            INIT_09 => X"000000190000000d000000380000002b0000003800000044000000200000004c",
            INIT_0A => X"00000029000000330000001c0000000b0000000d0000000b0000001700000044",
            INIT_0B => X"0000004a0000003500000011000000340000001d000000570000002b0000003e",
            INIT_0C => X"00000016000000320000001d0000003000000023000000230000002e00000020",
            INIT_0D => X"0000003600000034000000350000002a0000004000000032000000440000003c",
            INIT_0E => X"0000002300000040000000200000002f0000003f00000041000000370000002f",
            INIT_0F => X"0000003000000036000000430000003c000000380000002f0000003600000001",
            INIT_10 => X"0000002200000014000000280000002100000026000000290000002c0000002a",
            INIT_11 => X"0000002c00000048000000410000003f00000033000000360000002f00000032",
            INIT_12 => X"00000027000000190000001a0000002d0000002f0000002c000000300000002c",
            INIT_13 => X"000000180000001d0000003e0000003d0000003e0000003a0000002e00000032",
            INIT_14 => X"0000002c0000002b000000160000001a0000002b00000039000000360000002d",
            INIT_15 => X"00000036000000390000003d0000003a0000004000000042000000430000002b",
            INIT_16 => X"0000002c0000002e00000021000000180000002300000030000000310000003c",
            INIT_17 => X"0000002a0000002f00000032000000400000002a0000001a0000002600000038",
            INIT_18 => X"0000000d00000031000000220000001500000022000000230000003000000031",
            INIT_19 => X"0000002f000000240000003b0000002c000000230000002c0000001400000000",
            INIT_1A => X"0000001e000000000000000e000000160000000f00000021000000000000002e",
            INIT_1B => X"0000002e0000002800000019000000280000001e000000000000000000000006",
            INIT_1C => X"0000000400000011000000000000000000000019000000120000001200000030",
            INIT_1D => X"000000380000002000000011000000190000001e000000050000000000000000",
            INIT_1E => X"00000030000000370000001b000000200000000600000017000000030000000f",
            INIT_1F => X"0000001a00000045000000170000000f00000014000000380000005100000037",
            INIT_20 => X"0000003e0000002f00000013000000380000000c000000240000002500000000",
            INIT_21 => X"0000000d0000002a0000003600000000000000090000001b0000001d0000001b",
            INIT_22 => X"0000002b00000032000000580000004b000000480000003f0000001c00000041",
            INIT_23 => X"000000000000001f0000002a000000470000000b000000180000001d00000030",
            INIT_24 => X"0000001e00000020000000250000002f0000003f0000001c0000001a00000028",
            INIT_25 => X"0000000e00000027000000210000003f000000360000002a0000002b0000002c",
            INIT_26 => X"000000170000000f00000013000000150000001b0000002e0000003500000034",
            INIT_27 => X"00000029000000350000003000000036000000390000003b0000001f00000031",
            INIT_28 => X"000000180000001800000013000000200000001f0000002a0000004100000030",
            INIT_29 => X"0000003e0000002d000000230000002d0000003b000000270000003e00000032",
            INIT_2A => X"00000028000000340000003200000034000000360000003e0000003d00000043",
            INIT_2B => X"00000004000000170000000d0000000f00000011000000180000000000000000",
            INIT_2C => X"00000011000000120000000400000000000000000000000a0000001300000012",
            INIT_2D => X"000000020000000a000000100000000a0000000d000000060000000b00000019",
            INIT_2E => X"00000008000000170000000c0000000d000000140000001f0000000b00000001",
            INIT_2F => X"0000000000000015000000150000000b000000100000000d0000001300000007",
            INIT_30 => X"000000120000000f000000120000000b0000001e000000170000000800000000",
            INIT_31 => X"0000000000000019000000240000001e000000260000001d0000001700000011",
            INIT_32 => X"000000050000000d00000007000000220000000f000000010000000f00000009",
            INIT_33 => X"0000002b0000001f000000250000000b00000000000000100000001e00000011",
            INIT_34 => X"0000001c00000012000000000000000000000004000000130000001e00000015",
            INIT_35 => X"00000015000000260000001a0000000d000000370000004f0000000100000000",
            INIT_36 => X"00000007000000000000000d0000001700000023000000000000001000000013",
            INIT_37 => X"00000002000000000000000c0000001000000000000000000000000000000021",
            INIT_38 => X"000000090000001000000000000000200000001b000000070000000300000014",
            INIT_39 => X"0000000a00000000000000070000001f00000009000000070000001200000010",
            INIT_3A => X"00000047000000300000000c00000018000000220000000c0000000000000019",
            INIT_3B => X"0000000d0000000b000000000000000000000015000000670000006300000049",
            INIT_3C => X"0000000d0000000c000000420000002d00000066000000250000001100000000",
            INIT_3D => X"000000180000001c00000000000000000000000600000000000000000000001b",
            INIT_3E => X"0000001a0000006200000030000000360000002a000000000000003000000023",
            INIT_3F => X"00000017000000070000002f000000210000001a000000000000001f00000020",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE38;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE39 : if BRAM_NAME = "samplegold_layer0_instance39" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000b00000004000000000000001100000000000000000000000100000000",
            INIT_01 => X"0000003e0000000000000018000000140000002c000000210000000a00000006",
            INIT_02 => X"0000000000000000000000000000000000000000000000030000002300000023",
            INIT_03 => X"0000002d0000000900000030000000230000001f000000030000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000170000001000000000",
            INIT_05 => X"0000000a000000000000000d00000018000000000000000a0000002100000000",
            INIT_06 => X"0000000f0000000e000000100000000e00000015000000190000003100000021",
            INIT_07 => X"0000000200000006000000110000001200000015000000030000001a00000003",
            INIT_08 => X"0000000a00000007000000000000000000000005000000030000000b00000000",
            INIT_09 => X"0000000000000000000000100000001700000019000000140000003500000038",
            INIT_0A => X"0000003c00000008000000080000000b0000000a000000060000000000000000",
            INIT_0B => X"0000000d000000080000000f0000001900000024000000220000001e0000003b",
            INIT_0C => X"000000360000003e000000080000000d00000004000000000000000000000000",
            INIT_0D => X"0000001b0000001a0000000d0000001d0000001a0000002c000000270000002b",
            INIT_0E => X"0000002d00000036000000330000000e00000002000000040000000800000008",
            INIT_0F => X"0000001f0000001e000000150000002900000033000000270000002c00000026",
            INIT_10 => X"000000380000003a0000002d00000028000000110000000e0000000c0000001f",
            INIT_11 => X"0000001600000023000000260000003700000056000000510000004f0000002c",
            INIT_12 => X"0000003900000049000000570000004d000000070000000e0000000500000009",
            INIT_13 => X"00000000000000070000002a0000003b0000003100000038000000580000005a",
            INIT_14 => X"000000690000005f0000004c0000005800000035000000070000000a00000002",
            INIT_15 => X"00000018000000070000000d0000003c000000690000006e0000006500000038",
            INIT_16 => X"0000004f0000006000000073000000370000005f000000300000001200000003",
            INIT_17 => X"0000001d00000034000000000000000000000041000000550000005a0000004e",
            INIT_18 => X"0000002f00000048000000530000005f0000002f000000780000003600000013",
            INIT_19 => X"000000200000003f000000410000000000000000000000000000000300000008",
            INIT_1A => X"0000002b000000260000002600000024000000000000002e0000006b0000002f",
            INIT_1B => X"0000001d00000025000000640000003e00000000000000090000000700000000",
            INIT_1C => X"000000000000000000000000000000000000000000000000000000260000004a",
            INIT_1D => X"0000002200000029000000150000005500000011000000070000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000014000000170000002700000052",
            INIT_1F => X"000000110000002b000000280000001f0000001c000000000000000000000000",
            INIT_20 => X"00000000000000000000000000000009000000110000001d0000001100000030",
            INIT_21 => X"00000016000000130000001e000000150000001e000000150000000000000000",
            INIT_22 => X"0000001200000015000000090000000c0000000f0000001f000000160000001a",
            INIT_23 => X"000000000000000000000000000000000000000000000000000000070000000c",
            INIT_24 => X"0000000000000000000000000000000000000001000000070000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000130000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000019",
            INIT_28 => X"0000000100000000000000000000000300000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"00000000000000060000000000000000000000000000000b0000000000000000",
            INIT_2B => X"0000000000000016000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_2D => X"0000001c00000000000000020000003500000004000000000000001000000000",
            INIT_2E => X"000000000000000000000000000000000000000000000000000000000000002c",
            INIT_2F => X"0000000d00000018000000000000000000000000000000000000001300000000",
            INIT_30 => X"0000000000000001000000000000000000000004000000040000000000000000",
            INIT_31 => X"0000000000000017000000070000000000000000000000000000000000000000",
            INIT_32 => X"00000000000000030000002f0000000000000000000000000000001b00000000",
            INIT_33 => X"0000000000000000000000120000005e0000005a000000210000003900000030",
            INIT_34 => X"0000001c0000000f00000000000000570000000000000000000000000000001d",
            INIT_35 => X"0000000d00000000000000000000000000000000000000180000002f00000000",
            INIT_36 => X"0000003f00000021000000590000001400000026000000170000000000000001",
            INIT_37 => X"0000000000000000000000000000000000000000000000210000002100000035",
            INIT_38 => X"000000210000001c000000000000000000000000000000000000000000000000",
            INIT_39 => X"00000000000000000000000000000030000000000000001f0000000a0000000c",
            INIT_3A => X"0000000000000000000000000000000000000002000000000000000000000012",
            INIT_3B => X"0000000a00000000000000100000002700000000000000000000000000000000",
            INIT_3C => X"000000000000000000000000000000000000000000000000000000030000000c",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000020000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE39;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE40 : if BRAM_NAME = "samplegold_layer0_instance40" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"000000000000001e000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000220000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000100000000000000000000000000000004",
            INIT_0F => X"0000001a00000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"000000000000002000000000000000000000000c000000000000000000000003",
            INIT_11 => X"000000100000000d000000000000000000000000000000000000000000000000",
            INIT_12 => X"00000000000000190000001b0000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000021000000000000000000000008000000000000000000000004",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"00000000000000000000000a0000000f00000019000000090000000900000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"000000000000000000000006000000000000000e000000060000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000002200000015000000480000000000000000000000000000000000000000",
            INIT_1C => X"000000100000001600000015000000000000001e0000000b0000001a00000014",
            INIT_1D => X"0000001d0000001d00000014000000110000001f000000000000002a00000016",
            INIT_1E => X"00000020000000130000002500000005000000000000001c000000100000001b",
            INIT_1F => X"000000150000001e0000001c000000200000002c000000000000000d0000000d",
            INIT_20 => X"0000000f000000190000000a00000034000000000000000e000000200000000d",
            INIT_21 => X"0000000a000000150000001c000000260000001a000000290000000000000017",
            INIT_22 => X"00000016000000200000000b000000000000000a000000100000001e00000011",
            INIT_23 => X"0000001d0000000c000000180000001f0000001f000000200000002b0000000e",
            INIT_24 => X"0000005900000017000000160000002600000000000000170000002600000004",
            INIT_25 => X"000000000000001000000007000000380000000c0000001b0000002f0000000c",
            INIT_26 => X"000000320000008600000020000000180000002a00000000000000050000002e",
            INIT_27 => X"0000002e0000003c000000000000000000000031000000230000001000000013",
            INIT_28 => X"0000000900000068000000060000001900000021000000240000000000000000",
            INIT_29 => X"0000000000000010000000160000002c00000014000000090000004100000011",
            INIT_2A => X"00000000000000110000005c0000000300000000000000360000002700000000",
            INIT_2B => X"0000000000000000000000000000001400000014000000000000001700000047",
            INIT_2C => X"0000005200000000000000180000005a00000000000000000000004e00000049",
            INIT_2D => X"0000004300000015000000050000000000000000000000420000000000000034",
            INIT_2E => X"0000000e0000003e000000000000001000000038000000000000000000000069",
            INIT_2F => X"0000006700000035000000140000001200000000000000000000003100000000",
            INIT_30 => X"0000002a0000001b000000000000000000000013000000250000000000000000",
            INIT_31 => X"0000001100000033000000310000002b0000000e0000000b0000000000000000",
            INIT_32 => X"00000000000000170000000c000000000000001b000000180000000900000019",
            INIT_33 => X"000000080000003c0000000e0000003c000000270000000e0000000f00000001",
            INIT_34 => X"0000000c000000000000002b0000001d000000000000001c0000000000000021",
            INIT_35 => X"0000002e00000007000000030000002e000000160000002e000000110000000c",
            INIT_36 => X"000000050000000b0000000300000013000000180000000d0000001900000000",
            INIT_37 => X"000000000000001c000000000000001f000000020000000a0000001c0000001d",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"00000000000000000000001d0000001400000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE40;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE41 : if BRAM_NAME = "samplegold_layer0_instance41" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000002f00000006000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000c0000000a00000000000000000000000c000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000002c0000000e000000190000000000000000000000000000000000000000",
            INIT_0D => X"000000000000000000000000000000000000000000000000000000000000001e",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"000000000000000000000000000000260000001f000000200000001900000007",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"00000000000000000000000c0000001e00000025000000180000000800000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000002800000024000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000100000018000000220000002b00000035000000360000003400000031",
            INIT_15 => X"0000002e000000390000002e0000000a0000000d000000010000000a00000007",
            INIT_16 => X"00000001000000010000002a000000350000003d000000390000003a00000036",
            INIT_17 => X"00000038000000360000002b00000036000000090000001c000000170000000b",
            INIT_18 => X"0000001e00000018000000220000003700000033000000410000003f0000003c",
            INIT_19 => X"000000410000003600000036000000320000001f00000017000000140000001e",
            INIT_1A => X"00000012000000250000002e0000003700000035000000390000004300000045",
            INIT_1B => X"000000430000003c0000003c0000003900000029000000180000001700000011",
            INIT_1C => X"000000140000000b0000002e0000002d0000002e000000320000003400000031",
            INIT_1D => X"0000003900000025000000380000003f00000031000000340000000000000016",
            INIT_1E => X"000000130000000c000000000000000c0000002a000000200000002400000025",
            INIT_1F => X"0000002100000020000000420000001f00000039000000400000001d0000000d",
            INIT_20 => X"00000025000000110000000a000000000000000000000022000000280000001d",
            INIT_21 => X"000000300000003600000041000000380000002d000000270000003a00000013",
            INIT_22 => X"000000210000002e000000160000001000000000000000030000002e0000002e",
            INIT_23 => X"000000240000002800000033000000450000001b000000380000002b00000034",
            INIT_24 => X"0000002e0000001a000000350000001e0000001500000000000000000000000f",
            INIT_25 => X"0000000000000000000000440000002d0000002e000000300000000000000040",
            INIT_26 => X"0000001b0000002e000000230000003c00000033000000120000000000000003",
            INIT_27 => X"0000000000000000000000000000000800000021000000000000000000000000",
            INIT_28 => X"000000210000002000000018000000360000002b0000002e0000000e00000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000210000001e0000000b",
            INIT_2A => X"000000320000002c000000140000002e000000320000002e000000120000000d",
            INIT_2B => X"0000000000000000000000000000000000000000000000030000002100000020",
            INIT_2C => X"0000002b000000210000001800000022000000340000001f0000003600000018",
            INIT_2D => X"000000140000001700000014000000160000000f000000180000001700000032",
            INIT_2E => X"0000002a0000003400000038000000290000002e0000002f0000003600000024",
            INIT_2F => X"0000002500000015000000290000002c0000002b000000280000001e0000002b",
            INIT_30 => X"00000023000000080000000c000000100000000d000000040000000d00000017",
            INIT_31 => X"00000018000000090000001100000000000000040000000f000000020000000c",
            INIT_32 => X"000000250000002100000005000000160000000b000000070000000a00000009",
            INIT_33 => X"0000000c000000000000002b000000030000000c000000000000000000000000",
            INIT_34 => X"00000002000000230000000a00000008000000120000000d0000000700000006",
            INIT_35 => X"000000000000000a0000000d0000001300000002000000000000000200000014",
            INIT_36 => X"000000280000001000000000000000010000000d0000000b000000040000000c",
            INIT_37 => X"000000050000000a000000080000000000000005000000000000000000000006",
            INIT_38 => X"000000000000003b000000000000000000000022000000050000000700000010",
            INIT_39 => X"0000000000000016000000110000000000000013000000000000000000000005",
            INIT_3A => X"00000007000000000000002c00000016000000000000000c000000110000002e",
            INIT_3B => X"0000000200000018000000000000000f00000011000000000000000000000000",
            INIT_3C => X"000000070000000700000007000000210000002d00000011000000060000000f",
            INIT_3D => X"00000000000000130000000c00000000000000040000000c0000000000000016",
            INIT_3E => X"0000000300000032000000000000000000000029000000380000000500000006",
            INIT_3F => X"0000000000000000000000250000000000000000000000280000000500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE41;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE42 : if BRAM_NAME = "samplegold_layer0_instance42" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000900000048000000000000000000000013000000250000000e",
            INIT_01 => X"0000001200000040000000000000001800000000000000000000006200000000",
            INIT_02 => X"00000006000000000000000a0000005b00000000000000000000001c0000000b",
            INIT_03 => X"000000100000001e000000120000000000000000000000010000001000000046",
            INIT_04 => X"0000001600000000000000000000000000000035000000000000000000000000",
            INIT_05 => X"000000130000001b00000017000000240000002800000007000000000000002a",
            INIT_06 => X"00000025000000000000000b0000000000000000000000000000000000000000",
            INIT_07 => X"0000000d0000000f000000240000001e0000001e0000001a000000000000000f",
            INIT_08 => X"0000000000000009000000000000000a00000000000000050000000300000000",
            INIT_09 => X"0000000c0000001200000005000000070000000e000000000000000700000000",
            INIT_0A => X"000000000000000000000000000000000000000000000000000000000000000b",
            INIT_0B => X"000000000000000f000000040000000000000000000000000000000300000000",
            INIT_0C => X"000000110000000b0000001000000016000000130000000c0000000b00000000",
            INIT_0D => X"0000001300000000000000000000000000000003000000060000001b00000000",
            INIT_0E => X"0000000000000003000000000000000100000004000000070000000800000009",
            INIT_0F => X"0000000900000000000000000000000000000004000000000000000400000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000003",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000c00000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000090000000000000000000000120000001e00000003",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000010",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000042000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"000000400000000000000000000000000000000000000004000000000000000d",
            INIT_20 => X"0000000000000000000000000000001e00000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000f00000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000001c00000000",
            INIT_25 => X"000000000000000000000002000000000000002b000000000000000000000000",
            INIT_26 => X"000000000000000000000000000000020000000000000000000000000000000d",
            INIT_27 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000007",
            INIT_34 => X"000000000000000000000000000000160000001f000000340000002500000008",
            INIT_35 => X"000000000000000000000000000000000000000000000000000000000000000e",
            INIT_36 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"000000070000001b000000070000000900000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"000000000000000b0000000a000000040000000b000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000140000000000000000",
            INIT_3B => X"0000000000000000000000000000000100000007000000020000000000000020",
            INIT_3C => X"00000000000000000000002b00000007000000010000003a000000350000003b",
            INIT_3D => X"0000000100000000000000000000000500000003000000000000000000000002",
            INIT_3E => X"0000000d000000030000000000000000000000050000000e0000002800000000",
            INIT_3F => X"0000000000000003000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE42;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE43 : if BRAM_NAME = "samplegold_layer0_instance43" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001d0000001a0000000000000000000000030000000e0000002700000000",
            INIT_01 => X"0000000000000011000000180000002e0000005900000058000000570000003f",
            INIT_02 => X"0000000000000000000000020000000000000000000000070000000d0000002c",
            INIT_03 => X"0000000100000007000000060000001900000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"000000040000000e000000000000000100000001000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000090000000100000000000000120000000000000000",
            INIT_0A => X"00000002000000050000000b0000000500000004000000020000000400000005",
            INIT_0B => X"00000008000000070000000000000000000000050000000a0000000000000004",
            INIT_0C => X"000000210000001800000007000000000000000a000000090000000600000007",
            INIT_0D => X"0000000500000008000000090000000000000000000000060000000a0000000a",
            INIT_0E => X"000000150000000000000005000000120000002c0000001f0000000900000004",
            INIT_0F => X"0000000500000005000000080000000800000002000000000000000500000000",
            INIT_10 => X"000000000000004c000000390000000000000000000000000000000000000020",
            INIT_11 => X"0000000300000019000000120000000600000008000000000000000100000008",
            INIT_12 => X"0000000000000000000000350000005a00000048000000190000000000000012",
            INIT_13 => X"00000001000000000000000d0000000e0000000c000000090000002100000006",
            INIT_14 => X"000000440000002c00000000000000190000002c0000002b000000480000002b",
            INIT_15 => X"00000039000000130000000000000017000000000000004b0000000c0000002c",
            INIT_16 => X"00000017000000240000003300000014000000130000001d0000003200000034",
            INIT_17 => X"0000002f00000052000000170000000000000006000000000000000c00000031",
            INIT_18 => X"0000001400000000000000130000001700000037000000180000000000000011",
            INIT_19 => X"000000000000003000000047000000290000000b000000000000001500000015",
            INIT_1A => X"00000013000000100000000000000000000000210000002d000000070000000b",
            INIT_1B => X"0000001900000000000000300000004a0000003400000031000000010000001a",
            INIT_1C => X"0000000a000000170000000f00000002000000000000001d000000110000000c",
            INIT_1D => X"0000000000000016000000000000000000000002000000060000000b00000000",
            INIT_1E => X"0000000f0000000e000000060000000c00000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000180000000200000006000000090000000a00000009",
            INIT_20 => X"0000000000000000000000000000000000000000000000010000000000000000",
            INIT_21 => X"0000003200000003000000030000000d00000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000100000000000000000000000a00000000",
            INIT_23 => X"0000000000000026000000220000000000000000000000000000000100000000",
            INIT_24 => X"00000000000000000000000000000006000000030000000e0000000600000009",
            INIT_25 => X"00000015000000000000000d0000003c0000000f000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_27 => X"0000000000000009000000070000000200000000000000520000000000000000",
            INIT_28 => X"0000000000000000000000030000000300000000000000040000000000000000",
            INIT_29 => X"0000000100000000000000030000000a00000019000000040000003f00000027",
            INIT_2A => X"0000006100000053000000450000000a00000000000000000000000400000004",
            INIT_2B => X"0000000f00000004000000000000000a0000002f00000000000000a400000038",
            INIT_2C => X"00000000000000000000002000000044000000490000001b0000000000000000",
            INIT_2D => X"0000001a000000000000000700000001000000150000001300000024000000fb",
            INIT_2E => X"000000fd0000004e0000000000000000000000000000002f000000060000003a",
            INIT_2F => X"0000005c000000130000001d000000000000000700000000000000000000006c",
            INIT_30 => X"00000000000000ad000000960000005700000057000000000000000000000000",
            INIT_31 => X"000000000000005000000009000000b700000000000000000000001e00000000",
            INIT_32 => X"0000004c0000002f0000007a00000041000000980000004c0000003400000000",
            INIT_33 => X"00000000000000000000002400000040000000a4000000360000000000000074",
            INIT_34 => X"00000092000000800000007f000000000000000000000071000000c200000041",
            INIT_35 => X"00000051000000000000000000000000000000640000003e0000001000000000",
            INIT_36 => X"0000000000000013000000b40000002d000000000000002c0000000d0000010c",
            INIT_37 => X"000000f500000048000000000000000b000000000000004a000000220000000e",
            INIT_38 => X"0000000f00000001000000000000008f00000000000000110000004e00000000",
            INIT_39 => X"00000000000000900000004e000000420000003800000015000000410000003b",
            INIT_3A => X"0000000d0000001b0000000e0000000100000022000000050000004100000045",
            INIT_3B => X"00000041000000000000001600000016000000140000000f0000000f00000027",
            INIT_3C => X"0000000000000000000000100000003a00000000000000050000000700000034",
            INIT_3D => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000500000000000000070000000000000000",
            INIT_3F => X"000000000000001e0000000c0000000800000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE43;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE44 : if BRAM_NAME = "samplegold_layer0_instance44" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000200000000000000000000000000000000000000000000000e0000000d",
            INIT_01 => X"000000270000001a000000000000003200000011000000110000000b00000007",
            INIT_02 => X"0000001d0000000f0000000d0000000c0000000700000004000000000000000e",
            INIT_03 => X"0000000000000000000000010000000000000000000000240000002600000028",
            INIT_04 => X"0000000e00000006000000200000000900000009000000060000000a00000009",
            INIT_05 => X"0000000a000000000000000300000009000000290000004b0000008000000042",
            INIT_06 => X"0000000000000046000000820000003c0000000c000000070000000a0000000c",
            INIT_07 => X"000000090000000c000000000000000400000000000000440000006400000000",
            INIT_08 => X"000000000000000000000000000000000000000000000038000000040000000a",
            INIT_09 => X"000000220000000a0000000500000000000000000000002e0000004f00000025",
            INIT_0A => X"00000011000000fa000000f300000073000000030000000d0000000000000045",
            INIT_0B => X"00000000000000120000001800000006000000610000000c0000000000000000",
            INIT_0C => X"000000000000000000000000000000000000006b000000000000000000000000",
            INIT_0D => X"000000000000000000000030000000ab000000150000003b000000a80000002f",
            INIT_0E => X"0000008600000060000000000000000000000000000000000000000600000000",
            INIT_0F => X"0000002e00000000000000000000000000000000000000200000000000000018",
            INIT_10 => X"000000000000000000000000000000000000000000000000000000000000004c",
            INIT_11 => X"0000000f000000240000001b0000000000000000000000000000000300000000",
            INIT_12 => X"000000000000000000000000000000000000000400000009000000000000000c",
            INIT_13 => X"000000000000004d000000780000005f00000016000000000000000000000001",
            INIT_14 => X"0000000d00000000000000000000000000000008000000330000000f00000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000b0000000e000000000000000000000000000000000000000000000000",
            INIT_17 => X"000000000000000a000000110000001f00000026000000230000004a00000012",
            INIT_18 => X"000001450000013c0000012f0000000c00000008000000070000000000000000",
            INIT_19 => X"000000ba000000bb000000f00000010c0000011900000127000001410000014b",
            INIT_1A => X"000001170000012000000126000001340000008a0000003e0000005c0000009c",
            INIT_1B => X"000000840000009d000000b9000000ca000000db000000e4000000ec00000102",
            INIT_1C => X"000000cc000000d8000000de000000df000000e30000009c000000470000002d",
            INIT_1D => X"00000046000000290000006d000000b2000000bc000000c1000000c5000000c4",
            INIT_1E => X"000000c3000000c0000000bd000000bb000000b9000000b3000000a300000079",
            INIT_1F => X"000000a50000007e0000001700000047000000a8000000bc000000c2000000bf",
            INIT_20 => X"000000a3000000b9000000bd000000bf000000bf000000bd000000af000000a9",
            INIT_21 => X"000000a1000000a20000008a00000031000000290000008c0000008d000000a1",
            INIT_22 => X"0000003c0000004f0000006e000000a7000000bd000000bf000000be000000ba",
            INIT_23 => X"000000c0000000930000006f000000190000005500000000000000000000002e",
            INIT_24 => X"000000170000001c00000022000000380000007c000000a2000000be000000c0",
            INIT_25 => X"000000be000000be0000005f0000001f00000027000000330000000000000000",
            INIT_26 => X"0000000300000000000000000000000b0000001e000000310000007000000085",
            INIT_27 => X"0000005c00000090000000bd0000001100000000000000170000003500000000",
            INIT_28 => X"0000002000000000000000000000000000000000000000000000001100000006",
            INIT_29 => X"0000000000000034000000420000009800000000000000070000001300000045",
            INIT_2A => X"00000000000000000000001b0000000000000000000000000000000000000013",
            INIT_2B => X"0000000700000009000000000000000800000075000000220000000000000000",
            INIT_2C => X"00000000000000000000000e000000000000002a000000000000000000000000",
            INIT_2D => X"00000000000000000000000e00000000000000010000006b000000190000000a",
            INIT_2E => X"0000001f000000000000000000000009000000000000002a0000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000004e00000011",
            INIT_30 => X"0000001900000011000000000000000f0000000d000000000000002b00000000",
            INIT_31 => X"000000000000000000000000000000000000000000000000000000100000004c",
            INIT_32 => X"000000450000000a000000060000000100000017000000020000000000000000",
            INIT_33 => X"0000000600000000000000000000000000000000000000020000000000000018",
            INIT_34 => X"0000007800000082000000020000000600000007000000070000000600000000",
            INIT_35 => X"0000004a0000006e000000660000007900000075000000770000008300000088",
            INIT_36 => X"0000007300000078000000870000004400000041000000150000004600000051",
            INIT_37 => X"000000550000005a0000006100000062000000700000006d000000770000007a",
            INIT_38 => X"0000006b0000006e00000062000000650000004e0000004b000000080000002f",
            INIT_39 => X"000000010000003b0000005f0000005d0000006000000065000000660000006a",
            INIT_3A => X"0000006a00000063000000650000006900000063000000420000004f00000028",
            INIT_3B => X"000000490000003a00000000000000500000005d000000600000006b00000067",
            INIT_3C => X"000000660000006f000000660000006a0000006b000000650000005100000049",
            INIT_3D => X"0000005700000042000000290000000000000024000000570000005900000053",
            INIT_3E => X"0000004a000000630000006a00000064000000650000006a0000006900000053",
            INIT_3F => X"00000050000000280000003f0000000000000000000000000000001200000021",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE44;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE45 : if BRAM_NAME = "samplegold_layer0_instance45" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000230000005f000000640000005f000000690000006b",
            INIT_01 => X"0000006c0000003d00000022000000020000000000000036000000720000000e",
            INIT_02 => X"0000003b00000012000000000000002f000000050000003e0000006300000063",
            INIT_03 => X"0000006500000068000000360000001f00000000000000000000000000000044",
            INIT_04 => X"00000000000000000000003e0000005b00000017000000000000002000000022",
            INIT_05 => X"000000000000007c00000073000000180000004c0000003c0000000000000000",
            INIT_06 => X"0000000c0000000000000000000000060000007300000031000000000000001f",
            INIT_07 => X"0000000000000000000000180000009500000000000000000000000d00000000",
            INIT_08 => X"0000006900000021000000000000000000000000000000720000003000000000",
            INIT_09 => X"0000001e0000000000000000000000150000005d000000000000000000000000",
            INIT_0A => X"000000060000005d000000000000001200000000000000000000005600000033",
            INIT_0B => X"0000000b0000003b000000000000000600000018000000500000001500000000",
            INIT_0C => X"000000000000002f00000017000000000000002b00000000000000000000002f",
            INIT_0D => X"0000000300000008000000170000000000000000000000290000003e00000026",
            INIT_0E => X"0000001b000000020000001400000000000000000000002c0000000000000000",
            INIT_0F => X"0000000600000007000000080000000800000000000000060000000b00000035",
            INIT_10 => X"000000ac0000001a000000110000001000000000000000000000003400000007",
            INIT_11 => X"000000a7000000b1000000b6000000bf000000cc000000cd000000c4000000bf",
            INIT_12 => X"000000b1000000c40000006800000032000000410000007a000000880000008b",
            INIT_13 => X"000000860000008f0000009b000000a1000000a8000000b8000000c1000000ba",
            INIT_14 => X"000000a4000000aa0000009c0000007200000026000000320000005300000072",
            INIT_15 => X"0000003600000082000000830000008800000091000000900000009a000000a2",
            INIT_16 => X"0000008b0000008b0000008d0000008900000071000000400000002700000018",
            INIT_17 => X"00000018000000390000006f000000740000007a000000810000008d0000008c",
            INIT_18 => X"0000008d0000008f0000008f0000008f00000082000000820000007a00000055",
            INIT_19 => X"0000004e00000000000000000000001800000046000000680000006000000079",
            INIT_1A => X"00000042000000860000008d0000008d000000900000008e0000007800000073",
            INIT_1B => X"000000340000001f000000000000000000000000000000000000000000000000",
            INIT_1C => X"00000026000000310000003e000000860000008f0000008f000000900000006d",
            INIT_1D => X"0000004200000025000000000000000000000000000000000000003400000031",
            INIT_1E => X"000000000000000500000003000000120000002b00000068000000910000008f",
            INIT_1F => X"0000009000000000000000190000000a00000000000000000000000000000000",
            INIT_20 => X"00000000000000000000000000000011000000050000000f0000002e00000082",
            INIT_21 => X"00000000000000950000000000000000000000150000001f0000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000009000000120000000000000000",
            INIT_23 => X"0000000000000011000000680000000000000000000000000000000000000000",
            INIT_24 => X"000000120000002d000000000000000000000000000000000000001c00000000",
            INIT_25 => X"000000000000000000000000000000760000002f000000000000000000000000",
            INIT_26 => X"0000000000000001000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000100000059000000190000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"00000020000000080000000a0000000000000016000000440000002100000018",
            INIT_2A => X"0000002200000021000000110000000c000000000000002e0000002700000022",
            INIT_2B => X"00000000000000000000000000000000000000000000001e0000003500000017",
            INIT_2C => X"0000000a00000010000000120000001c0000000c0000000b0000000b00000002",
            INIT_2D => X"0000004a0000004c0000005100000059000000550000004c0000003f00000026",
            INIT_2E => X"0000004c0000001a0000001b0000002f000000300000002b0000004200000040",
            INIT_2F => X"000000320000003b0000003f000000460000004f000000530000004f00000045",
            INIT_30 => X"00000053000000570000001c000000000000000a0000001a0000001400000029",
            INIT_31 => X"0000001f00000023000000240000002b0000002c000000340000004100000047",
            INIT_32 => X"000000290000002a0000002b000000250000000100000000000000250000002c",
            INIT_33 => X"000000290000001e00000015000000120000001c000000280000002600000028",
            INIT_34 => X"0000002e0000002d0000002b000000250000002b000000270000001000000000",
            INIT_35 => X"000000000000000000000000000000000000001300000028000000300000002c",
            INIT_36 => X"000000200000002c0000002b0000002c0000002a00000027000000260000001a",
            INIT_37 => X"0000002e0000000000000000000000970000008a000000540000000a00000000",
            INIT_38 => X"0000003a0000002700000025000000320000002d0000002b000000230000000f",
            INIT_39 => X"0000003200000000000000000000000000000000000000130000002400000029",
            INIT_3A => X"0000000000000007000000060000000a0000001e0000002e0000002e00000022",
            INIT_3B => X"00000000000000000000000e0000006b00000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000030000002500000021000000010000001600000031",
            INIT_3D => X"0000001d0000000000000000000000000000000600000000000000130000001f",
            INIT_3E => X"0000000300000000000000000000000f00000014000000000000000000000000",
            INIT_3F => X"000000860000002f000000220000000000000000000000000000008c0000006d",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE45;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE46 : if BRAM_NAME = "samplegold_layer0_instance46" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003100000030000000000000000000000000000000060000000000000023",
            INIT_01 => X"00000000000000000000002900000056000000370000002e0000005300000001",
            INIT_02 => X"0000000000000000000000300000000000000000000000000000000000000004",
            INIT_03 => X"0000000000000000000000030000001d00000001000000270000000f00000006",
            INIT_04 => X"0000000000000000000000000000001200000000000000000000000000000000",
            INIT_05 => X"0000004f000000470000003e0000001f0000000900000007000000350000002c",
            INIT_06 => X"00000012000000050000000e000000000000007a000000900000008b0000007e",
            INIT_07 => X"0000000000000000000000000000000000000000000000130000000000000010",
            INIT_08 => X"00000000000000000000000e0000003300000010000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"00000000000000000000000000000000000000000000001c0000000700000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000200000012",
            INIT_11 => X"0000001e0000000b000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"000000020000009d000000ab0000008600000063000000490000000000000000",
            INIT_14 => X"000000000000000000000000000000000000000000000000000000000000001c",
            INIT_15 => X"0000000000000078000000d9000000400000002d000000410000006400000036",
            INIT_16 => X"000000240000002c000000000000000000000000000000000000000000000022",
            INIT_17 => X"0000000000000016000000ba000000e8000000760000002f0000001f00000030",
            INIT_18 => X"000000450000002000000036000000490000000500000000000000000000001f",
            INIT_19 => X"0000007e000000220000001600000051000000e100000102000000ee000000bf",
            INIT_1A => X"000000df00000053000000090000000c000000270000003e0000003c00000000",
            INIT_1B => X"00000000000000910000009f0000007900000098000000f1000000d6000000e6",
            INIT_1C => X"000000c5000000d6000000560000000a000000000000001c0000008700000098",
            INIT_1D => X"000000290000000000000052000000a5000000c7000000ce000000370000005f",
            INIT_1E => X"0000001700000093000000d80000009800000040000000000000001600000077",
            INIT_1F => X"000000750000002e00000000000000000000005b000000a80000002c00000012",
            INIT_20 => X"000000230000002e0000007e000000d70000009e000000670000003400000022",
            INIT_21 => X"0000003b000000540000001c0000000000000000000000320000007500000000",
            INIT_22 => X"00000000000000430000003100000072000000a20000009d0000008d00000056",
            INIT_23 => X"000000000000000800000019000000030000000000000000000000000000000e",
            INIT_24 => X"0000000000000000000000290000001600000000000000000000000000000004",
            INIT_25 => X"0000001500000016000000110000000000000000000000000000000000000000",
            INIT_26 => X"0000000100000039000000000000000c0000002600000017000000110000000f",
            INIT_27 => X"0000000a0000000e000000120000001600000018000000050000000800000000",
            INIT_28 => X"0000000000000000000000000000002700000000000000000000000300000007",
            INIT_29 => X"000000000000000000000000000000020000000d0000000d0000002800000026",
            INIT_2A => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000004800000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_2F => X"000000000000001f0000003b0000000000000000000000000000000000000000",
            INIT_30 => X"000000000000000000000000000000000000000300000000000000000000005d",
            INIT_31 => X"0000000000000000000000000000002d00000074000000600000004f00000000",
            INIT_32 => X"0000001a00000000000000000000000000000000000000090000000e00000031",
            INIT_33 => X"000000000000006e000000000000000000000000000000000000000000000000",
            INIT_34 => X"00000018000000390000000c0000003d00000000000000000000000000000000",
            INIT_35 => X"00000000000000000000003e0000002d00000000000000100000000000000000",
            INIT_36 => X"00000000000000000000002a0000000500000039000000000000000000000000",
            INIT_37 => X"0000004200000000000000000000000000000000000000810000000000000000",
            INIT_38 => X"000000000000000000000000000000060000001e000000020000007700000000",
            INIT_39 => X"000000140000007a0000004c000000290000000000000075000000590000007a",
            INIT_3A => X"0000005d00000000000000000000000000000000000000250000000000000000",
            INIT_3B => X"00000000000000090000000000000061000000000000002b0000000100000000",
            INIT_3C => X"000000000000003b000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000003900000002000000000000000500000040000000180000002500000000",
            INIT_3E => X"000000190000000000000048000000a50000009d000000930000006900000038",
            INIT_3F => X"0000000000000000000000000000000000000000000000070000003f00000021",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE46;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE47 : if BRAM_NAME = "samplegold_layer0_instance47" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000b000000200000001e0000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000017000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000180000000000000000",
            INIT_0D => X"0000004600000069000000230000001d0000001c0000000d0000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000130000000b00000000",
            INIT_0F => X"000000000000001f0000003b0000001100000012000000020000001100000000",
            INIT_10 => X"000000010000001d0000000000000000000000000000000d0000001b00000000",
            INIT_11 => X"0000000e00000000000000020000001a0000001c0000003c000000460000002e",
            INIT_12 => X"000000350000000000000030000000000000000d00000000000000140000001d",
            INIT_13 => X"0000001800000014000000000000002700000016000000280000003700000076",
            INIT_14 => X"00000078000000360000000d00000014000000000000002c000000040000000a",
            INIT_15 => X"000000000000001100000016000000810000005500000005000000060000002e",
            INIT_16 => X"00000022000000690000004b00000025000000000000001f0000002800000000",
            INIT_17 => X"00000000000000080000000000000035000000690000000b0000002400000000",
            INIT_18 => X"000000000000002b000000530000002600000042000000000000003100000026",
            INIT_19 => X"0000002000000000000000150000000000000052000000260000000000000031",
            INIT_1A => X"0000004600000000000000490000004f0000005100000054000000250000002d",
            INIT_1B => X"0000001c0000000b000000000000001900000012000000310000000600000010",
            INIT_1C => X"000000170000003900000013000000180000001a0000001c0000001d00000010",
            INIT_1D => X"0000000b00000019000000130000002b0000001a000000150000001400000002",
            INIT_1E => X"00000005000000000000000000000008000000000000000c0000000200000000",
            INIT_1F => X"0000000000000000000000000000000200000006000000080000001400000000",
            INIT_20 => X"0000000000000000000000140000000700000005000000000000000700000000",
            INIT_21 => X"000000040000000300000000000000000000000000000004000000070000003d",
            INIT_22 => X"000000340000000900000000000000300000000f0000000c0000000900000007",
            INIT_23 => X"0000000e0000000a0000000a0000000300000006000000060000000400000005",
            INIT_24 => X"000000000000000a000000190000002000000000000000150000001200000011",
            INIT_25 => X"0000000e0000001c000000170000000c0000000300000004000000060000000b",
            INIT_26 => X"0000000900000008000000040000000d0000002b00000000000000040000001a",
            INIT_27 => X"0000002c000000330000004c0000002a00000012000000040000000400000004",
            INIT_28 => X"0000000200000005000000050000000800000025000000000000003c00000000",
            INIT_29 => X"000000600000000000000000000000000000000e000000340000000b00000000",
            INIT_2A => X"000000160000000000000003000000070000001c00000000000000000000006c",
            INIT_2B => X"0000001f0000009c0000005f0000002e00000000000000250000000000000019",
            INIT_2C => X"00000009000000030000000e00000001000000510000001b0000000000000000",
            INIT_2D => X"0000000000000000000000060000002200000095000000410000001f00000000",
            INIT_2E => X"000000000000002300000000000000800000000c000000430000005100000022",
            INIT_2F => X"00000039000000000000000b0000000000000010000000370000008600000036",
            INIT_30 => X"000000470000000000000007000000000000000e000000450000000000000015",
            INIT_31 => X"0000000000000000000000610000002b00000000000000000000002000000093",
            INIT_32 => X"0000007c000000600000002800000000000000250000000e0000001a00000000",
            INIT_33 => X"00000002000000000000002000000067000000000000001e0000000000000017",
            INIT_34 => X"000000090000006a0000003a0000005a00000000000000320000001e00000012",
            INIT_35 => X"000000160000002200000000000000530000001c000000000000003900000000",
            INIT_36 => X"0000000000000000000000000000000800000030000000000000001e00000022",
            INIT_37 => X"000000030000001300000022000000000000002100000000000000000000004d",
            INIT_38 => X"0000003d0000001000000012000000180000001c000000190000001200000009",
            INIT_39 => X"000000000000000000000000000000270000001c0000001a0000000000000004",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_3E => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000011",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE47;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE48 : if BRAM_NAME = "samplegold_layer0_instance48" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"000000000000000000000000000000270000002b0000002b0000001900000000",
            INIT_03 => X"000000000000003b000000150000000000000000000000000000000000000000",
            INIT_04 => X"00000000000000000000000000000000000000020000002a0000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"000000000000000000000000000000000000000f000000020000000000000000",
            INIT_07 => X"0000006e000000d10000006d0000000000000000000000000000000000000000",
            INIT_08 => X"000000000000000000000000000000510000000c000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000f0000000d000000000000000000000000",
            INIT_0A => X"0000000000000000000000450000000000000010000000680000003100000000",
            INIT_0B => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"000000000000000000000000000000000000000000000000000000000000002a",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000001f00000030",
            INIT_0E => X"000000040000001f000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000600000000000000000000000000000000",
            INIT_10 => X"000000000000004e000000500000001100000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000019000000110000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000003000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000f000000120000001e0000002400000025000000380000001d00000000",
            INIT_15 => X"0000008400000080000000130000000f0000000f000000000000000000000000",
            INIT_16 => X"0000003c0000005a000000640000006d00000074000000850000008900000089",
            INIT_17 => X"00000076000000760000007b0000001f000000000000000e0000002800000038",
            INIT_18 => X"0000002d00000036000000430000004b0000005200000055000000610000006c",
            INIT_19 => X"000000490000004900000050000000560000002c000000000000000000000021",
            INIT_1A => X"0000000000000024000000370000003c0000003f000000420000004100000043",
            INIT_1B => X"0000003f0000003c0000003d0000003900000033000000360000001c00000000",
            INIT_1C => X"00000018000000000000000c0000003a00000040000000440000004200000042",
            INIT_1D => X"000000410000003e0000003f0000003f0000003d000000360000002e00000032",
            INIT_1E => X"0000002b000000270000000000000000000000380000002e000000380000003f",
            INIT_1F => X"0000002400000020000000330000003e0000003f0000003f0000003c0000002c",
            INIT_20 => X"000000250000002600000000000000190000000d0000000d0000003800000035",
            INIT_21 => X"000000000000000000000019000000280000002e000000400000004000000040",
            INIT_22 => X"0000003f00000008000000000000000000000024000000150000000000000000",
            INIT_23 => X"000000000000000000000000000000000000000c00000028000000210000003f",
            INIT_24 => X"000000280000003f0000000000000000000000000000002a000000200000001a",
            INIT_25 => X"0000001b0000002e0000001d0000000000000000000000000000000000000012",
            INIT_26 => X"0000001c00000025000000240000001400000000000000000000000000000035",
            INIT_27 => X"00000000000000210000000a0000001500000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000110000001c000000170000000f0000001a00000015",
            INIT_29 => X"000000000000000000000000000000300000000a000000000000000000000000",
            INIT_2A => X"000000000000000000000000000000000000001a00000000000000090000000c",
            INIT_2B => X"0000000000000000000000000000000000000022000000100000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000040000000000000005",
            INIT_2D => X"0000000000000000000000000000000000000000000000100000000300000002",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000004",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000004000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000029000000000000000300000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000190000002700000000",
            INIT_36 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"000000000000000000000000000000000000000600000000000000160000001b",
            INIT_38 => X"000000000000003e000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000b000000140000002f0000002400000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000001",
            INIT_3C => X"0000000f000000000000008a00000000000000000000000b0000001200000000",
            INIT_3D => X"0000000a00000005000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000300000000000000440000006000000000000000000000000000000017",
            INIT_3F => X"0000000000000019000000000000001f0000000e000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE48;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE49 : if BRAM_NAME = "samplegold_layer0_instance49" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000020000001d0000005d000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000200000033000000000000002500000000",
            INIT_02 => X"00000000000000000000000000000000000000000000003f0000001a00000000",
            INIT_03 => X"0000002200000000000000000000000000000000000000320000000000000078",
            INIT_04 => X"0000001e00000000000000000000001f00000008000000100000000100000000",
            INIT_05 => X"0000000900000013000000400000000000000000000000000000001900000028",
            INIT_06 => X"0000004200000000000000000000000000000039000000190000000800000000",
            INIT_07 => X"0000000000000020000000040000007800000000000000000000000000000003",
            INIT_08 => X"000000000000002c000000000000000000000000000000030000005900000000",
            INIT_09 => X"000000000000001e00000030000000000000006d000000000000000000000000",
            INIT_0A => X"00000000000000000000000c0000000d00000000000000000000000a0000003c",
            INIT_0B => X"00000010000000140000003100000012000000000000000b0000000000000000",
            INIT_0C => X"000000200000001c0000001e0000002c00000011000000130000000000000012",
            INIT_0D => X"000000130000001c0000001d000000210000001200000003000000200000001e",
            INIT_0E => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"000000000000000b000000100000000100000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000008000000250000001c00000017000000140000000000000000",
            INIT_13 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"000000000000001100000015000000140000001d000000210000001f00000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000006",
            INIT_16 => X"000000170000001c0000001e0000002000000014000000040000000500000007",
            INIT_17 => X"0000000c00000000000000070000000000000000000000000000000000000000",
            INIT_18 => X"00000002000000210000001f0000001b0000001b000000220000001300000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"000000000000000d000000180000001f00000015000000140000001f00000011",
            INIT_1B => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"000000000000000a0000001d0000001c00000021000000130000000a0000000a",
            INIT_1D => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"00000000000000000000000000000019000000220000001c0000001b00000014",
            INIT_1F => X"0000001300000018000000000000000c00000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000001600000019000000220000001600000016",
            INIT_21 => X"000000110000000b00000010000000140000002c000000070000002b00000011",
            INIT_22 => X"0000000000000013000000000000000000000004000000180000002900000016",
            INIT_23 => X"00000009000000200000001700000000000000100000001c0000000c00000000",
            INIT_24 => X"0000000000000000000000000000000000000001000000000000001100000014",
            INIT_25 => X"0000001300000000000000070000000300000018000000000000000000000000",
            INIT_26 => X"0000000800000000000000000000000000000000000000000000000000000016",
            INIT_27 => X"000000170000001c000000120000000000000001000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000a00000000000000000000000000000005",
            INIT_29 => X"000000000000000e000000000000000000000000000000000000000600000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000050000000000000000",
            INIT_3E => X"000000200000000c000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE49;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE50 : if BRAM_NAME = "samplegold_layer0_instance50" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000020000000800000000000000020000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000003000000000000000100000000",
            INIT_09 => X"0000000500000008000000050000000200000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000100000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000001a00000015000000000000000000000001000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000012000000150000000000000003000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"00000000000000080000000d0000000e00000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"00000000000000000000000e000000140000000e000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000008",
            INIT_15 => X"00000000000000000000001a000000210000001c000000120000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"000000000000000000000000000000000000001d000000330000003800000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000001f0000002c",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000002000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000500000003",
            INIT_1E => X"0000000000000003000000010000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"000000150000002600000011000000220000001f000000000000000000000000",
            INIT_23 => X"000000170000001e0000001c0000001d0000001f0000001b0000001e0000000c",
            INIT_24 => X"00000000000000160000000e00000018000000250000001f000000100000000a",
            INIT_25 => X"0000000d0000000800000008000000090000001100000011000000090000000e",
            INIT_26 => X"000000000000000000000005000000050000002f0000001f0000001d00000018",
            INIT_27 => X"00000025000000270000001d0000001a000000170000000d0000000000000000",
            INIT_28 => X"00000000000000000000000000000000000000000000002b0000001000000016",
            INIT_29 => X"000000000000001500000020000000150000001d000000080000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000240000006600000008",
            INIT_2B => X"0000002e00000021000000110000001400000005000000000000000000000000",
            INIT_2C => X"000000000000000000000001000000020000000000000000000000230000007b",
            INIT_2D => X"0000003a000000320000002f0000002000000013000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000010000000000000000000000060",
            INIT_2F => X"000000310000003b0000001d0000001d0000002f0000000d0000000000000000",
            INIT_30 => X"00000000000000000000000d00000000000000000000000d0000000000000053",
            INIT_31 => X"0000003c0000003e0000001e0000000800000015000000110000000000000000",
            INIT_32 => X"0000000000000000000000000000000400000000000000080000000d00000052",
            INIT_33 => X"000000690000001f000000a300000065000000380000001b0000002900000004",
            INIT_34 => X"0000001600000000000000000000000000000000000000000000001700000000",
            INIT_35 => X"000000000000001d0000001400000033000000970000007b000000510000000d",
            INIT_36 => X"0000001800000005000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000001900000000000000000000002d0000003800000051000000610000007d",
            INIT_38 => X"000000340000002c000000000000000300000005000000000000000000000000",
            INIT_39 => X"00000000000000160000000000000018000000330000001c0000002100000029",
            INIT_3A => X"00000015000000140000000400000000000000120000000c0000000a00000000",
            INIT_3B => X"000000000000000000000004000000000000000e0000000a0000002700000025",
            INIT_3C => X"0000000b0000001e0000002700000000000000030000000c0000000100000000",
            INIT_3D => X"0000000000000000000000000000000f0000001100000002000000000000000b",
            INIT_3E => X"0000000000000000000000000000000000000007000000000000000b00000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000040000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE50;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE51 : if BRAM_NAME = "samplegold_layer0_instance51" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000002000000000000000000000000000000000000000d0000000300000000",
            INIT_01 => X"000000350000002a000000150000000300000000000000030000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000002a00000036",
            INIT_03 => X"0000000000000005000000180000002100000032000000180000000000000000",
            INIT_04 => X"0000000f00000005000000000000001b0000001b000000030000000000000000",
            INIT_05 => X"0000000b00000007000000000000000000000000000000000000000000000008",
            INIT_06 => X"00000014000000270000000700000005000000070000004f000000640000004e",
            INIT_07 => X"0000001b000000210000001b0000000600000000000000000000000000000004",
            INIT_08 => X"000000070000000000000000000000250000001a000000120000000000000003",
            INIT_09 => X"0000000000000000000000050000000200000000000000000000000500000008",
            INIT_0A => X"000000100000000d000000000000000000000000000000000000003b00000000",
            INIT_0B => X"0000000f00000011000000000000000000000000000000000000000000000005",
            INIT_0C => X"000000050000000b0000000d0000000f0000001f000000480000005400000000",
            INIT_0D => X"0000006b0000005e00000025000000140000000b000000000000000000000004",
            INIT_0E => X"0000000b0000000f00000000000000000000001b000000150000003f00000031",
            INIT_0F => X"000000000000000000000000000000580000007b000000000000000000000000",
            INIT_10 => X"00000000000000080000000b0000000000000005000000050000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000300000000000000000000000000000000000000000000000000000015",
            INIT_14 => X"0000001000000000000000000000000b0000001200000000000000000000000d",
            INIT_15 => X"0000000000000000000000230000001300000001000000000000000000000000",
            INIT_16 => X"00000000000000000000000100000008000000000000001d0000000a00000013",
            INIT_17 => X"00000000000000000000000f0000000400000000000000000000000000000005",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000200000000000000000000000000000000",
            INIT_1A => X"0000000a0000000c000000080000000000000000000000000000000000000000",
            INIT_1B => X"0000000f00000012000000100000001100000025000000250000001b00000010",
            INIT_1C => X"00000011000000110000000c000000080000000e0000000b0000000d0000000e",
            INIT_1D => X"0000001b0000001b000000130000001f0000003300000033000000350000002d",
            INIT_1E => X"00000033000000150000001e0000000a0000000a0000001d0000001a0000001a",
            INIT_1F => X"0000002a0000002b000000250000002100000032000000510000004c00000041",
            INIT_20 => X"00000042000000330000002d0000001b0000000c0000000d0000002900000027",
            INIT_21 => X"00000029000000290000003a0000002d0000003b0000005f0000005e0000004f",
            INIT_22 => X"0000003f00000028000000390000002e000000370000000e0000000b00000030",
            INIT_23 => X"00000047000000430000003900000047000000520000005f000000620000005a",
            INIT_24 => X"0000004b000000420000002e0000002a00000032000000270000001b00000017",
            INIT_25 => X"000000160000004e000000510000004f0000004e000000670000006100000052",
            INIT_26 => X"00000044000000470000004300000028000000380000003d0000001500000018",
            INIT_27 => X"00000019000000130000003c0000004400000056000000510000005d00000050",
            INIT_28 => X"00000045000000400000004f0000004c00000030000000370000001d0000002c",
            INIT_29 => X"0000001b00000015000000180000003600000039000000470000005900000055",
            INIT_2A => X"0000004c0000003d0000003d000000580000003a000000550000003300000049",
            INIT_2B => X"000000370000002d000000210000001900000052000000490000004100000055",
            INIT_2C => X"00000053000000460000003a0000003e0000005700000038000000480000002e",
            INIT_2D => X"0000003e00000034000000440000002d0000001a000000500000005300000049",
            INIT_2E => X"00000052000000510000004b000000450000004400000042000000480000003f",
            INIT_2F => X"0000003b0000003c0000002000000022000000150000001e0000005a0000004c",
            INIT_30 => X"0000004f000000600000004c0000003d0000003b00000037000000400000002e",
            INIT_31 => X"0000003800000034000000290000002500000017000000140000001a0000005d",
            INIT_32 => X"0000004f000000620000006000000045000000340000002a0000002f00000039",
            INIT_33 => X"000000490000003c000000400000003f0000004000000035000000260000001c",
            INIT_34 => X"000000350000005a000000600000005b0000003b0000002b0000003e00000043",
            INIT_35 => X"0000005b0000005a00000051000000490000004f00000053000000470000003e",
            INIT_36 => X"00000000000000000000005f00000063000000580000004e0000004800000051",
            INIT_37 => X"000000000000000000000000000000000000000000000000000000000000000a",
            INIT_38 => X"000000050000000000000000000000050000000b000000010000000000000000",
            INIT_39 => X"0000000600000003000000000000000000000000000000020000000000000005",
            INIT_3A => X"00000009000000000000000000000000000000090000000f0000000d0000000a",
            INIT_3B => X"0000000600000005000000030000000a00000000000000000000000000000000",
            INIT_3C => X"000000000000000f000000000000000000000000000000060000000700000008",
            INIT_3D => X"0000000d00000000000000000000000800000000000000060000000000000000",
            INIT_3E => X"0000000a0000000000000000000000000000000e000000100000000c00000006",
            INIT_3F => X"0000001300000011000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE51;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE52 : if BRAM_NAME = "samplegold_layer0_instance52" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000015000000000000000000000000000000000000000600000015",
            INIT_01 => X"00000012000000190000001a0000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000100000001800000000000000000000000000000000",
            INIT_03 => X"0000000100000003000000180000000000000005000000000000000000000000",
            INIT_04 => X"0000000000000002000000000000002400000000000000000000000000000007",
            INIT_05 => X"0000000f00000007000000100000000900000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000900000000000000000000000000000000",
            INIT_07 => X"0000000000000008000000140000000600000005000000000000000000000000",
            INIT_08 => X"000000000000000000000000000000000000000f000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000022000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000170000000e00000000",
            INIT_0C => X"0000000000000000000000000000000000000007000000000000000a00000000",
            INIT_0D => X"000000000000000000000009000000000000000000000000000000000000002c",
            INIT_0E => X"0000002300000000000000000000000000000009000000000000000000000007",
            INIT_0F => X"0000000f000000130000001400000001000000010000000c0000000800000020",
            INIT_10 => X"0000002a0000001c000000000000000000000000000000060000000100000004",
            INIT_11 => X"000000120000000e00000022000000340000001a000000160000000900000003",
            INIT_12 => X"00000000000000270000002600000009000000120000001a000000170000001e",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000040000000400000003000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"000000000000000000000000000000000000000c000000010000000000000000",
            INIT_19 => X"0000000000000000000000030000000500000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000080000000000000003",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000700000007",
            INIT_1D => X"0000001200000006000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000010",
            INIT_1F => X"0000001300000013000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000006000000080000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"00000000000000000000002b0000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000003300000016000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000100000000000000010000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000026000000100000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000200000001d0000000c",
            INIT_2A => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"000000130000002b0000001d0000000000000000000000000000002200000024",
            INIT_2C => X"0000002e00000001000000000000000000000000000000080000000300000006",
            INIT_2D => X"000000110000001d0000002c0000002b0000002e000000270000000a0000002e",
            INIT_2E => X"0000003b00000036000000280000001e0000001a000000210000002f00000029",
            INIT_2F => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000030000000a00000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000700000012",
            INIT_34 => X"0000000000000000000000000000000d0000000e000000050000000000000000",
            INIT_35 => X"0000000000000008000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000001e000000030000000000000000000000090000000d0000000c00000008",
            INIT_3B => X"0000001800000002000000000000000000000000000000000000000000000006",
            INIT_3C => X"0000000000000000000000000000001d0000000000000000000000000000001c",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000027000000080000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE52;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE53 : if BRAM_NAME = "samplegold_layer0_instance53" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000000000000210000001a000000350000003d00000000",
            INIT_01 => X"0000001e000000030000000e0000000200000000000000000000000000000000",
            INIT_02 => X"00000000000000000000001a000000060000002500000018000000130000001b",
            INIT_03 => X"00000021000000430000006a0000000200000000000000000000000000000000",
            INIT_04 => X"000000000000000000000000000000000000000000000000000000000000000f",
            INIT_05 => X"0000000000000000000000130000001d000000000000000f0000000000000000",
            INIT_06 => X"00000000000000000000000000000000000000000000000b0000000000000012",
            INIT_07 => X"0000001300000025000000170000000000000000000000120000000300000000",
            INIT_08 => X"0000000500000000000000190000000800000002000000020000000000000001",
            INIT_09 => X"0000000b0000000a0000000a0000000f00000022000000200000001100000013",
            INIT_0A => X"0000001100000012000000140000000300000001000000070000000e00000003",
            INIT_0B => X"0000003c00000042000000400000004900000046000000440000004a00000015",
            INIT_0C => X"00000002000000080000000f00000019000000240000002a0000002f0000003b",
            INIT_0D => X"0000002a00000038000000350000003100000030000000400000004200000048",
            INIT_0E => X"000000430000001400000012000000110000001300000019000000220000002a",
            INIT_0F => X"000000280000001c0000001700000016000000210000001f0000003300000042",
            INIT_10 => X"0000003a00000039000000250000003100000031000000340000003500000033",
            INIT_11 => X"0000004200000019000000110000000c00000011000000120000000000000022",
            INIT_12 => X"0000005900000055000000450000001600000024000000320000003b00000043",
            INIT_13 => X"0000002a0000001700000016000000160000002d0000002c0000000d00000006",
            INIT_14 => X"0000000b000000880000008f000000810000001900000020000000330000003a",
            INIT_15 => X"0000002b0000001100000011000000220000002d0000003c0000002700000013",
            INIT_16 => X"0000001c00000022000000860000008b0000008f0000002c0000003000000035",
            INIT_17 => X"000000340000001c000000180000002400000032000000280000003800000038",
            INIT_18 => X"0000000e000000270000007300000081000000800000007e000000340000003c",
            INIT_19 => X"0000002b00000031000000160000001d0000003b000000410000001f00000020",
            INIT_1A => X"000000480000005000000087000000650000009b000000910000008300000023",
            INIT_1B => X"000000170000002a000000290000001d0000002900000044000000430000001d",
            INIT_1C => X"0000002f000000490000008500000093000000c6000000e0000000ce000000b3",
            INIT_1D => X"000001010000000000000016000000230000002300000036000000440000003c",
            INIT_1E => X"0000003700000034000000420000005b000000620000008900000094000000fb",
            INIT_1F => X"000000cb000000e800000000000000140000001a000000240000003300000040",
            INIT_20 => X"00000033000000230000000c0000003300000019000000220000005600000082",
            INIT_21 => X"0000005c00000065000000750000000600000017000000110000002d00000037",
            INIT_22 => X"0000004f000000380000001b0000002e00000023000000100000003b0000004d",
            INIT_23 => X"0000002f0000003d0000003e000000450000001a000000040000001e0000003f",
            INIT_24 => X"000000370000004b000000220000000c00000019000000070000001e0000001c",
            INIT_25 => X"00000000000000000000000c0000001e0000002e000000010000000200000026",
            INIT_26 => X"000000030000000d000000000000000000000000000000020000001000000013",
            INIT_27 => X"0000000000000003000000070000000000000002000000000000000000000000",
            INIT_28 => X"0000000000000000000000040000000400000001000000000000000000000005",
            INIT_29 => X"000000000000000c000000000000000900000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000009000000000000000400000000000000220000000000000004",
            INIT_2C => X"000000000000000c000000070000000000000000000000000000000000000000",
            INIT_2D => X"0000000c000000000000000000000000000000000000000d0000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000060000000000000001",
            INIT_2F => X"0000000100000000000000000000000000000000000000010000000900000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000400000000000000000000000000000011000000000000000000000015",
            INIT_32 => X"0000000000000000000000070000000a00000000000000000000000000000000",
            INIT_33 => X"0000000000000001000000000000000000000000000000020000000b00000019",
            INIT_34 => X"00000000000000000000000000000000000000000000001d0000000800000005",
            INIT_35 => X"0000000000000003000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000001",
            INIT_37 => X"0000000b00000000000000000000000000000000000000000000000500000000",
            INIT_38 => X"000000000000000300000018000000040000002d000000000000000000000025",
            INIT_39 => X"0000000000000013000000050000000000000000000000000000000000000002",
            INIT_3A => X"000000120000001a0000002c0000002e000000460000007b0000001b00000000",
            INIT_3B => X"0000007300000002000000000000000000000000000000090000000200000000",
            INIT_3C => X"0000000a0000001a000000000000000f0000002500000000000000020000005e",
            INIT_3D => X"000000190000001f00000000000000000000000a000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000b00000000000000000000000000000005",
            INIT_3F => X"0000001600000000000000000000000000000007000000000000000200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE53;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE54 : if BRAM_NAME = "samplegold_layer0_instance54" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000150000002300000009000000080000000000000000000000110000002a",
            INIT_01 => X"0000000000000009000000250000001e0000000a000000070000001000000003",
            INIT_02 => X"000000140000000d000000000000000100000004000000010000000000000000",
            INIT_03 => X"000000060000000e000000160000000d00000010000000070000000300000007",
            INIT_04 => X"0000000d0000000b0000000c00000009000000090000000d0000000300000000",
            INIT_05 => X"00000000000000000000000a000000120000000b000000100000000a00000011",
            INIT_06 => X"0000000000000000000000010000000300000007000000090000000000000000",
            INIT_07 => X"0000000000000000000000000000000d000000040000000e0000001200000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000003000000000000000f0000000e",
            INIT_0A => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000003",
            INIT_0C => X"0000000800000009000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_0E => X"000000000000000a0000000e0000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_10 => X"0000000000000000000000090000000d00000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_12 => X"0000000000000000000000000000000a00000008000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000f0000000e",
            INIT_19 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000020000000b00000010",
            INIT_1B => X"0000000200000007000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000001700000025000000180000001c00000000000000000000000000000000",
            INIT_20 => X"00000010000000140000001a00000016000000190000001a0000002700000028",
            INIT_21 => X"0000002d0000001300000026000000170000001b000000130000001b00000014",
            INIT_22 => X"00000024000000200000001c0000001b00000017000000290000002b0000003d",
            INIT_23 => X"0000003d0000002a0000002b0000000f0000001a0000001c0000001c00000026",
            INIT_24 => X"00000012000000180000002300000026000000330000003a0000003f00000040",
            INIT_25 => X"00000044000000420000003a0000002b00000003000000210000001e0000000b",
            INIT_26 => X"0000001600000011000000150000001600000032000000360000004000000047",
            INIT_27 => X"0000003200000047000000580000003f00000000000000150000003e00000036",
            INIT_28 => X"0000002e0000001e000000190000002700000032000000480000004400000043",
            INIT_29 => X"0000004400000031000000330000006400000033000000000000000000000021",
            INIT_2A => X"0000001200000019000000110000001b0000003500000046000000420000003d",
            INIT_2B => X"00000035000000480000003f0000002a00000047000000340000000000000008",
            INIT_2C => X"0000001e00000026000000240000000200000023000000330000005100000037",
            INIT_2D => X"00000034000000300000004d000000470000002b000000450000000000000004",
            INIT_2E => X"0000001600000023000000300000002e00000015000000240000003b00000045",
            INIT_2F => X"0000003a0000003900000033000000490000002a000000330000001300000028",
            INIT_30 => X"00000026000000000000000e0000003e00000043000000050000002a00000048",
            INIT_31 => X"0000003f000000320000003d0000003f00000049000000190000003c00000000",
            INIT_32 => X"000000180000002a000000030000000000000001000000180000000d0000000b",
            INIT_33 => X"00000022000000310000002e000000300000003e000000440000002400000037",
            INIT_34 => X"00000047000000350000000a0000000c0000000000000000000000000000000a",
            INIT_35 => X"00000001000000330000001a0000002f00000041000000410000003f00000015",
            INIT_36 => X"0000001d0000003e000000270000000b0000001d000000100000001200000005",
            INIT_37 => X"000000180000001e000000280000001d00000030000000400000005800000046",
            INIT_38 => X"0000002d00000026000000240000001e0000000c000000090000001d00000026",
            INIT_39 => X"00000008000000130000002600000016000000230000002d000000320000003f",
            INIT_3A => X"00000021000000170000000e0000001f0000002900000026000000110000000d",
            INIT_3B => X"000000000000000000000000000000160000001c00000011000000220000002c",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_3E => X"0000001900000009000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000110000001d00000023",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE54;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE55 : if BRAM_NAME = "samplegold_layer0_instance55" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000d00000004000000000000000000000000",
            INIT_01 => X"0000000000000000000000010000000a00000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000004",
            INIT_03 => X"000000080000000000000000000000000000000a000000340000002d00000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"00000000000000000000000c0000000900000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"000000000000000000000000000000000000002d0000001b0000000000000000",
            INIT_0A => X"0000002300000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000012",
            INIT_0C => X"0000000000000000000000000000002400000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000001",
            INIT_12 => X"0000000000000003000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000005000000000000000000000008000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000002200000000000000000000000000000000",
            INIT_20 => X"0000000800000004000000010000000000000001000000040000000200000002",
            INIT_21 => X"000000000000000000000000000000000000001800000011000000100000000b",
            INIT_22 => X"0000001200000016000000060000000000000007000000040000000100000000",
            INIT_23 => X"0000000000000000000000000000000000000009000000060000000900000009",
            INIT_24 => X"00000002000000050000000a0000000c00000000000000030000000000000000",
            INIT_25 => X"00000001000000000000000b0000000000000018000000000000001700000008",
            INIT_26 => X"000000100000000d000000000000000000000000000000000000000000000001",
            INIT_27 => X"00000000000000000000000b0000000700000029000000230000002200000017",
            INIT_28 => X"000000360000003c000000260000000d00000003000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000800000002000000240000001400000030",
            INIT_2A => X"000000000000001b0000003b0000003400000000000000040000000000000000",
            INIT_2B => X"0000000000000002000000000000000000000000000000000000000000000000",
            INIT_2C => X"00000000000000060000000000000009000000240000000a0000000600000000",
            INIT_2D => X"0000000600000007000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000500000000000000000000000000000000000000000000001200000007",
            INIT_2F => X"0000000d0000000c000000000000000400000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000400000005000000000000000000000007",
            INIT_31 => X"0000000c0000000a0000000a0000000000000000000000000000000000000000",
            INIT_32 => X"0000000900000008000000090000000000000000000000000000000000000002",
            INIT_33 => X"000000180000000b000000080000000600000001000000000000000000000006",
            INIT_34 => X"0000001f000000180000002a000000210000001c000000140000000c0000001c",
            INIT_35 => X"0000001d000000190000001c000000160000001e000000200000001e0000001f",
            INIT_36 => X"000000190000002200000036000000310000002e0000002f0000001800000015",
            INIT_37 => X"00000029000000190000001a0000001c000000180000001a0000001a0000001d",
            INIT_38 => X"0000001d0000001c000000200000003e00000046000000410000003900000013",
            INIT_39 => X"0000003200000026000000170000001a0000001900000018000000190000001c",
            INIT_3A => X"0000002b0000001e000000200000004200000045000000440000004600000041",
            INIT_3B => X"0000004700000040000000450000000d0000000a00000017000000170000000e",
            INIT_3C => X"00000014000000310000003a0000004a0000004d000000580000004100000025",
            INIT_3D => X"0000002900000034000000410000003600000009000000070000001600000012",
            INIT_3E => X"0000000c000000180000003c0000005400000051000000460000004d0000004d",
            INIT_3F => X"000000450000001d000000280000004a0000000b000000060000000600000015",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE55;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE56 : if BRAM_NAME = "samplegold_layer0_instance56" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001c0000000e0000003300000041000000550000004d0000003c00000044",
            INIT_01 => X"0000003b00000044000000200000004a00000008000000170000000200000006",
            INIT_02 => X"000000030000001300000023000000390000005300000057000000500000003c",
            INIT_03 => X"0000003f00000051000000120000004000000019000000410000000000000000",
            INIT_04 => X"00000000000000000000001f000000320000003f0000005c0000005200000049",
            INIT_05 => X"00000044000000430000004e0000001f000000390000001d0000002b0000000e",
            INIT_06 => X"0000004c00000009000000000000000d000000360000004b000000600000004b",
            INIT_07 => X"00000045000000430000003f0000002e00000039000000370000002e00000023",
            INIT_08 => X"000000290000000b000000040000000f00000025000000190000004500000053",
            INIT_09 => X"0000004d00000038000000350000002e00000049000000230000004200000053",
            INIT_0A => X"000000220000000f0000000a0000000f0000000d00000026000000090000003f",
            INIT_0B => X"000000400000004b000000400000002c0000003b000000360000002900000038",
            INIT_0C => X"0000000e0000000a0000001d00000020000000120000000f000000080000001d",
            INIT_0D => X"0000001c00000045000000410000002600000030000000340000003000000028",
            INIT_0E => X"000000220000000d00000008000000170000000f000000160000001e00000010",
            INIT_0F => X"0000001200000015000000230000002200000023000000200000001d0000001f",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000008",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000003000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000040000000200000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000400000001",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000003",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE56;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE57 : if BRAM_NAME = "samplegold_layer0_instance57" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000200000007000000030000000900000026000000000000000000000000",
            INIT_09 => X"000000060000000a000000130000002300000000000000000000000600000000",
            INIT_0A => X"0000000b0000001200000019000000100000000d000000170000000200000003",
            INIT_0B => X"0000000a0000000c0000000c0000000f00000039000000000000000e0000000b",
            INIT_0C => X"000000110000000a000000060000002f0000001c000000170000000700000002",
            INIT_0D => X"000000070000000f000000140000001100000012000000250000000c00000000",
            INIT_0E => X"000000140000000a000000150000001700000028000000010000002d00000027",
            INIT_0F => X"00000018000000010000000f0000000c0000002200000029000000140000002e",
            INIT_10 => X"000000230000001500000000000000150000002100000030000000000000000d",
            INIT_11 => X"000000020000000e000000070000000b0000000000000017000000210000001b",
            INIT_12 => X"0000001b000000280000001d0000000e000000090000001d0000002400000004",
            INIT_13 => X"0000000e00000000000000090000000200000000000000000000001000000023",
            INIT_14 => X"00000021000000230000001a000000160000001f000000140000002400000014",
            INIT_15 => X"000000190000002a000000000000000a00000000000000000000000800000015",
            INIT_16 => X"00000009000000100000000d0000001c0000000e000000200000001800000016",
            INIT_17 => X"000000220000001b00000030000000180000000a000000000000000800000009",
            INIT_18 => X"000000000000001b000000000000000f00000008000000210000000800000024",
            INIT_19 => X"0000001c0000001f0000001d000000140000001a0000000d000000000000000f",
            INIT_1A => X"0000000c0000000c000000150000000a000000010000001d0000001300000016",
            INIT_1B => X"0000002100000021000000080000001c0000001d0000001a0000000300000005",
            INIT_1C => X"000000070000000c00000006000000120000001500000007000000040000000d",
            INIT_1D => X"000000130000001a0000001d0000000c0000001a0000001f0000002300000000",
            INIT_1E => X"0000000000000001000000020000000b000000140000000e0000001800000000",
            INIT_1F => X"00000000000000050000000f0000001b0000001c000000090000001c00000013",
            INIT_20 => X"0000000a000000000000000000000009000000050000000d0000000a0000000f",
            INIT_21 => X"0000000d0000000000000003000000060000000a000000270000000c0000001c",
            INIT_22 => X"0000001e0000000800000000000000000000001000000011000000030000000a",
            INIT_23 => X"0000000c000000080000000d0000000000000003000000000000000e00000012",
            INIT_24 => X"0000002800000025000000060000000000000014000000080000001100000005",
            INIT_25 => X"0000002000000019000000000000005800000037000000100000001e0000000e",
            INIT_26 => X"000000370000002f00000003000000000000000000000011000000230000001d",
            INIT_27 => X"000000270000002e0000002e00000000000000790000003a0000001a00000020",
            INIT_28 => X"0000002c0000008600000016000000010000000000000000000000110000002c",
            INIT_29 => X"0000003500000031000000350000001c000000000000000b0000003d00000017",
            INIT_2A => X"000000420000004b00000062000000020000004b000000000000000000000035",
            INIT_2B => X"0000004a0000001d0000006300000049000000000000003c0000000000000017",
            INIT_2C => X"0000001b0000006a0000005e0000003c000000000000005d0000003100000001",
            INIT_2D => X"0000002300000035000000090000006800000046000000090000001600000000",
            INIT_2E => X"00000002000000270000003a0000006500000044000000140000003f0000003e",
            INIT_2F => X"0000005000000022000000330000001f00000064000000440000000000000016",
            INIT_30 => X"000000140000001b0000004f000000100000006300000018000000310000001e",
            INIT_31 => X"000000000000007100000023000000410000003a0000004f0000003700000002",
            INIT_32 => X"00000011000000450000001f0000001f0000004d000000480000004100000054",
            INIT_33 => X"0000003f0000000a0000003c000000140000005a000000250000005900000014",
            INIT_34 => X"00000000000000340000003a0000003300000000000000780000004a0000003e",
            INIT_35 => X"000000440000002b0000003c0000003200000022000000490000000000000038",
            INIT_36 => X"000000340000000e0000001f00000050000000130000004b0000004f00000046",
            INIT_37 => X"00000014000000650000003700000036000000130000004f000000360000000a",
            INIT_38 => X"0000002d000000400000002800000016000000180000005f0000005c00000032",
            INIT_39 => X"0000003400000026000000500000005600000042000000000000005c00000032",
            INIT_3A => X"000000390000003600000042000000280000002e00000000000000610000004d",
            INIT_3B => X"000000500000003900000025000000100000007d0000003f0000000000000045",
            INIT_3C => X"000000400000003f0000002c0000002700000033000000290000000b00000044",
            INIT_3D => X"0000002100000040000000320000004600000029000000670000003000000000",
            INIT_3E => X"0000000000000030000000360000002100000000000000390000002200000012",
            INIT_3F => X"0000001900000000000000450000002700000052000000570000004c0000001c",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE57;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE58 : if BRAM_NAME = "samplegold_layer0_instance58" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000010000000000000000000000000000001e00000016000000280000001f",
            INIT_01 => X"00000029000000000000002b0000002c000000140000000d0000000000000004",
            INIT_02 => X"0000002500000000000000000000000000000001000000140000001a0000001f",
            INIT_03 => X"000000150000001a000000500000000700000002000000090000000000000013",
            INIT_04 => X"0000000e0000000a000000180000000000000000000000030000000b00000010",
            INIT_05 => X"0000001700000005000000000000003a00000000000000000000000000000000",
            INIT_06 => X"0000004e0000001200000000000000000000008d0000007d000000970000001f",
            INIT_07 => X"00000000000000010000001f0000000e000000000000000a0000000800000021",
            INIT_08 => X"0000000000000001000000000000000600000000000000120000005c00000034",
            INIT_09 => X"0000000800000000000000000000000b00000013000000000000000000000000",
            INIT_0A => X"00000027000000000000000000000000000000120000000a0000000000000005",
            INIT_0B => X"0000000000000000000000050000000e00000000000000000000000000000017",
            INIT_0C => X"0000000b00000018000000090000000700000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000002200000014000000000000000100000007",
            INIT_0E => X"0000000000000000000000000000002000000000000000000000001500000008",
            INIT_0F => X"0000002400000012000000000000000200000000000000000000000000000000",
            INIT_10 => X"000000120000000a000000000000000000000008000000310000003a00000008",
            INIT_11 => X"000000000000000e000000060000001c00000008000000000000000000000000",
            INIT_12 => X"0000002200000000000000000000001b0000004c000000180000000000000000",
            INIT_13 => X"00000000000000180000000e0000000000000002000000000000000000000010",
            INIT_14 => X"0000000000000009000000160000000000000000000000000000000000000000",
            INIT_15 => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000006000000000000000000000016000000000000000000000006",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000004000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000005400000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000005500000007000000060000000000000011000000030000000000000000",
            INIT_1D => X"00000007000000580000004e00000059000000670000005d000000530000005c",
            INIT_1E => X"0000003f000000400000000d00000008000000740000006f0000006e00000054",
            INIT_1F => X"000000490000000f000000470000004f000000410000003d000000450000001d",
            INIT_20 => X"0000000e0000004f000000180000000d0000000c0000006c000000660000005e",
            INIT_21 => X"0000003f0000003200000026000000170000003e0000003e0000003800000039",
            INIT_22 => X"0000002000000007000000550000002a00000001000000380000004600000040",
            INIT_23 => X"0000003c0000002d0000001d0000002200000015000000280000003800000031",
            INIT_24 => X"000000310000001d000000140000004f000000370000002c0000003a00000027",
            INIT_25 => X"0000003a0000004d000000360000002700000018000000140000002000000039",
            INIT_26 => X"0000002600000031000000220000001f000000450000003e000000350000003c",
            INIT_27 => X"00000046000000470000004c00000032000000210000001d000000140000001e",
            INIT_28 => X"000000210000000f000000340000001b00000031000000370000005b0000003e",
            INIT_29 => X"0000003e0000004a0000003e0000003300000031000000210000001a00000014",
            INIT_2A => X"0000002c00000014000000360000001800000020000000320000002000000066",
            INIT_2B => X"0000003f0000003a0000004c0000002a000000410000001b000000350000002f",
            INIT_2C => X"000000390000003b0000002d00000033000000280000001b0000001a00000032",
            INIT_2D => X"0000003000000030000000370000003d000000260000003b0000003d0000004f",
            INIT_2E => X"0000004300000048000000380000004a0000001a00000015000000290000002b",
            INIT_2F => X"0000002f000000320000001b000000430000003400000042000000490000003b",
            INIT_30 => X"0000003c0000003c00000031000000530000002e00000029000000240000003e",
            INIT_31 => X"0000003800000037000000290000001d00000041000000360000004600000043",
            INIT_32 => X"00000045000000340000003c00000035000000490000003d0000003300000030",
            INIT_33 => X"000000390000003e0000004d0000002600000025000000430000003a0000003c",
            INIT_34 => X"00000040000000320000003e0000003b00000036000000460000004600000041",
            INIT_35 => X"000000490000004800000046000000390000001f0000002c000000490000003e",
            INIT_36 => X"0000003b00000039000000310000003f0000003b00000039000000380000004c",
            INIT_37 => X"0000004b000000410000004c000000460000002e00000010000000380000003f",
            INIT_38 => X"0000007e0000000e000000350000003d000000380000003a0000003600000034",
            INIT_39 => X"00000000000000000000001b0000001500000024000000120000000c00000031",
            INIT_3A => X"00000049000000500000001100000014000000170000001a0000001d00000065",
            INIT_3B => X"0000006c0000000000000003000000160000001b000000050000000600000026",
            INIT_3C => X"0000002b00000067000000240000001200000012000000120000000900000004",
            INIT_3D => X"0000000b000000230000001a00000004000000260000000b0000000000000027",
            INIT_3E => X"0000003200000000000000430000004200000000000000000000000500000000",
            INIT_3F => X"0000000000000026000000000000004a00000018000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE58;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE59 : if BRAM_NAME = "samplegold_layer0_instance59" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000070000003c000000000000000000000019000000000000000800000000",
            INIT_01 => X"0000000000000000000000160000001b00000034000000190000000000000000",
            INIT_02 => X"00000000000000020000001f000000000000000000000002000000000000000c",
            INIT_03 => X"0000000000000000000000000000002300000019000000290000000d00000000",
            INIT_04 => X"000000280000000000000016000000000000000c000000000000000100000000",
            INIT_05 => X"00000000000000000000000000000000000000200000001b0000001000000000",
            INIT_06 => X"00000013000000000000000000000000000000000000004b0000000000000006",
            INIT_07 => X"000000090000000000000000000000000000000f0000002b0000000000000012",
            INIT_08 => X"000000000000003e00000000000000000000000000000000000000300000000b",
            INIT_09 => X"0000000700000000000000000000002700000000000000410000000000000005",
            INIT_0A => X"0000000000000024000000000000000000000000000000020000000500000000",
            INIT_0B => X"000000000000001500000000000000000000001b000000060000001e00000016",
            INIT_0C => X"0000001b0000001300000000000000000000000d0000001d0000000000000002",
            INIT_0D => X"00000000000000010000002500000000000000000000000f0000000000000011",
            INIT_0E => X"000000130000000a0000002f0000000000000000000000080000000f00000000",
            INIT_0F => X"0000002f00000000000000000000001500000000000000000000000000000000",
            INIT_10 => X"0000000d0000000c0000000b000000210000000000000000000000050000001c",
            INIT_11 => X"0000000000000022000000000000000500000016000000000000000000000007",
            INIT_12 => X"0000001500000027000000000000000f0000001b0000000a0000000000000006",
            INIT_13 => X"00000011000000000000000000000000000000130000000f0000000000000000",
            INIT_14 => X"0000000d000000120000001d0000000600000013000000130000002700000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000050000000000000001",
            INIT_16 => X"000000040000000f000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000300000000000000000000000000000000000000000000000c00000009",
            INIT_18 => X"000000000000000b000000110000000000000000000000000000000000000000",
            INIT_19 => X"00000000000000000000000d0000000500000001000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000018",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"000000000000000000000000000000000000000a000000030000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000c00000007",
            INIT_31 => X"00000002000000060000001200000003000000130000000b0000000000000000",
            INIT_32 => X"0000000000000003000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000e00000007000000210000000000000000000000160000001600000000",
            INIT_34 => X"00000000000000000000000a0000000000000000000000000000000000000010",
            INIT_35 => X"000000010000003b0000002b0000000f00000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000700000000000000000000000000000000000000000000001300000017",
            INIT_38 => X"000000080000000000000000000000000000000c000000150000000200000000",
            INIT_39 => X"0000000000000006000000000000000300000016000000110000000800000000",
            INIT_3A => X"0000000300000000000000070000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000001000000017",
            INIT_3C => X"0000000000000000000000000000001e00000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000f00000002",
            INIT_3E => X"00000010000000010000000b0000000900000010000000100000000500000000",
            INIT_3F => X"0000000000000012000000290000005f000000110000000b0000001400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE59;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE60 : if BRAM_NAME = "samplegold_layer0_instance60" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000200000000000000010000000000000000",
            INIT_01 => X"000000000000001a000000390000001500000000000000090000000900000009",
            INIT_02 => X"00000000000000000000001b0000001f00000000000000000000000000000000",
            INIT_03 => X"00000000000000000000000b00000007000000000000000d0000001c00000000",
            INIT_04 => X"00000018000000190000000f0000000300000000000000000000000000000000",
            INIT_05 => X"000000000000000000000000000000140000000c00000001000000000000000e",
            INIT_06 => X"00000000000000160000000b00000003000000000000002b000000100000000c",
            INIT_07 => X"00000000000000000000000900000000000000010000000a0000000b00000010",
            INIT_08 => X"00000011000000070000001800000021000000180000000f0000001700000010",
            INIT_09 => X"0000000800000002000000000000000400000005000000000000001b00000022",
            INIT_0A => X"0000000d0000000500000003000000130000001e000000170000001600000000",
            INIT_0B => X"0000000d000000040000000a0000000700000000000000170000000600000000",
            INIT_0C => X"0000000100000000000000050000000900000000000000190000002100000031",
            INIT_0D => X"0000005e000000620000006100000065000000620000000e0000000000000010",
            INIT_0E => X"0000006b0000006e0000006e000000750000004c000000230000006200000064",
            INIT_0F => X"0000007f0000007d0000006c000000880000006b0000005f0000000000000000",
            INIT_10 => X"000000000000008100000087000000910000009d0000005c0000005500000088",
            INIT_11 => X"00000080000000760000005d00000087000000ae0000005f0000004900000000",
            INIT_12 => X"0000000a00000000000000a6000000b1000000b6000000b80000008b00000070",
            INIT_13 => X"0000006e000000530000004f00000062000000ab000000b00000007600000057",
            INIT_14 => X"000000a1000000730000008e000000c3000000c3000000ca000000c0000000b1",
            INIT_15 => X"000000aa00000071000000600000006d000000a2000000b40000009000000071",
            INIT_16 => X"0000007d000000ac000000a2000000a8000000a7000000b4000000da000000cb",
            INIT_17 => X"000000d80000009800000072000000690000006900000096000000aa00000098",
            INIT_18 => X"0000008a0000009100000088000000a0000000a900000098000000bb000000e3",
            INIT_19 => X"000000e5000000cb000000990000008b000000870000007b0000009000000097",
            INIT_1A => X"0000009f000000a80000009500000070000000a3000000a9000000a3000000da",
            INIT_1B => X"000000e1000000e0000000ae00000097000000840000009400000072000000a3",
            INIT_1C => X"0000009c000000b2000000c2000000870000009300000091000000a7000000ca",
            INIT_1D => X"000000bb000000b700000080000000470000008d00000075000000660000008d",
            INIT_1E => X"000000a6000000cd000000cb000000b4000000a7000000af00000096000000b8",
            INIT_1F => X"000000c4000000760000006e0000005c0000006b0000007a0000007d00000062",
            INIT_20 => X"000000b1000000b2000000a80000009e000000b3000000af000000ba000000a6",
            INIT_21 => X"000000ae000000c000000065000000720000007c0000006d0000006b0000007a",
            INIT_22 => X"0000006e0000009d000000a0000000960000009d000000be000000ca000000b2",
            INIT_23 => X"000000ad000000a9000000b70000005d00000071000000890000007800000060",
            INIT_24 => X"00000067000000630000008d000000990000009e00000063000000ae000000c8",
            INIT_25 => X"000000cc0000009c00000095000000ae0000006000000072000000760000006d",
            INIT_26 => X"0000005f0000005d000000500000006b0000007a0000008300000069000000af",
            INIT_27 => X"000000b5000000c700000083000000900000009f0000006d0000005500000056",
            INIT_28 => X"000000520000005e00000056000000430000004f00000064000000730000009b",
            INIT_29 => X"0000000000000001000000000000000000000000000000000000006700000053",
            INIT_2A => X"000000000000000000000000000000000000002d000000000000000000000000",
            INIT_2B => X"0000000000000012000000000000000000000000000000050000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000002c0000002c000000100000000000000000000000000000000500000000",
            INIT_2E => X"000000000000000000000000000000000000000000000000000000000000002b",
            INIT_2F => X"0000000000000000000000000000000000000000000000210000000000000000",
            INIT_30 => X"0000000000000000000000000000001100000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000180000000000000000000000000000001100000000",
            INIT_32 => X"0000000000000000000000000000000400000013000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000017000000060000000000000000",
            INIT_34 => X"0000000000000036000000000000000000000001000000000000000000000000",
            INIT_35 => X"00000000000000000000000000000000000000000000000a000000000000000b",
            INIT_36 => X"000000000000000000000011000000000000000c000000000000000000000000",
            INIT_37 => X"0000000000000043000000100000000700000000000000130000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000070000000000000015",
            INIT_39 => X"0000002d000000430000000100000000000000000000000a0000000000000000",
            INIT_3A => X"000000000000001e0000000c0000000000000000000000000000000000000000",
            INIT_3B => X"0000002b00000000000000000000000000000020000000000000000000000000",
            INIT_3C => X"0000000600000000000000180000000000000000000000000000001100000000",
            INIT_3D => X"0000000000000009000000070000000000000000000000000000002d00000000",
            INIT_3E => X"0000000400000000000000000000000000000007000000000000000000000000",
            INIT_3F => X"000000070000000100000000000000000000000000000004000000000000000f",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE60;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE61 : if BRAM_NAME = "samplegold_layer0_instance61" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000d000000180000000e0000000000000021000000290000000000000000",
            INIT_01 => X"000000000000000e000000070000000000000000000000220000000300000000",
            INIT_02 => X"00000000000000080000001a000000110000001b000000000000000000000000",
            INIT_03 => X"0000000000000014000000000000001900000000000000000000000a00000000",
            INIT_04 => X"0000000000000000000000000000001c00000006000000250000001400000000",
            INIT_05 => X"0000000000000000000000000000004900000013000000030000000000000000",
            INIT_06 => X"00000000000000000000002e0000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000800000038000000140000000000000000",
            INIT_08 => X"0000000000000000000000000000003a00000000000000000000000000000000",
            INIT_09 => X"00000003000000000000001d0000000000000027000000220000001200000000",
            INIT_0A => X"000000000000000000000000000000000000001700000000000000000000000e",
            INIT_0B => X"0000000000000000000000000000002b00000000000000190000001a00000000",
            INIT_0C => X"0000000000000004000000000000000000000013000000000000002c00000005",
            INIT_0D => X"0000000d00000000000000000000000900000030000000000000000000000001",
            INIT_0E => X"00000000000000000000000800000000000000000000000f0000000a00000024",
            INIT_0F => X"0000001d00000007000000000000000000000005000000130000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000001800000012",
            INIT_11 => X"0000001200000016000000000000001000000000000000150000000300000000",
            INIT_12 => X"0000001a00000000000000000000000000000000000000000000000000000014",
            INIT_13 => X"0000001600000000000000050000000700000000000000000000000500000000",
            INIT_14 => X"0000000000000010000000000000000000000000000000000000000000000009",
            INIT_15 => X"0000002b00000000000000000000000000000018000000000000000000000000",
            INIT_16 => X"0000000e0000000d000000000000000000000000000000000000001300000000",
            INIT_17 => X"0000000000000000000000000000000000000001000000000000000000000005",
            INIT_18 => X"000000170000000000000000000000000000000d000000000000000000000009",
            INIT_19 => X"000000000000000000000000000000000000000000000000000000000000000c",
            INIT_1A => X"00000000000000000000000000000000000000000000001e0000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000080000000000000000",
            INIT_1C => X"0000000000000000000000010000000500000000000000040000001400000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000800000013",
            INIT_1F => X"0000000c00000000000000000000000000000008000000000000000000000000",
            INIT_20 => X"0000000000000005000000000000000000000000000000000000000000000018",
            INIT_21 => X"0000000f000000440000007b0000001400000000000000000000000000000000",
            INIT_22 => X"00000036000000620000000000000001000000260000001c000000240000001b",
            INIT_23 => X"0000001d000000160000006200000053000000160000001b0000002300000021",
            INIT_24 => X"00000019000000240000009c00000000000000150000002c0000002400000010",
            INIT_25 => X"000000000000003900000028000000800000002e00000014000000170000001c",
            INIT_26 => X"000000210000001a000000270000006100000013000000020000002600000006",
            INIT_27 => X"00000002000000000000004700000000000000910000004f000000050000001b",
            INIT_28 => X"000000290000000c0000001a0000004800000027000000530000001c00000000",
            INIT_29 => X"0000000000000000000000120000005700000000000000290000005600000006",
            INIT_2A => X"0000001b0000003e000000000000001a00000053000000370000003900000020",
            INIT_2B => X"000000280000000000000000000000110000003e000000000000001a00000029",
            INIT_2C => X"0000001d0000001c0000002a000000000000001d000000560000003300000039",
            INIT_2D => X"0000002d000000100000001e00000000000000150000000f0000002d00000000",
            INIT_2E => X"0000000000000021000000120000000c00000011000000240000005800000030",
            INIT_2F => X"0000001c0000001d000000210000001b0000000000000019000000070000005f",
            INIT_30 => X"00000042000000040000001f0000000000000024000000140000003d00000034",
            INIT_31 => X"0000000400000022000000010000003b00000000000000080000001e00000012",
            INIT_32 => X"000000200000001500000028000000240000000c0000004f0000000a00000048",
            INIT_33 => X"0000002500000019000000000000003100000009000000000000000d00000014",
            INIT_34 => X"000000000000001d0000001800000033000000070000001c000000320000001a",
            INIT_35 => X"00000000000000230000002c0000000f00000000000000000000001800000032",
            INIT_36 => X"00000031000000000000000d000000160000004c000000000000002200000017",
            INIT_37 => X"0000000200000007000000260000001300000043000000000000000c00000017",
            INIT_38 => X"0000000f00000030000000000000000000000019000000420000000d0000001c",
            INIT_39 => X"00000013000000110000000b000000150000000e000000330000000000000000",
            INIT_3A => X"000000000000000c0000000b000000270000000000000029000000410000000f",
            INIT_3B => X"0000001d0000000c000000200000002f00000000000000150000002a00000000",
            INIT_3C => X"0000002e00000000000000140000000000000006000000050000003b0000002f",
            INIT_3D => X"0000000000000000000000020000001b0000002c0000000b0000001f0000001b",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000200000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE61;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE62 : if BRAM_NAME = "samplegold_layer0_instance62" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000e000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"00000000000000000000000000000037000000730000005e0000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000009",
            INIT_05 => X"0000000000000000000000000000000000000000000000020000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000001b0000002b000000290000003000000025000000250000002c0000002a",
            INIT_1B => X"0000001d00000000000000000000003d0000003b0000003c0000003600000000",
            INIT_1C => X"000000020000001600000032000000290000001e000000230000001800000016",
            INIT_1D => X"0000001e0000000000000000000000000000003c0000003a0000003900000033",
            INIT_1E => X"0000002100000025000000000000001b000000120000000d0000002800000015",
            INIT_1F => X"000000120000002e0000001f000000000000000b00000034000000310000002e",
            INIT_20 => X"000000360000001e000000240000000200000005000000190000001c0000001c",
            INIT_21 => X"0000001b0000000f000000210000002800000022000000200000001e00000039",
            INIT_22 => X"0000003000000030000000310000001300000001000000030000001b00000024",
            INIT_23 => X"00000024000000200000001d0000001d0000002b000000230000002700000020",
            INIT_24 => X"0000002200000032000000330000002600000013000000060000001000000002",
            INIT_25 => X"000000000000002100000004000000200000002300000030000000230000002b",
            INIT_26 => X"0000002b0000002900000033000000320000002b0000000c0000000f00000021",
            INIT_27 => X"0000000a000000250000000c000000230000002a0000001e0000003800000023",
            INIT_28 => X"000000170000002f0000001b0000003c00000028000000180000002600000012",
            INIT_29 => X"000000160000000900000022000000220000002a0000001c0000002e00000024",
            INIT_2A => X"0000002b0000001f0000002a000000160000001b0000000f0000002000000024",
            INIT_2B => X"0000002c000000160000002a0000001c0000001b000000240000002300000026",
            INIT_2C => X"0000002b000000180000002a000000280000002200000028000000160000001b",
            INIT_2D => X"000000200000000800000036000000230000001d000000170000003000000027",
            INIT_2E => X"000000360000002a000000180000002a000000270000001b0000001d00000024",
            INIT_2F => X"0000001f0000001e000000130000001e0000002c000000260000002a00000021",
            INIT_30 => X"000000060000003a000000270000001900000025000000260000001800000021",
            INIT_31 => X"000000100000001d000000150000001500000016000000260000002700000027",
            INIT_32 => X"00000032000000230000002b0000002200000011000000230000002600000019",
            INIT_33 => X"000000160000000b000000110000001200000014000000060000001b00000021",
            INIT_34 => X"000000190000001e0000002f000000230000001b000000100000001b00000019",
            INIT_35 => X"0000001600000015000000150000000f000000130000000f0000000100000017",
            INIT_36 => X"00000018000000060000001000000000000000100000000d0000000000000000",
            INIT_37 => X"00000000000000140000000b0000000a0000000600000003000000000000004b",
            INIT_38 => X"0000002f0000000c00000000000000000000001f000000000000000000000000",
            INIT_39 => X"00000000000000090000001500000008000000080000000c0000000700000000",
            INIT_3A => X"000000000000000000000000000000000000000e0000002e0000000000000001",
            INIT_3B => X"0000002d0000000000000000000000510000000b000000020000000200000000",
            INIT_3C => X"00000000000000000000000000000000000000230000001c0000000000000000",
            INIT_3D => X"000000000000003500000011000000090000001f000000000000001900000000",
            INIT_3E => X"0000000100000000000000000000000000000000000000250000000900000000",
            INIT_3F => X"00000000000000000000001900000013000000090000000f0000000700000034",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE62;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE63 : if BRAM_NAME = "samplegold_layer0_instance63" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003500000008000000000000000000000000000000010000000700000012",
            INIT_01 => X"0000001a000000000000000e00000000000000290000000a0000001b00000027",
            INIT_02 => X"0000002f00000010000000000000000000000000000000000000001300000000",
            INIT_03 => X"0000001500000000000000020000001300000000000000240000000300000026",
            INIT_04 => X"0000003600000000000000160000000000000000000000090000000600000000",
            INIT_05 => X"00000000000000210000000f0000000000000000000000000000000000000007",
            INIT_06 => X"0000001500000024000000000000000000000000000000210000000100000007",
            INIT_07 => X"000000000000002a000000020000000000000000000000000000000000000000",
            INIT_08 => X"000000000000002a00000011000000030000001400000000000000000000001d",
            INIT_09 => X"000000000000002a000000010000000000000000000000240000000000000002",
            INIT_0A => X"00000000000000000000002a000000110000000d0000000f0000000000000000",
            INIT_0B => X"0000000600000000000000220000000a00000000000000000000000000000005",
            INIT_0C => X"0000002100000000000000000000002900000019000000110000001100000000",
            INIT_0D => X"000000080000000500000000000000140000000e000000010000000000000000",
            INIT_0E => X"000000000000001400000000000000000000002f0000001e0000000c00000000",
            INIT_0F => X"0000000000000014000000050000000100000009000000110000000500000016",
            INIT_10 => X"0000001900000018000000050000000000000015000000200000001a00000000",
            INIT_11 => X"00000000000000080000000c0000000300000006000000000000001e00000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"000000000000000000000000000000000000000f000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000001500000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"000000250000001e000000190000001200000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000015",
            INIT_32 => X"000000180000000100000000000000090000001b000000000000000000000000",
            INIT_33 => X"000000000000000000000000000000000000000000000000000000000000001e",
            INIT_34 => X"00000000000000080000001c0000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000003",
            INIT_36 => X"0000000a00000016000000180000001d0000001d000000240000001a0000000d",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000002800000029000000280000003000000028000000160000001f00000035",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"000000180000000d000000090000000d0000000e000000150000001a00000012",
            INIT_3B => X"0000002100000022000000000000000000000000000000000000000000000003",
            INIT_3C => X"00000029000000450000002f0000001f000000330000002a0000001000000018",
            INIT_3D => X"00000000000000000000000a0000001700000000000000000000000000000000",
            INIT_3E => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"000000120000002a000000170000002700000000000000110000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE63;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE64 : if BRAM_NAME = "samplegold_layer0_instance64" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000150000001e000000160000002d0000002c0000002700000029",
            INIT_01 => X"0000002f00000000000000000000001700000005000000000000000000000000",
            INIT_02 => X"0000000000000000000000060000000000000003000000060000001400000009",
            INIT_03 => X"000000050000000f0000001a000000310000000900000000000000000000000b",
            INIT_04 => X"0000000000000000000000040000001a000000320000000b0000000000000000",
            INIT_05 => X"00000000000000000000000d0000000b00000006000000000000000000000003",
            INIT_06 => X"000000000000000000000000000000000000000a0000000c0000000100000000",
            INIT_07 => X"0000000400000026000000350000000000000000000000000000000000000005",
            INIT_08 => X"0000000a0000000a00000000000000040000000a000000160000000a00000000",
            INIT_09 => X"000000000000000e000000180000000d00000005000000000000000000000000",
            INIT_0A => X"000000280000001d000000120000002500000022000000220000000c0000000c",
            INIT_0B => X"00000019000000160000001e000000190000001c000000270000002b00000023",
            INIT_0C => X"0000002b0000002c0000001f0000000b000000230000002b0000002b00000009",
            INIT_0D => X"00000015000000040000001c000000240000000f0000000f0000002200000021",
            INIT_0E => X"0000004a0000005100000050000000480000000c0000001f0000002e0000002d",
            INIT_0F => X"0000002d0000000f000000000000001b000000270000002b0000003e00000048",
            INIT_10 => X"0000004d0000004d000000420000004a000000600000000e0000002800000028",
            INIT_11 => X"000000270000002c0000000800000011000000190000002c0000003400000054",
            INIT_12 => X"0000004e00000051000000500000003a0000004d0000004f000000180000001b",
            INIT_13 => X"0000002200000020000000320000002f000000180000002b000000440000003e",
            INIT_14 => X"00000040000000470000003d000000420000004c000000460000003f00000020",
            INIT_15 => X"000000220000002400000015000000340000002e0000002c0000004300000035",
            INIT_16 => X"0000003500000025000000370000004a0000003e0000003e0000004d0000004a",
            INIT_17 => X"000000340000001b000000310000000b000000210000002c0000002c00000031",
            INIT_18 => X"0000002f0000001e00000028000000200000002200000033000000400000002f",
            INIT_19 => X"000000380000003800000003000000330000000a0000002a0000004700000043",
            INIT_1A => X"0000004300000051000000330000002300000047000000400000001f0000002a",
            INIT_1B => X"0000002b0000001d000000290000000d0000001a000000070000002300000048",
            INIT_1C => X"0000005700000020000000320000002e0000002b0000003d0000001f00000045",
            INIT_1D => X"000000240000003700000025000000190000001300000023000000000000002f",
            INIT_1E => X"000000340000004e0000003c000000300000003e00000032000000320000002f",
            INIT_1F => X"0000003e0000000000000026000000150000000d000000310000002000000000",
            INIT_20 => X"000000200000003c000000530000001e00000000000000340000002700000013",
            INIT_21 => X"0000004e00000020000000110000000b0000000d00000014000000290000003d",
            INIT_22 => X"0000002700000032000000450000005b000000200000000a0000000e0000002c",
            INIT_23 => X"000000330000002d00000022000000190000000f000000050000002500000020",
            INIT_24 => X"0000001b0000002b0000003a0000003e000000530000002d0000000600000008",
            INIT_25 => X"00000014000000320000002a0000002000000019000000140000001000000020",
            INIT_26 => X"0000003d00000060000000550000003a0000004600000062000000250000000b",
            INIT_27 => X"00000052000000390000004a0000004c000000340000002b000000330000003a",
            INIT_28 => X"000000490000005a00000099000000740000004d000000500000004000000035",
            INIT_29 => X"0000005d000000440000002f00000036000000380000004f0000005600000046",
            INIT_2A => X"000000460000004500000025000000c700000075000000520000005300000016",
            INIT_2B => X"000000000000005e0000005d0000003500000000000000320000004b0000005b",
            INIT_2C => X"0000006c000000930000005600000012000000da000000560000006300000052",
            INIT_2D => X"0000004d0000002d000000650000004c000000100000004d000000550000006a",
            INIT_2E => X"0000005e0000005e0000007c0000004b0000002d000000ab000000860000006c",
            INIT_2F => X"0000008300000031000000300000006700000035000000100000007300000055",
            INIT_30 => X"00000048000000590000005d000000680000004500000018000000b500000071",
            INIT_31 => X"0000004a00000080000000360000005100000054000000010000001f00000051",
            INIT_32 => X"0000005e000000690000004b0000005e0000007d0000005c0000003a0000006e",
            INIT_33 => X"0000008d00000000000000800000005f0000004300000031000000250000001f",
            INIT_34 => X"0000003a0000004d0000003600000047000000630000003c0000004e00000057",
            INIT_35 => X"0000001e000000830000000e0000008700000062000000000000001e00000006",
            INIT_36 => X"0000000800000023000000610000000c00000019000000520000004900000041",
            INIT_37 => X"00000049000000180000005500000025000000af000000690000000000000056",
            INIT_38 => X"000000670000004f000000460000005c0000003a00000069000000040000001e",
            INIT_39 => X"000000060000000b000000310000004400000031000000bd0000005500000000",
            INIT_3A => X"000000000000002b0000005a00000005000000390000004e0000000000000071",
            INIT_3B => X"000000690000000900000019000000690000003c00000002000000d100000068",
            INIT_3C => X"000000570000000000000027000000850000004a000000410000004e00000000",
            INIT_3D => X"00000000000000100000001c0000004b000000600000005e0000002900000093",
            INIT_3E => X"0000007a00000050000000000000000000000056000000ba0000006000000000",
            INIT_3F => X"000000060000000a0000000d0000001500000068000000460000006600000080",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE64;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE65 : if BRAM_NAME = "samplegold_layer0_instance65" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000080000000610000006600000000000000000000003f000000bf00000028",
            INIT_01 => X"000000220000001e000000190000001d00000020000000460000003d00000063",
            INIT_02 => X"0000000000000017000000210000001c00000000000000000000004200000077",
            INIT_03 => X"0000000000000004000000070000003000000061000000360000001d00000000",
            INIT_04 => X"0000000000000000000000020000000d0000000d000000130000002e00000026",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000003200000000000000010000000000000000000000000000000100000000",
            INIT_07 => X"00000000000000000000000a00000000000000000000000e0000003d0000003a",
            INIT_08 => X"0000000700000000000000120000000000000000000000000000000000000000",
            INIT_09 => X"000000000000002a0000000000000000000000020000001d0000000600000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"000000000000006a000000210000000c00000007000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000020000000600000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"00000000000000040000000000000000000000000000004a0000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000020",
            INIT_11 => X"00000000000000090000000d0000001f00000000000000000000000000000000",
            INIT_12 => X"000000bd000000ab000000b5000000b80000003a000000060000000500000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000002e000000a0",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000f00000001000000000000000000000000",
            INIT_16 => X"0000001f000000000000001e0000000000000004000000000000001c0000002e",
            INIT_17 => X"00000000000000000000001f0000004300000000000000000000000000000007",
            INIT_18 => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_19 => X"00000000000000000000001a0000000a000000000000006b0000005300000000",
            INIT_1A => X"000000060000001d00000000000000000000003a0000005b0000006200000000",
            INIT_1B => X"0000001a00000014000000130000000400000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000700000000000000000000000000000000",
            INIT_1D => X"00000000000000040000000f0000001100000000000000000000000000000002",
            INIT_1E => X"00000027000000220000001d0000001b000000000000000c0000000000000000",
            INIT_1F => X"000000290000001b000000140000000c000000060000000d0000001b00000032",
            INIT_20 => X"00000028000000250000001700000016000000220000002a000000200000001b",
            INIT_21 => X"0000001f0000001f000000040000000000000000000000000000000000000000",
            INIT_22 => X"00000000000000310000001d0000001700000017000000220000003a00000024",
            INIT_23 => X"000000390000001b000000000000000000000000000000000000000000000000",
            INIT_24 => X"00000000000000000000001c000000160000001e00000017000000240000003c",
            INIT_25 => X"0000003d0000001b0000000c0000000000000000000000000000000000000000",
            INIT_26 => X"00000000000000000000000000000000000000220000001f0000001500000034",
            INIT_27 => X"00000024000000200000000b0000000000000000000000000000000000000000",
            INIT_28 => X"00000000000000000000000000000000000000030000000a0000002900000011",
            INIT_29 => X"0000001d00000017000000160000000000000000000000000000000000000000",
            INIT_2A => X"000000000000000000000000000000000000000000000000000000210000002d",
            INIT_2B => X"0000003800000033000000040000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000002f00000000",
            INIT_2D => X"00000014000000270000002c0000000000000000000000000000000000000000",
            INIT_2E => X"000000000000000000000000000000000000000000000000000000000000001a",
            INIT_2F => X"0000000f000000020000003a0000001f00000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000400000000000000070000002700000018000000000000000000000000",
            INIT_32 => X"0000000f00000000000000000000000000000000000000190000000000000000",
            INIT_33 => X"000000040000000d000000000000000000000033000000040000000000000000",
            INIT_34 => X"00000000000000040000000b0000000000000000000000000000000000000000",
            INIT_35 => X"000000000000000f000000000000000000000005000000000000000000000000",
            INIT_36 => X"0000000000000000000000090000001800000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000700000015000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_3B => X"000000000000000000000007000000050000000d000000020000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"00000000000000080000000f0000000a00000014000000120000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000008000000000000000000000009",
            INIT_3F => X"000000020000003e0000001900000006000000000000000e0000000c00000022",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE65;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE66 : if BRAM_NAME = "samplegold_layer0_instance66" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004a000000000000000000000000000000000000001a0000000000000000",
            INIT_01 => X"000000000000002d000000000000000d00000000000000000000000000000019",
            INIT_02 => X"000000160000002a000000000000000000000000000000000000000000000000",
            INIT_03 => X"000000000000000b0000003c000000000000000c0000000c0000000a00000000",
            INIT_04 => X"00000007000000110000002b0000000000000000000000000000001700000005",
            INIT_05 => X"0000000000000000000000390000001b0000000f000000130000000400000008",
            INIT_06 => X"00000005000000000000000f0000001900000000000000080000000000000019",
            INIT_07 => X"0000000100000003000000240000002a0000002d00000000000000060000001f",
            INIT_08 => X"0000000e00000004000000120000000000000006000000000000004a00000000",
            INIT_09 => X"000000000000000000000050000000330000002e000000160000000c0000000f",
            INIT_0A => X"000000270000001c00000000000000050000001f0000002a0000000000000035",
            INIT_0B => X"0000002300000000000000000000005b0000000f0000002f0000000900000000",
            INIT_0C => X"000000000000001c000000000000004f0000001f000000000000002500000000",
            INIT_0D => X"000000000000000a00000000000000010000008100000000000000130000000a",
            INIT_0E => X"000000290000000a0000000000000039000000000000002b000000290000000d",
            INIT_0F => X"0000000000000009000000340000000000000000000000630000002000000000",
            INIT_10 => X"0000000000000019000000080000000000000065000000000000003500000019",
            INIT_11 => X"0000000000000000000000000000001d00000000000000060000008500000018",
            INIT_12 => X"000000290000000000000000000000000000006a0000002d0000001a00000011",
            INIT_13 => X"000000120000000000000007000000000000000000000000000000110000007a",
            INIT_14 => X"000000650000003e0000000000000000000000230000002e0000002d0000001f",
            INIT_15 => X"000000140000000e000000000000000900000000000000000000000000000000",
            INIT_16 => X"000000000000007200000032000000000000000000000027000000200000001b",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_25 => X"0000000000000000000000000000000d0000000d000000030000001b00000014",
            INIT_26 => X"00000000000000000000000000000000000000000000002a0000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000600000000000000030000000000000007",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"00000000000000000000000700000000000000000000000e0000000700000000",
            INIT_2B => X"0000000000000009000000010000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000022000000150000000700000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000001200000012",
            INIT_2E => X"00000006000000000000000000000000000000010000000a0000000c00000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000003",
            INIT_30 => X"000000000000000f000000000000000000000000000000000000000000000003",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_33 => X"000000000000000000000005000000120000000e000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000003000000000000000500000000",
            INIT_35 => X"00000066000000630000004a0000004100000041000000460000000f00000000",
            INIT_36 => X"000000030000000200000000000000060000000800000000000000170000003e",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000017",
            INIT_38 => X"0000000600000004000000010000000c0000001300000007000000000000000b",
            INIT_39 => X"00000000000000020000000200000014000000120000002e0000001100000031",
            INIT_3A => X"0000003d0000004100000009000000050000000400000000000000010000001b",
            INIT_3B => X"0000000600000009000000130000001600000012000000310000001400000009",
            INIT_3C => X"000000130000000c0000000b0000002400000016000000000000000000000001",
            INIT_3D => X"000000000000000100000029000000020000001b0000001f0000000800000004",
            INIT_3E => X"00000014000000000000000b0000002100000033000000090000000100000002",
            INIT_3F => X"000000530000003e000000260000002600000040000000240000001300000028",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE66;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE67 : if BRAM_NAME = "samplegold_layer0_instance67" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000160000001a0000000e00000037000000280000000e",
            INIT_01 => X"0000000a0000000e00000029000000410000002200000029000000360000000b",
            INIT_02 => X"000000000000001a000000340000000000000051000000000000001b00000008",
            INIT_03 => X"00000007000000180000000f0000000000000000000000000000000000000000",
            INIT_04 => X"0000001f00000030000000070000000a0000001e00000008000000350000001d",
            INIT_05 => X"000000220000000e000000000000001c000000340000001b0000002700000014",
            INIT_06 => X"0000000000000000000000000000000000000010000000000000000400000000",
            INIT_07 => X"000000230000002d0000001c0000000000000000000000000000000000000000",
            INIT_08 => X"0000000a0000003e0000002a000000390000002f000000010000000000000000",
            INIT_09 => X"0000000e00000000000000000000000f00000000000000220000003600000036",
            INIT_0A => X"0000000e00000002000000000000000000000000000000060000000000000000",
            INIT_0B => X"0000000e0000001f000000090000001f00000006000000000000000000000013",
            INIT_0C => X"0000000b00000026000000290000001b0000000a000000000000000000000003",
            INIT_0D => X"000000090000000b0000001d0000000400000009000000170000000000000000",
            INIT_0E => X"0000000000000000000000290000001100000000000000000000000000000000",
            INIT_0F => X"000000a9000000a2000000b0000000a8000000d6000000cb000000d500000000",
            INIT_10 => X"000000b0000000b3000000c7000000e0000000d7000000e2000000cf000000af",
            INIT_11 => X"000000ca000000b2000000b5000000a8000000a5000000ee000000f0000000f2",
            INIT_12 => X"000000fb000000cd000000c3000000e1000000da000000d8000000d7000000e1",
            INIT_13 => X"0000008c000000880000008d0000008e0000008c0000008a000000ef000000fc",
            INIT_14 => X"000000f8000000fa000000b7000000b1000000ce000000de000000bb0000008d",
            INIT_15 => X"000000b9000000be000000c9000000c0000000d2000000ab000000ae000000dd",
            INIT_16 => X"000000cb000000f7000000f80000008d000000ae000000d5000000de0000009b",
            INIT_17 => X"000000c9000000c1000000be000000b5000000c4000000ad000000a1000000a8",
            INIT_18 => X"00000078000000b0000000ef000000eb000000ab000000d9000000e1000000bf",
            INIT_19 => X"000000ac000000b10000009e0000009800000096000000930000009800000078",
            INIT_1A => X"0000006a0000008500000097000000c1000000c6000000fb000000fc000000e8",
            INIT_1B => X"000000cc0000008e00000078000000970000008400000076000000990000008a",
            INIT_1C => X"000000690000008800000081000000870000007b000000b2000000ff000000f2",
            INIT_1D => X"000000920000007a000000520000004d00000055000000560000005b00000066",
            INIT_1E => X"0000007b00000075000000700000006c0000006f00000062000000aa000000e9",
            INIT_1F => X"000000c100000088000000540000003000000050000000410000003800000055",
            INIT_20 => X"0000007e000000530000004f00000052000000300000007200000064000000c2",
            INIT_21 => X"000000c90000009800000077000000ad0000009a000000a00000009b0000009d",
            INIT_22 => X"0000006e000000350000004f000000400000001d0000003d000000390000006f",
            INIT_23 => X"00000060000000cb0000007b0000007400000057000000700000006400000063",
            INIT_24 => X"00000081000000470000004b0000004b000000140000001d000000560000005d",
            INIT_25 => X"0000003e0000007c000000c20000007d0000005d000000500000008c0000007a",
            INIT_26 => X"0000009c000000850000001c0000000f000000080000000d0000004700000086",
            INIT_27 => X"0000007d00000089000000bd000000bb000000690000002e0000001d00000083",
            INIT_28 => X"00000090000000ac000000730000002b0000001100000005000000250000005b",
            INIT_29 => X"000000500000005800000092000000ad000000be0000007b0000002c00000016",
            INIT_2A => X"0000000c0000007900000067000000460000002b000000200000001800000031",
            INIT_2B => X"00000000000000000000001e000000000000000000000000000000830000002d",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"00000054000000310000003d0000005200000001000000000000000000000000",
            INIT_2E => X"00000000000000110000000000000000000000080000001c0000004700000069",
            INIT_2F => X"000000000000000000000000000000000000003a000000010000000000000000",
            INIT_30 => X"00000000000000020000001c0000001600000000000000000000002900000000",
            INIT_31 => X"00000000000000000000001900000000000000000000003d0000000500000000",
            INIT_32 => X"00000000000000000000001a0000000000000000000000000000002900000000",
            INIT_33 => X"000000040000000300000000000000160000002300000000000000310000005d",
            INIT_34 => X"000000000000001b000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000001b0000000c0000001c0000001a0000001800000000000000190000003e",
            INIT_36 => X"000000000000002c000000360000000a00000000000000000000000000000003",
            INIT_37 => X"000000240000001e000000040000000000000000000000000000000e00000000",
            INIT_38 => X"000000210000001d000000000000006500000013000000000000002900000047",
            INIT_39 => X"000000140000003a000000310000002400000038000000320000001e0000000e",
            INIT_3A => X"00000000000000000000006e000000000000001300000000000000000000001c",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"00000037000000170000001c0000000e00000013000000540000000000000000",
            INIT_3D => X"000000000000003d000000250000003600000046000000390000003a00000009",
            INIT_3E => X"0000004800000000000000000000002000000000000000030000001e00000000",
            INIT_3F => X"0000000f00000000000000000000004300000000000000000000001300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE67;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE68 : if BRAM_NAME = "samplegold_layer0_instance68" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001400000014000000530000001f0000001000000000000000000000006f",
            INIT_01 => X"0000000000000000000000000000004800000037000000380000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000010000000000000000200000000",
            INIT_03 => X"00000009000000160000000000000000000000000000002b0000000000000000",
            INIT_04 => X"0000001d00000043000000000000000000000000000000040000000000000009",
            INIT_05 => X"0000002d00000004000000000000000e0000000000000000000000080000003b",
            INIT_06 => X"000000030000001a000000050000000000000000000000000000000000000002",
            INIT_07 => X"000000040000000000000000000000010000000000000000000000000000000f",
            INIT_08 => X"0000000000000004000000000000000000000006000000000000000000000000",
            INIT_09 => X"0000003a00000024000000000000000000000004000000040000000000000000",
            INIT_0A => X"00000000000000010000000c00000007000000190000002e0000002f00000037",
            INIT_0B => X"00000044000000420000004f00000000000000000000000b0000000a0000000a",
            INIT_0C => X"0000001400000000000000000000000b00000030000000430000004200000039",
            INIT_0D => X"0000004d0000002a00000031000000610000000000000008000000060000000a",
            INIT_0E => X"0000000c0000000000000000000000000000002b0000002f0000004200000043",
            INIT_0F => X"0000005000000054000000390000005c0000005f000000030000000a00000000",
            INIT_10 => X"000000000000001b000000000000000000000010000000350000003300000051",
            INIT_11 => X"0000005a00000051000000520000004500000052000000610000000000000000",
            INIT_12 => X"0000001300000000000000190000000b000000090000003f0000005300000054",
            INIT_13 => X"0000002500000038000000480000003b0000003d000000450000003e00000002",
            INIT_14 => X"00000000000000290000000000000000000000150000002e0000004200000046",
            INIT_15 => X"0000004700000038000000480000004300000032000000420000003900000043",
            INIT_16 => X"00000042000000000000002e00000000000000000000004d0000005a00000065",
            INIT_17 => X"0000002e0000000000000000000000110000000a00000004000000220000002c",
            INIT_18 => X"0000002700000048000000030000002900000000000000000000005b0000002d",
            INIT_19 => X"0000001f0000003c00000040000000380000004b000000270000005a0000004a",
            INIT_1A => X"0000003b0000003d00000022000000140000001700000000000000090000007c",
            INIT_1B => X"00000062000000380000002000000045000000380000002c0000005800000016",
            INIT_1C => X"00000007000000560000002e0000000000000014000000350000000000000015",
            INIT_1D => X"0000002d0000008200000040000000000000003000000020000000140000005d",
            INIT_1E => X"00000033000000260000001d00000003000000060000001e0000002000000000",
            INIT_1F => X"0000001b0000002d0000007b000000330000000800000000000000000000004b",
            INIT_20 => X"000000530000002f00000022000000180000000000000025000000160000000f",
            INIT_21 => X"0000000c0000002b0000002f00000074000000460000000a0000000000000043",
            INIT_22 => X"00000045000000350000002a0000001f000000180000000f0000002700000011",
            INIT_23 => X"000000000000001000000020000000170000007d0000003e0000000600000008",
            INIT_24 => X"0000001e0000001b0000001d0000004200000044000000250000001c00000015",
            INIT_25 => X"0000000000000000000000020000001700000015000000080000002d00000005",
            INIT_26 => X"0000001800000031000000140000001d0000000e000000000000000000000009",
            INIT_27 => X"0000000a00000013000000000000000000000013000000110000003900000001",
            INIT_28 => X"00000000000000090000002c0000004700000015000000000000000000000000",
            INIT_29 => X"00000000000000140000005500000000000000000000000a0000001000000043",
            INIT_2A => X"0000001f00000004000000010000003d00000022000000030000000000000000",
            INIT_2B => X"00000000000000000000000d0000003100000000000000000000000200000014",
            INIT_2C => X"000000230000001f000000000000002d00000048000000000000000000000003",
            INIT_2D => X"0000000000000000000000000000000000000015000000000000000000000000",
            INIT_2E => X"000000000000001f00000013000000100000004f000000210000000000000007",
            INIT_2F => X"000000080000000f000000000000000000000000000000120000000000000000",
            INIT_30 => X"00000032000000000000000200000026000000140000002e0000002a00000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"00000000000000540000000000000000000000600000001a0000001e0000000e",
            INIT_33 => X"00000026000000020000003c0000003000000000000000060000001700000028",
            INIT_34 => X"0000002000000000000000210000000000000000000000640000001100000051",
            INIT_35 => X"00000000000000000000000000000000000000000000002a0000000c00000000",
            INIT_36 => X"0000001100000000000000000000001900000000000000000000007700000000",
            INIT_37 => X"0000002600000000000000260000000000000000000000270000000000000023",
            INIT_38 => X"0000002a00000017000000000000001a0000002000000000000000000000005a",
            INIT_39 => X"0000006600000012000000000000002e00000014000000000000006900000000",
            INIT_3A => X"000000170000001100000000000000000000000a000000270000000000000000",
            INIT_3B => X"0000000d0000007a0000001f00000000000000000000001d0000009400000020",
            INIT_3C => X"0000003100000021000000140000000000000000000000000000000000000000",
            INIT_3D => X"00000000000000000000005b0000003f0000000000000000000000020000003b",
            INIT_3E => X"0000001800000016000000130000000d00000000000000050000000000000000",
            INIT_3F => X"000000000000000000000000000000790000003100000000000000000000001c",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE68;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE69 : if BRAM_NAME = "samplegold_layer0_instance69" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000700000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000050000000700000006",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000001a00000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000006a0000007a000000830000002400000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000005400000088",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_14 => X"00000000000000000000001a0000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000006000000000000000000000026000000200000000000000000",
            INIT_17 => X"000000000000000000000000000000000000000a000000350000000000000000",
            INIT_18 => X"0000000c0000000e000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000002000000060000000000000000000000000000000000000000",
            INIT_1B => X"0000002c00000027000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000002b00000034000000250000001a0000001800000017000000200000002d",
            INIT_1D => X"0000003a00000031000000300000001e0000002a00000026000000270000002f",
            INIT_1E => X"0000001b0000000e000000100000000600000000000000020000000f0000001c",
            INIT_1F => X"000000220000002e000000300000002f0000001c0000002a0000002b0000002a",
            INIT_20 => X"0000002e00000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"000000000000001b0000001e000000360000002f000000140000002800000036",
            INIT_22 => X"000000220000000f000000150000000000000000000000000000001300000000",
            INIT_23 => X"00000000000000000000000000000022000000360000002e0000002600000032",
            INIT_24 => X"0000002f0000002a0000000b0000000000000000000000000000000000000000",
            INIT_25 => X"000000000000000000000000000000070000000b0000003a0000002300000024",
            INIT_26 => X"00000030000000300000000d0000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000130000002500000029",
            INIT_28 => X"000000310000002a000000080000000c00000000000000000000000000000000",
            INIT_29 => X"00000000000000000000000000000000000000000000002f0000000000000012",
            INIT_2A => X"000000090000002c000000070000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000019",
            INIT_2C => X"000000000000000f00000027000000000000000100000006000000000000000d",
            INIT_2D => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000001000000070000002200000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"000000000000000000000000000000080000001e000000000000000000000000",
            INIT_31 => X"0000000000000012000000000000000000000000000000000000000000000000",
            INIT_32 => X"00000000000000000000000a0000000400000000000000070000000000000000",
            INIT_33 => X"00000000000000000000002a0000002300000000000000000000000000000000",
            INIT_34 => X"00000000000000000000000000000006000000000000000f0000000c00000000",
            INIT_35 => X"0000000000000000000000000000001500000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000060000000000000004",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"00000000000000000000000000000000000000000000001a0000000000000001",
            INIT_39 => X"0000000000000000000000150000001400000009000000000000000900000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000002f00000008",
            INIT_3B => X"000000000000000000000000000000000000001f000000000000000000000000",
            INIT_3C => X"000000000000000000000000000000000000000000000000000000000000004a",
            INIT_3D => X"0000003d000000000000000000000000000000000000001d0000000f00000000",
            INIT_3E => X"0000000000000001000000000000000000000000000000010000000000000000",
            INIT_3F => X"0000000000000004000000170000000000000000000000190000002300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE69;


    MEM_SAMPLEGOLD_LAYER0_INSTANCE70 : if BRAM_NAME = "samplegold_layer0_instance70" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000310000000000000006000000000000000000000006",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000070000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000026000000000000002000000000",
            INIT_06 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"000000000000000000000000000000000000000000000026000000000000002a",
            INIT_08 => X"00000049000000000000000000000000000000000000000f0000001900000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_0A => X"0000000a0000003f000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000002000000000000003500000000000000000000000e00000003",
            INIT_0C => X"0000000000000000000000510000000000000000000000000000001c00000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000b00000032",
            INIT_0E => X"0000000800000000000000100000000700000000000000000000000000000015",
            INIT_0F => X"0000002600000038000000050000000000000000000000010000000c0000002c",
            INIT_10 => X"0000002200000000000000000000000100000000000000000000000000000000",
            INIT_11 => X"000000000000001300000028000000000000000000000000000000020000000e",
            INIT_12 => X"0000000c00000009000000000000001300000003000000000000000000000000",
            INIT_13 => X"0000000000000000000000240000000000000000000000000000000000000004",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYER0_INSTANCE70;

    MEM_EMPTY_18Kb : if BRAM_NAME = "default" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 36, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 36, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST"      -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate;


end a1;