library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 4000000) of integer;

  constant input_wght : mem := (
    -- bias
    -12555, 5187, 421, -594, 6712, -7672, 9532, 3569, -7946, 2656,

    -- weights
    -- filter=0 channel=0
    -2, -4, -11, -10, -7, -4, -9, -2, -5, -5, -4, -4, -9, -10, -8, -4, -11, -6, -10, -10, -7, -4, -11, -4, -9, -10, -5, -5, -2, -9, -5, -7, -1, -1, -4, -1, -5, -7, -1, -2, -5, -7, -8, -2, -1, -4, -9, -3, -9, -5, -10, -3, -8, -10, -1, -5, -8, -3, -3, -8, -6, -8, -7, -7, -5, -3, -5, -9, -5, -1, -7, -9, -8, -8, -7, -3, 0, -6, 0, -7, -1, -7, -8, -8, -8, -6, -1, 0, 0, -8, -2, -7, -7, -7, -9, 0, -6, -7, -5, -8, -3, -2, -7, -3, -9, -9, -10, -5, -1, -5, -8, -4, -9, -5, -4, -8, -9, -6, -7, -1, -7, -1, -2, -5, -3, -8, -8, -3, -4, -6, -2, -1, -8, -9, -4, -5, -5, -4, -4, -5, -1, -1, -1, -7, -1, -1, -9, -2, -5, 0, 0, 0, -5, -5, -3, -5, -4, -1, -2, 0, -3, 0, -8, 0, -2, -7, -6, -6, -4, -3, -4, -3, -3, -3, 0, -5, -3, -5, -9, -3, -2, 0, -6, -3, -6, -5, -6, -2, 0, -7, 0, -3, -5, -2, 0, -7, -5, -2, 0, -4, -1, -6, -7, 0, 0, -4, -2, -4, -4, -3, -1, -6, -6, -1, -6, -7, 0, -1, -8, -4, -4, -5, -6, -2, 0, -4, 0, -4, -1, -3, 0, 0, 0, 0, -6, -8, -6, -6, -2, -6, -10, -10, -3, -3, -3, -2, -6, -4, -6, -2, 0, -1, -9, -2, -1, 0, 1, -4, -3, -1, 0, -2, -6, -3, 0, -3, -5, -1, -6, -4, -8, -9, -7, -6, -10, -5, -6, -4, -10, -7, -1, -1, -4, 0, -1, -5, -4, 1, -3, -2, -4, -7, -3, -3, -4, -3, 1, -5, -3, -4, -6, -8, -5, -3, -12, -6, -3, -7, -9, -10, -7, -8, -7, -9, -7, -5, -8, -2, -3, 2, -2, -1, -3, -7, -6, 0, -7, -5, -7, -5, -7, -3, -11, -4, -4, -10, -5, -4, -9, -3, -9, -6, -1, -8, -2, -4, -6, -4, -7, -4, -2, -1, -5, -3, 0, -4, -4, -7, -8, -8, -2, -8, -3, -8, -7, -6, -6, -7, -13, -4, -5, -9, -4, -3, -8, -5, -2, -7, -3, -9, -10, -4, 0, 0, 3, 1, -3, -4, -8, -7, -10, -9, -9, -6, -9, -12, -10, -9, -14, -14, -13, -10, -10, -11, -5, -3, -8, -4, -9, -9, -2, -2, -6, -3, -5, 3, 0, -4, -2, -2, 1, -4, -5, -7, -4, -4, -13, -14, -9, -14, -17, -13, -13, -15, -12, -7, -4, -6, -5, -2, -8, -3, -2, -1, -2, 0, -4, 1, 0, -2, -1, -3, -2, -7, -3, -7, -9, -10, -9, -9, -14, -12, -12, -17, -11, -9, -14, -11, -13, -6, -10, -9, -7, -3, -2, -3, -3, 0, -3, 1, -3, -2, -2, -2, 0, -4, -1, -6, -9, -11, -11, -14, -15, -11, -13, -14, -15, -12, -15, -5, -6, -9, -5, -7, -9, -10, -8, 1, 0, -5, 2, 0, 0, 2, 1, -3, -5, -1, -5, -3, -11, -10, -7, -6, -8, -10, -15, -16, -17, -17, -16, -8, -10, -6, -8, -5, -12, -7, -5, 1, 3, -4, 0, 0, 0, 1, -1, 2, -1, -4, -7, -3, -8, -6, -11, -11, -16, -14, -20, -14, -17, -21, -15, -11, -9, -5, -8, -10, -6, -8, -1, 0, -4, -3, 1, -6, 0, -4, -2, 3, 1, 0, -4, -2, -4, -12, -7, -9, -11, -12, -16, -16, -18, -23, -16, -11, -11, -11, -12, -11, -8, -2, 0, 2, -5, -5, 1, 1, -5, -2, -2, 3, 0, 1, -5, 0, -5, -10, -12, -16, -17, -17, -14, -14, -19, -15, -18, -11, -9, -4, -10, -4, -9, 0, 1, 0, -6, -1, -4, -3, -4, 3, -1, 0, -3, -1, 1, -1, -8, -12, -11, -7, -8, -12, -13, -17, -14, -21, -10, -13, -6, -5, -3, -1, -7, -6, -4, -3, -3, 1, -5, 0, -6, 0, 0, -3, 3, 4, -3, -5, -2, -8, -10, -11, -5, -9, -13, -12, -12, -18, -12, -8, -8, -12, -3, -7, 1, 1, -1, -2, -2, -3, -7, -7, -3, -5, -3, -2, 2, 0, -4, -3, 0, -7, -5, -3, -5, -11, -7, -8, -9, -12, -8, -4, -7, -4, -3, -6, -4, -3, 1, 0, 0, -5, -5, -4, -2, 0, -2, 3, -3, 0, 1, -1, 0, -7, -7, -5, -10, -7, -9, -8, -4, -3, -7, -7, -7, -4, -6, -6, -4, -5, 3, 0, 2, -5, -3, 0, -2, -7, 1, 0, -2, 0, 1, -1, -5, 0, -6, -2, -7, -9, -3, -7, -5, 0, -5, -2, 0, -5, -4, 0, -3, 1, -4, 3, -2, 1, -2, -6, -2, -3, 0, 1, -1, -5, -2, -4, 3, -4, 1, 0, -7, -7, -6, -1, -6, -5, 0, -2, 0, 1, -6, 1, 0, 2, -4, -4, 0, -4, -1, -5, -5, 0, 0, -5, 0, -5, -4, 3, 1, 1, -1, -3, -5, -4, -3, -4, -1, 1, -3, -3, -2, -2, -6, -1, 2, 1, 0, 0, -3, 1, 0, -6, -2, -7, -4, 0, 0, -5, 0, 0, 1, -3, 2, 0, -1, -4, -1, -6, -4, -2, -4, -1, 0, 0, -3, 0, 1, 0, -3, -4, -1, -1, -6, 0, -7, -8, 0, 1, 1, 0, 3, 0, -1, 0, 2, -2, 0, 0, 2, 1, -2, 5, -2, 3, -5, -3, 1, -6, 0, -4, -2, -1, -1, -3, -6, -6, -8, -4, -4, -4, -5, 0, 2, -3, -2, -3, 0, 0, -3, -1, 0, 1, 2, 0, -3, -2, -1, 0, -1, -4, 1, -4, 0, 0, -4, -8, -9, -8, -4, 0, -4, 0, -5, -1, 1, 0, 0, -3, 2, 1, 2, 0, 0, 2, 3, 0, -4, -2, -2, 0, -5, 0, -2, -2, -3, 0, -7, -3, -1, 0, -9, -6, -7, -5, -5, -6, -8, 0, -6, -5, -8, 0, -5, -5, -1, -1, 0, 0, -1, -2, -6, -6, -7, -3, -6, -1, -2, -2, -4, -9, -2, -9, -2, -1, -9, -7, -4, -5, -1, -1, -4, -6, -3, -1, -4, -4, -8, -4, -6, -4, -6, -10, -4, -8, -4, -1, -6, -6, -6, -8, -7, -9, -4, -7, -1, -1, -7, -3, 0, -6, -1, -4, -8, -8, -8, -5, 1, -2, -3, -1, -3, -2, -1, -1, -1, 0, -3, -8, -3, -8, -8, -1, -6, -6, -3, 0, -3, -7, -9, -3, -7, -1, -3, -1, -6, -1, -7, -2, -1, -4, -5, 1, -3, 0, 0, -6, 0, 1, 2, 0, -3, 0, 0, -1, -8, -2, -2, 0, -6, -5, -8, -7, -8, 0, -3, 0, -3, -6, -2, -6, -4, -4, -5, 1, 1, 0, 0, 0, -3, -5, -3, 0, -4, -2, 0, -5, -8, -6, -6, 0, -6, 1, 0, -4, -9, -1, 0, -2, -5, 2, -2, -2, 0, 0, 0, -3, -2, 2, -1, 2, -2, 1, -4, -4, -5, -1, -2, 0, -4, -6, -5, -1, -1, -7, 0, 1, -7, -1, -2, -1, -5, -5, 2, -2, 5, 1, -3, -1, -4, 0, -1, 3, 4, 0, -5, -2, -5, 0, 0, -2, -5, 0, 1, -3, -2, -6, 0, 0, -3, 0, -1, 4, -1, -2, 2, -1, 5, 1, -1, 2, 4, -3, 3, 3, 4, 4, 1, 0, 4, -2, -4, -5, 0, -2, -6, 0, -4, -6, -1, -5, -5, -4, 0, 0, 4, 3, -4, 4, 2, 0, 4, 4, -4, 3, -1, 4, 2, 3, -1, 0, -3, 0, 2, -2, 1, -4, -3, 0, -3, -4, -6, -2, -2, -3, 2, 0, 1, 0, -3, -2, 0, 0, 1, 0, 1, 4, 2, 3, -1, -2, -3, -3, 0, 2, 0, 0, -7, -5, 0, 1, -5, 1, -2, 0, -2, 0, 1, -1, 2, 0, 3, -1, 3, -1, -2, 0, 0, 4, -3, -1, 4, 0, -4, 1, -3, 0, -1, -7, -1, 0, 1, 2, -4, 2, -1, -5, -7, -7, -4, -1, -3, 0, 3, 4, -2, 1, 0, 0, -2, -3, 5, -1, 4, 3, -2, -1, 0, -3, -5, -3, -6, -5, -3, -1, -2, -3, 0, -6, -4, -2, -5, -4, -2, 4, 1, -1, 0, -3, 0, -4, -2, 2, 0, -1, 0, 0, 3, 1, 2, -4, -2, -3, -9, -3, 0, 2, -2, -2, -3, -4, -1, -7, -7, 0, -3, 0, 1, -4, -7, 0, -6, -1, -7, 0, 0, -3, 0, 2, 1, -1, -2, -7, -5, -6, -5, -7, -3, 2, 4, -2, -3, -4, -1, -5, -3, -1, -3, -1, -2, 0, -6, -3, 0, -4, 0, 0, -4, -1, 1, -6, -3, 0, -1, -5, -6, -8, -5, -2, 4, -1, 0, -2, 3, 0, -2, -6, 0, -2, -8, 1, -2, -7, -4, -1, -1, 0, -5, 1, 2, 0, -1, -4, 3, 1, -4, -4, -5, -3, -7, 0, -5, -2, 0, 4, 0, 1, -3, -6, -1, 0, -6, -2, 0, -3, -7, -4, -4, -7, -5, -10, -1, -4, 1, -3, -3, -3, -3, 1, -2, 0, -6, -1, -5, -4, -2, 3, 3, 0, 1, -4, -6, 0, -3, 2, -3, -3, -3, -10, -4, -4, -11, -11, 0, -1, 0, -1, 0, -2, -3, -4, -3, -1, 3, -1, 0, 2, 3, -2, -1, 4, 0, 1, 2, 3, -5, -5, -2, -5, -5, -4, -8, -6, -10, -8, -8, -8, 0, 0, 0, 0, -4, -3, 3, -1, 2, 2, -3, 1, -4, -2, 0, 2, -1, 4, 2, -1, -3, -4, 0, -4, 0, -9, -8, -8, -6, -14, -7, -3, -6, 0, 0, -3, -2, 0, 0, 5, 4, 2, -5, -4, -2, -2, -2, 2, 2, 7, 3, 1, -4, -4, -1, -7, -5, -2, -7, -13, -9, -7, -6, -2, -4, -3, 2, 2, 1, 0, 0, 2, 6, 1, -2, -5, -4, 3, 2, 2, 5, 1, 7, 5, -2, 3, 0, -3, -5, -7, -7, -11, -9, -5, -9, -6, -4, -4, 0, -1, 5, 3, 8, 5, 1, -1, 2, 0, 0, 0, 6, 6, 6, 5, 4, 1, -1, 0, 0, -1, 0, -3, -5, -6, -3, -3, -2, 0, 1, 4, 5, 3, 1, 8, 10, 9, 4, -1, 0, -6, -1, -1, -1, 7, 8, 2, 2, 5, 5, 1, 1, 0, 3, -1, 1, -3, -3, -2, 0, -3, 0, 0, 2, 0, 1, 0, 6, 2, 8, 5, -4, -5, -2, -1, 4, -1, 0, 1, 2, 3, 0, 4, 4, 5, 3, 0, 6, 3, 3, -3, -2, 0, -2, -1, 0, 7, 6, 7, 1, 1, 4, 0, -2, -3, -3, 0, -3, -3, 1, -1, 7, -1, 2, 4, 3, 2, 1, 4, 3, 4, 1, 2, 5, -1, 3, 1, 1, 5, 7, 3, 0, 2, 0, 1, -3, -3, -2, -8, -1, 1, 0, 2, 4, 0, 3, 3, 6, 5, 1, -1, 4, 0, 5, 7, 2, 2, 0, 0, 0, 0, 5, 2, 2, -2, 2, -2, -4, -5, -7, -7, -1, 0, -2, -5, 0, 6, 2, 0, 0, 5, 1, -2, 4, 3, 3, 2, 3, 5, 4, 2, 5, 3, 4, -2, 0, 2, 3, -3, -1, -4, -6, -3, -5, -6, 0, -4, 5, 0, 6, 1, 2, 1, 0, 5, 3, 4, 4, 0, 7, 0, 1, 0, 0, -1, -1, -4, -3, -1, 0, -3, -4, -11, -3, -7, -5, -6, -1, 1, -1, -1, 3, 3, 1, 2, 7, 6, 0, 1, 2, 7, 7, 0, 2, 0, 1, 2, -1, -3, -3, -6, -6, -8, -11, -7, -12, -5, -9, -5, -2, -5, 0, 1, 1, 4, -1, 4, 1, 3, -1, 0, 5, -1, 1, -3, 0, -1, -4, -3, -3, 0, -4, -1, -7, -3, -3, -4, -10, -4, -5, -7, -5, -4, 0, -2, 0, -1, -6, 1, 0, 3, 4, -2, 4, 1, 2, -4, -1, 0, 0, -2, 1, -3, -7, -10, -6, -6, -12, -11, -8, -3, -11, -5, -6, -7, -8, -4, -6, -3, -7, -3, -6, 0, -7, 0, -2, -6, -4, -7, -5, -3, -2, 0, -6, -3, -9, -6, -3, -7, -6, -10, 7, 4, 8, 8, 6, 3, 5, 8, 2, 3, 7, 5, 6, 8, 8, 6, 6, 4, 7, 6, 4, 1, 0, 3, 1, 5, 0, 4, 5, 3, 2, 7, 6, 9, 6, 9, 2, 7, 5, 4, 3, 8, 11, 9, 4, 4, 10, 7, 6, 10, 8, 4, 2, 5, 3, 2, 4, 2, 11, 4, 1, 2, 6, 9, 5, 6, 3, 6, 8, 9, 6, 8, 4, 7, 3, 6, 5, 4, 10, 7, 5, 4, 7, 4, 3, 5, 12, 9, 9, 8, 10, 11, 3, 9, 10, 8, 8, 8, 2, 7, 3, 11, 5, 8, 13, 12, 9, 6, 7, 11, 10, 9, 5, 7, 12, 9, 12, 12, 13, 7, 12, 8, 11, 10, 10, 10, 4, 4, 6, 4, 2, 4, 4, 3, 5, 5, 11, 10, 5, 5, 5, 12, 11, 10, 8, 12, 5, 11, 5, 8, 13, 10, 5, 5, 5, 4, 10, 5, 8, 5, 9, 3, 10, 10, 10, 10, 8, 11, 7, 13, 8, 10, 8, 9, 8, 8, 13, 7, 6, 9, 15, 13, 11, 12, 7, 7, 7, 10, 7, 7, 11, 14, 13, 6, 7, 7, 9, 6, 9, 14, 6, 15, 6, 9, 11, 15, 9, 9, 12, 13, 9, 11, 9, 10, 9, 11, 8, 11, 5, 11, 4, 7, 11, 10, 14, 13, 11, 6, 5, 6, 8, 11, 12, 10, 12, 11, 8, 13, 6, 13, 7, 11, 13, 8, 13, 12, 5, 7, 12, 7, 7, 12, 8, 5, 15, 13, 8, 5, 9, 7, 1, 5, 8, 6, 12, 12, 11, 11, 8, 11, 12, 12, 9, 13, 13, 9, 10, 12, 6, 10, 7, 12, 10, 9, 5, 6, 15, 9, 7, 7, 10, 2, 6, 6, 11, 5, 11, 9, 9, 6, 11, 13, 10, 14, 10, 11, 7, 6, 11, 6, 9, 10, 5, 12, 3, 6, 10, 8, 11, 16, 6, 6, 2, 4, 7, 8, 3, 9, 12, 8, 4, 9, 9, 5, 8, 6, 9, 14, 12, 13, 10, 12, 9, 12, 4, 5, 9, 3, 4, 4, 15, 10, 14, 8, 6, 2, 7, 0, 6, 9, 12, 10, 7, 7, 2, 8, 3, 6, 5, 8, 6, 11, 7, 8, 5, 11, 7, 2, 7, 0, 4, 3, 6, 17, 10, 7, 8, 8, 5, 6, 5, 8, 5, 6, 5, 3, 4, 7, 6, 2, 0, 7, 0, 6, 5, 5, 1, 5, 5, 6, 0, 7, 1, 10, 11, 15, 11, 12, 6, 9, 2, 4, 5, 7, 2, 1, 1, 3, 2, 2, 2, 0, 0, 0, 3, 1, 3, -1, 4, 9, 6, 3, -2, 7, 5, 8, 9, 13, 11, 11, 13, 3, 3, 4, 1, 6, 1, 2, 4, 3, 2, -3, -3, 2, -3, 3, -1, 5, 5, 1, 4, 1, 3, 2, -2, 3, 4, 9, 9, 14, 16, 13, 11, 7, 7, 0, 3, 6, -1, 0, 2, -4, -5, 0, -6, -6, -5, -5, -5, 2, -1, 6, 1, 5, -1, 5, 5, 6, 1, 6, 8, 15, 8, 11, 9, 4, 8, 2, 7, 4, 5, 3, 6, -1, 0, -1, -8, -6, -7, -7, 0, 0, 0, 3, 5, -1, 1, 4, 7, 7, 5, 13, 7, 12, 10, 8, 12, 5, 5, 9, 2, 3, 6, 4, -1, 0, -3, -10, -3, -8, -5, -9, -7, 0, -3, 6, 3, 3, 3, 3, 10, 5, 5, 13, 11, 6, 9, 13, 10, 13, 7, 8, 5, 12, 1, 4, -2, 3, -1, -3, -7, -5, -5, -3, -3, -1, 5, 3, 2, 10, 6, 12, 13, 10, 12, 8, 10, 8, 11, 6, 8, 12, 13, 8, 8, 8, 4, 0, 5, 2, -2, 0, -5, -5, -4, -6, -7, 4, 5, 5, 4, 9, 7, 7, 8, 11, 14, 7, 5, 13, 11, 9, 13, 12, 11, 9, 13, 7, 4, 7, 8, 6, 5, -3, 1, -8, -3, -5, 0, 3, 4, 4, 7, 11, 14, 9, 11, 11, 10, 11, 11, 3, 3, 11, 15, 9, 13, 13, 15, 8, 9, 4, 6, 2, 10, 2, 3, 2, 1, 0, -1, 8, 6, 11, 9, 9, 18, 13, 18, 19, 17, 12, 4, 3, 6, 8, 9, 16, 13, 16, 15, 10, 8, 14, 11, 7, 3, 11, 5, 4, 0, 8, 7, 9, 10, 10, 9, 9, 12, 14, 19, 18, 14, 9, 11, 2, 2, 4, 7, 10, 14, 11, 9, 9, 13, 13, 15, 10, 11, 7, 10, 13, 5, 9, 6, 8, 13, 11, 8, 12, 17, 19, 16, 16, 10, 10, 11, 2, 7, 10, 7, 14, 8, 11, 16, 8, 10, 14, 10, 7, 9, 7, 7, 14, 8, 11, 9, 13, 13, 10, 16, 9, 16, 14, 14, 16, 7, 9, 3, 6, 6, 9, 8, 11, 11, 12, 9, 9, 10, 15, 11, 9, 7, 12, 9, 11, 11, 17, 13, 10, 15, 14, 9, 13, 14, 7, 10, 7, 14, 3, 8, 6, 4, 5, 1, 8, 8, 7, 8, 12, 11, 17, 13, 14, 15, 8, 12, 16, 8, 12, 13, 11, 12, 12, 11, 15, 10, 13, 14, 8, 13, 7, 2, 6, -2, 4, 3, 2, 6, 13, 7, 13, 17, 7, 8, 10, 16, 11, 8, 8, 12, 11, 15, 16, 11, 15, 11, 11, 12, 6, 10, 10, 7, 8, 2, 5, -3, 0, 6, 2, 6, 6, 8, 8, 8, 8, 11, 11, 14, 9, 13, 9, 13, 11, 12, 12, 12, 9, 7, 9, 10, 5, 8, 3, 7, 3, 4, 2, 0, 5, 0, 4, 10, 9, 10, 7, 13, 9, 6, 15, 8, 12, 13, 14, 16, 11, 8, 14, 5, 6, 4, 8, 7, 6, 1, 2, 3, -2, -1, -1, 1, -4, 3, 2, 8, 8, 4, 9, 7, 10, 11, 8, 9, 8, 11, 12, 10, 6, 13, 10, 10, 9, 3, 11, 10, 5, 5, 6, 0, -1, -1, -2, -3, -3, 1, 1, 0, 3, 0, 5, 7, 3, 3, 2, 8, 4, 3, 9, 3, 4, 5, 0, 8, 7, 3, 6, 0, 1, -1, 0, 2, -1, -1, 1,
    -- filter=0 channel=1
    0, 1, 6, 4, 1, 8, 1, 7, 6, 6, 4, 5, 9, 6, 7, 3, 8, 8, 8, 8, 4, 5, 6, 8, 4, 7, 9, 4, 3, 8, 4, 6, 0, 5, 8, 3, 6, 3, 2, 5, 2, 3, 3, 10, 6, 3, 6, 1, 1, 6, 5, 5, 2, 7, 7, 3, 2, 2, 3, 8, 8, 6, 4, -2, -2, 2, 1, 7, 7, 7, 1, 7, 7, 5, 10, 8, 5, 0, 7, 7, 5, 2, 0, 5, 3, 9, 1, 3, 1, 8, 8, 5, 5, 6, 7, 0, -5, 1, 3, 1, -2, 5, 3, 3, 4, 5, 7, 6, 2, 1, 3, 2, 4, 6, 0, 2, 3, 7, 1, 8, 0, 1, 3, 5, 5, -1, 4, -1, 1, 5, 1, 3, -1, 6, 6, 1, 4, 4, 3, 0, 4, 0, 2, 5, 0, -2, 0, 7, 4, 2, 6, 4, 4, 2, 1, 2, 7, 6, 2, 0, -1, -1, 2, 3, -1, -1, -2, -2, 0, 3, 0, 5, -3, 0, 0, -5, 1, -1, -3, 4, 2, -2, 5, 0, 5, 0, -2, -2, 2, -1, 0, 0, 5, -1, 6, 0, 3, -1, 1, -4, 3, 0, -3, -2, -5, -4, -1, -8, -5, -4, -7, -5, -4, -3, -3, 0, -3, 2, 2, 0, 3, -1, 0, 1, 1, 6, 3, 2, 4, -2, 3, -4, 0, -1, -7, -8, -2, -7, -8, -3, -5, -6, -10, -7, -9, -6, 0, 0, -1, 0, 2, -2, 2, -2, 4, 2, 4, 5, 5, 5, -1, -4, -6, 0, -7, -6, -6, -13, -10, -13, -12, -10, -7, -13, -7, -9, -11, -7, -10, -2, -2, 0, -6, 4, 1, 5, 0, 3, -1, 0, 9, 8, 1, 2, -2, 0, -2, -8, -8, -9, -8, -16, -16, -17, -16, -15, -9, -7, -7, -6, -9, -3, -6, -6, -1, -1, 7, 2, 2, 2, 0, 0, 9, 2, 0, -3, 1, -5, -4, -7, -5, -11, -7, -11, -16, -13, -10, -9, -14, -13, -6, -8, -3, -1, 0, -2, 0, 2, 9, 5, 3, -2, 3, 7, 9, 2, 4, 0, 1, 1, -2, -4, -7, -3, -7, -12, -10, -7, -3, -7, -3, -2, -8, -3, -3, -2, 4, 0, 2, 8, 6, 2, 6, 0, 6, 2, 10, 3, 9, 5, 6, 9, 5, 2, 2, -1, -6, -2, -4, -6, -1, 0, -1, -4, 0, -3, -2, 1, 3, 11, 11, 10, 11, 10, 7, 3, 6, 1, 8, 7, 4, 6, 13, 9, 10, 7, 7, 2, 1, 3, 4, 0, 6, 4, 4, 4, 5, 5, 2, 4, 4, 7, 5, 8, 5, 8, 7, 1, 0, 3, 2, 10, 7, 13, 16, 9, 11, 9, 12, 13, 4, 5, 9, 12, 5, 9, 8, 4, 9, 11, 8, 10, 13, 7, 9, 5, 5, 10, 3, 4, 2, 6, 0, 5, 6, 12, 12, 14, 13, 16, 12, 6, 7, 11, 10, 7, 14, 14, 11, 6, 9, 9, 12, 12, 7, 11, 13, 8, 4, 3, 9, 3, 6, 5, 4, 9, 8, 13, 5, 15, 15, 10, 7, 7, 11, 13, 12, 10, 8, 5, 8, 9, 9, 6, 5, 4, 4, 8, 7, 4, 3, 0, 3, 7, 2, 4, 3, 5, 1, 0, 2, 7, 8, 11, 5, 3, 9, 11, 7, 3, 6, 7, 4, 9, 5, 6, 5, 0, 3, 3, 1, 2, 5, 4, 1, 4, 11, 1, 5, 0, -4, 2, -3, -1, 1, 4, 5, 8, 2, 6, 4, 0, 5, 2, -1, 2, 0, 0, -2, 4, 4, 0, -1, 0, -2, 1, 1, 2, 6, 2, 4, 0, -7, -5, 1, 2, -4, 2, 0, 1, 3, 5, -1, -2, -2, 4, 1, 5, 3, 2, 3, 1, 0, -5, -4, -4, -4, 4, 8, 4, 13, 10, -1, 1, -1, -5, -3, -3, 0, -3, -2, 1, 2, 2, -2, -1, 0, -5, -4, -4, -4, -3, -7, -3, -7, -10, -8, -2, -5, -3, 5, 12, 15, 5, 1, -1, -1, -2, -1, -7, -6, -6, -3, 0, 0, -6, -9, -6, 0, -7, -7, -1, 0, -7, -7, -7, -3, -11, -11, -7, -6, -1, 7, 13, 9, 11, 1, 0, -9, -7, -5, -7, -7, -5, -3, -8, 0, 0, -7, -4, -5, -5, -1, 0, -7, -9, -7, -9, -12, -8, -4, -10, 0, 5, 2, 10, 17, 3, 0, 1, -8, -6, -2, -9, -8, -6, -12, -4, -5, -2, -12, -11, -4, -6, -10, -7, -3, -10, -8, -13, -12, -9, -5, -7, -4, 2, 4, 11, 14, 6, 0, 0, -7, -11, -12, -9, -11, -8, -9, -10, -5, -13, -5, -5, -13, -11, -9, -12, -14, -14, -16, -13, -7, -14, -5, -7, -4, 0, 8, 10, 18, 8, 6, -1, -2, -5, -3, -7, -14, -8, -6, -12, -14, -14, -13, -14, -11, -8, -15, -14, -10, -16, -12, -8, -12, -7, -6, -8, 0, 4, 11, 13, 12, 7, 3, -6, -9, -6, -7, -12, -6, -6, -11, -12, -11, -14, -14, -13, -11, -14, -16, -11, -16, -13, -8, -4, -4, -8, -7, -6, -1, 2, 4, 12, 16, 12, 5, 3, -4, -6, -2, -8, -4, -6, -9, -8, -16, -18, -10, -12, -14, -16, -16, -12, -9, -6, -3, -2, -4, -8, -7, -6, 1, 0, 10, 12, 7, 7, 3, 3, 1, -5, -3, -2, -3, -5, -5, -6, -11, -11, -10, -13, -16, -8, -6, -5, -9, -7, -1, 0, -2, 1, 0, 1, 6, 7, 10, 15, 11, 12, 11, 8, 3, 1, 2, 2, -4, -5, -1, -7, -7, -5, -5, -6, -7, -6, -5, -8, -8, 2, 3, -1, 0, 5, -1, 5, 3, 13, 10, 14, 12, 6, 8, 10, 2, 8, 5, 3, 6, 2, 0, -1, -2, 1, -3, 1, -1, -3, -1, 0, 4, 3, 4, 2, 8, 2, 10, 9, 9, 14, 10, 16, 12, 13, 7, 5, 11, 11, 2, 3, 8, 6, 6, 6, 0, 3, 2, -2, -1, 3, 0, 2, 5, 3, 6, 8, 2, 11, 7, 13, 11, 5, 14, 6, -6, 0, -2, 0, -4, 0, -5, 2, -1, 0, -1, 0, 1, -1, 1, 0, -4, -2, -1, -1, -2, 0, 0, -2, -1, 0, 2, -4, -1, -2, -1, 0, -2, 0, -4, 1, -3, -3, 3, 0, 2, -3, -1, 5, 1, 0, 0, -3, 1, -6, 0, -4, 1, 2, 0, -1, 3, -1, 2, 0, -4, -4, 0, -2, -7, -6, 1, 1, -2, -5, -6, -5, -3, 5, 4, -2, 3, -2, -3, 1, -3, -2, 0, -4, -2, -1, 0, 3, -5, 3, -1, -1, -5, -2, 1, -7, -4, -1, 0, -1, 0, -4, -6, 1, -3, 2, 4, -1, -2, -3, -1, 0, 0, 0, 3, -1, -4, 1, 1, 0, -6, -2, -2, -1, 1, -1, 0, -5, -2, -2, -6, 1, -6, -3, -5, -2, 0, 2, 0, -2, 2, -5, -4, 1, 1, -3, -2, -2, 3, -4, 2, 0, -1, 0, 1, -7, 0, -5, -2, -8, -9, 0, -6, 1, -5, -2, -7, -6, -6, 0, 0, -5, 0, -3, 0, 2, -1, 3, -5, 1, 0, 0, -1, 0, 2, -2, -6, -3, -2, 0, -7, -1, -6, -2, 2, -4, 2, -1, -1, -2, 0, -6, -3, -4, -4, -1, 0, -1, 1, -5, -1, -5, -3, -5, -4, -4, 0, -1, -7, -4, 0, -7, -5, 0, -6, -3, 0, 2, -4, -2, -5, 0, -5, -7, -5, -3, -4, -5, -4, 0, -6, -1, -3, -4, -4, -3, -5, 1, -3, -6, -9, -4, 0, 0, 0, -8, -4, -5, 3, 3, -2, -2, -4, -7, -8, -3, -3, -5, -2, -5, -7, -3, -7, -4, -9, -2, -8, 0, -7, -7, -8, -1, -6, -2, -3, -5, 0, -7, -4, 2, 0, 4, -2, -5, 0, -5, -4, -4, -8, -9, -1, -7, -9, -5, -8, -2, -1, -8, -7, -4, -6, -3, -5, 0, -1, -3, -3, 3, -4, -4, -4, -1, 4, 0, 1, 0, 1, -4, 0, -5, -5, -2, -5, -9, -1, -8, 0, -1, 1, -4, -4, -4, -6, -5, -5, 3, -1, 1, 2, 1, -1, -8, -2, 1, -1, 2, 0, -4, -3, -4, 0, 1, -6, 1, -3, 0, 1, -3, 2, -4, 3, -3, 0, 3, 2, 0, 0, 0, 6, 0, 0, 3, 0, -5, 0, -1, 4, 2, 1, 1, 1, 7, 4, -2, 5, 3, 2, 2, 5, 0, -1, 1, 6, 2, 3, 2, 2, 7, 3, 3, 2, 6, 4, 0, 2, -1, -6, -6, -4, 2, 1, 3, 2, 9, 8, 7, 7, 7, 8, 10, 7, 5, 11, 4, 4, 3, 10, 10, 4, 10, 9, 3, 3, 6, 3, 3, 0, 1, 1, -6, -1, 2, 1, 2, 6, 10, 3, 9, 4, 11, 5, 11, 10, 6, 11, 12, 8, 4, 4, 11, 3, 1, 3, 2, 4, 3, 0, 3, 0, 0, 1, 1, 0, 3, 1, 7, 1, 10, 7, 10, 4, 8, 11, 5, 8, 14, 8, 14, 5, 12, 12, 1, 9, 0, 5, 2, 4, 0, 0, 4, -5, -2, 2, 3, 1, 0, 2, 5, 6, 2, 8, 0, 2, 1, 8, 9, 7, 4, 6, 5, 4, 6, 8, 1, 4, -2, -2, -1, 0, -3, -3, 2, 0, 0, 0, 1, 2, 0, 0, -7, -4, 0, 1, 3, 2, 6, -1, 6, 1, 4, 5, 1, -2, 0, -2, -2, -6, -2, -5, -3, -1, -4, -7, 0, 0, 0, 2, 5, 0, -4, -8, -8, -5, -8, -3, -4, 0, -3, 4, 0, 0, -1, -4, -2, 0, 0, 1, -6, 0, 0, -7, -8, -6, -10, -3, -5, 0, 0, 5, 0, 1, -7, -12, -12, -10, -6, -11, -7, -6, -7, -5, -6, -1, -1, -5, -5, -1, -4, -5, -5, -10, -7, -7, -6, -12, -12, -5, -1, 0, 8, 4, 1, 1, -7, -8, -12, -10, -6, -8, -12, -7, -7, -10, -11, -8, -10, -10, -11, -4, -4, -6, -7, -11, -11, -11, -11, -6, -11, -4, -2, 2, 9, 10, 0, -3, -4, -8, -12, -13, -13, -11, -12, -10, -8, -6, -11, -8, -8, -11, -6, -8, -3, -3, -3, -7, -8, -9, -15, -10, -4, -9, -5, 2, 9, 8, 0, 2, -6, -3, -9, -5, -6, -7, -10, -10, -5, -12, -11, -8, -8, -11, -8, -5, -5, -2, -11, -7, -13, -6, -11, -8, -5, -10, 0, 2, 9, 10, 1, -1, -8, -6, -7, -7, -5, -13, -12, -12, -12, -7, -4, -12, -12, -7, -7, -8, -5, -9, -13, -11, -8, -9, -8, -7, -11, -7, -1, 1, 3, 6, 2, 2, -2, -8, -11, -11, -13, -14, -7, -14, -13, -11, -9, -9, -11, -10, -9, -11, -9, -14, -13, -17, -15, -14, -14, -7, -10, -7, 4, 9, 9, 7, 5, 4, -4, -10, -6, -10, -6, -9, -9, -7, -9, -15, -10, -12, -12, -11, -12, -11, -12, -15, -13, -14, -9, -9, -10, -6, -10, -7, 3, 1, 14, 6, 11, 5, -2, -8, -9, -8, -9, -6, -11, -6, -6, -14, -16, -11, -11, -17, -12, -14, -17, -17, -13, -12, -6, -4, -4, -3, -2, -3, 4, 7, 9, 9, 10, 2, -6, -7, -11, -4, -11, -9, -6, -11, -12, -12, -9, -10, -15, -11, -18, -11, -9, -8, -10, -5, -7, -2, -5, -7, 1, -3, 0, 8, 6, 6, 8, 6, 2, -2, 0, -1, -7, -7, -8, -10, -8, -14, -11, -15, -8, -10, -13, -8, -10, -3, -2, -1, 1, 2, -4, -4, 3, 0, 5, 6, 13, 12, 9, 8, 5, -3, 3, 1, 0, -5, -3, -2, -1, -4, -5, -4, -5, -10, -7, -7, -1, -1, -2, 1, 0, 5, 2, 0, 1, 4, 8, 10, 6, 11, 5, 9, 1, 0, 4, 0, 4, -1, 3, 3, 0, -2, 0, -4, -5, -6, 0, 0, 0, 3, -2, 0, 4, 4, 4, 10, 4, 8, 10, 5, 13, 8, 5, 3, 10, 5, 5, 1, 7, 0, 2, 0, 6, 7, 0, 6, 4, 5, 0, -1, 0, 3, 7, 1, 5, 1, 6, 9, 10, 3, 12, 7, 6, -9, -5, -10, -3, -5, -3, -9, -5, -10, -2, -3, 0, -2, -5, -3, -8, -6, -2, -3, -8, -8, -1, -6, -1, -7, -1, -3, -8, -2, -10, -6, -10, -9, -6, -8, -5, -5, -6, -2, -2, -5, -9, -1, -5, -7, -7, -1, -6, -2, -8, -10, -4, -8, -3, -5, -7, -2, -4, -2, -4, -4, -10, -7, -8, -6, -12, -11, -3, -3, -9, -7, -6, -7, -6, -6, -7, -8, -2, -10, -3, -5, -5, -11, -6, -3, -8, -8, -2, -8, -7, -5, -9, -7, -2, -7, -10, -7, -7, -6, -9, -5, -10, -4, -6, -1, -1, -3, -3, -2, -1, -5, -7, -1, -4, -9, -2, -10, -8, -9, -5, -2, -8, -10, -6, -4, -8, -6, -8, -8, -9, -5, -9, -5, -11, -3, -7, -6, -7, -2, -5, -3, -5, -6, -6, -5, -5, -2, -2, 0, -7, -1, -4, -4, -7, -6, -10, -8, -11, -10, -10, -8, -11, -3, -9, -4, -10, -6, -1, -8, -5, -1, -4, -5, -6, -2, 1, -1, 0, 1, -5, -6, -6, -4, 0, -4, -6, -3, -10, -4, -8, -7, -13, -8, -9, -6, -1, -5, -6, -3, -3, -3, -6, -5, -5, 0, -2, 1, 0, -1, 0, 0, -5, 1, -6, -6, -3, -4, -6, -10, -1, -11, -12, -10, -4, -6, -11, -4, -8, -5, -6, -7, -3, -5, -3, -5, 2, 1, -3, -3, 5, 0, 0, 3, -2, 2, 1, -2, 0, -7, -10, -9, -3, -6, -7, -10, -5, -7, -1, -8, 0, -7, -2, 0, -5, -8, -5, 2, 3, -1, 0, 5, 0, -1, 6, 1, 4, 3, 2, -5, -5, -5, -3, -1, -6, -2, -5, -4, -10, -8, 0, -4, -4, -2, -6, 2, 0, -3, -6, 1, 0, -1, 3, 2, 5, 5, 2, 3, 1, 0, 6, 5, 1, 3, 0, 2, 2, 0, -2, 0, -7, -3, 0, -2, 0, 0, 1, 0, 4, -1, 0, 2, 5, 6, 9, 3, 8, 7, 8, 8, 7, 3, 2, 3, 2, 6, 2, 3, 6, 1, 0, -2, -6, -6, -5, -2, -3, -1, 0, 0, 4, 4, 1, 5, 11, 11, 11, 11, 7, 14, 8, 9, 9, 11, 14, 4, 6, 4, 3, 6, 2, 3, -2, -5, -9, -8, -2, 0, 1, 1, 7, 9, 12, 7, 9, 13, 16, 15, 17, 15, 18, 13, 15, 17, 16, 13, 15, 14, 11, 11, 11, 13, 7, 9, 0, 1, -9, -5, -1, 2, 2, 5, 9, 9, 15, 13, 19, 15, 18, 16, 23, 23, 22, 25, 18, 20, 19, 21, 18, 17, 12, 12, 19, 17, 10, 6, -1, 2, -8, -7, -1, -2, 6, 8, 13, 13, 19, 13, 17, 21, 22, 26, 27, 22, 29, 24, 22, 21, 22, 23, 21, 16, 19, 20, 12, 11, 9, 11, 0, 3, -7, -2, -3, 1, 7, 10, 11, 10, 16, 14, 14, 17, 16, 20, 25, 26, 23, 21, 23, 21, 22, 21, 15, 17, 13, 14, 10, 16, 12, 7, 8, -1, -5, -4, 2, 4, 5, 2, 6, 15, 17, 12, 18, 21, 20, 15, 20, 17, 19, 24, 23, 26, 19, 22, 14, 15, 15, 7, 12, 13, 7, 4, 8, 0, 0, 4, 0, 3, 2, 8, 3, 8, 7, 11, 10, 14, 13, 14, 19, 13, 12, 14, 17, 15, 15, 12, 14, 11, 4, 6, 11, 2, 3, 9, 7, 0, -1, 0, 3, 3, 4, 5, 0, 5, 2, 6, 9, 9, 7, 8, 14, 16, 13, 12, 12, 10, 13, 10, 5, 4, 7, 4, 0, 1, 2, 4, 5, 3, 6, 5, 8, 6, 4, -4, 2, 2, 0, 1, 3, 5, 4, 8, 9, 12, 4, 6, 3, 6, 8, 6, 5, 6, 6, 3, 0, -3, 2, 0, 6, 6, 1, 4, 1, 0, 2, 0, 0, 5, -1, 3, 2, 0, 6, 0, 3, 1, 1, 0, 2, 2, 4, 0, 2, 0, 2, 0, -4, 0, 0, -3, 0, 10, 7, 9, 1, 2, 0, 0, 0, 2, 1, 3, 3, 4, 5, 5, 0, -4, -2, 2, 6, 1, 4, 1, 0, 4, 1, 0, -3, -4, -3, -3, 0, 4, 8, 13, 3, 4, -4, -5, 2, 1, 0, 1, 0, -4, -3, -1, -3, 1, -5, -2, 0, 1, -1, 0, 0, -6, -1, -2, -1, -5, -1, 0, 1, 10, 6, 12, 7, 6, 0, 0, -5, -2, -4, -3, 0, -2, -5, -3, 2, 0, -4, 0, -1, -1, -1, -2, -4, -2, -1, -6, -9, -3, 1, -6, 0, 7, 14, 9, 6, 2, -1, -4, -3, -1, -7, -2, -3, -7, -5, -7, -1, -5, -4, 1, 0, -5, -2, 0, -8, -4, -7, -4, -6, -8, -6, -3, 2, 11, 15, 12, 4, 5, -3, 0, -6, -6, -4, -10, -6, -6, -7, -6, -4, -2, -7, -7, -8, -3, -9, -9, -6, -10, -6, -1, -2, -1, 0, 0, 6, 9, 8, 15, 10, 2, -1, 0, -7, -6, 0, -1, -2, -6, -5, -10, -6, -8, -7, -6, -9, -12, -9, -4, -2, -7, -5, -7, -2, -6, -3, 4, 2, 8, 9, 12, 6, 5, 1, -2, 0, -5, -5, -4, -5, -7, -8, -6, -9, -7, -10, -4, -8, -13, -5, -3, -4, -2, -1, 2, 2, 0, -3, -1, 3, 11, 15, 15, 13, 3, 0, 1, 0, 0, -1, 0, -2, -4, -1, -8, -10, -10, -10, -3, -4, -6, -3, -3, 1, 0, 1, 0, 2, 4, 7, 3, 11, 11, 15, 12, 9, 4, 8, 1, 0, 4, 3, 6, -2, -1, 0, 1, -7, -7, -2, -6, -3, -4, -2, -3, 0, 3, 3, 8, 2, 8, 2, 8, 7, 11, 15, 6, 6, 8, 9, 4, 7, 10, 8, 6, 7, 5, 1, 1, 2, 4, -1, 5, 0, 3, 5, 8, 4, 9, 3, 11, 6, 12, 7, 6, 9, 9, 15, 9, 9, 11, 8, 11, 5, 12, 9, 7, 9, 3, 3, 3, 2, 5, 6, 2, 2, 1, 4, 7, 12, 5, 12, 5, 13, 6, 11, 13, 8, 11, 9,
    -- filter=0 channel=2
    3, 0, 0, 4, 4, 0, -1, 0, 3, 0, 3, -1, -2, 0, 2, -4, -1, 0, 0, 0, -3, 3, 1, 1, 4, -2, -1, 0, 0, -2, 1, 0, -1, -1, 1, -3, 0, -2, 3, 0, -2, 1, 2, -4, 0, 0, -2, -1, 0, 3, 0, -3, -3, 0, -3, -4, 2, -2, -1, 0, 0, 0, -3, 3, 4, 3, 1, -3, 0, -1, -2, 1, -1, 3, -2, 0, -3, 3, -3, -4, 1, 3, 3, 4, 3, -2, -1, 0, 0, -1, 1, 0, 3, 3, 1, 1, 0, 2, 4, 1, -2, 1, 0, 4, 1, -2, -2, 1, 1, 0, 3, -3, 3, -1, 1, 0, -1, 3, 0, 0, -3, -4, 0, 0, -3, 4, -1, -1, 4, -2, 3, 4, 1, 0, 1, 2, 2, 3, -1, -1, 0, 0, 4, 0, 2, 3, -1, -4, 0, 2, 0, 2, 0, 0, -2, 0, 1, 2, 2, -2, -2, 4, -3, -3, -1, 0, 4, 0, -3, -2, -1, 0, 0, -4, 0, -3, -1, 3, 4, 0, -3, -2, -3, 0, 1, -4, 0, -1, 1, 1, 0, -1, 0, -1, 2, -3, -3, 3, 4, 0, 0, 0, 4, -3, -3, 1, 3, -2, 0, 4, 3, -1, 0, 3, 2, 3, 2, -1, -3, 0, -2, 1, 0, -1, 0, -1, 0, 1, 0, -1, 1, 0, -2, 0, -3, 0, 3, 0, -1, 2, 4, 4, -2, 1, -2, 3, -4, -3, -4, 4, -3, 3, 5, 5, -1, 2, 0, 1, 1, 3, -3, -3, 1, 2, -1, -4, 1, 3, -1, -2, -2, -2, 3, -4, 3, -3, -1, 3, -4, 2, 0, 2, -2, -3, -2, -1, 0, 3, -1, 3, 1, 0, 4, 5, 0, 1, 3, 1, -2, -3, -4, 0, -1, 0, 0, -2, -1, 3, 0, 0, 4, -3, 0, -1, 0, 4, 0, 0, 0, 4, -2, -2, 0, -2, 0, -1, -3, 1, 4, -1, -3, -2, -2, -2, 0, -2, 2, 3, 3, 0, -3, 0, -1, 4, 0, 3, -2, -3, -3, 0, -1, 0, 4, -2, 4, 5, -3, 2, 0, 4, -4, 2, -1, 0, -1, -5, -5, 0, 3, 3, 0, 0, -5, -2, -3, 0, -3, -3, -3, 3, 5, 1, 0, 0, -2, 4, -3, 1, 2, 0, -3, -3, -2, 1, 3, 0, -4, -3, -2, 1, -3, 0, -4, -4, 2, 0, -2, 0, 3, 3, -2, -3, 4, -1, -1, -3, 1, 5, 4, 0, 1, 2, 4, 3, 2, -5, 0, -2, 2, -2, 0, -6, -6, -5, 0, 0, -1, 0, 0, -1, -1, -3, -4, -3, -1, 3, 1, -2, 1, -2, -3, 0, -2, 0, -2, -1, -2, -3, -1, 0, -5, -3, -2, 1, -5, -5, -3, 1, 0, -5, 2, 0, -3, -1, 3, 0, -1, -2, 2, 0, 0, 3, 2, -3, 4, 0, 0, -1, 0, -4, -5, -6, -2, -4, -5, -1, -2, 1, -4, -4, 1, 1, 0, 0, 0, 3, 0, 4, 0, 4, -1, 4, 1, 1, 2, -3, 0, -1, -1, -2, 2, -1, 2, -3, 0, -6, -1, -4, -2, 0, 0, 0, -1, -1, 2, -4, 2, 2, 2, 0, 1, -3, -1, 2, 3, 0, -2, -2, -1, -2, -3, -2, 0, 0, -4, -4, 0, 0, -2, -3, 0, -4, -5, 0, -5, -3, -3, -2, 2, 0, 1, 0, 3, -1, 0, 0, 1, 4, -2, 2, 5, 0, 3, 1, -2, 1, 2, 2, -5, -3, -7, -5, 0, -5, 0, 2, 0, -4, -1, -4, 0, -4, -1, 0, 3, -2, -3, 1, -2, 4, 5, 0, -2, 0, -2, -4, -3, -4, -2, -5, 0, -5, 0, -5, 0, 0, 0, -6, -6, -3, -2, 2, -3, 3, 4, 4, 0, 0, -1, -3, 3, -2, 4, 3, 1, 4, 1, 0, 1, 1, 3, -1, 2, -1, -5, 1, -5, 1, -4, 0, -4, -4, 0, 1, -3, -1, -2, -1, -3, 3, -2, 0, -1, 0, -1, -2, -1, -3, 0, 1, -4, 0, -1, -5, -4, -1, 1, -5, -1, 2, 0, 1, 2, 0, 3, 0, 0, -2, 0, 0, 4, 4, 4, 4, 3, 0, 3, 1, -3, -2, 0, 0, 2, 2, 0, 0, -5, 1, 1, -6, -3, 0, -1, 2, -1, 3, 2, -2, -1, 1, 0, -3, 2, -2, -2, -2, -4, 0, 2, 1, 0, 3, -3, 1, -4, 4, 4, -5, 1, -3, 0, 2, 0, -4, -4, 0, 2, 1, 1, 1, 2, -3, -1, 3, -1, 1, 3, 2, 0, 1, 1, -1, 4, -3, 2, 1, 4, 2, -2, -4, 1, -2, 4, -3, -3, -2, 1, 1, -3, 0, 1, 4, 0, 0, -3, 0, 3, -2, -2, 1, 1, 0, 3, 1, -1, 0, -3, -3, 1, 2, 3, 2, 0, 3, 0, -4, 0, 2, -1, 2, 2, 0, 2, 3, -2, 3, 2, 0, -2, 0, -1, 3, -3, -1, -2, 0, 1, -2, 3, 0, -2, 2, 2, -2, 1, 3, 0, 0, 4, -1, -1, 0, 2, -3, 2, 0, 1, 3, 2, 1, 0, -1, -4, 1, 3, 0, 3, 3, -1, 4, 2, 1, 0, 3, 3, -2, 3, 3, 2, 0, 2, 3, 3, 0, 0, 1, -4, 0, -2, -3, 0, 1, 1, -3, 1, 2, -2, 2, -2, 1, 3, 1, 2, -1, -2, 4, -1, 4, 4, 0, 2, -2, 3, -1, 1, -2, 1, 3, 4, -2, -3, 0, -3, -4, 0, -1, 2, -1, 1, 2, -1, -3, -2, 0, 3, -3, -1, -2, 0, 4, 0, -2, 3, -3, -1, -3, 3, -2, -2, 0, 2, -1, -1, -2, 4, -1, 3, 0, 0, 3, -3, 0, 1, -3, -4, -4, -1, -1, -2, -3, -4, -4, 2, 1, -3, 0, 0, 0, 1, -1, 2, 3, -4, -4, -3, 0, 0, 0, 0, -1, 0, 0, 0, -5, -4, -4, 0, 0, 3, -4, -5, -2, -1, -1, 3, 2, 1, 3, -3, -4, 0, 0, 0, -2, -4, 0, -3, -4, -5, 2, 3, -3, 1, 0, -3, -2, -3, 3, 4, 0, 0, -1, 3, -1, 1, 2, 2, -1, -3, 3, -3, -3, 2, -3, -3, 4, -1, 3, -3, 3, 0, 3, 0, -2, -1, 3, 0, 1, 1, -1, 2, 1, 3, -1, -2, -1, -3, -2, 0, -2, 3, 1, 0, 2, -1, 1, -2, -1, -2, 2, -1, 1, 4, 4, 4, 4, 0, -1, 0, -2, 1, 3, -2, 0, 0, 1, -2, 3, 2, 2, 3, 2, -1, -1, -2, 2, 0, 4, 2, 1, 2, -1, 1, -2, 0, -1, 1, 0, 2, -2, 1, 4, 2, 0, -1, 0, -3, 3, 3, 1, -3, 2, -1, 0, 2, 0, 1, -1, 0, -3, 4, -2, 2, 0, 1, 1, 0, 3, 1, 2, -2, -1, 1, 1, 0, 1, 3, 0, 0, 4, -2, -3, 1, 1, 0, 3, -1, -2, 2, -3, -2, -1, 1, 1, 2, 0, -1, 4, 2, -1, 0, 3, 4, 0, -3, -3, -1, 0, 1, -2, 2, 2, -1, 4, -2, -1, 0, -3, 0, 1, 1, 2, -3, -1, 1, -1, 0, -4, -1, 3, 0, -1, 0, -3, 3, 0, 0, 4, -2, 3, 2, 4, 1, -3, 4, 1, 3, 0, 3, 0, -1, -4, 1, -3, 4, -2, -1, 0, -2, 3, -1, 3, 3, 5, 4, 0, 3, -2, -2, 4, -1, 2, -3, 1, 0, 4, -1, 3, 0, -1, 4, 0, 0, 0, 0, -3, -3, 0, 3, 2, 4, 2, 4, -1, 4, 0, 1, 3, 2, 1, 5, 5, 2, 4, 0, 4, 5, -1, 0, -1, -1, -2, 4, -2, 4, 2, 0, 4, 0, -3, 3, 3, 3, 0, 0, -3, -2, 5, 2, -2, 0, 0, 5, 3, -1, 2, 5, 0, 3, 0, 0, 3, 5, 1, 1, 1, 3, 0, -2, 2, 2, 2, -1, 0, 3, 0, 3, 3, 2, -1, -1, -2, 0, 3, 3, 5, 6, 0, -1, 2, -1, -1, 0, -1, 0, 2, 2, -1, 3, -1, -4, -1, -1, -3, -1, 2, 2, -1, -1, -1, 0, 2, 1, 0, -3, 1, 0, -1, -1, 5, -2, 3, -2, 0, 3, -3, -3, -1, -1, -2, -5, -3, 2, -2, 0, 2, 2, 2, -2, -2, 3, 1, -3, 1, 3, -2, 1, -2, 2, 0, 5, 0, 4, 5, 4, -3, -1, -2, 1, 3, 1, -4, 2, 0, -1, -2, -4, 1, -3, 2, 3, 2, 5, -1, 1, 0, 3, 2, 2, 2, -2, 3, 1, -1, 3, 0, 0, -3, 2, 3, -1, 2, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -3, 4, -1, 0, -1, 1, 1, 2, 3, 3, -1, 0, 5, 4, 4, -1, 5, 3, 5, -2, -3, 0, -4, -4, -4, 0, -3, -6, 0, 0, 3, -3, 0, 2, 3, -1, 0, 5, 6, -2, 3, 5, 4, 3, 0, -1, 2, 2, -1, -2, 5, 1, 3, -1, 0, 2, 0, -4, -6, 2, 0, -4, -2, 0, 2, 2, 4, 2, 5, 1, 3, 2, 1, 0, 5, -1, 0, 1, 1, 0, 0, 0, 2, -1, 1, -5, 0, -2, 2, 2, -3, -4, -2, -4, -4, -2, 4, -2, 4, 1, -2, 5, 1, 1, 1, 5, 3, -2, -2, 0, 0, 5, -1, 0, -3, 0, 3, -1, -2, -2, 2, -5, -2, -4, 0, 0, 2, -2, 2, 0, 0, -3, 3, 3, 2, 0, 3, 3, 5, 4, 0, 1, 5, 0, -1, 4, 0, 2, -2, 1, -5, 0, -1, -4, -2, -4, -4, -4, -3, 2, -2, 3, -3, -1, -2, 3, 4, 2, 2, 0, -1, 3, 1, 6, 2, 4, 4, 2, 3, 0, 3, 0, -2, -3, 2, -5, 0, 0, 1, -1, -3, 1, -2, 1, 5, 4, 4, 0, 0, 4, 2, -2, -3, -3, -2, 2, -1, 2, 1, 1, 2, 3, -3, 2, 1, -2, -1, -5, 0, -2, -4, 3, 1, -3, 0, -2, -2, 0, 0, -2, -2, 1, 0, 4, 1, 3, -2, 2, 3, 1, 4, -2, 5, 1, 0, 0, 3, -1, 2, -4, 2, -1, -3, -1, 0, 0, 4, -3, 5, 2, -3, -2, 4, 0, 4, 1, 1, 0, -1, 4, 0, 1, 0, -1, 1, 0, -1, 2, -3, -3, 0, 0, -3, 1, 3, 0, -1, 0, 2, 4, 0, 2, -2, 4, 5, 3, 0, 2, 0, 0, 4, 2, 4, 2, 3, 0, 2, 0, -3, -1, 1, 1, 0, 3, 0, -3, 4, 0, 3, 3, 2, 0, 0, 2, 2, 0, -2, 4, 0, 4, 1, 2, -2, -3, 5, 1, -2, 4, 1, -2, 2, 4, 0, 2, -4, -2, 0, 0, 0, -1, -1, 0, -2, 0, -1, -1, -2, 5, 4, 4, 0, 2, 4, -2, -2, -2, 1, 3, 0, 0, 0, 0, 4, -2, 0, -2, 3, 0, 1, -1, 1, -1, 2, 1, 0, 0, 0, 1, 3, 3, 0, -2, 4, -3, 0, -1, 2, 0, -3, 5, -1, 0, 2, -3, 0, -4, -2, -1, 2, -3, 3, 1, 3, 1, 1, -1, 4, 1, 1, -1, -3, 3, -2, 3, -2, 4, 4, 0, -3, 0, 1, 2, -3, 3, -2, 0, 2, 4, 0, 2, 4, 3, 3, -3, 1, 3, -3, 1, 2, -3, -2, 0, -2, -3, 4, -3, -1, -1, 0, 3, 0, 2, -1, 3, -3, 3, 4, -3, 2, -1, -3, -3, 0, 1, -1, -3, -1, -1, 3, 0, 2, 0, -2, 0, -3, -4, 0, 4, 2, 1, -1, 3, -4, -1, 0, -2, 3, 2, 0, 1, -2, 2, -3, -2, -4, 2, 0, -4, -3, 2, -2, -1, 0, -3, -4, 2, -3, -4, 0, 1, 0, -1, -1, -1, 0, -1, 2, 2, 0, 0, 0, 4, -2, -1, 3, 3, 1, 2, -1, -1, -2, -4, -1, 3, 3, -3, -1, 2, 3, -1, 1, 1, -3, -3, -1, -1, 0, -1, -4, -2, 0, -3, 3, 3, 3, 0, 3, -1, -4, 0, 2, -3, 1, 3, -1, 0, 0, -2, -5, -4, -1, -1, 1, -1, 0, -1, -3, -3, -2, -3, 0, -5, -4, 1, 0, -4, 0, -3, -6, -6, 0, -6, -4, -3, 0, 0, 0, 0, -3, -3, -1, -6, -2, 0, -3, -2, -2, 1, -3, 0, -1, -3, -3, 0, -3, 0, -3, -1, -5, -1, 0, 1, 0, 0, 0, 2, -4, -2, -1, -4, -3, -5, -2, -4, -6, 0, -2, -5, 1, 0, 0, -4, -6, -5, -3, -3, -1, 0, 0, 1, -2, -1, -5, -2, 0, -4, -3, -5, -3, -4, -4, -5, 1, -1, -1, -1, -5, -6, -2, 0, -6, 0, -5, -1, -5, -3, 2, 2, 1, 2, -3, 1, 0, 2, -3, -2, -2, 0, -5, 1, 0, -2, -4, 0, -6, 0, -4, -4, 0, -3, 0, 1, -3, 0, -1, 1, -2, 0, -1, 1, 1, -3, 0, -2, 0, -4, 0, 0, -3, 0, -2, 1, 0, 0, -1, -4, -4, -1, -5, -5, 2, 0, 2, -5, 1, -2, -5, -4, 0, -3, -1, -4, -1, -3, -4, -3, 3, 2, 2, 0, 1, 0, -5, 0, -3, -4, 0, 0, -5, -4, 2, 0, 0, 0, -4, -1, 1, 3, 2, -2, 0, -3, 0, 3, -4, 0, 0, -1, -5, -2, -3, 0, -5, 0, -3, 0, -4, -4, -2, 2, -3, 1, -4, -2, -2, -3, -5, -2, 0, 1, 0, 3, 0, -2, -4, 1, 3, 1, -1, -2, 3, -2, -1, -1, -2, 1, -4, 0, 0, 1, -3, 3, 3, 0, 0, 2, 3, -4, 2, -1, 3, 1, -4, 0, 0, -2, -4, 2, 1, -3, -1, -3, 0, 1, -3, 2, 3, -1, -4, -4, 0, 1, -3, -2, 0, 0, 2, 0, -5, 0, 0, 0, -3, 2, -1, 0, 2, 1, 0, 3, 3, 0, 4, 0, 0, -1, 1, 1, 3, -1, 3, 2, -1, 1, -3, 3, -3, -1, -2, 2, 1, 1, 1, 0, -1, -4, -4, 3, 1, -4, 2, -2, 0, -3, -2, -2, 1, 0, -3, 0, 0, -3, 2, -4, 3, -2, -2, 3, 0, -4, -2, -1, 0, -3, 2, -3, -2, -3, -1, -4, 0, 0, 4, 1, -1, -2, -2, 1, 0, -4, 3, 1, -1, -2, 0, -3, 0, -2, -3, -4, 2, -2, 4, -4, -2, -2, 0, -4, -2, 2, -3, 2, -1, 1, 0, 4, -1, -2, -1, 1, 3, 2, 3, -4, -5, 1, -2, -4, 1, 0, 3, 3, -2, -1, 2, -3, 3, 0, 0, 3, 4, -1, -3, -3, 3, 0, 0, -3, 3, -3, -3, 0, 0, -2, 2, -2, 2, 0, 0, -4, -2, -2, -3, 2, -3, 2, 4, -2, 4, -2, 4, 0, 1, 3, 0, 2, -1, 3, 0, 3, -4, 4, -3, 1, 3, 1, 3, -3, -4, -5, -3, -3, 0, -3, -4, -2, 2, -2, 0, 3, 3, -4, 0, 0, -2, -4, -2, -3, -3, -2, 1, -1, 0, 2, -1, 0, 3, 1, -3, 3, 1, -4, -3, 2, 0, 1, -3, -5, -1, -4, -3, -2, 4, -3, 3, -1, 3, 0, 1, 1, -2, 1, -3, 0, -2, -2, -2, 0, 1, -5, 2, -1, -5, -1, 0, -3, -3, 2, -1, 3, 0, -3, -1, -2, 2, 0, -1, 2, 2, 2, -2, -1, -1, -4, 4, 2, -2, 2, 2, 0, -1, 2, -1, 1, -3, 1, -3, -4, 2, -2, 0, 0, -2, 2, 1, 4, -1, -2, -4, 3, 0, 2, 1, 3, -2, 0, 0, 2, 0, 0, -4, 1, -1, -1, 0, -2, 1, -5, 0, -2, -4, 0, -2, 2, -2, 0, 0, 3, 2, 4, 3, 2, -2, -3, 1, 0, 1, 2, -2, 1, -4, 3, -1, 2, -2, -3, 2, 0, 1, -1, -3, 1, -5, 0, -3, -4, 0, -1, 0, 1, -1, 3, -3, 0, 0, -4, 1, 2, -3, 0, -1, 1, 4, -1, -2, 0, -4, 0, 1, 0, 1, 0, 2, -2, -1, -5, -2, -1, -3, 0, 1, -2, 0, 4, 3, 0, 2, 0, -4, -2, 0, -3, 0, -1, -1, 3, -3, -3, 0, 0, -1, -4, -4, 0, -4, -4, 3, 2, -1, 4, -3, -3, -1, -3, 4, 4, -2, 0, 3, -4, -2, 4, -3, 3, 2, 0, 0, -3, -2, 4, 0, -3, -4, 2, 3, -2, 1, -3, 3, 0, -1, -1, -2, -1, -1, -1, 1, -3, 2, 4, 0, -3, -2, -3, -2, 0, -1, -2, 3, 0, 1, -3, -1, 4, 0, -4, -4, 0, 3, 3, -3, 0, 2, 1, 2, 1, -2, 0, 3, -3, -4, -1, -3, 1, -2, -2, 3, -2, -3, 0, -3, 0, -2, 1, -2, 0, -4, 3, 0, -1, -2, 3, -2, 4, 0, -3, -2, 3, 0, 0, -3, 0, 2, -4, 3, 0, -3, 0, -4, -2, 2, 3, 3, 0, -3, 0, 2, -3, 0, 0, -2, -2, 1, 0, 1, -2, 0, -2, -4, 0, 0, 2, -2, 1, 0, -2, -4, 1, -1, 0, 0, -2, -2, 3, 4, -2, 1, 1, 0, -3, 0, -1, 3, -2, -1, -4, 4, 0, 3, 3, 1, 0, -4, -2, -2, 0, 4, -5, -4, -3, 2, 1, 0, 1, -1, 3, 2, 2, 0, 0, 0, -4, -3, 0, 0, -2, 0, 1, 0, 3, -2, -3, -3, -2, -2, 1, 3, -2, -4, -4, -1, 0, -2, -4, -3, 0, 0, 1, 0, 0, -4, -1, 1, -3, -2, -1, 3, 0, 0, 3, 1, -3, -1, 2, -4, -2, 2, 2, 0, 3, -5, -3, 3, 2, -4, 0, -4, 0, 0, 2, -1, 3, 2, -3, 0, 2, 0, 0, -2, 2, -3, 1, -2, 1, 0, 3, -1, -2, 0, 2, -5, 0, -2, 1, -4, 0, 2, -3, 1, 0, -5, 2, 1, -2, 0, 1, 0, 2, -4, 1, 0, 0, -2, 1, 1, 2, 2, -4, -1, -4, -3, 1, 3, -2, -3, 2, -4, -3, 1, -3, -5, -2, 0, 2, -4, 1, 1, 0, -1, -4, -1, 0, 1, 0, -4, 0, -3, -1, 0, -1, -1, -5, 1, 0, 0, -4, -1, 0, -4, 1,
    -- filter=0 channel=3
    0, 0, 4, 5, 3, 0, 2, 4, 4, 4, 2, 0, 1, 4, 0, 1, 4, -3, 1, 3, -1, 0, 4, 0, 0, 4, 0, 0, 2, 1, 3, -2, 5, 4, -1, 0, 5, 5, 3, 1, -2, 3, -3, 2, 4, 1, 1, 0, 1, -3, -3, 5, 1, -2, -1, -1, 1, 1, 6, 4, 2, 1, -1, 3, 0, 2, 3, 2, 1, 4, 2, 4, 5, -1, -2, 2, 2, 0, 0, 1, -3, -1, -3, -2, 1, -2, 1, 4, 5, 5, 3, 7, 3, 1, 0, 4, -2, -1, 2, -1, 6, 6, 5, 4, 4, 0, 3, 0, -3, 0, 2, -2, 2, -4, 1, 1, -3, 3, 2, 0, 1, 0, 4, 2, 2, 1, -1, 4, 0, 6, 1, 5, 2, 5, 0, 0, -1, -2, 0, 0, -3, -1, -3, -2, -1, -5, -3, 0, -3, 3, 4, 1, 2, 3, 0, 2, 2, 0, 7, 3, 1, 7, 0, 4, 4, -1, 5, 1, 2, -1, 3, -2, -2, 0, -2, -5, -2, -1, -6, 0, 0, 0, -1, -2, 0, 1, 8, 0, 2, 2, 0, 6, 4, 5, 6, 3, 3, 5, 0, 4, 0, 2, -4, 1, 0, -6, -2, -2, 0, -4, -1, 0, 0, 0, 0, -2, 3, 1, 7, 1, 0, 2, 7, 2, 0, 6, 0, 2, 0, 2, 4, 3, 2, 0, 0, 3, 0, 0, -6, -4, -3, 0, 0, -2, -3, -5, 1, 0, 0, 6, 0, 7, -1, 1, 0, 6, 0, 5, 0, 2, 0, 0, 3, -1, 2, 1, 2, 2, 1, -5, -3, -5, 1, 0, 0, -5, -3, 0, 1, -2, -1, 0, 5, 2, 1, 1, 1, 3, 6, 3, 3, 0, 0, 5, 5, -1, -2, 2, 0, -2, -6, -1, -3, -3, -6, -6, -5, 0, -4, 2, 0, 3, 2, 0, 1, 4, 7, -1, 7, 4, 7, 4, 5, 1, 6, 0, 1, -2, 1, 0, -4, 0, 1, -2, -4, 0, -4, -5, 0, 0, 2, -5, -1, 0, 0, -2, 4, 2, 0, 2, 0, 5, 5, 1, 0, -1, 4, 2, 0, 0, 1, 0, 0, 2, 0, -1, -1, -4, -4, -2, -3, -4, -1, 0, 2, -3, 0, 3, 2, 6, 0, 0, 2, 2, 3, 4, 6, 0, 0, 2, 2, -1, 0, -1, -1, -5, 2, -4, -2, -3, -6, -5, -2, -4, -3, 0, 1, -2, 1, 0, 3, 2, 6, 6, 1, 6, 3, 0, 2, 0, 3, 1, -1, -4, -4, 2, 2, -5, -3, 0, 0, -4, -2, 0, -4, 2, 0, 2, 1, 2, 1, 4, 1, 4, 4, 3, 0, 0, 3, 4, -1, 0, -3, -3, 3, 2, -4, -5, -5, -4, 2, 0, 0, -1, -4, 2, -3, 1, 2, 3, -3, 0, -4, 3, 0, 0, 4, 0, 3, 3, 4, 1, 5, 4, -4, 0, -3, -2, 1, 0, 1, 1, 0, -3, 2, -2, 1, -3, -4, 1, -4, -2, 1, 0, 1, -2, 1, 2, -1, 5, 0, 3, 1, 0, 0, 1, 0, -2, 0, 0, 1, 3, -1, 0, 0, -3, -3, -1, 0, 2, 0, -1, 0, 2, -1, 2, 3, 1, -1, 5, 2, 1, 4, 2, -2, -2, 4, 0, 2, 0, 0, -2, 0, -4, 1, 0, -1, 1, 3, 0, 3, 1, 0, -4, -3, 0, -3, 1, 1, 0, -1, 0, 2, 6, -1, -3, 0, 1, 1, 0, -2, 3, 0, -1, 0, 1, -4, 0, 0, -3, 0, 1, 3, -4, -1, 3, -2, 0, 0, 2, -1, 0, 5, -2, 0, 0, 0, 0, 0, -3, 2, 1, 4, 3, 3, 1, -1, -3, 2, 0, 0, 2, 0, 0, -1, 4, 4, -1, 2, 0, -3, 4, 0, 0, 5, 1, 4, 4, 4, -3, 3, 4, -2, -3, 3, 1, 0, 0, 4, 1, -3, 0, 1, 2, 0, 6, 2, 0, 3, 0, 0, -3, -2, 4, -3, 0, 3, -2, 2, 5, -1, -3, 2, -2, -3, -2, 0, -3, 2, 1, -1, 2, 4, 2, 0, -1, -1, 0, 2, -2, 1, 2, 0, 0, -3, 3, -1, -1, 0, 1, -2, 0, -1, 1, -3, 4, 4, -2, 2, 2, 4, 4, -3, 5, -2, 2, 2, -2, 4, 5, 5, 3, 4, 3, 0, 0, -2, -2, 2, 5, 4, 1, -1, 4, 2, -1, 4, -1, 0, 0, 2, 1, 3, 0, 4, 5, 1, 0, 5, 4, -1, 0, 6, 7, 4, 2, -2, 2, -3, -1, 4, 1, 0, 2, 2, 0, 0, -3, 1, 1, 1, -1, 3, -2, 1, 0, 3, -1, 4, 4, -1, 4, 5, 2, 5, 0, 5, 3, 2, 4, 3, 6, 2, 5, -1, 0, 3, 1, 5, -2, 2, 1, -2, -3, 4, 0, 4, 6, 5, 0, 3, 4, 0, 5, 2, 4, 8, 2, 0, 1, -1, 0, -1, -2, 6, 0, 0, 1, 2, 2, -1, 2, 2, 3, 2, 0, 2, 3, -1, -2, 5, 4, -1, 2, 7, 6, 4, 3, 0, 4, 4, 6, 7, 1, -1, 4, -2, -2, 1, 0, -2, 3, -3, 0, 0, 3, 1, 5, -2, 4, 5, 2, 5, 0, -2, 4, 3, 1, 2, 5, 8, 4, 4, 7, 3, 6, 1, 2, 3, -1, -1, 1, 5, 5, 0, 0, 4, 3, -3, 4, -1, 5, 0, 6, 6, 1, 6, 2, 0, 6, 6, 7, 5, 6, 2, 3, 1, 3, -1, 3, 4, 0, 4, 1, 3, -2, 2, 0, 0, 3, -3, 4, 0, -2, 1, 6, 0, 6, 2, 0, 0, 2, 7, 2, 2, 3, 0, 4, 1, 1, 0, 0, 0, 3, 0, -2, 5, -1, 2, 2, 3, 1, 0, -1, 3, 1, 4, -1, 1, 0, -1, 2, 0, -1, 2, 4, 6, 3, 2, 6, -1, 0, 0, 1, 3, 0, -2, -1, -1, -3, -3, 0, 0, 0, -4, 3, 4, -2, 0, -1, 5, 1, 0, 2, 0, -1, 0, 4, 0, 4, 0, 5, 4, 5, 5, 0, -2, 1, 1, -1, -1, 2, 2, 0, -3, -3, 2, 3, -5, -1, 1, -4, 1, 0, -4, -3, -5, -4, 0, 0, -1, -3, -3, 0, -4, -1, -6, -5, -1, 2, -2, -2, -2, 0, -2, 0, 1, 2, -3, 0, -1, 3, -1, 0, -1, -5, -1, -3, 1, -1, -1, -6, -2, -6, 1, -1, 2, 1, 1, -5, 0, -2, 0, 0, 0, -2, 1, -3, 2, -4, -2, 0, 3, 2, 2, 0, 1, -1, -2, -5, -5, -7, -4, -5, 0, -1, -5, -6, 0, -2, -3, -3, 1, 0, -1, -1, 0, 1, 1, -4, 3, -4, -2, 0, 2, 0, -2, -2, 2, -2, -3, -1, -2, -6, -6, -6, -2, 0, 0, 0, -4, -1, 0, -4, 1, 3, 2, 0, 3, -2, -3, -3, 0, 1, 1, 2, 1, 1, 2, -5, -3, 0, -2, 0, -3, -5, -4, 0, -7, -5, -4, -6, -7, 0, -2, -1, -2, 2, 2, -3, 2, 1, 1, -1, 3, 1, 0, -1, -3, 2, 0, 3, 1, 0, -7, -4, -7, -8, -7, -6, -2, -1, -1, -1, -7, -7, -3, 1, -2, 0, 0, -2, -2, 0, 0, 0, 4, 1, 0, 2, 0, -1, 0, 3, -4, 1, 0, -6, -4, 0, -2, -4, -8, -1, -8, -5, -6, -5, -4, -2, 2, 2, 3, -1, -3, 1, 0, 2, 2, -1, -3, 2, -3, -2, 1, 0, -4, -6, -5, -7, -8, -7, -2, -4, -7, -7, -5, 0, -7, -6, -6, 0, 1, 3, 2, -1, -3, 1, 1, -3, 1, -2, -3, 0, -1, -4, 0, 0, 2, -3, 0, -2, -8, -1, -5, -4, -6, -3, -4, -1, -5, 0, -6, 0, -5, 0, -1, 2, 3, -2, 0, 3, 3, -3, 2, -3, 4, 2, -3, 3, 2, -6, 1, 0, -4, -4, -2, -4, -4, -8, -6, -5, -4, -1, -3, 1, -5, 0, 4, 0, -3, -1, -1, 1, 2, 0, 5, 1, 1, -2, 0, -4, 0, -5, 1, -7, -6, -1, 0, -5, -3, -6, -4, 0, 0, -5, -1, 0, 2, -3, 0, 2, 4, 4, 0, 3, 0, 3, 3, 0, 3, -2, -1, 2, -3, 0, -5, 0, -1, -4, -7, -3, -4, -6, -7, -4, -3, -3, -1, 0, 0, 1, 0, -2, -2, 2, 1, -2, -3, -2, 0, 2, -3, 0, -1, 0, -2, -4, -6, -3, -5, -2, -6, -4, -3, -4, 0, 0, -6, 0, -3, -5, 0, -4, -3, 0, 0, 3, 0, 4, 4, 0, 1, 3, -3, -3, -3, -3, 1, 0, -5, 0, -6, -2, 2, 0, 2, 0, 0, -3, -5, -3, 0, -1, 2, -4, 0, -2, 3, 0, 4, 0, 1, -4, 0, -3, -1, -4, -2, -1, 1, -5, 2, -3, -4, 0, -1, 2, 0, 1, 0, -4, -3, 2, 1, 0, 1, 0, -1, -1, 0, -1, 2, 3, 3, 3, 2, 0, -3, -2, -2, 0, 2, -5, 2, -1, 2, 0, 1, 3, -2, -4, -4, -3, 1, 3, 0, -5, 2, -1, 0, 0, -4, 0, 3, -3, -3, 3, -1, 3, 3, -4, -1, -4, -1, 0, 2, -3, -4, 3, -4, -4, 2, -3, 1, 1, -4, -2, 0, 3, 1, 0, 3, 3, 4, 3, -4, 0, 1, 1, 0, -4, -4, 1, 1, -4, 0, 0, 0, -4, -1, -2, 4, 2, 4, 1, 0, 3, -4, -1, -5, 0, -1, 0, 2, 2, 3, -3, 3, -5, -1, 0, -5, 1, 0, -4, 2, -2, 1, -4, -3, -5, 4, 4, 0, -3, 5, 2, 0, 3, 1, 0, 4, -3, -3, -2, -1, 1, 2, 2, -4, 0, -1, 0, 3, -3, -3, -3, 1, -3, -1, -1, -3, -3, 3, -3, 5, 4, 0, 5, 5, 4, -2, 2, -1, -2, 5, -3, 0, -2, -4, 0, 3, -5, -2, 0, -1, 1, -1, -1, 1, 4, 1, 0, -3, 0, 2, 3, -2, 1, 3, 5, 5, 2, -3, 4, 4, -2, -1, -2, -3, -3, 4, 2, -4, 0, 0, -3, -1, -2, 2, 0, -4, 0, -1, 2, 3, -1, 3, -2, 4, 1, 4, -1, 2, 5, 0, 0, 4, 0, -1, -4, -2, -2, 2, 1, -3, -1, -5, -4, -2, 1, -4, 4, 3, 3, -3, -3, 0, 2, 5, 5, 5, -2, 0, 6, -1, 5, -1, 1, 4, 1, 3, 0, 4, 1, 0, 2, -4, -1, 2, -1, 0, 2, 2, 4, 2, -2, 0, 1, 5, -3, -1, 0, 5, 0, 6, 1, 0, -1, 3, 0, 3, 0, 0, -4, 0, 3, -2, 2, -1, 2, 1, 2, -3, 1, -2, -1, -2, 0, -2, 3, -3, 0, 0, 0, 1, 4, 0, 1, 3, 4, -2, 4, 4, 0, 0, -2, 3, -2, 0, 0, 0, 2, 2, 0, 0, -4, -2, 3, -1, 3, 1, 1, -3, 0, 4, 6, 5, 0, 5, 0, 0, -1, 2, 3, 1, 1, 4, 4, 1, -2, 3, -1, -1, -4, 0, -1, 2, -4, -4, -4, 4, 3, -3, -2, 0, 4, -1, 5, 0, 3, 0, 0, 3, -1, -1, -3, 2, 2, 0, 0, -1, 4, 0, 0, -5, 2, 1, 2, 0, -5, -4, 1, 0, 4, 2, -2, 3, 1, 6, 0, 5, -1, 3, 6, -1, 1, -2, 1, 0, 5, 2, 4, -1, 1, 0, 3, 1, -1, 2, 2, -3, -4, -4, -3, 2, 2, -3, -1, -3, -1, 5, 4, 6, 3, 5, 0, 1, 5, -2, 3, 0, -1, 0, 4, 1, -4, 0, 3, -4, -1, 0, 1, 1, -1, -4, 1, 3, 0, 4, -2, -2, 4, 4, -2, 4, 0, 6, 2, 1, -1, 5, 0, -1, 1, 0, 0, 4, 4, -2, -4, -2, -3, -2, 0, -1, -5, -2, 3, -2, 4, -1, -1, 5, 4, 5, 4, 3, 0, 0, 1, 4, 1, -3, 0, -1, -1, -1, 2, -1, 3, -4, -4, 2, -1, 1, 0, -4, 1, -3, 0, 1, 3, 3, -1, -1, 1, 4, 0, 0, 3, 3, 0, -1, -2, -2, 0, 3, 4, -3, -3, -4, -4, -3, 0, 2, -4, 2, -5, -4, 0, -3, -1, -2, 1, -4, -4, -6, -5, -1, 0, 1, -4, -4, 1, 0, -5, -6, 1, -2, 1, -5, -3, -1, -1, 1, -3, -4, 0, 3, -1, -3, -4, -2, 0, 2, -5, -5, -2, 0, -3, -5, 0, 1, 0, -6, 0, -6, -6, -1, -6, 0, -6, 0, 0, 1, 0, 3, -3, -2, 0, 0, -3, -1, 0, 1, -4, -5, 1, -1, -4, -1, -5, -1, -1, 0, -6, -6, -4, -3, -4, -1, 0, 0, 0, 2, -1, 3, 2, -2, -2, 0, -1, 0, -4, 2, 0, 0, 1, 3, 0, -3, -3, -6, 1, 0, 0, -1, 0, -2, -4, 0, 0, -7, 0, 1, -3, 0, -3, -2, -1, 1, -3, -2, 3, -1, 0, -4, 0, -2, 4, -2, 0, -3, 0, -3, -3, -2, -4, -1, -6, -7, -3, -1, -7, -6, -5, -1, -4, 0, 0, 0, 2, -1, 0, 0, 0, -3, -1, 2, 1, 3, -3, -3, 0, -1, -3, -1, -3, -4, -5, -3, -3, -3, -8, -8, -8, 0, -7, -1, 2, 0, 1, 0, 3, 1, -1, 4, -3, 2, -3, 2, 0, 3, -3, 1, 0, -5, 0, -5, -4, -6, -4, -7, -8, -8, -9, -9, -2, -3, -6, 0, 1, 3, -2, -3, -3, 4, 1, 0, -3, 5, -2, 3, -3, 0, 2, 3, 3, -3, -6, -1, 0, -6, -8, -1, -5, -1, -6, -6, -3, -2, 1, 1, -5, 0, 2, 4, 0, 0, 5, 0, 5, 0, 1, -3, 2, 0, -3, -1, -1, -2, -3, 0, -7, 0, -6, -3, -8, -4, -1, -8, -6, -5, -3, -5, 1, 3, 4, -1, -3, 3, -1, 2, 4, 0, 3, -1, 0, 0, -2, 4, 2, 0, -1, 0, -7, -2, -3, -7, 0, -5, -9, -6, -3, -2, -5, -2, 1, 1, 1, -3, 0, -1, 2, -2, -1, 0, 1, -1, -2, 2, 2, 2, 3, -1, -6, -6, -7, -1, -2, -2, -7, -5, -6, -5, -5, -4, -6, -5, -6, 1, 2, 0, 1, 0, -2, 4, 1, 5, 0, -2, -3, -3, -2, 0, -5, -5, -5, -2, -4, -2, -4, -7, -4, -4, -5, 0, 1, -1, -6, -2, 0, -2, 0, 0, 4, -3, 3, 2, 4, 1, 4, -1, 4, -1, 1, 0, -4, 1, 1, -4, -4, -3, -1, -6, 0, -4, -5, -3, -5, -6, 0, 1, 2, 3, 4, -3, 3, -1, 0, -1, 2, 2, 5, 1, 3, 2, -2, -3, -3, -4, 2, 0, 0, -3, 0, -3, -1, 1, 0, 0, -3, 1, -2, -1, -1, 1, -3, 1, 4, 0, 2, 4, 5, 2, 0, 0, -2, 3, -3, -2, -4, -2, -3, -1, 0, -4, -2, 3, -5, 2, 0, 0, -4, 1, 1, 3, 0, -3, 0, -2, 0, 0, 0, 0, 0, 0, 0, 3, 3, -1, 2, 1, -4, -3, 0, -3, 0, -2, 1, -2, 2, 0, -1, -4, -2, 0, -2, 1, 2, 2, 2, 0, -1, -1, -2, 0, -2, 0, 3, 4, -2, -1, -2, -3, -4, -5, -1, -2, 3, 1, -4, 0, 1, -3, 0, 4, 1, 0, 2, -3, 0, -4, 1, -1, 4, -1, 2, 0, -1, -2, 5, 2, -1, -4, -3, -1, -3, 3, 1, -4, 2, -2, -2, -1, 1, 4, -1, 3, 0, 2, -3, 2, 3, -2, 0, 2, 0, 0, 2, 5, -3, 2, 0, -2, 3, 0, -1, -2, 0, -3, -4, 0, 2, 1, 1, -1, 4, 0, 3, -3, 0, 3, 0, -4, 0, 5, 1, 2, 3, 1, -1, -3, 4, -2, 0, 0, -1, -3, 2, 3, 2, 2, -3, 1, 0, 5, 0, -2, 0, 3, 0, 4, 0, -2, 2, -1, -2, 1, -1, 5, 4, 0, -2, -2, 2, -2, 1, 3, -3, 3, 3, -1, 2, -2, -3, -3, 0, 0, -1, 0, -2, -2, 3, 1, 0, -1, 0, 3, 0, -1, 4, 3, 3, -1, 0, 1, 1, 4, -3, -1, 0, 0, -3, 4, 4, -2, -1, 4, -3, 1, 0, 6, 0, 4, 0, 6, 4, 0, 1, 5, 4, 2, 3, 2, 2, 3, 0, 4, 4, 0, 4, 0, 4, -1, -3, -2, 1, 0, -2, 1, 0, 1, 4, 2, 0, 3, 6, 3, 4, -1, 0, 2, 3, 0, 0, 5, 3, 3, 5, 1, 0, 0, 4, 0, 5, -1, -1, 0, -2, 1, -1, 0, 4, 4, 5, 0, 2, 2, 7, 7, 2, -1, 1, 3, -1, 5, 1, 2, -2, 5, 3, 1, 0, -2, 0, -1, 2, -3, 2, 5, 2, 1, 0, 4, 2, 4, 0, 7, 0, 4, 1, 8, 7, 5, 0, 0, 4, 6, -2, 1, 5, 5, -1, -2, 1, 0, 0, 2, 0, 0, 0, -2, 4, 6, 6, 0, 6, -1, 6, 8, 8, 8, 5, 0, 0, 5, 2, 6, 1, 4, 3, 0, 3, 5, 5, 1, 3, 4, 1, 1, 0, 1, 1, 0, 4, 3, -2, 6, 7, 0, 6, 8, 1, 7, 3, 7, 1, 3, 2, 1, 4, 0, 0, 2, 4, 3, -2, 1, 2, 3, -2, 2, 3, 3, 6, -2, 0, 0, 5, 0, 0, 6, 2, 5, 4, 3, 8, 5, 5, 6, 1, 0, 0, 3, 6, -1, 0, 4, 4, -1, 0, 3, -3, 4, 4, 2, 0, 6, 6, 6, 5, 2, 1, 1, 7, 0, 1, 1, 2, 2, 5, 6, 5, 2, 1, 5, 6, 0, 6, 1, 2, 1, 2, -1, 2, 1, -1, 4, -1, -1, -1, 0, -1, 6, 6, 1, 8, 6, 5, 8, 6, 5, 8, 4, 0, 0, 7, 7, -1, 0, 5, 4, 3, -1, -2, 5, 4, 0, 3, 0, 0, -1, 5, 3, 4, 6, 0, 0, 0, 1, 8, 8, 2, 8, 3, 3, 0, -1, 0, 6, 0, 3, 2, 1, 1, 5, 3, 1, 0, 1, 2, 4, 4, 6, 4, 4, 2, 2, 1, 2, 4, 3, 3, 8, 5, 6, 1, 1, -1, 1, 1, 4, -1, -2, -1, -2, -2, 3, 2,
    -- filter=0 channel=4
    -9, -9, -11, -5, -9, -2, -7, -2, -5, -6, -2, -1, -8, -9, -7, -8, -2, 0, -4, -4, -7, -3, -6, -9, -6, -9, -3, -4, -7, -5, -9, -8, -9, -2, -1, -4, -8, -7, -7, -9, -1, -8, -5, -4, -7, -3, -7, -5, -4, 0, -6, -6, -7, -9, -6, -5, -7, -9, -9, -2, -9, -11, -10, -14, -4, -10, -2, -6, 0, -7, -6, -7, 0, -5, -3, -2, -7, -3, -7, -5, 0, -1, -2, 0, -5, -6, -4, -6, -5, 1, -1, -6, 0, -5, -3, -10, -5, -2, -8, -1, 0, -3, -5, 0, -4, 2, -2, -5, -5, -3, -4, 0, -1, -5, -2, -3, -4, 1, 1, -4, 1, -1, -6, 0, -4, -2, -3, -2, -10, -3, -6, 0, 0, -2, -2, 1, 4, -2, -6, 1, -2, -4, 0, 0, -4, 0, -1, -2, 0, 0, -1, -3, -1, 2, -1, 0, 0, 0, -7, -3, -4, -4, -7, -4, -6, -2, -4, 1, -1, 1, -2, -6, -8, -3, -8, -5, 0, -3, -6, 0, -5, -5, 0, 1, 3, 5, 0, 2, 1, -4, -3, -5, -9, -7, -9, -4, -2, 0, 1, 0, 2, 0, 0, -3, -3, -1, -5, -3, -9, -4, -6, -4, 0, 1, 1, 0, -3, 4, 3, 0, -6, -4, 0, -2, -7, -7, -3, -7, 0, -2, -4, 2, 2, 1, -2, -2, -3, -5, -5, -7, -4, -1, 1, -2, -4, -4, -4, 2, -4, 1, -3, 2, -5, -8, 0, -3, -2, 0, -3, -5, -1, 0, -1, 0, 6, 0, 1, 0, -2, -7, 0, -3, -5, 0, -4, -8, -7, -1, -4, 0, -2, 0, 1, -1, -3, -6, -7, -7, -4, -1, -4, -1, -3, -3, 5, 5, 4, 0, -1, -3, 0, -7, -7, -2, -5, -7, -5, -6, -1, 0, -2, -7, -2, -1, -6, -1, -4, -1, -7, -5, 0, 1, 0, -5, -3, -2, -1, -1, -3, 2, 0, -4, -3, 0, -1, 0, 0, -2, 0, -5, -3, -5, -2, 0, -6, 0, 0, -4, -2, -4, -3, -2, -3, -1, -6, 0, -6, -2, -4, 4, 0, 5, 4, 2, -5, -2, 0, 0, -5, -3, 0, -2, -3, -6, -5, -5, 0, -6, -1, -5, -2, -4, -6, -4, -3, -6, -2, -3, -1, 0, -5, 0, 3, 3, 3, -4, -4, -3, -7, 0, 3, -1, -4, 0, -4, 2, -5, -6, -1, -6, -2, -7, -6, -1, -3, -3, -4, -4, -7, 1, -1, -4, -1, 1, -4, -3, 1, -3, -6, -8, -4, 0, -5, 2, 2, -1, 0, 4, 2, -2, 1, -3, -5, -1, -3, -1, -5, -3, -1, 0, -6, 2, 0, -5, -3, 3, 1, -5, -6, 1, -1, -3, -3, 2, 3, 0, 0, -2, 2, -3, 0, 1, -3, -2, 1, -2, -5, -2, 0, -8, -9, -3, -6, -4, -1, -1, -1, -1, -1, -1, 0, 1, 0, -4, -1, 1, -1, 5, 2, 0, 0, -1, 0, 0, 4, -3, 0, 0, -2, -1, 0, -9, -4, -7, -3, 0, 2, -3, 0, -3, -2, 1, 0, 3, -2, 0, 1, 0, -2, 3, -2, -3, 0, 1, 5, -1, 0, 4, 1, 0, -3, 3, -4, -5, -3, -5, -3, -3, -4, 2, 3, 1, -1, -1, -1, -1, 0, -4, 2, 0, 5, 3, -2, 6, 5, 3, 3, 0, 4, 2, 5, 2, 2, -3, -1, -5, -5, -5, -4, -1, -2, 1, 0, 0, 5, 0, 5, 0, -1, 2, 2, 0, -1, -1, 2, 3, 5, 3, 4, 9, 6, 7, 4, 1, 5, 0, -3, -9, -3, 4, 2, 4, -1, 1, 6, 4, 1, -1, -1, 1, 4, -2, -2, -8, -4, -3, 0, -2, 6, 0, 0, 2, 8, 1, 8, 2, 5, 4, 0, -9, 1, 4, 0, 6, 4, 3, 0, 2, 0, 2, 4, -1, -2, 2, -3, -12, -6, -2, 1, -1, -2, -3, 0, 4, 6, 2, 8, 1, 6, 5, 2, -7, -3, -2, 2, 4, 5, 1, 5, 2, 5, 1, 0, 4, 2, 0, -6, -7, -6, -6, -3, -3, 1, 1, -4, 2, 7, 1, 1, 6, 0, 0, -1, -1, 0, -1, 6, 5, 2, 6, 5, 0, 6, 1, 3, 6, 4, 0, -3, -5, -6, -6, 1, 2, 0, 3, -2, 5, 8, 7, 8, 4, 0, 5, 0, -8, -1, 6, -2, 1, 2, 3, 1, 4, 3, 4, 3, 0, 5, -1, -3, -4, -3, -3, -1, -1, 1, 0, 4, 3, 3, 2, 1, 5, 6, 0, 0, 0, -3, -2, 0, 5, 6, 6, 2, 2, 1, 6, 2, 8, 6, 4, -2, -2, 0, -3, 3, 6, 5, 3, 4, 0, 3, 0, 5, 0, 6, -1, 1, -5, 1, -3, 5, 2, 3, 0, 2, 0, 0, 3, 5, 6, 8, 4, 4, 6, 1, -4, -2, 2, 0, 1, 2, 2, 9, 2, 1, 7, 3, 3, -6, -2, -3, 0, 3, 5, 2, 3, 1, 0, -2, 0, 7, 4, 2, 6, 4, 6, -1, 2, 0, 0, 6, 1, 8, 0, 6, 6, 3, 0, 1, -5, 0, 0, 2, -3, -2, 1, 6, -1, 0, 1, 0, 5, 6, 6, 9, 9, 2, 2, 5, 5, 1, 3, 4, 4, 4, 5, 3, 1, 2, 2, 1, 2, -2, -5, 0, -1, -2, -2, 0, 6, 5, 3, 3, 4, 7, 2, 2, 9, 7, 8, 1, 9, 4, 4, 1, 4, 4, 5, 3, 7, 6, 1, -2, 0, -4, -5, 0, 2, 0, -1, 5, 3, 4, 4, 8, 7, 3, 4, 3, 2, 9, 2, 5, 8, 1, 2, 2, 3, 9, 6, 1, 0, 2, 3, 0, 0, 3, 0, -2, 0, 3, 3, 6, 5, 4, 1, 5, 5, 6, 7, 5, 6, 8, 1, 4, -1, 3, 7, 3, 3, 0, 4, 0, 3, 0, 2, 2, -1, -4, -1, -1, 5, 0, 3, -1, -1, 3, 0, 0, -1, 5, 2, 5, -1, 4, 5, 4, 0, 3, 0, 2, -2, 3, 0, -2, 1, 0, 4, -2, 0, -1, -6, -9, -4, 1, -3, -2, -2, -3, 3, 2, 1, 0, 1, 1, 2, 0, 5, 3, 5, 5, 5, 5, 3, 0, 0, -1, 3, -4, -5, -1, 0, -2, -7, 0, -2, -4, 0, 0, -2, -1, 0, -2, 5, 4, 2, 0, 5, 3, 1, 3, 7, 4, -1, 3, -2, 3, 0, -1, -3, 0, 0, -3, 1, -6, -3, -6, -1, -4, -3, 4, 4, 3, -1, 5, 0, 0, 3, 5, 0, 5, 1, 6, 7, 0, 6, 5, 4, 7, 0, 5, 3, 0, 5, 4, 1, -4, -2, -4, 1, -2, 3, 2, 0, 1, 4, 1, 6, 7, 9, 4, 2, 4, 0, 8, 6, 6, 0, 8, 7, 3, 6, 6, 7, 3, 5, 4, 5, 1, 1, -5, 2, 1, 4, 6, 2, 5, 1, 4, 7, 1, 8, 8, 7, 1, 1, 3, 0, 1, 0, 4, 6, 8, 4, 6, 3, 6, 3, 5, 4, 6, -1, 2, -1, 4, 2, 2, 2, 5, 3, 6, 4, 5, 7, 1, 5, 7, 7, 1, 2, 3, 1, 6, 6, 4, 4, 7, 13, 2, 6, 3, 0, 1, 5, -3, 3, 4, 0, 5, 10, 7, 9, 4, 3, 9, 0, 3, 1, 5, -1, 9, 7, 9, 2, 3, 8, 7, 4, 11, 6, 6, 2, 8, 5, 3, 0, 4, 1, 5, 1, 8, 6, 6, 7, 5, 10, 6, 4, 6, 0, 2, 2, 3, 8, 11, 6, 8, 6, 7, 8, 4, 12, 8, 8, 6, 5, 2, -1, 3, 6, 0, 8, 11, 10, 8, 11, 8, 12, 11, 8, 3, 8, 7, 9, 9, 10, 6, 5, 4, 11, 9, 5, 11, 5, 8, 4, 5, 6, 6, -1, 4, 8, 4, 5, 5, 9, 9, 14, 10, 9, 5, 5, 7, 8, 3, 6, 3, 3, 2, 2, 4, 4, 7, 8, 6, 6, 4, 9, 3, 2, 5, 2, 6, 10, 4, 9, 3, 1, 8, 7, 12, 14, 12, 9, 8, 10, 7, 3, 6, 0, 1, 6, 7, 8, 8, 6, 10, 5, 3, 2, 10, 9, 2, 3, 6, 4, 8, 4, 6, 1, 5, 11, 12, 10, 10, 2, 0, 7, 2, 3, 7, 1, 1, 4, 10, 10, 6, 8, 10, 4, 10, 6, 10, 2, 3, 4, 1, 5, 10, 9, 6, 3, 4, 5, 8, 4, 7, 6, 3, -3, 0, 4, 3, 7, 6, 1, 1, 8, 12, 11, 7, 8, 3, 8, 3, 6, 7, 3, 2, 5, 4, 5, 11, 5, 7, 9, 4, 7, 0, 3, 3, 0, -5, 0, -4, 0, -3, 1, 1, 10, 10, 11, 3, 10, 10, 6, 10, 6, 11, 5, 3, 4, 9, 6, 9, 4, 6, 4, 8, 4, 0, 1, 2, -2, -4, -2, 0, -1, 3, 0, -1, 4, 7, 6, 10, 10, 6, 7, 6, 8, 4, 8, 7, 7, 13, 8, 9, 7, 3, 4, 0, 4, 0, 0, 0, -2, -8, -6, 0, -1, -3, -1, -3, 0, 8, 7, 3, 5, 7, 9, 12, 9, 10, 6, 2, 12, 7, 7, 7, 5, 11, 7, 8, 0, 1, -3, 1, -4, -2, -3, -6, -3, -6, 1, 0, 0, 0, 4, 6, 6, 10, 9, 12, 7, 4, 0, 2, 9, 11, 8, 13, 14, 13, 4, 5, 9, 3, -1, 2, -6, -7, -2, -1, -6, 0, -2, 2, 4, 1, 11, 7, 11, 11, 16, 8, 8, 6, 3, 2, 12, 8, 9, 12, 15, 9, 5, 7, 9, 7, 0, 4, 0, -5, -10, -9, -6, -8, 0, 2, 4, 8, 11, 11, 9, 13, 15, 12, 15, 9, 3, 10, 10, 12, 7, 16, 9, 7, 5, 9, 9, 7, 6, 1, 1, -5, -11, -12, -4, -9, -5, -1, 3, 5, 12, 14, 16, 17, 13, 9, 9, 9, 6, 8, 6, 15, 14, 15, 13, 11, 13, 11, 8, 8, 3, 4, -1, -9, -6, -11, -12, -6, -5, 2, 0, 1, 8, 6, 9, 13, 11, 12, 11, 10, 1, 6, 11, 12, 14, 16, 12, 12, 6, 12, 9, 6, 4, 0, 2, -6, -6, -5, -9, -7, 0, 6, 6, 1, 7, 5, 7, 14, 10, 8, 10, 12, 1, 9, 11, 12, 12, 12, 10, 17, 15, 15, 9, 5, 11, 4, 0, 0, -2, -9, -2, -2, 6, 9, 8, 8, 8, 10, 7, 16, 10, 8, 13, 11, 0, 6, 12, 8, 12, 15, 13, 15, 15, 15, 7, 14, 9, 9, 4, 2, -1, -1, 1, 0, 1, 10, 11, 11, 11, 11, 13, 13, 15, 15, 8, 6, 6, 2, 9, 12, 14, 13, 12, 12, 11, 12, 13, 11, 11, 5, 8, 1, 0, -2, 5, 8, 11, 8, 8, 10, 14, 11, 7, 15, 13, 9, 7, 6, 5, 7, 6, 13, 7, 10, 11, 11, 13, 13, 15, 15, 12, 8, 7, 5, 8, 4, 1, 7, 5, 12, 11, 9, 13, 12, 13, 15, 9, 8, 9, 5, 0, 3, 6, 7, 12, 10, 14, 10, 7, 13, 8, 15, 8, 11, 13, 14, 13, 3, 8, 11, 8, 14, 7, 11, 13, 10, 10, 14, 9, 6, 9, 2, 4, 5, 9, 7, 5, 8, 13, 6, 10, 13, 14, 15, 11, 16, 15, 7, 14, 14, 11, 15, 16, 14, 15, 12, 8, 13, 13, 9, 10, 6, 11, 6, 7, 4, 5, 6, 14, 5, 13, 10, 9, 15, 14, 17, 12, 12, 11, 14, 16, 15, 10, 12, 14, 12, 9, 13, 12, 11, 14, 9, 10, 6, 5, 8, 10, 3, 5, 10, 12, 7, 8, 14, 11, 15, 14, 16, 15, 9, 15, 14, 12, 10, 17, 11, 12, 16, 13, 9, 10, 14, 9, 12, 10, 6, 8, 9, 8, 4, 8, 11, 12, 6, 7, 14, 12, 13, 14, 15, 9, 12, 11, 9, 9, 10, 9, 13, 8, 7, 9, 12, 12, 6, 13, 5, 10, 6, 10, 12, 7, 6, 12, 5, 12, 7, 9, 13, 7, 8, 10, 14, 7, 6, 9, 13, 10, 4, 10, 11, 10, 8, 10, 12, 7, 12, 7, 6, 6, 5, 6, 10, 2, -13, -9, -11, -10, -9, -6, -12, -11, -6, -10, -6, -12, -9, -8, -10, -5, -10, -9, -12, -13, -7, -12, -6, -9, -10, -14, -8, -7, -9, -14, -16, -16, -14, -11, -8, -5, -12, -5, -9, -10, -5, -5, -10, -7, -12, -7, -10, -12, -2, -7, -8, -4, -8, -9, -10, -12, -4, -10, -12, -8, -12, -11, -10, -11, -10, -9, -11, -7, -2, -6, -7, -3, -9, -5, -4, -9, -5, -3, -9, -9, -4, -8, -9, -9, -4, -7, -3, -5, -7, -1, -6, -8, -5, -10, -6, -8, -17, -13, -10, -10, -2, -6, -6, 0, 0, -3, -4, -2, -2, -6, -7, -4, -6, -3, -7, -5, -4, -3, -8, 0, -6, -1, -1, -8, -8, -8, -9, -9, -8, -9, -4, -8, -5, 0, -5, -5, 0, -3, -5, 0, -2, -6, -2, -3, -3, -1, -7, -3, -5, -2, -1, 0, 0, -1, 1, -3, -2, -8, -4, -8, -7, -8, -11, -10, -6, -7, -4, 0, 2, 0, -4, -7, -8, 0, -7, -9, -9, -1, 0, 0, -7, -5, 0, -2, -2, -3, 0, -2, -9, -6, -6, -7, -11, -12, -11, -1, -5, 1, 1, -2, -1, 0, -7, -2, -7, -6, -6, -7, -3, -5, -1, -6, -3, 0, 0, -3, 0, 2, -5, 0, -7, -4, -9, -11, -10, -2, -8, -1, 0, -2, -5, -2, -4, -4, 2, 2, -7, -6, -8, -6, -3, 0, 2, -6, -3, -6, -4, 0, 0, 0, 1, 1, -2, -6, -9, -12, -3, -8, -7, -2, -1, 3, 0, -2, -1, 1, 0, 3, -3, -5, -6, 0, -2, -1, -7, -5, -6, -3, -4, 1, -1, -5, 0, 0, -1, -4, -3, -8, -6, -5, -5, -2, -4, -3, 2, -1, -2, -2, 1, 4, 2, -4, -7, -3, -7, -8, -2, -2, -1, -2, 1, 1, -1, -1, -5, -1, 0, 0, -6, -5, -8, -4, -1, -6, 0, -7, 2, -2, -2, 2, 0, -1, -3, -4, -9, -8, -6, -6, -2, -1, -6, -3, -3, -1, -3, -2, -4, -2, 0, -5, -2, -8, -5, -2, 0, -5, -4, -1, -6, 0, 4, 0, 1, -4, -4, -7, -8, -5, -2, -6, -3, -1, 0, -3, -6, -5, -6, -2, 0, -4, -5, -4, -3, -5, -8, -3, -3, 0, -7, -3, -4, -5, -1, -3, -1, -6, -3, -5, -5, -9, -5, -4, -7, -5, -2, -4, 0, 0, -5, -5, -9, -3, -3, -8, -2, -8, -5, -8, -7, -1, -7, -7, -6, 0, -1, -2, 0, -2, -4, -4, -2, -3, -4, -2, -8, -3, -7, -5, -1, -1, -2, -7, -9, -5, -9, -7, -1, -5, -4, -9, -4, -6, -2, -4, -5, 1, -8, -9, 0, -6, -5, -11, -9, -9, -4, -5, -9, -6, -4, -1, 0, -3, -6, -5, -9, -4, -8, 0, -7, -8, -3, -5, 0, -6, 0, -6, 0, -7, -4, -3, -7, -2, -3, -8, -9, -8, -4, -2, -4, -5, -3, -5, -1, -7, -6, -4, -1, -2, -1, -2, -3, -2, -4, -3, -2, -5, -6, -3, 0, -2, -4, -2, -7, -9, -2, -6, -13, -9, -11, -5, -3, -8, -3, 0, -3, -4, 1, -4, -6, -7, -3, -4, -3, -12, -11, -7, 0, 0, -4, 1, 0, -1, -7, -8, -6, -5, -6, -3, -7, -6, -3, -6, -5, -7, -8, -7, 0, -7, 0, -6, -2, 0, -6, -3, -2, -12, -5, -1, -7, -7, -3, -2, -5, -5, -8, -5, 0, -4, -2, -9, -13, -8, -13, -5, -11, -6, 0, -8, -6, -5, -4, -3, -4, 3, -3, -5, -1, -3, -6, -7, -2, 0, -1, 0, -2, -8, -7, -8, -6, -6, -8, -10, -14, -12, -12, -12, -8, -4, -8, -6, 0, -5, -1, -6, 0, 0, -4, 2, 0, -6, -9, -4, -3, -2, -3, -5, -4, -8, -8, -2, 0, -5, 0, -4, -6, -17, -14, -16, -6, -7, -8, -8, -8, 0, -4, -1, -3, 1, -4, 0, -2, -4, -4, -2, -7, -1, -1, 0, 0, -2, -5, -3, 0, -6, -7, -10, -12, -18, -11, -16, -6, -5, -5, -3, -2, 0, -3, 1, -5, 0, 0, 0, 0, -5, -4, -6, -8, 0, 1, -2, 0, -1, 0, -3, 0, -5, -4, -4, -9, -12, -10, -7, -8, -1, -2, -1, -4, -6, 0, -3, -1, -4, -7, -1, -3, -12, -6, -2, -5, -8, -1, -3, -3, -1, -1, -2, -3, -2, -7, -9, -5, -7, -9, -5, -8, -4, -7, 0, 0, -1, -4, -3, 0, 0, -7, -2, -3, -8, -9, -8, -8, -5, -6, -8, -2, -9, -6, -7, -3, 0, -3, -4, -5, -7, -10, -7, -9, 0, -4, -3, 1, -1, -1, -1, 0, -4, -3, -8, -10, -8, -5, -3, -8, -7, -8, -1, -3, -8, -5, -6, 0, 0, -8, 0, -4, -5, -7, -4, -1, -6, -3, 1, -1, -2, -8, -1, -1, -5, -9, -4, -7, -10, -10, -4, -12, -12, -7, -8, -11, -4, -12, -6, -1, 0, -6, -6, -5, -2, -3, -3, -4, -8, -3, -6, -7, -3, -9, -7, -7, -5, -4, -4, -7, -11, -11, -5, -7, -8, -4, -7, -3, -12, -12, -3, -5, -2, -7, -4, -1, -9, -8, -11, -4, -6, -8, -11, -10, -6, -5, -10, -10, -6, -6, -3, -7, -9, -10, -9, -12, -10, -9, -8, -8, -7, -7, -7, -3, -6, -5, -2, -8, -10, -9, -3, -9, -5, -3, -8, -7, -5, -3, -10, -3, -12, -10, -8, -12, -9, -11, -13, -4, -5, -2, -2, -5, -4, -7, -8, -5, -4, -9, -9, -1, -5, -8, -3, -2, -3, -2, -7, -7, -11, -8, -7, -11, -11, -7, -6, -11, -5, -11, -10, -12, -4, -10, -8, -2, -3, -12, -7, -4, -10, -9, -6, -10, -5, -5, -4, -12, -6, -5, -4, -6, -10, -9, -11, -11, -5, -6, -6, -6, -10, -8, -12, -4, -10, -11, -10, -8, -10, -11, -8, -10, -12, -11, -12, -10, -7, -9, -7, -9, -6, -7, -11, -13, -9, -5, -12, -7, -12, -9, -13, -9, -9,
    -- filter=0 channel=5
    -1, -8, -3, -3, -1, -2, -4, -6, 0, -5, 3, 0, -2, 1, -3, -2, 0, 1, 0, 0, -1, -3, 3, 0, -4, -7, -4, -1, 0, -4, 1, -5, -1, -5, 2, -3, -3, -4, -4, -3, -1, 1, -1, 6, 8, 9, 8, 8, 6, 7, 2, 9, 10, 6, 0, 0, -4, 0, 1, -6, 0, -2, -6, 0, 2, -1, -2, 1, 0, 3, 3, 0, 6, 4, 8, 4, 13, 6, 12, 13, 12, 14, 16, 16, 6, 8, 9, 5, 0, -1, -5, -1, 1, 1, 1, -5, 3, 2, -4, 3, 5, 2, 4, 6, 5, 4, 11, 12, 8, 15, 11, 13, 15, 12, 15, 17, 8, 10, 8, 5, 5, 0, -1, -2, -3, -2, -5, -1, 2, 1, -3, -3, 4, 1, 1, 6, 9, 6, 14, 13, 18, 22, 20, 15, 17, 14, 20, 11, 17, 14, 11, 10, 7, 5, -3, -4, 1, -2, -3, -3, 1, 3, 2, 4, 5, 3, 9, 3, 7, 11, 10, 18, 17, 22, 20, 21, 17, 14, 19, 13, 11, 14, 14, 8, 8, 4, 0, -2, -3, -4, -4, 1, -1, 3, -1, 6, 3, 1, 4, 5, 11, 11, 15, 18, 17, 19, 20, 19, 16, 22, 17, 15, 15, 16, 10, 11, 7, 2, 6, 4, -1, -2, -2, -2, -1, -2, 2, 0, 5, 5, 1, 7, 5, 6, 9, 13, 17, 12, 20, 16, 18, 16, 18, 15, 18, 12, 15, 11, 7, 3, 8, 4, 2, -3, 1, -4, -2, -3, 0, 5, 6, 4, 9, 5, 3, 6, 7, 6, 14, 14, 17, 12, 16, 17, 12, 16, 10, 15, 11, 8, 9, 8, 2, 4, 1, 0, -1, -4, 0, 2, 2, 0, 6, 5, 7, 8, 10, 8, 10, 4, 4, 8, 8, 12, 9, 6, 9, 14, 9, 13, 12, 5, 3, 6, 2, 0, 0, -3, 0, -1, -3, -3, 1, 0, 0, 5, 5, 4, 1, 6, 3, 1, 6, 2, 6, 11, 5, 5, 10, 8, 4, 9, 7, 8, 3, 7, 2, 5, 4, 4, -4, -3, 0, 1, 2, 5, 2, 7, -1, 1, 6, 6, 0, 5, 2, 4, 5, 5, 6, 7, 4, 10, 7, 6, 0, 4, 1, 0, 5, 5, 0, -2, 5, -1, 1, 2, -2, 3, 4, 0, 2, 4, 0, 0, -1, 1, -2, -1, -3, 1, -2, -4, 0, 3, 2, -2, 0, 1, 3, 7, 6, 0, 3, 2, 0, 3, 1, 4, 5, 4, 2, 0, 0, 5, -1, 0, 2, -2, 1, 0, 0, -5, 1, 0, -3, 1, -2, -1, 3, -1, 6, 6, 0, 0, 0, 3, 2, -1, -1, -2, 3, -3, 1, 0, 1, -1, 2, 0, 2, -3, 1, -2, -6, -2, -3, -5, -4, -7, -4, -5, -3, -1, 0, -2, 1, 2, 1, -2, 1, 0, -4, 2, -3, 0, 3, -3, 0, -2, 0, -4, -3, 0, 2, 0, -4, -7, -3, -8, -1, -3, -4, -5, 1, -2, 4, 2, 2, 6, 1, 0, -1, 3, -1, 3, -2, -1, -3, 0, 3, 1, -1, 4, -3, 3, -3, -5, -3, -1, -5, -2, -2, -7, -5, 1, -3, 1, 0, 0, -1, 4, -2, -2, 3, -1, 2, 4, 0, -3, -1, -3, 1, 0, 4, 4, 2, 0, 3, -2, -2, -3, -1, -3, 1, 0, 0, 2, 4, 7, 6, 7, 6, -2, 0, 0, -4, -1, -2, -4, -4, -3, -2, 5, 3, 0, 0, 4, 9, 0, -1, 2, 5, 4, -1, -4, -5, -1, 0, 1, 8, 2, 6, 1, 5, 0, 0, -2, -4, -2, 0, -2, -5, -4, 4, -1, 5, 1, 2, 6, 4, 2, 8, 5, 1, 3, 0, 3, -3, 2, 5, 2, 8, 1, 9, 6, 0, 2, -3, 3, 0, -2, 0, -4, -2, 2, 0, -3, 1, 0, 4, 2, 9, 8, 3, 7, 2, 1, -1, 3, 3, 4, 4, 7, 9, 8, 10, 1, 7, 6, 0, 0, -6, -9, -7, -6, -3, -5, -3, 4, 5, 0, 5, 4, 5, 13, 8, 3, 1, 6, 3, 2, 1, 7, 3, 4, 8, 1, 2, 7, 4, 4, -4, -5, -4, -7, -10, -4, -3, -5, 0, -1, 0, 6, 6, 6, 6, 11, 6, 7, 11, 5, 2, 2, 10, 2, 2, 9, 4, 9, 6, 5, 0, -1, 1, -2, 0, -11, -12, -3, -4, -2, 1, 0, 3, 3, 5, 6, 9, 11, 7, 11, 9, 2, 7, 3, 5, 10, 9, 3, 6, 11, 9, 2, 7, 2, 0, -2, 1, -5, -4, -3, 0, -3, 2, 0, -1, 1, 8, 4, 6, 9, 7, 11, 5, 3, 8, 11, 6, 12, 10, 8, 2, 10, 11, 3, 7, 8, 1, 0, -1, -9, -5, -3, -1, 0, -2, -1, 4, 7, 3, 3, 11, 11, 11, 9, 3, 11, 13, 8, 7, 10, 6, 2, 7, 8, 9, 6, 7, 7, 3, -5, -1, -6, -11, -11, -3, 0, 2, 2, 4, 6, 10, 6, 10, 14, 9, 13, 4, 5, 6, 13, 13, 8, 9, 4, 8, 5, 6, 4, 0, 6, 4, -2, -1, -12, -4, -5, -1, -6, -3, 5, 6, 0, 10, 12, 13, 11, 11, 8, 12, 8, 9, 12, 9, 13, 12, 4, 3, 1, 3, 1, 4, 2, 1, 0, -2, -11, -11, -3, -9, 2, -3, 5, 4, 5, 6, 6, 9, 5, 7, 10, 12, 4, 4, 8, 7, 11, 5, 7, 2, 2, 3, 5, -1, 3, -1, 0, -9, -8, -5, -11, -2, -3, 2, -3, 4, 6, 9, 1, 7, 7, 6, 5, 9, 9, 2, 7, 4, 5, 6, 5, 1, 0, 4, 5, 5, -3, 1, -3, -8, -5, -4, -10, -3, -3, -1, 0, 3, 5, 7, 7, 6, 4, 3, 5, 5, 2, 4, 6, 2, 8, 0, 2, 1, 6, 2, -2, 0, 1, -3, 0, -2, -5, -7, -6, -5, -1, -1, 0, -1, 4, 3, 2, 0, 4, 6, 0, 1, 5, -1, 2, -2, 0, 1, -1, 0, 0, 0, -1, 0, -1, -3, -7, -7, -5, -6, -10, -11, -14, -12, -12, -13, -8, -16, -9, -14, -12, -12, -4, -8, -7, -5, -8, -8, -7, -12, -5, -7, -8, -11, -14, -9, -11, -11, -7, -11, -9, -13, -14, -6, -12, -11, -11, -13, -5, -5, -5, -4, -6, -1, -7, -7, -3, -6, -3, 0, 1, 0, -5, -10, -10, -4, -11, -8, -11, -13, -7, -7, -8, -4, -12, -10, -9, -4, -8, -4, -7, -7, -2, -1, -6, -4, -1, 0, 0, 5, -1, 0, 0, -2, -4, -7, -5, -11, -6, -13, -9, -6, -6, -13, -5, -3, -6, -11, -8, -2, -1, -7, -1, -4, 0, 2, 0, -2, 4, 1, 6, 7, 2, 2, 4, 0, 2, -5, -2, -9, -6, -11, -6, -7, -6, -7, -6, -2, -6, -11, -3, -3, -1, -1, -1, -4, -3, 0, -1, 1, 9, 4, 8, 4, 5, 9, 7, 5, 5, 2, -4, -2, -9, -5, -11, -3, -10, -13, -7, -6, -6, -9, -9, -9, 0, 1, -3, -3, 0, 0, 7, 2, 10, 5, 10, 5, 5, 8, 3, 4, 0, -1, 0, -6, -3, -1, -7, -4, -7, -7, -8, -7, -1, -2, -3, -3, -6, -4, -7, -2, 3, 3, 7, 6, 6, 4, 4, 8, 2, 5, 1, 5, 4, 2, -3, -4, -1, 0, -5, -7, -3, -4, -3, -4, -10, -2, -3, -5, 0, -4, -2, 0, 1, 0, 6, 2, 2, 5, 5, 2, 8, 3, 4, 6, 1, -1, -3, -2, -3, 1, -2, -5, -1, -3, -8, -10, -2, -6, -9, -8, -5, -2, -7, 0, -3, -1, 2, 3, 3, 8, 1, 4, 3, 6, 0, 0, 0, 1, -3, 2, 0, -6, -5, -1, -6, -3, -6, -8, -10, -7, -6, -3, -3, 0, -1, 1, -2, 2, -5, 0, 3, -1, 2, 0, 1, 3, 0, 0, 1, 2, 0, 0, -2, -6, 0, -1, -1, -5, -10, -6, -6, -10, -9, -4, -7, 0, -1, -2, -1, -3, -3, -8, -5, 4, -4, -2, 0, -1, -3, -4, 0, 1, 0, -3, -8, -10, -6, -8, -9, -4, -5, -7, -7, -4, -9, -2, -2, -1, -3, -5, -2, -8, -2, -6, -4, -3, 1, -2, 0, 0, -1, 1, 0, -1, -1, -7, -8, -4, -4, -5, -7, -7, -10, -3, -3, -8, -7, -1, -8, 0, 1, -4, -3, -7, -6, -1, -7, -6, -3, -3, -6, -8, -4, -2, 0, -7, -5, 0, -2, 0, 0, -8, -9, -3, -7, -2, -4, -2, -5, -9, -4, -1, -4, -2, -8, -1, -2, -9, -8, -7, -2, -5, -8, -5, -7, -7, -3, -2, 0, -7, 0, -1, -7, -2, -4, -3, -1, -4, -5, -9, -5, -8, -5, -8, -7, -2, -2, -2, -8, -3, -6, -3, -1, -3, -8, -3, -9, -2, -7, -5, -6, 0, -4, -1, -6, -1, -7, -5, -3, -10, -7, -11, -10, -7, -6, -3, -2, -2, -8, -3, -1, -3, -7, -5, -4, -2, -3, -8, -2, -11, -3, -5, -3, -4, -3, -2, 1, -8, -4, -2, -6, -9, -5, -5, -4, -2, -9, -6, -4, 0, -2, -2, -3, -5, 0, -3, -4, 0, 0, 0, -8, -5, -7, 1, -3, 2, -6, 1, -5, -6, -3, -3, -8, -10, -3, -10, -5, -7, -3, 0, -4, 2, 4, 4, 0, -2, 4, 0, 0, 0, -3, 0, -6, -3, 0, 4, -1, 3, 3, 0, -1, -6, -2, -6, -4, -10, -4, -5, -7, -4, 0, 0, -4, 3, 1, 4, 5, -1, 1, 3, -2, 3, 0, -4, 1, -5, 1, 0, -4, 2, -3, 2, -2, -3, -3, -4, -11, -9, -8, -1, -6, -7, 0, 0, 0, 3, 4, 1, 5, 1, 0, 3, 0, 2, -6, 0, 0, 3, 0, 2, -1, 0, 0, -2, -4, -6, -7, -6, -10, -13, -2, -7, -7, -3, -5, 1, -2, -1, 6, 1, 7, 1, 3, 2, -2, 0, 1, -3, -2, -1, 5, 3, 0, 1, 5, 0, -3, -2, -7, -3, -9, -13, -8, -6, -10, 0, 0, 0, 3, 4, 4, 5, 4, 7, 6, 5, 1, 2, 4, -2, 0, 0, 2, 3, 0, 4, -2, -1, -4, -4, -5, -10, -11, -14, -8, -6, -9, -1, -5, 0, 3, 0, 2, 4, 8, 7, 7, 7, 2, 1, 6, 4, 0, 5, 0, 3, 7, 0, -1, 0, 0, -7, -5, -5, -9, -11, -14, -12, -8, -7, -7, -1, -5, 1, 4, 0, 3, 1, 5, 5, -1, 4, 0, 2, 8, 3, 7, -2, 1, 0, 3, 3, -1, -6, -7, -10, -7, -15, -10, -6, -10, -7, -4, 0, 2, 2, -1, 0, 5, 2, 3, 4, 5, 5, 1, 1, 1, 2, 0, 5, 0, 0, 6, 3, -3, 0, -2, -5, -13, -15, -13, -5, -2, -6, -6, -6, -3, -3, 0, 5, 2, 0, 1, 5, 7, 2, 3, 8, 7, 3, 2, 3, -1, -2, 5, 4, 1, 0, -4, -8, -15, -10, -11, -10, -11, -5, -8, -3, 0, -1, 4, 3, 0, 8, 9, 0, 0, 6, 2, 0, 2, 1, 2, 4, 1, 0, 0, 0, -5, -1, -3, -11, -15, -15, -14, -9, -4, -7, -2, -5, 1, 0, 0, 6, 0, 2, 4, 3, 4, 0, 0, 0, 3, 1, 4, 4, 0, 2, -5, -3, -7, -5, -10, -6, -10, -10, -10, -8, -8, -10, -7, -5, 1, 1, 1, 1, 2, 2, 0, 5, 0, 1, 0, -3, 4, 0, -2, -4, 1, 2, 1, -5, 0, -6, -13, -11, -11, -15, -10, -10, -7, -8, -1, -2, -3, 4, -4, -3, 3, -3, 2, -1, 3, -1, 0, 3, 1, 0, 1, -2, -3, 0, -1, -5, -1, -4, -6, -12, -17, -12, -14, -9, -12, -11, -6, -1, 0, 1, 1, 0, 0, 4, 2, -5, 0, 0, -5, -1, -1, -2, -4, -5, -1, -3, -6, -7, -8, -8, -9, -14, -9, -13, -14, -10, -13, -13, -3, -6, -5, -4, -1, -2, 0, 0, -8, -3, -8, -1, -2, 0, -1, 1, 0, -7, -3, -9, -5, -10, -9, -9, -12, -8, -14, -11, -16, -14, -10, -13, -17, -9, -13, -19, -13, -11, -8, -12, -11, -11, -8, -8, -8, -13, -10, -12, -13, -8, -11, -8, -16, -14, -17, -17, -18, -18, -12, -10, -13, -16, -12, -8, -14, -9, -13, -7, -10, -6, -10, -8, -9, -9, -5, 0, -7, -8, -7, -4, -10, -10, -10, -12, -9, -17, -12, -13, -12, -11, -15, -7, -8, -12, -11, -10, -13, -11, -11, -3, -8, -2, -8, 0, 1, 2, 0, -4, 3, -3, -2, -5, -3, -1, -11, -11, -7, -14, -8, -7, -7, -8, -8, -13, -8, -5, -6, -7, -6, -8, -10, -9, -2, -5, 0, -3, 4, 3, 4, 1, 2, 0, 6, -1, 1, -2, -2, -11, -3, -11, -13, -9, -10, -11, -7, -8, -7, -13, -14, -12, -10, -2, -3, -1, -5, 0, 1, 7, 9, 4, 9, 3, 5, 9, 7, 6, 1, -5, -1, -8, -6, -10, -12, -5, -13, -15, -7, -9, -11, -5, -11, -8, -3, -3, -5, -1, -2, 5, 7, 7, 10, 12, 7, 12, 8, 4, 9, 2, 3, 0, 0, -3, -2, -8, -10, -9, -10, -7, -6, -7, -8, -7, -3, -7, -4, -5, -1, 0, 1, -1, 8, 11, 4, 4, 6, 6, 9, 2, 7, 2, 4, 6, 1, -1, 1, -3, -7, -10, -11, -5, -5, -11, -12, -11, -8, -6, -2, -1, -1, -2, 3, 4, 6, 2, 10, 4, 2, 11, 6, 4, 6, 7, 4, 4, -1, 0, -2, 1, -9, -1, -10, -9, -12, -8, -3, -3, -10, -2, -6, 0, 0, 0, -3, 1, 2, -2, 6, 8, 5, 4, 10, 9, 3, 2, 7, 3, 0, 0, -6, -2, -8, -8, -7, -8, -3, -9, -8, -7, -7, -2, -1, -1, 1, 0, -2, 3, -1, 0, 8, 3, 2, 3, 4, 7, 7, 1, 4, 5, -1, -5, 0, -7, -1, -8, -10, -3, -7, -3, -9, -2, -1, -10, -3, -5, 2, 0, 2, -2, -1, -2, 0, 2, 9, 7, 2, 8, 6, 0, 2, 0, 0, -4, -1, -4, -8, -4, -5, -10, -6, -9, -9, -1, -3, -6, -4, -1, -3, -1, 2, 0, 0, 1, 0, 0, 3, 2, 3, 0, 4, 1, 1, 0, 2, 0, -2, -4, -2, -5, -9, -8, -9, -1, -7, -4, -5, -8, 0, -6, 0, 1, 1, -3, -1, 4, 4, 3, 1, 5, 4, -2, 0, 3, -1, -1, 2, -1, -4, 1, -1, -3, -7, -3, -5, -1, -6, -4, -8, -1, -4, -5, -3, -3, -3, 0, 3, 1, 0, 3, -1, 3, 1, 3, -2, -3, -3, 2, -1, 0, 2, -2, -2, -3, -5, -1, -2, -1, -1, 0, -1, -3, -2, -2, -3, -3, -4, -3, 1, 0, 1, -1, 2, 2, 3, 5, 2, -3, -4, 1, -3, 3, -3, -3, -2, 0, -7, -5, -1, -1, -2, -2, -1, 0, -2, 3, 0, -2, 1, -2, 0, 3, 0, -1, 2, 0, 4, -1, 0, -3, 0, 0, 0, 2, 3, -3, -1, -7, -8, 0, 0, -1, -2, -5, -5, -4, -1, 0, 3, 3, 0, 0, 5, 2, 6, 2, 7, 0, 9, 0, -1, 2, 4, 3, 6, 0, 1, -3, -3, -5, -9, -8, -6, -4, -8, -8, -7, 0, -1, 4, 1, 8, 8, 6, 6, 7, 2, 11, 9, 9, 6, 1, 0, 0, 3, 0, 3, 2, 2, 1, 1, -1, -7, -6, -6, -7, -1, -9, -6, -5, 0, 0, 0, 6, 9, 13, 4, 5, 10, 9, 9, 11, 8, 6, 8, 9, 9, 8, 4, 8, 1, -2, -3, -2, -3, -9, -10, -3, -7, -6, -2, 1, -1, 0, 5, 3, 4, 12, 8, 7, 9, 7, 11, 5, 5, 1, 4, 9, 4, 6, 2, 8, 2, 3, 1, -2, -7, -1, -11, -9, -2, -4, 0, -1, -1, 0, 7, 2, 9, 7, 14, 9, 6, 9, 12, 7, 5, 9, 5, 9, 5, 9, 10, 6, 3, -1, 0, 0, -6, -7, -9, -3, -9, -3, -5, -4, -3, 2, 8, 7, 10, 6, 11, 17, 7, 12, 12, 6, 5, 6, 6, 11, 7, 9, 5, 5, 9, 4, -1, 2, -3, -10, -9, -8, -5, -9, 0, -5, 1, 0, 2, 9, 11, 13, 14, 9, 12, 10, 9, 9, 8, 8, 13, 5, 8, 7, 7, 7, 3, 4, 0, 2, -6, -5, -7, -10, -10, -4, 0, 0, 0, 2, 6, 8, 7, 10, 8, 14, 12, 10, 11, 14, 13, 12, 15, 16, 10, 11, 4, 5, 9, 5, -1, 1, -5, -1, -4, -10, -3, -2, -2, -2, -2, 0, 6, 3, 9, 6, 6, 6, 12, 10, 9, 5, 11, 11, 8, 13, 13, 9, 3, 6, 6, 4, 0, 0, 1, -7, -6, -9, -7, -5, -2, 0, -2, 1, 7, 2, 3, 5, 9, 13, 12, 5, 10, 7, 11, 7, 8, 8, 12, 2, 4, 9, 8, 11, 0, 2, -4, -10, -7, -13, -7, -2, 1, -2, -1, 6, 5, 7, 8, 15, 12, 7, 14, 5, 13, 10, 15, 12, 12, 7, 6, 8, 10, 8, 4, 3, 2, 0, 0, -9, -14, -11, -2, -6, -2, 3, 0, 5, 9, 9, 8, 13, 7, 11, 12, 7, 9, 12, 9, 8, 6, 6, 5, 10, 7, 11, 0, 6, 2, 0, 1, -2, -5, -11, -9, -1, 0, 4, 4, 1, 5, 4, 11, 6, 14, 6, 6, 7, 7, 10, 9, 9, 9, 4, 3, 8, 9, 5, 3, -1, -1, 0, -2, -9, -9, -3, -8, -7, -3, -1, 2, -1, 5, 6, 2, 7, 4, 10, 7, 11, 6, 3, 7, 5, 2, 8, 3, 6, 3, 6, 7, 5, 4, 0, -3, -4, -9, -7, -7, -6, -2, 0, 3, 1, 8, 4, 8, 10, 7, 5, 5, 10, 4, 1, 1, 7, 7, 8, 9, 2, 6, 5, 0, 3, 0, 0, -5, -8, -4, -8, -8, -3, 1, -5, -5, 3, 5, 3, 6, 5, 7, 2, 0, 4, 6, 6, 4, 6, 1, 1, 6, 1, 6, 0, 2, -2, 2, 1, -5, -9, -9,
    -- filter=0 channel=6
    3, 4, 7, 0, 3, 2, 7, 5, 8, 0, -1, -1, 2, 6, -3, -1, 0, 0, 2, -3, -2, -3, -2, 0, -1, 0, 2, 5, 3, 8, 7, 8, 6, 9, 7, 5, 2, 5, 9, 3, 1, 2, 3, 0, 7, 4, 4, -3, 0, 1, -1, 3, -1, 6, 6, 5, 5, 6, 6, 3, 1, 10, 6, 9, 4, 6, 3, 7, 8, 7, 9, 3, 1, 7, 4, 6, 4, 2, -1, 4, 2, 2, 1, 1, 3, 2, 6, 5, 2, 3, 10, 4, 2, 4, 0, 7, 6, 6, 5, 11, 2, 6, 5, 1, 1, 5, 0, 2, -2, 0, 4, 0, 0, -4, -2, -4, 0, 2, 3, 4, 1, 1, 3, 6, 4, 4, 6, 8, 4, 9, 3, 9, 2, 9, 9, 7, 0, -2, 6, 2, -3, 4, -2, -2, -1, 1, 0, -1, 4, 1, 0, 4, 6, 0, 3, 1, 2, 0, 4, 6, 10, 8, 9, 2, 6, 6, 8, 8, 6, 0, 7, 4, 0, 5, -3, 3, -2, 0, 3, 4, 8, 6, 6, 3, 6, 2, 6, 1, 2, 7, 10, 4, 6, 9, 7, 5, 2, 0, 6, 10, 7, 7, 6, 6, 2, 6, -1, 8, 5, 4, 6, 1, 8, 1, 8, 1, 6, 6, 1, 2, 8, 8, 4, 3, 11, 4, 7, 7, 2, 2, 6, 9, 1, 10, 0, 2, 7, 8, 7, 6, 3, 8, 4, 10, 2, 3, 2, 9, 5, 3, 4, 5, 8, 7, 5, 2, 10, 6, 4, 3, 8, 1, 8, 8, 6, 7, 6, 8, 6, 12, 9, 2, 7, 10, 13, 8, 11, 9, 7, 8, 10, 10, 4, 7, 1, 9, 8, 9, 8, 4, 5, 5, 4, 4, 0, 5, 1, 3, 9, 8, 15, 7, 8, 8, 12, 16, 10, 11, 12, 9, 11, 2, 9, 3, 1, 8, 3, 2, 0, 9, 8, 0, -1, 5, 7, 0, 0, 0, 0, 6, 6, 6, 8, 16, 13, 8, 17, 17, 12, 15, 12, 7, 12, 4, 2, 4, 1, 3, 2, 2, 3, 2, 5, -1, 0, -2, 0, 2, 6, 6, 0, 3, 4, 5, 11, 9, 9, 11, 16, 11, 13, 14, 14, 14, 10, 9, 5, 0, 0, 0, 2, -1, 3, 4, 1, 7, 2, 4, -1, 0, 3, -1, 4, 8, 3, 11, 16, 12, 19, 10, 9, 16, 12, 14, 5, 5, 6, 2, 6, -3, 0, 0, -5, -2, 3, 5, 3, 4, -4, -3, 0, 0, 2, -2, 0, 9, 9, 14, 12, 10, 13, 15, 16, 15, 12, 7, 11, 4, 3, 0, 1, -1, -3, 0, -5, 0, 4, 5, 2, 0, 0, -7, 1, -5, -9, 0, 3, 1, 9, 9, 12, 11, 10, 12, 12, 14, 16, 15, 10, 4, 3, 3, -2, -3, -1, -2, -5, 0, -1, 0, 2, -1, 0, -3, 0, -10, -3, -3, 1, 1, 1, 12, 13, 14, 19, 14, 12, 15, 7, 6, 5, 2, 0, -5, -10, -7, -7, -11, -6, 1, -3, -3, 0, -1, -3, -2, -6, -5, -5, -6, -10, -5, 5, 2, 8, 17, 16, 17, 15, 9, 13, 14, 7, 7, 4, -6, -5, -7, -6, -10, -3, -2, -2, 3, 0, -1, -2, -7, -7, 0, -11, -4, -4, -5, 1, 7, 7, 14, 17, 16, 19, 14, 19, 12, 4, -1, -6, -7, -7, -8, -7, -5, -7, -2, 3, 3, 3, 0, -2, -5, -5, -3, -9, -6, -1, -1, 1, 0, 8, 8, 16, 14, 12, 16, 13, 12, 3, 0, -4, -6, -11, -7, -2, 2, -2, 2, -3, 0, -2, 0, -2, 4, 0, 3, -3, 0, -1, -1, -4, 0, 7, 6, 16, 15, 11, 15, 15, 12, 1, -4, -8, -1, -3, -8, 0, -2, -1, -3, -4, 7, 1, -5, 1, 2, -2, 2, 0, -3, -7, -4, -1, -2, 7, 3, 14, 15, 14, 16, 10, 9, 3, 1, 0, -1, -5, 1, 0, 0, 1, -2, 0, 7, 0, 0, 0, -2, 0, 1, 2, -3, 1, -4, 0, -2, -2, 0, 5, 4, 8, 10, 4, 0, -1, -1, -2, -2, 0, 4, 0, 3, 3, 1, 1, 5, 3, 0, -2, 1, 2, 8, 5, 4, 2, 0, -3, 1, -2, 0, 0, 4, 4, 0, 4, -4, -1, 2, 0, -4, -1, -1, 0, 5, 0, 6, -2, 3, 0, -2, 0, 4, 0, 1, 1, 0, 2, 3, 1, 5, -2, -2, 0, -2, -2, 3, -5, -3, -2, 3, 0, -1, 2, 2, 7, 4, 7, 1, 4, 4, -2, 6, 2, -1, -1, 8, 6, 3, 3, 0, 5, 6, 3, 0, 2, 0, -1, 4, 1, 3, 0, 0, -1, -2, 3, 1, 2, 5, 3, 2, 4, 7, 3, 0, 0, 2, 4, 7, 8, 8, 6, 2, 6, 3, 4, 5, 3, -3, 3, 3, 4, 0, 5, 7, 5, -1, -1, -2, 6, 1, 2, 0, 3, 4, 3, 0, 5, 5, 1, 6, 9, 7, 5, 8, 3, 1, 0, 2, 1, 2, 2, 6, -1, -1, 2, 1, 6, 0, -1, 6, 1, 5, 5, 2, 9, 12, 2, 2, 7, 4, 5, 8, 1, 3, 5, 0, 4, 4, 0, -1, 3, -1, 7, 1, 1, 3, 1, 4, 5, 2, 1, 6, 2, 3, 6, 4, 5, 8, 4, 1, 3, 4, 3, 8, 0, 2, 2, 4, 0, 1, -1, 0, 0, 1, 3, 1, 8, 8, 2, 3, 2, 4, 6, 3, 3, 12, 10, 7, 2, 7, 0, 3, 1, 4, 6, 3, 2, 3, 1, 4, 0, 1, 0, 2, 0, 2, 2, 2, 6, 0, 3, 4, -1, 4, 3, 7, 10, 10, 4, 0, 6, 2, 4, 0, 5, 2, 0, 0, 0, -2, 1, 4, 1, 4, -4, 3, 4, 3, -2, 1, 3, 0, 3, -3, 0, 7, 4, 3, 5, 1, 3, 5, 10, 8, 5, 1, -1, 0, 4, 6, 0, 2, 3, -3, 0, -3, 2, -1, 0, 0, -4, 1, 4, -3, 1, 5, 1, 1, 6, 5, 8, 0, 5, 10, 6, 9, 8, 1, -1, 2, -2, 1, -1, 2, -1, -2, -5, 1, 1, 0, -3, 0, -1, -3, -7, 2, 0, 0, 0, -1, 2, 2, 3, 3, -3, 3, 3, 5, 2, 3, -2, 3, 4, -1, 0, -3, 3, 4, 0, 3, 3, -1, -1, 0, -2, 0, -2, 0, -4, -5, -5, 0, 2, 0, 1, 3, 3, 0, 5, 1, 6, 0, 0, 2, -1, 0, 3, 3, 3, -1, 3, 0, -5, 3, -2, 0, -5, -2, -3, 0, -4, -1, 0, 2, 5, 1, 0, 5, 4, 1, 5, 2, 2, 2, 5, 4, 5, 4, 5, -1, 2, 1, 3, 1, 0, 2, -3, -2, 1, 1, -7, 0, -4, 0, -2, 2, -1, 6, 4, 0, -3, -1, 0, 0, 1, 5, 7, 6, 2, 6, 6, 0, 3, -2, -1, 3, -3, 0, -2, -3, -4, -1, -2, -3, 0, -3, -4, -2, -1, 2, 1, 1, 3, 3, -1, 3, 7, 6, 0, 6, 3, 6, 0, 6, 0, -1, 2, 0, 2, 1, -5, -2, -6, -1, -1, -2, 3, -2, 0, 0, 0, -1, 3, 6, -1, -1, -1, 4, 1, 1, 6, -1, 0, 1, 3, 2, 6, 0, 6, 0, -1, 0, -4, 4, -5, 1, 4, 2, -1, 0, 0, 1, 2, 6, 6, 0, 0, 7, 4, 7, 8, 7, 5, 4, 5, 6, 5, 8, 0, 7, 5, 3, 6, 3, -2, 4, -5, 1, 1, 4, 1, -1, 4, 6, 7, 0, 3, 5, 4, 1, 0, 8, 0, 4, 5, 3, 5, 1, 1, 5, 0, 9, 3, 1, 9, 0, 4, 6, -1, 0, 6, 2, 8, 5, 2, 7, 2, 4, 6, 7, 8, 0, 0, 0, 3, 2, 4, 4, 2, 3, 4, 3, 2, 4, 3, 7, 8, 8, 8, 11, 8, 6, 5, 12, 4, 6, 3, 5, 6, 4, -1, 1, 6, 2, 3, 3, 8, 1, 1, 1, 2, 6, 6, 5, 3, 1, 4, 12, 14, 13, 15, 9, 15, 8, 10, 9, 7, 8, 10, 9, 1, 3, 5, 5, 3, 6, 3, 2, 3, 3, 1, -2, 5, 3, 4, 5, 8, 7, 7, 7, 12, 11, 17, 9, 9, 12, 14, 11, 7, 7, 4, 8, 1, 6, 0, 3, -2, 0, 0, 3, 8, 2, 2, -4, 1, 0, 7, 2, 3, 5, 8, 16, 13, 12, 16, 12, 13, 17, 12, 7, 14, 7, 5, 5, 6, 5, -3, 1, 3, 2, 3, 2, 2, 2, -5, 1, 0, 0, 0, 0, 1, 9, 12, 14, 18, 22, 15, 16, 17, 17, 20, 19, 10, 11, 7, 1, 2, 2, 1, -2, -4, 0, 4, 3, 0, -4, 0, -4, -5, -1, 0, 3, 8, 7, 14, 12, 17, 23, 19, 19, 25, 17, 17, 13, 13, 14, 4, 4, 2, -6, 1, -1, 0, -3, -3, 3, 0, -3, 0, -1, -6, -4, 0, -5, 0, 11, 9, 19, 18, 19, 24, 20, 16, 25, 16, 17, 18, 13, 12, 4, -4, -8, -2, -5, -2, -5, -3, -1, 4, -4, -2, -1, -3, -6, -6, 0, 0, 9, 15, 15, 16, 19, 23, 20, 22, 18, 20, 24, 20, 11, 8, 6, -5, 0, -1, -2, 0, 1, 2, 0, 4, -4, -6, 0, 0, 0, -7, -2, -1, 6, 8, 11, 18, 22, 21, 21, 22, 30, 20, 24, 21, 7, 3, 1, -3, -2, -7, -2, -1, -4, 3, -2, -1, 0, -4, 2, -4, -2, -3, -1, 0, -2, 6, 7, 16, 24, 25, 18, 25, 20, 23, 16, 16, 7, 3, 2, -1, 0, -1, -3, -1, -4, 0, -2, 0, -5, 1, -4, -2, 3, 0, -6, 1, -2, 2, 4, 12, 17, 16, 18, 21, 18, 17, 10, 12, 6, 0, 0, -3, 1, 0, 0, 2, -4, -4, 2, -4, 0, -4, -4, 4, 4, -3, 4, 1, 0, 4, 1, 10, 10, 10, 12, 20, 16, 16, 8, 1, 0, 5, 0, -2, 0, 3, 0, 1, -3, -4, 2, -4, 2, -2, 3, 0, -1, 3, -1, 3, 1, -4, 4, 6, 3, 5, 12, 7, 11, 10, 2, 2, 3, -1, 5, 2, 5, 2, 6, 0, 0, -4, 2, -1, 0, 0, 1, 4, 3, 0, -3, 1, 0, -2, -3, -2, 2, 3, 7, 7, 0, 2, 0, -2, 0, 4, 2, 3, 5, 7, 2, 6, -3, 0, 7, 1, -3, -1, 0, 4, 1, 2, 0, 0, 2, 2, 3, 4, 0, 0, -2, 2, -2, -2, -6, -4, 3, -2, 1, -3, 1, 4, 0, 2, 1, 0, 0, 3, 2, 4, -3, 3, -2, 2, -1, 2, 0, 4, -3, -4, 0, -2, -4, 0, 0, -5, -1, -4, 1, -3, 3, 2, 1, 6, 0, 7, 3, -1, 7, 0, 4, -2, -2, 1, 0, 5, 1, 3, 3, 1, 0, 0, -6, -8, -4, -2, -4, -7, 0, -1, -4, -4, -2, 2, 0, 1, 0, 3, 2, 3, 9, 3, 3, 0, 1, 2, 1, 5, -3, 4, -4, 2, -3, -5, -2, -2, -3, -4, 0, -5, 0, -4, -4, -3, 0, 0, -1, 2, 5, 0, 3, 3, 2, -1, -2, 3, 7, 0, 6, -2, -4, -2, 2, 0, 1, -2, -3, -4, -2, 2, -4, -5, -6, 0, 0, -3, 0, -2, -2, 6, 2, 0, 0, 5, 8, -1, -1, 6, 3, 7, 2, 1, 0, -4, 0, -4, 2, -4, -1, -3, -1, 1, 2, 0, 2, 2, -2, 0, -4, 2, 1, 1, 3, 0, 0, -1, 0, 4, 4, 3, -1, 2, 0, 4, -4, 0, -4, 0, -3, 0, 0, -7, 0, -6, -3, 0, -5, 1, 0, 0, -2, 0, 5, 6, 0, 2, 6, 5, 2, 3, -1, 1, 1, 4, 0, 0, -4, -4, -2, -7, 0, -1, -1, -5, -3, -4, -4, -6, -6, 0, -7, 2, -4, 4, 1, 0, 3, 0, 1, 0, 4, -1, 0, 0, 1, -1, 0, 1, 0, 0, -2, -9, -3, -6, -7, -3, -5, -6, -5, -1, -8, -5, 1, 0, -3, -2, 1, 3, 0, 2, 8, 2, 7, -5, -8, -6, -12, -10, -16, -10, -14, -11, -11, -9, -12, -8, -17, -12, -11, -12, -13, -14, -14, -13, -11, -8, -9, -14, -10, -13, -8, -8, -13, -9, -11, -11, -12, -9, -7, -9, -6, -8, -8, -12, -6, -10, -8, -13, -15, -10, -9, -10, -8, -11, -12, -9, -13, -7, -14, -14, -13, -10, -5, -7, -4, -4, -5, -3, -4, -10, -9, -12, -7, -13, -12, -13, -12, -10, -9, -9, -14, -14, -12, -9, -14, -16, -11, -12, -13, -15, -5, -11, -5, -3, -5, -9, -5, -6, -5, -5, -8, -5, -9, -10, -5, -12, -6, -9, -10, -15, -8, -10, -16, -13, -12, -11, -17, -15, -15, -15, -14, -10, -8, -5, -3, -2, -7, -6, -8, -3, -8, -2, -7, 0, 0, -7, -11, -7, -9, -10, -12, -7, -12, -11, -10, -12, -15, -11, -17, -15, -18, -10, -8, -7, -6, -9, -11, -10, -6, -4, -10, -8, -3, -5, -7, -4, -5, -8, -6, -4, -13, -7, -11, -14, -14, -10, -18, -19, -17, -17, -19, -18, -19, -10, -11, -14, -12, -11, -7, -10, -10, -10, -7, -2, -6, -5, -3, -3, -6, -7, -10, -7, -4, -11, -11, -10, -8, -10, -17, -17, -16, -18, -23, -15, -13, -14, -10, -10, -13, -12, -8, -7, -7, -7, -1, 0, 0, -5, 0, -7, -4, -9, -5, -11, -4, -5, -10, -16, -12, -10, -18, -14, -19, -18, -15, -18, -14, -18, -15, -9, -12, -8, -3, -5, -9, -10, -7, -2, 0, 0, 0, -1, -2, -5, -6, -5, -11, -7, -9, -11, -12, -12, -15, -19, -16, -22, -18, -21, -17, -12, -13, -16, -11, -8, -3, -9, -9, -1, 0, -7, 0, -1, 1, -9, -1, -1, -2, -7, -13, -5, -11, -14, -9, -16, -17, -18, -14, -13, -12, -18, -16, -9, -8, -15, -17, -7, -9, -8, -8, -4, -1, -5, -5, -3, -3, -3, 0, -7, -2, -5, -12, -8, -11, -10, -9, -12, -17, -11, -12, -13, -18, -16, -10, -13, -8, -10, -11, -10, -5, -7, -8, -3, -2, -3, -1, 4, 0, -2, 0, -8, -2, -12, -7, -8, -11, -15, -9, -9, -16, -17, -17, -15, -16, -14, -9, -15, -12, -10, -6, -9, -10, -8, -9, -2, -5, 0, -2, -1, -5, -7, -5, -3, -12, -4, -6, -9, -14, -8, -6, -8, -7, -14, -9, -9, -9, -8, -11, -9, -14, -9, -11, -13, -10, -5, -11, -2, -7, 1, -1, 2, -5, -7, -8, -9, -9, -14, -9, -11, -9, -10, -13, -4, -9, -14, -7, -6, -11, -9, -8, -7, -7, -14, -12, -9, -9, -6, -8, -6, -2, -2, -3, 5, 0, -8, -12, -9, -12, -8, -11, -10, -7, -6, -7, -11, -8, -11, -9, -9, -13, -10, -10, -12, -6, -12, -12, -10, -16, -14, -9, -8, -3, -6, 0, 0, 2, -3, -9, -5, -10, -10, -11, -15, -14, -11, -3, -3, -2, -1, -9, -8, -6, -3, -8, -10, -5, -6, -11, -9, -13, -7, -13, -10, -6, -4, 2, 0, -2, -7, -10, -12, -6, -14, -18, -15, -10, -11, -10, -3, 0, -5, 0, -4, -4, 0, 0, -8, -12, -6, -10, -15, -9, -12, -10, -7, -3, -6, 0, 0, -4, -7, -10, -10, -5, -13, -13, -9, -8, -9, -4, -5, -2, -3, -6, -5, 0, -2, 2, -4, -8, -11, -10, -10, -9, -5, -10, -7, -5, 1, -1, 2, 0, -5, 0, -5, -6, -12, -6, -12, -10, -6, -3, -4, -1, -4, -4, -3, 1, -3, 2, -6, -8, -13, -7, -15, -8, -12, -6, -6, -3, -2, -3, -1, -4, -2, -6, -1, -9, -12, -6, -11, -9, -10, -13, -5, -1, 2, 0, 0, 3, -5, -7, -5, -6, -11, -12, -9, -7, -4, -7, -5, -7, -4, 0, -2, -3, 0, -6, -7, -7, -3, -5, -7, -10, -11, -6, -3, -5, -7, -5, -2, -2, -1, -3, -6, -12, -13, -3, -5, -9, -5, 0, -4, 0, -2, 1, -2, -2, -2, 2, -1, 0, -8, -6, -10, -12, -11, -10, -10, -11, -11, -4, -5, 1, -7, -6, -6, -12, -12, -3, -3, -3, -2, -5, -5, -2, -3, -2, 1, 3, 3, 1, 0, 3, 0, -1, -7, -7, -8, -9, -8, -8, -9, -7, -4, -6, -11, -17, -12, -10, -5, -11, -4, -2, -5, -2, -2, -4, -2, 7, 3, 1, 0, 3, 0, 1, -3, -5, -2, -2, -7, -9, -7, -9, -8, -13, -7, -14, -11, -12, -9, -5, -8, -2, -2, 0, -2, -5, -3, -1, -3, -2, -2, 4, 0, 1, -1, 1, 2, 1, -4, -3, -3, -4, -5, -6, -13, -13, -8, -12, -8, -15, -12, -11, -9, -5, -5, -1, -7, -1, -3, -1, 1, 4, 0, 5, 0, -2, 0, 1, 2, -3, -2, 0, 0, -3, -5, -9, -6, -13, -12, -6, -9, -14, -11, -9, -10, -3, -5, -4, -4, 0, -1, 5, 4, 0, 1, 5, 0, 0, 2, 1, 1, -1, -1, -5, 0, -3, -6, -10, -3, -11, -8, -9, -11, -6, -4, -9, -1, -2, -7, -5, 0, 2, -1, -3, 4, 2, 0, 5, 1, 2, 0, 5, -3, 3, -6, -1, -3, -3, -9, -2, -9, -9, -3, -8, -4, -5, -1, -3, 0, -7, -3, 0, -2, 2, 3, -4, 0, 7, 0, 0, 6, 4, 2, -2, 4, 2, -2, -6, -5, -1, -4, -9, -9, -1, 0, -7, 1, -2, 1, -2, -4, -4, -2, 3, 3, 7, 0, 0, 3, 0, 3, 5, 7, 1, 3, -4, 0, 2, 2, -1, -2, -6, 1, -3, -1, -2, -6, -2, -7, 1, -2, -8, -5, -1, -1, 0, 1, 0, -2, 3, 2, 0, -1, 3, 0, 3, 2, 0, -3, -2, -4, 0, -1, -3, -4, 0, -4, -5, -1, -1, -2, -4, -5, -1, -1, 0, -1, 4, 2, 4, 0, -2, 1, 1, 1, 1, 4, 4, -2, -2, 1, 1, -3, 2, -3, -2, -5, -4, -5, -4, -3, -5, 1, 0, -2, 3, -4, -2, -2, 5, 0, 1, 6, 5, 0, 7,
    -- filter=0 channel=7
    -1, 6, 6, 1, 0, 1, 3, 1, 5, 1, 4, -1, -1, -1, 3, 2, -1, 1, 4, -1, 3, 3, 2, 3, 0, 3, 8, 0, 6, 1, 9, 5, 1, 0, 0, -3, -4, 1, -4, 3, -3, -3, 1, -1, 1, 2, -5, 3, -4, -4, 0, 3, 3, 0, -3, 0, -1, -4, -5, -1, 2, 3, -1, 0, 2, -2, -3, 1, -2, 0, -5, -2, -5, -5, 2, -4, 0, 0, -3, -3, -3, 1, -3, -3, 3, -3, -2, 1, 1, -2, -8, -7, -4, -1, 2, 0, -1, 0, -1, -7, 0, -1, -8, -3, -1, -5, -2, -3, 0, -1, -6, -3, 0, -6, -3, -3, -3, -3, -7, -7, -6, -2, -5, -9, -1, 1, 4, -1, 1, -3, -3, -7, -3, -6, -10, -4, -9, 0, -5, 2, -7, 0, 0, -6, 1, 0, 3, -2, -2, 0, -8, -5, -8, -5, -6, -3, 0, -3, -1, 0, -3, -5, -5, -1, -3, -6, -5, -7, -3, -3, -6, 2, -3, 2, -3, 0, -3, -3, -1, 0, -3, -1, -5, -9, -6, -3, -7, -6, 3, 2, -4, 0, -1, 0, -7, 0, -7, -5, -12, -3, -1, -7, 0, -2, -1, 5, 1, -1, 6, -2, 2, 0, -4, -2, 0, -3, -6, -9, 0, 0, -3, 2, -3, -4, -2, -3, 0, -7, -8, -9, -9, -11, -6, -1, -2, 2, 1, 4, 3, 7, 0, 0, 0, 3, 1, -4, 1, -7, -1, -4, -8, -8, -2, -3, -2, 0, -3, 0, -2, -2, -2, -5, -2, -4, -3, -6, -4, 2, 2, 0, 5, 8, 5, 2, 6, 4, -3, 1, 1, -6, -8, -8, -4, 0, -3, -3, 0, 1, 0, -5, -5, -7, -4, -5, 0, -1, -5, -4, 0, 4, 7, 0, 7, 6, 8, 3, 5, 2, 4, 3, 2, 1, -6, -3, -2, 0, -5, 1, -1, 0, -3, -5, 0, -3, -4, 0, 0, 0, -3, -2, -1, 6, 3, 7, 0, 7, 5, 4, 4, 0, 1, 0, 0, 2, 2, 1, 0, -2, 1, 4, 3, 2, 3, 0, 2, 0, -1, 0, 5, -2, -2, -4, 1, 1, 7, 3, 4, 6, 6, 5, 0, 6, 7, -1, 5, 1, -1, 6, 0, 5, 0, -2, -1, 3, 6, 2, 6, 0, 1, 4, 5, 0, -2, 3, 3, 7, 5, 0, 2, 5, 3, 7, 4, 6, 4, 3, 0, 1, 5, 2, -1, 5, 7, 2, 3, 6, 2, 2, 5, 5, 0, 6, 2, 5, -3, -4, 3, 2, 4, 4, 1, 0, 0, 1, -1, 2, 2, -2, -1, -2, 2, 4, 0, 0, 3, 8, 1, 2, 4, 10, 5, 8, 5, 2, 0, 1, 1, 0, -1, -2, -1, 2, 2, 0, 2, 1, -4, -3, 1, -5, -7, -3, -3, 3, 2, 6, 4, 9, 7, 9, 11, 7, 2, 8, 6, 0, 4, 3, -2, -4, 0, -2, -6, -7, -9, -3, -4, -5, -9, -4, -8, -4, -4, 2, 0, -1, -1, 0, 1, 2, 10, 12, 14, 9, 12, 3, 2, 1, 3, 4, 0, -2, -10, -9, -4, -13, -8, -12, -7, -15, -10, -14, -5, -11, -8, -5, -3, 0, 2, 0, 3, 4, 11, 6, 11, 13, 11, 6, 2, 8, 6, 0, -1, -1, -8, -8, -15, -14, -18, -15, -19, -16, -13, -12, -7, -10, -3, 2, 2, 2, -2, 0, 2, 6, 4, 13, 11, 10, 7, 10, 8, 6, 3, 3, -2, -5, -6, -10, -11, -13, -16, -12, -11, -20, -15, -13, -6, 0, 0, 0, 2, 0, 3, 7, 5, 4, 5, 7, 11, 11, 3, 7, 6, 0, 4, 6, 3, -2, -5, -2, -6, -10, -9, -3, -1, -10, -10, -5, -3, -2, 1, 4, 0, -2, 1, 6, 1, 6, 11, 11, 9, 4, 5, 2, 7, 1, 4, 6, 6, 1, -4, 2, -3, 2, 1, 8, 7, 3, 3, 0, -1, 2, 0, 6, 3, 4, 5, 5, 3, 7, 8, 13, 10, 7, 1, 4, 3, 8, 2, 2, 7, 3, 2, 5, 4, 3, 8, 15, 14, 9, 4, 1, 0, 7, 4, 7, 1, 4, 1, 2, 6, -1, 2, 7, 10, 9, 9, 9, 5, 3, 9, 10, 10, 8, 9, 3, 3, 4, 7, 17, 17, 15, 7, 7, 9, 8, 5, 10, 9, 0, 1, 5, 4, 4, 7, 5, 7, 7, 8, 0, 6, 1, 3, 5, 5, 9, 3, 7, 7, 5, 12, 16, 9, 9, 7, 12, 10, 5, 9, 3, 2, 7, 5, 0, 1, 3, 8, 10, 10, 6, 3, 4, 1, 8, 8, 11, 4, 8, 6, 7, 6, 11, 9, 8, 8, 9, 8, 11, 9, 11, 13, 9, 5, 5, 3, 4, 1, 0, 6, 4, 10, 2, 6, 5, 8, 12, 5, 5, 6, 5, 8, 6, 3, 7, 2, 10, 7, 12, 11, 10, 6, 8, 13, 8, 9, 5, 6, 2, 2, 4, 9, 7, 4, 2, 2, 1, 10, 8, 4, 7, 9, 2, 8, 1, 6, 1, 6, 12, 5, 4, 4, 4, 7, 7, 6, 6, 7, 4, 5, 3, 0, 3, 7, 8, 10, 5, 6, 4, 9, 6, 10, 4, 8, 3, 9, 5, 1, 5, 8, 7, 7, 7, 6, 7, 8, 2, 2, 1, 3, 6, 5, 0, 8, 1, 1, 9, 8, 0, 1, 5, 2, 4, 6, 8, 9, 5, 5, 0, 7, 7, 1, 4, 0, 3, 5, 4, 4, 10, 9, 5, 4, 9, 0, 2, 0, 6, 6, 1, 3, 1, 1, 8, 7, 2, 6, 6, 0, 7, 4, 1, 2, 7, 5, 1, 5, 8, 4, 2, 4, 5, 8, 7, 1, 0, 4, 6, 0, 3, 1, 9, 5, 4, 7, 7, 4, 7, 2, 0, 7, 3, 6, 2, 6, 1, 8, 5, 5, 0, 1, 6, 9, 8, 4, 3, -1, 5, 0, 2, 0, 6, 0, 3, 7, 7, 6, 4, 2, 4, 2, 10, 11, 9, 4, 8, 10, 10, 10, 5, 11, 9, 12, 11, 5, 3, 7, 7, 2, 7, 9, 2, 2, 3, 7, 10, 8, 3, 6, 11, 6, 6, 9, 6, 6, 9, 10, 8, 10, 4, 4, 8, 4, 7, 5, 9, 7, 12, 8, 6, 9, 13, 9, 11, 11, 12, 8, 8, 5, 7, 2, 7, 8, 8, 6, 9, 6, 5, 11, 7, 5, 2, 6, 8, 3, 3, 6, 8, 8, 8, 6, 4, 3, 9, 8, 5, 3, 5, 9, 9, 8, 9, 5, 0, 4, 3, 0, 3, 4, 3, 8, 6, 6, 2, 3, 5, 7, 0, 2, 6, 9, 3, 6, 5, 2, 1, 2, 0, 3, 5, 3, 4, 2, 1, 4, -3, 3, -5, 0, 1, 0, 3, 0, 4, 0, 4, -1, 2, 4, 7, 5, 4, 9, 0, -3, 0, 2, -3, -2, 3, -1, 3, 1, 9, 0, 2, 5, -2, 0, -5, -1, -1, 0, 1, 2, 1, -1, 0, 2, 3, 0, 5, 0, 6, 2, 2, -7, -4, -1, -4, -4, -3, 0, 6, 0, 0, 7, 1, -2, 0, 1, -1, -4, -4, -6, 0, 3, 3, 0, -1, 0, 0, 4, 2, 1, -3, -2, -6, -9, -9, -3, -6, -5, 0, 2, 6, 2, 3, 3, 2, 1, 0, -8, -12, -5, -8, -7, -3, -7, -4, -1, 5, 5, 6, 4, 3, 1, 1, -2, -9, -10, -7, -6, -9, -9, -6, -4, -1, 2, 0, 3, 4, -4, -7, -5, -9, -7, -9, -12, -8, -5, -1, -4, -1, 0, 1, 1, 4, -3, 1, -2, -10, -3, -6, -13, -4, -3, -5, -4, 5, 0, -1, 7, -1, -1, 0, -10, -5, -7, -10, -13, -11, -6, -9, -4, -4, -7, 0, -5, -3, -6, -1, -9, -8, -12, -6, -12, -9, -7, -4, -7, 0, 1, 6, 3, -2, -4, -3, -3, -1, -9, -8, -8, -13, -8, -9, -8, -3, -11, -6, -4, -4, -8, -1, -4, -10, -4, -9, -12, -9, -3, -3, -6, 3, -3, 0, 6, 0, -4, -5, -3, 1, -6, -7, -13, -15, -5, -10, -10, -12, -8, -10, -9, -6, -4, -12, -5, -7, -12, -6, -6, -6, -3, 1, -2, -1, 1, 3, 5, 2, 5, -1, -2, -3, -6, -11, -10, -8, -14, -11, -12, -9, -6, -14, -11, -7, -5, -6, -7, -11, -12, -8, -7, -6, -1, 2, 0, 0, 6, 6, 5, 3, 6, -1, 0, 6, 0, -9, -6, -15, -9, -10, -10, -7, -9, -15, -7, -12, -13, -10, -8, -11, -11, -10, -7, -7, 1, 1, 5, 4, 6, 0, 8, 5, 9, 5, 2, 0, 2, 0, -10, -7, -6, -13, -12, -7, -7, -14, -11, -15, -9, -8, -14, -15, -11, -10, -5, -6, -3, 4, 1, 9, 2, 4, 10, 5, 4, 6, 8, 4, 1, -4, -10, -4, -13, -10, -14, -13, -17, -11, -11, -11, -9, -16, -14, -9, -10, -10, -3, 1, 0, 5, 8, 3, 9, 10, 11, 10, 6, 4, 3, 7, 4, 2, 0, -6, -15, -9, -16, -14, -14, -20, -12, -15, -19, -16, -9, -13, -9, -10, -5, 3, -1, 5, 4, 10, 10, 14, 9, 10, 11, 12, 5, 6, 3, 0, -3, -7, -9, -17, -12, -16, -20, -19, -20, -19, -21, -19, -10, -15, -14, -9, -6, 1, 0, 4, 6, 6, 9, 10, 15, 12, 11, 6, 11, 2, 6, 1, -1, 0, -6, -12, -15, -15, -16, -19, -16, -20, -17, -20, -9, -6, -2, 0, 2, 0, 5, 8, 3, 9, 12, 9, 15, 14, 6, 11, 9, 7, 5, 6, 2, 0, -8, -8, -12, -18, -9, -10, -11, -14, -12, -16, -8, -7, -2, 3, -3, -2, 0, 2, 6, 3, 6, 11, 9, 9, 8, 7, 8, 3, 3, 10, 6, 4, 0, 0, -1, -7, 0, -3, -2, -4, 0, -5, -1, 0, 3, 1, 4, 0, 1, 7, 8, 10, 10, 12, 8, 6, 8, 4, 3, 2, 9, 7, 9, 3, 4, 3, 0, 3, 11, 12, 13, 6, 4, 6, 4, 7, 8, 8, 2, -1, 3, 3, 7, 7, 11, 13, 8, 8, 5, 9, 5, 6, 8, 10, 10, 9, 9, 11, 5, 12, 20, 16, 20, 15, 16, 11, 12, 10, 8, 5, 10, 1, 3, 2, 4, -1, 7, 10, 12, 6, 9, 0, 0, 1, 2, 11, 13, 13, 12, 12, 9, 14, 18, 20, 20, 21, 13, 10, 15, 10, 11, 12, 11, 1, 5, 4, 1, 0, 8, 3, 11, 6, 3, 7, 5, 4, 9, 9, 14, 8, 8, 11, 12, 13, 19, 15, 19, 18, 12, 10, 11, 15, 16, 6, 9, 5, 4, -1, 3, 5, 1, 7, 9, 1, 5, 0, 1, 2, 3, 6, 12, 14, 7, 7, 3, 9, 16, 14, 18, 10, 12, 13, 10, 7, 8, 7, 5, 7, 6, 0, 2, -2, 0, 2, 5, -1, 0, 0, 2, 5, 11, 9, 8, 4, 5, 7, 10, 8, 10, 12, 7, 15, 9, 4, 12, 8, 7, 15, 8, 6, 5, 4, -2, 4, 2, 4, 4, -2, -2, 6, 6, 6, 11, 11, 3, 4, 8, 6, 4, 2, 11, 14, 8, 4, 11, 7, 9, 3, 5, 7, 10, 3, 1, -3, -2, 0, 6, 1, 0, -1, 3, -2, 6, 0, 1, 5, 3, 9, 5, 8, 0, 5, 11, 5, 5, 8, 1, 5, 3, 4, 11, 1, 8, 2, 3, -1, 0, 0, 0, 4, 0, 6, 0, -1, 3, 5, 0, 7, 8, 3, 2, 5, 3, 5, 1, 9, 3, 4, 8, 6, 3, 7, 0, 5, 7, 0, 0, 1, -1, -1, 0, 2, 7, 1, -1, 4, 4, 0, -2, 3, 0, 3, 3, 0, 5, 0, 7, 7, 6, 3, 0, 6, 0, 3, 0, 5, 1, 0, 5, -3, 2, -2, 4, 0, 5, -2, 3, 0, 2, 5, 3, 1, -1, 4, 0, 4, 4, 4, 2, 3, 4, 2, 2, 4, 0, 0, 1, 2, 3, 1, 0, 0, -1, 0, -1, 5, 2, 0, 2, 0, 7, 7, 3, 1, 3, 5, 6, 2, 8, 2, 10, 4, 2, 3, 7, 7, 2, 7, 1, 2, 4, 1, 3, 0, 4, 2, 3, 5, 9, 13, 14, 17, 12, 15, 15, 17, 13, 13, 14, 13, 10, 14, 11, 9, 9, 11, 16, 17, 12, 9, 13, 11, 18, 16, 18, 11, 16, 11, 12, 20, 14, 8, 10, 7, 10, 14, 9, 12, 12, 15, 11, 16, 7, 8, 12, 13, 12, 7, 11, 6, 12, 6, 7, 15, 12, 10, 7, 7, 13, 8, 15, 15, 7, 8, 4, 7, 7, 8, 7, 11, 7, 9, 13, 8, 7, 6, 10, 10, 7, 4, 3, 13, 6, 7, 6, 8, 10, 3, 5, 5, 3, 5, 10, 8, 6, 11, 5, 0, 5, 0, 1, 2, 5, 7, 8, 7, 3, 4, 8, 5, 3, 6, 3, 5, 6, 3, 7, 3, 3, 1, -1, 3, 2, 5, 11, 7, 9, 6, 2, 5, -2, 3, -6, -2, 1, 6, 5, 4, 4, 5, 9, 6, 4, 7, 3, 2, 6, 6, 3, 3, 0, 1, -4, 0, 6, 0, 6, 7, 7, 5, 1, 0, 1, -6, 0, -3, 1, 0, 6, 4, 9, 5, 4, 5, 3, 4, 6, 4, 3, 5, -3, -1, 0, 1, -4, 4, 5, 7, 1, 3, 5, 4, 0, 3, -2, -6, -10, -4, -6, 0, 4, 0, 6, 1, 9, 10, 10, 2, 7, 3, 2, -2, 0, -1, -8, -5, -5, -3, 0, 3, -2, 6, 5, 0, -1, -3, -1, -4, -7, -12, -4, -1, -5, -3, 5, 3, 1, 5, 7, 3, 5, 0, 0, -4, 0, -4, -11, -8, -1, -8, 0, 3, 4, 0, -3, -1, -7, 0, 0, -6, -8, -12, -5, -12, -1, 0, 0, 3, 0, 0, -1, 4, 0, 2, -5, 0, -9, -8, -6, -2, -3, -7, -2, -4, -1, 0, 0, -4, -7, 0, -6, -3, -6, -10, -6, -7, -8, 0, -4, 1, 1, -4, 0, 1, -1, 0, -2, -2, -7, -3, -11, -5, 0, 1, 0, -4, -3, 0, 0, -3, -5, -7, -5, -2, -4, -7, -10, -5, -1, 0, -5, -5, -6, -2, -6, 0, -6, -3, -4, -10, -7, -5, -7, -1, -2, 3, -5, -4, -2, -1, 0, 0, 0, -3, -2, -4, -5, -6, -14, -8, -10, -9, -8, -4, -3, -5, -7, -2, -8, -2, -4, -4, -10, -7, -3, -3, 0, -2, -5, -4, 0, -4, -4, -4, -4, -2, -4, -1, -4, -5, -11, -7, -10, -7, -3, -4, -5, -6, -3, -8, -2, -7, -3, -11, -7, -11, -2, -1, -2, 2, 1, 1, -3, -3, 2, -1, 3, 0, 3, 3, -4, -4, -10, -5, -3, -7, -9, -2, -7, -9, -11, -10, -4, -8, -12, -9, -14, -15, -10, -3, 2, 0, 0, -3, -5, 1, 3, -1, -1, 1, -3, 0, 1, -5, -9, -9, -11, -12, -12, -10, -7, -9, -7, -12, -11, -12, -11, -12, -11, -6, -8, -4, 0, 3, -1, 2, 0, 2, 4, -3, -4, 0, -1, -3, -2, -7, -8, -8, -13, -13, -15, -9, -14, -17, -12, -12, -14, -15, -14, -10, -16, -4, -9, -3, -5, -4, 2, 1, -1, -2, 0, -3, 0, 4, 3, -2, -4, -2, -1, -4, -12, -14, -16, -21, -17, -19, -13, -15, -12, -19, -15, -11, -12, -11, -6, -9, -1, 1, 0, 1, -2, 5, 0, 0, -2, -3, -1, -1, 0, -4, -8, -8, -15, -15, -16, -16, -20, -21, -15, -21, -18, -20, -18, -8, -8, -8, -4, -1, -8, -3, 0, -3, -4, -1, 0, -1, -6, -3, 0, -1, -1, -3, 1, -3, -13, -11, -11, -13, -15, -12, -13, -15, -14, -10, -12, -5, -6, -6, -2, -1, -6, -6, -3, -4, 0, -5, -3, -4, -4, -3, -3, -1, 0, -2, 2, 0, -3, -4, -10, -9, -9, -3, -11, -8, -5, -6, -7, -5, -4, -6, -8, -9, 0, -1, -6, -8, -5, 3, -7, -9, -6, -8, -3, -2, 0, 1, 3, -2, -2, -2, -2, -1, -4, 1, 3, 0, 2, 0, -2, 0, -1, -6, -8, -5, -2, -7, -5, -9, -9, -5, -6, -4, -7, -10, -1, 0, -6, -4, -4, -2, -1, 0, -4, 0, 1, 5, 4, 0, 0, -5, 0, -2, 0, -4, -6, -4, -10, -4, -8, -8, -6, -3, -1, -9, -8, -11, -4, -2, -7, 0, 1, -4, -1, 0, -5, 2, 5, 7, 3, 6, 5, -3, -4, 0, -1, 1, -5, -1, -6, -10, -12, -9, -5, -3, -10, -7, -6, -13, -5, -2, -1, -5, 0, -4, -1, -2, -7, 1, -1, 1, 0, 0, 3, 3, -5, 0, 0, -3, -4, -9, -12, -10, -15, -14, -9, -10, -11, -12, -13, -14, -12, -2, -5, -4, 1, -1, -8, -2, -6, -3, -5, 3, -5, 0, -5, -5, -3, -1, -2, -7, -2, -4, -8, -11, -13, -11, -10, -5, -7, -13, -9, -9, -7, -8, -2, -3, -2, -1, -10, -7, -2, -7, 0, -4, -3, -6, -5, -2, -2, -5, 0, 0, -3, -9, -11, -16, -9, -16, -9, -8, -7, -14, -10, -15, -6, -5, -9, -5, -4, -9, -4, -10, -6, -4, -8, -1, -2, -7, -8, -5, -10, -9, -7, -6, -8, -4, -6, -13, -15, -14, -13, -14, -9, -18, -10, -15, -9, -8, -10, -8, -11, -3, -5, -6, -7, -9, -8, -7, -8, -5, -4, -5, -6, -9, -9, -6, -5, -5, -12, -7, -15, -16, -18, -16, -13, -10, -12, -16, -7, -13, -14, -6, -11, -12, -9, -6, -7, -10, -12, -8, -7, -10, -14, -11, -12, -12, -12, -14, -11, -5, -16, -8, -16, -11, -13, -9, -16, -10, -16, -15, -11, -12, -8, -11, -11, -12, -9, -6, -15, -14, -12, -11, -7, -8, -15, -16, -15, -8, -8, -12, -13, -8, -15, -15, -11, -14, -16, -10, -12, -15, -19, -16, -16, -13, -11, -16, -11, -13, -9, -10, -9, -15, -8, -14, -7, -7, -15, -17, -11, -14, -14, -15, -17, -10, -17, -17, -12, -16, -18, -16, -11, -15, -16, -13, -15, -13, -7, -13, -7, -13, -14, -6, -14, -6, -10, -4, -6, -12, -6, -14, -14, -8, -15, -13, -8, -8, -9, -9, -11, -14, -14, -11,
    -- filter=0 channel=8
    -1, 2, -4, 0, -1, -1, -2, -2, 0, -6, -2, -5, -6, 1, 0, 0, 0, -2, -4, -2, -2, 0, -2, -6, 0, 1, 1, -2, -3, 2, 0, 4, 3, 3, 0, -4, -5, -7, -5, -2, 0, -4, -5, -5, -3, -4, -4, -2, -2, -3, -6, -5, -3, -2, -5, 0, -6, -5, -1, -1, 2, -2, -1, 0, 1, -3, 1, 0, -3, -2, -2, 1, -4, 0, -8, 0, -5, 0, -4, -1, -4, -2, -2, -4, -1, -2, 0, -4, -2, -4, 1, -2, -5, 3, 3, 2, -5, -3, -3, 0, -6, -5, 0, -1, -3, 0, -8, 0, 0, -5, -6, -2, -4, 0, -3, 0, -6, -2, -5, 0, -2, -7, 0, 1, 2, 2, -5, -3, -1, -2, -7, -1, 0, -5, 0, -5, -4, -8, -2, -3, -4, -8, -6, -7, -6, -1, 1, 0, -2, -6, -4, 0, -5, 0, -5, -1, -6, 0, -2, 1, -5, -8, -6, -2, -1, 1, 0, -2, -5, -1, -4, -6, -6, -9, -5, 1, -5, 0, -1, -5, -2, -1, -5, -7, 0, -5, -2, -4, -6, -4, -2, -2, -2, -3, -4, -1, -4, -3, 0, 0, -2, -7, -8, -2, -5, -7, -3, -3, -5, -1, 0, -6, -5, -6, -7, -1, -1, -4, -3, -4, -6, 0, -4, -3, -5, -3, 0, -6, -3, 0, 0, -5, 0, -8, 0, 0, 1, -1, -5, -2, -3, -1, 2, 3, -4, 0, -1, -4, -1, -7, -5, -2, -8, 0, -6, -4, -7, -10, -9, -3, -8, -1, 0, 1, 0, -6, -5, -5, -6, 0, -2, 4, 0, 1, 3, -2, 4, -4, 1, 0, -5, -3, 0, -3, 0, -1, -1, 0, -6, -10, -2, -4, -2, -1, -6, 1, 0, 3, 1, 0, 0, 4, 1, 6, 1, 1, 0, -3, -1, -3, 2, -2, -3, -5, -7, -1, -4, -2, -5, -3, -9, -11, -10, -8, -2, -5, -7, -4, 0, -2, 0, 0, 6, 3, 3, 0, 5, -1, 3, 4, 3, -3, -1, -4, 0, -6, -8, -3, -4, -7, -4, -1, -12, -10, -6, -4, -4, -1, -2, -4, -2, 2, 0, 1, 3, 0, 4, -1, 0, 3, 0, -2, 2, -2, -1, -5, 0, -5, -3, -4, -2, -8, -2, -2, -5, -13, -10, -12, -9, -5, -2, -4, 4, 0, 1, 4, 3, 0, 3, -3, -2, 5, -2, -1, -3, -3, -3, -3, -4, -6, -2, -6, -11, -11, -4, 0, -8, -6, -9, -8, -5, -3, -1, 0, 4, -3, 5, 6, 0, -1, 5, -4, 0, 3, -2, 3, -3, 0, 0, 1, -5, -8, -2, -6, -7, -6, -7, -5, -3, -3, -8, -9, -8, -5, -1, 2, -1, 0, -4, 2, 0, -2, -5, 0, 0, 0, 1, -3, -6, 0, 2, -1, -6, -5, -4, -4, -8, -10, -6, -7, -8, -5, -2, -3, -5, -8, -2, 0, -3, -2, 1, -2, -1, -5, -6, -6, -3, -2, -4, -7, -4, 1, -1, -1, 0, -6, -4, -7, -10, -4, -9, -8, -10, -12, -12, -3, -6, -5, 0, 2, -1, 0, -2, -4, -5, -4, 0, -1, 0, 0, 1, -2, -3, -1, -2, -2, -2, -2, -8, -10, -6, -11, -8, -3, -7, -10, -4, -3, -3, -6, 1, -2, 0, 2, 3, 1, -4, -3, -4, 2, 2, 4, 0, 1, 6, 1, -3, 0, -1, -5, -1, -4, -3, -2, -3, -1, -8, -4, -7, -7, 0, 0, 0, 4, 4, 5, 5, 0, 0, 0, 2, 3, 5, 10, 2, 7, 0, -1, 4, 3, -1, -2, 1, 0, -7, -7, -6, -2, -7, -9, 0, -1, -2, 0, -3, -2, 4, 1, -1, 3, -3, -1, 2, 5, 5, 10, 9, 7, 6, 0, -1, -1, 0, 0, -3, -1, -4, -4, -4, -2, -4, -3, -8, -2, -4, 0, -2, 2, -3, 3, 1, 0, 1, -2, -2, 6, 1, 1, 0, 5, 5, 2, 3, 3, 3, 0, 3, 3, -2, -4, -3, -4, -13, -2, -6, -4, -1, -1, 0, 0, 3, 0, 1, 2, 0, 6, 0, 7, 8, 5, 6, 0, 1, 4, 5, 2, -2, 0, -2, 4, -3, 0, -8, -4, -7, -8, -4, -6, -1, 0, -2, 2, -3, 4, 0, -2, 1, 1, -1, 6, 5, 3, 5, 2, 1, -1, 3, -1, 0, -2, -4, -2, 1, -6, -5, -13, -15, -4, -2, -4, 0, 0, 1, -4, 2, 0, 3, -2, 0, 2, 0, 0, 0, -5, -1, 0, -3, 2, -5, -1, -5, -5, 0, -3, -6, -7, -11, -11, -11, -11, -6, 0, -2, 2, -2, 0, -2, 0, -2, -1, 4, 1, -4, 0, -6, 0, 0, -1, -6, -2, -1, -4, 0, -4, -4, -6, -9, -11, -12, -12, -16, -16, -4, -3, -3, 2, 0, -5, 0, 0, 1, -1, 0, -2, -2, -3, -1, -1, 0, -7, -3, -1, -9, -7, -4, -10, -6, -5, -8, -13, -17, -13, -19, -17, -12, -3, -1, -5, -7, -8, -3, -3, -8, -5, 0, 0, -2, -6, -7, 0, -6, -6, 0, -7, -6, -7, -5, -11, -6, -7, -7, -10, -17, -15, -22, -20, -15, -11, -10, -10, -8, -10, -5, -4, -11, -11, -8, -9, -3, -8, -5, -11, -7, -7, -6, -7, -7, -9, -10, -11, -9, -14, -13, -11, -15, -15, -20, -17, -15, -9, -14, -7, -8, -13, -7, -9, -13, -12, -5, -6, -9, -8, -11, -8, -6, -8, -5, -8, -10, -14, -9, -11, -9, -16, -12, -20, -18, -19, -23, -22, -14, -16, -20, -13, -12, -12, -16, -10, -13, -15, -13, -12, -16, -17, -15, -9, -10, -9, -8, -13, -12, -18, -12, -15, -22, -18, -16, -24, -25, -26, -22, -27, -21, -17, -24, -22, -20, -17, -13, -22, -18, -18, -15, -18, -21, -15, -17, -12, -15, -19, -15, -18, -19, -23, -21, -20, -25, -20, -19, -25, -21, -21, -27, -24, -30, -21, -28, -20, -22, -28, -19, -24, -27, -26, -23, -25, -26, -27, -19, -20, -27, -27, -27, -22, -22, -29, -28, -26, -31, -30, -31, -22, -23, -23, 2, -2, 5, 0, 3, 4, 3, -2, 3, 1, 2, -3, 0, 2, 3, -1, 1, 0, 0, -2, 0, 1, -3, 0, 0, -1, 2, -2, 2, 3, 3, 0, -1, -2, 0, -2, 5, 0, -2, -2, -3, 0, 1, 0, -5, 1, -1, 3, -3, 1, 1, 0, 0, -2, 1, -4, -3, 3, -4, 0, 0, 0, 6, 0, 1, -1, 3, 3, 3, 5, 4, 1, 2, 0, -1, -2, 0, -3, -2, -3, 2, 3, 0, 0, 4, 5, 0, 1, 2, 2, 3, 1, 2, 5, 5, 0, 0, 2, -2, 3, -2, 5, 2, -2, 3, 1, 4, 0, 5, 1, 0, 1, -2, 2, 0, 3, 2, 1, -2, 1, 3, 3, 0, 4, 2, 0, -1, 5, 3, 3, -4, 0, 0, 4, 0, 1, 0, 0, -4, -1, 2, 3, 1, 5, 2, 4, -2, -2, 1, 2, 2, -2, -1, 4, 0, -2, -1, 0, 4, 2, 0, -1, 1, 0, -1, -1, 6, 0, 0, -1, 1, -4, 0, 4, 2, 0, 0, 1, 5, 0, -1, 2, -4, 2, 1, 1, 1, 0, 0, -3, -2, 1, -2, -4, 0, -2, 2, 6, 0, 5, 3, 4, -4, 2, 5, 5, 5, 3, -2, 0, 2, 3, 2, 4, 1, 1, -1, 1, 2, -1, 0, -4, -2, 2, 2, 0, 3, 1, 1, -1, 1, 3, 1, 0, 1, -2, 0, 7, 8, 1, 6, 0, 3, 1, 1, 1, -1, 3, 0, -2, -2, -1, 1, -1, 2, 2, -6, 2, -4, 4, 1, 2, 0, 3, 3, -1, -1, 5, 6, 1, 6, 0, 4, 1, 7, 8, 3, 6, 0, 5, -1, 5, 3, -2, 2, -3, -2, 0, -1, -5, 0, -1, 2, -2, 4, 5, 7, 8, 1, 5, 2, 2, 10, 2, 0, 4, 7, 4, 2, 6, 4, 4, 3, 4, 3, 0, -2, 2, 4, -1, 0, 0, -2, 3, 2, -3, 1, 0, 6, 2, 4, 8, 10, 9, 9, 5, 0, 5, 6, 1, 4, 5, -3, 3, 0, 5, 0, 2, -3, 0, -2, -3, -5, -4, -1, -2, 0, 3, 0, 6, 4, 2, 5, 9, 10, 3, 2, 3, 3, 2, 2, -3, 3, 3, 1, 4, 6, -2, -1, -1, 4, 0, 1, 0, -4, -8, 0, -3, -2, 1, -2, 0, 6, 2, 4, 4, 6, 2, 4, 0, 5, 7, 1, 4, -1, -2, -2, 1, 0, 4, -3, -4, -3, -3, -2, 4, -2, 2, 2, 1, -1, 2, -1, 6, 3, 6, 1, 4, 4, 2, 0, 2, 1, 5, 2, 6, 3, -2, 4, 0, 5, 2, 0, -3, 0, -2, 0, 4, 2, 0, -2, 2, 3, 1, 3, 2, 3, 4, 1, 2, 4, -2, -2, -3, -2, -2, -1, 2, 0, 0, 4, 1, 1, -1, -3, 0, 0, -3, -3, -2, -1, 1, -4, -3, 0, 3, -2, 6, -1, 3, 5, 6, 0, -3, 0, -1, -4, -4, 3, -5, 3, -2, 2, 6, 0, 0, 0, 0, -6, 2, -3, 2, 3, -2, 2, -1, 2, 3, -1, -3, 4, -1, -4, -3, -4, -3, 1, 0, 1, 5, 1, 1, 1, -2, 2, 2, 0, -2, -3, -3, 0, 3, 1, 2, 1, 1, -6, -5, 0, 0, 0, 0, -3, 2, 1, 0, 3, 0, 3, 0, 1, 4, 2, 4, -1, -2, 0, 0, 0, 0, -2, 0, -2, 0, 2, 7, -1, 0, -3, 3, -3, 4, 2, -1, -2, 6, -2, 2, -3, 0, 4, 1, 9, 1, 3, 7, 8, -1, 5, 0, 0, 3, 3, -1, -2, -2, 0, 0, 5, -4, 2, 2, 1, -4, -2, 0, 0, 2, 3, 1, 1, 3, -4, -1, 5, 8, 2, 5, 4, -5, 2, -3, 3, -1, 1, 2, -3, 0, -2, 8, 6, 0, 0, 3, -2, -1, -1, 1, 0, 1, 2, 0, 1, -4, -4, 4, 1, -1, 4, 4, 0, 1, -2, -2, -5, 2, 0, 5, 0, 5, 4, 6, 3, 3, 0, 1, -5, -2, -7, -3, -4, -4, 1, 1, -3, 4, 2, -2, 6, 5, 0, 3, -2, -3, 0, 4, -3, 3, 1, -1, 3, 6, 6, 5, -3, 4, 7, 2, -4, -7, -4, -1, -2, -3, -2, 0, -2, 1, 0, 1, 1, 1, 1, 0, -2, -1, 4, 0, -3, 0, -2, 1, 3, 4, 0, 1, 1, -1, 0, 0, 1, 1, 0, 0, -3, -5, 0, 1, -6, 2, -4, 0, -1, -2, -2, -5, -4, -2, -3, -1, 1, 1, 2, 0, 5, -1, 3, 3, -6, 3, 5, 4, 4, -2, -4, 3, -3, 0, -3, -4, 2, 2, 1, -7, -4, -5, -5, -6, -7, -6, -7, -6, 1, -1, -5, -5, 0, -4, -1, 0, -3, 0, 5, 0, 4, 3, 3, -4, 0, -1, -4, 1, -3, -4, -4, -5, -4, 1, -5, -1, -4, -4, -7, -2, -1, 0, -4, 3, 4, -3, -3, 0, -6, 0, 4, 1, 5, 6, 5, 2, 0, 2, 0, -6, -5, 3, 0, -2, -4, 2, -3, -1, 0, -5, -3, 0, 1, -5, -2, -2, 2, 1, 0, -4, -10, -1, 0, 0, 0, -2, 4, 2, -1, 1, -1, -3, -3, -2, 0, 0, -3, 0, -6, 1, -3, 0, -1, -2, -4, 0, 2, 0, -2, 0, -9, -3, -7, 0, -4, 0, 0, 4, 3, 0, -5, -2, 0, -3, -5, -7, 0, -1, -5, 0, 0, -5, 0, -4, 0, -6, -5, -2, -5, 1, -2, -6, -3, -10, -10, -2, -4, -2, -7, -1, -7, 0, -6, -8, -7, -6, -7, -1, -3, -7, 0, -7, -6, -3, -2, -8, -2, -7, -5, -5, -11, -4, -7, -2, -3, -3, -12, -5, -3, -5, -10, -4, -9, -7, -7, -8, -7, -9, -5, -11, -8, -11, -6, -3, -3, -4, -8, -5, -5, -9, -7, -5, -4, -5, -8, -9, -8, -7, -9, -6, -6, -13, -8, -13, -9, -11, -8, -13, -13, -15, -10, -10, -11, -14, -10, -9, -14, -9, -13, -10, -12, -13, -9, -12, -13, -13, -12, -11, -10, -7, 5, 13, 8, 8, 9, 9, 3, 6, 8, 10, 10, 6, 2, 9, 7, 9, 6, 8, 3, 2, 2, 5, 4, 5, 9, 6, 8, 4, 6, 9, 9, 15, 9, 11, 12, 14, 12, 5, 5, 10, 3, 3, 2, 4, 7, 9, 6, 9, 4, 5, 5, 3, 5, 9, 7, 5, 10, 4, 10, 9, 10, 7, 6, 6, 5, 4, 7, 12, 9, 12, 5, 11, 4, 8, 2, 5, 4, 10, 11, 7, 11, 6, 12, 5, 12, 10, 2, 11, 5, 4, 8, 5, 8, 11, 5, 10, 8, 8, 7, 8, 10, 13, 7, 11, 4, 9, 10, 10, 9, 6, 4, 10, 12, 8, 10, 8, 11, 8, 9, 3, 7, 2, 5, 8, 9, 8, 10, 8, 11, 4, 4, 5, 9, 13, 10, 7, 6, 7, 10, 5, 6, 8, 8, 8, 3, 8, 10, 11, 7, 2, 3, 10, 8, 4, 3, 10, 11, 8, 7, 7, 3, 4, 4, 13, 6, 7, 5, 8, 11, 5, 2, 3, 3, 8, 5, 9, 7, 11, 8, 2, 7, 8, 4, 5, 9, 3, 8, 12, 4, 5, 3, 8, 11, 12, 4, 6, 11, 7, 6, 9, 9, 5, 8, 3, 8, 6, 4, 2, 6, 3, 8, 7, 8, 8, 3, 6, 3, 10, 8, 4, 5, 7, 9, 2, 11, 3, 9, 8, 7, 7, 11, 5, 8, 4, 5, 6, 5, 6, 10, 8, 4, 5, 8, 10, 4, 9, 10, 10, 8, 3, 7, 3, 6, 2, 7, 5, 7, 4, 5, 7, 13, 10, 12, 14, 9, 6, 6, 7, 9, 7, 3, 8, 3, 8, 3, 9, 3, 5, 9, 8, 11, 7, 10, 6, 3, 9, 9, 7, 5, 4, 5, 6, 9, 5, 13, 7, 11, 8, 11, 13, 12, 3, 8, 4, 5, 3, 3, 7, 10, 8, 11, 9, 10, 4, 8, 6, 3, 4, 10, 12, 9, 3, 6, 8, 6, 5, 4, 11, 6, 5, 13, 15, 6, 11, 3, 9, 8, 4, 8, 1, 8, 3, 8, 10, 4, 10, 7, 9, 9, 5, 12, 5, 8, 5, 2, 8, 5, 4, 7, 12, 10, 8, 7, 13, 13, 5, 8, 4, 9, 3, 9, 1, 5, 1, 8, 7, 4, 2, 2, 2, 10, 4, 9, 7, 4, 4, 2, 8, 11, 9, 5, 7, 12, 11, 5, 11, 6, 9, 0, 5, 5, 2, 2, 7, 3, 5, 1, 8, 4, 8, 6, 1, 7, 3, 6, 7, 9, 11, 9, 6, 7, 6, 4, 8, 4, 10, 7, 7, 10, 8, -1, 1, -3, 0, 4, 7, 3, 0, 3, 8, 5, 5, 6, 7, 8, 7, 9, 13, 8, 8, 6, 7, 10, 5, 1, 3, 8, 1, 6, 8, 5, -1, -1, -1, -3, 4, 2, 1, 7, 6, 6, 4, 9, 6, 1, 9, 2, 6, 6, 9, 15, 8, 4, 6, 8, 1, 1, 5, 5, 8, 6, 2, 0, 1, 0, -2, -4, 0, 0, 1, -1, 0, 1, 7, 1, 2, 1, 3, 2, 8, 8, 14, 14, 6, 5, 2, 3, 9, 5, 4, 3, -2, 1, 0, -1, 2, 2, 2, 3, 5, 0, 0, 0, 2, -1, 4, 7, 2, 2, 0, 3, 2, 13, 13, 16, 6, 4, 5, 2, 0, 3, 4, 4, 5, 3, 3, 5, -1, 6, 0, 3, 2, 2, 4, 0, -2, -1, 1, 1, -3, 2, 5, 8, 5, 7, 12, 14, 9, 7, 10, 1, 0, 7, 3, 0, 3, 5, 3, 0, 4, 0, 3, 8, 7, 3, 0, 0, -1, 4, -3, 2, 2, 0, 0, 4, 10, 15, 12, 15, 14, 11, 9, 0, 4, 4, 3, 0, 3, -4, 2, -1, -1, -3, 0, 5, 2, 3, 0, -2, 1, -1, 0, -3, -1, 4, 5, 8, 9, 15, 13, 13, 17, 10, 5, 0, -2, 2, 1, 2, 2, -2, -1, 0, 2, 0, 2, 3, 2, 1, 4, 1, 0, 0, 2, 2, 1, 6, 0, 6, 11, 15, 18, 14, 9, 10, 4, 1, 4, -3, -3, -6, 0, -4, -3, -3, -4, -1, 3, 3, 2, 0, 0, -1, -5, 1, -4, -2, 3, 0, 6, 6, 7, 9, 17, 18, 10, 13, 7, 0, -2, -3, -1, 1, -5, 1, 2, 0, -4, 1, 1, 2, 1, 2, -1, -3, -3, -1, -3, 0, -1, -2, 4, 10, 13, 16, 14, 10, 16, 14, 9, 10, 2, -1, 1, 3, -1, 0, 2, -1, 2, 0, -1, -6, -8, -7, -6, 0, 0, -1, 0, 4, 1, 4, 5, 6, 10, 14, 9, 11, 15, 11, 9, 13, 5, 0, 6, 2, 0, 0, 2, 0, -3, -1, 0, -8, 0, -1, -4, -5, 0, 0, 0, 3, 4, 4, 9, 4, 10, 12, 11, 12, 12, 9, 9, 14, 11, 3, 4, 0, 3, 3, -1, 2, 1, 0, 4, 1, -1, -4, 0, -1, 2, 1, -2, -2, 6, 5, 10, 7, 8, 9, 16, 12, 14, 12, 12, 10, 10, 6, 6, 4, 4, -1, -1, -1, 0, 0, 1, 3, 2, 1, 3, 4, -1, 0, 3, 4, 5, 10, 9, 9, 7, 10, 14, 10, 10, 12, 16, 13, 6, 4, 5, 8, 1, -3, -2, 4, 3, 0, -1, 0, -1, 6, 3, 5, 2, 6, 0, 7, 9, 4, 10, 11, 12, 13, 6, 7, 10, 8, 13, 15, 12, 5, 6, 5, 2, -1, 4, 5, 6, 4, 0, 0, 1, 4, 3, 0, 2, 7, 1, 0, 1, 2, 8, 7, 15, 7, 7, 10, 9, 14, 5, 10, 4, 2, 7, 6, 4, 0, 5, -1, 0, 0, 3, 2, 6, 2, 1, 6, -1, 1, 4, -1, 7, 2, 4, 11, 9, 8, 6, 6, 3, 12, 4, 8, 2, 3, 3, 5, 2, -2, -1, -3, -2, 1, 2, -3, -1, 4, 0, 0, 5, 5, 2, 1, 0, 4, 7, 4, 9, 9, 4, 4, 5, 3, 1, 3, 0, 0, 3, 2, -4, -6, 0, -5, -2, -6, -3, -4, -6, -3, -2, -2, -2, -1, -5, -3, -2, 0, -1, 2, 2, 3, 2,
    -- filter=0 channel=9
    1, 3, 0, 5, 6, 8, 0, 8, 8, 3, 5, 3, 0, 3, 6, 3, 8, 8, 2, 5, 7, 4, 6, 1, 5, 1, 0, 6, 5, 0, 5, 2, 4, 3, 0, 3, 5, 5, 0, 0, -1, 2, 2, 0, 1, -3, 3, 2, 2, 1, -1, 4, 5, 0, 1, 2, 0, 3, 6, 4, 0, 3, 4, -2, 2, -1, 6, 0, 0, 5, 5, 0, -4, -1, -2, -8, -6, 0, -6, 0, -1, 3, -5, 1, -3, -5, 0, -5, 2, 4, 3, 1, 2, -1, 0, 0, 6, 4, 4, 6, -1, 3, -3, -2, -2, -1, -8, -2, 0, -7, -5, 0, -3, -3, -9, -3, 0, -9, -6, -4, 1, -1, 3, 2, 0, 0, 5, 2, 1, 5, 4, 0, 0, -1, 0, 0, 3, -4, -7, 0, -1, -5, -4, -4, 0, -4, -1, -6, -7, -1, -5, -1, -2, 0, 2, -1, -2, 5, -3, 1, 7, 0, -2, -2, 2, 5, 0, 4, 3, 2, 2, -5, -1, -7, 0, 1, 0, 0, -8, -5, -1, -8, -4, -4, 1, -4, -2, 1, -4, -2, 0, 2, 2, 2, 4, 3, 3, 2, 0, -1, 0, -3, 1, 0, -3, -5, -6, -6, -1, -1, -8, -8, 0, -1, -3, -2, 4, 2, 2, 2, 3, -4, 1, 2, 3, -1, 0, -2, -2, 0, 1, 2, -3, 0, -1, -1, 0, -1, -3, 0, -4, -3, -7, -8, 0, 2, -2, 1, 5, 4, 3, -2, 0, -3, -1, -3, 1, 1, 2, -2, 1, 2, 6, 1, 2, -4, -1, 0, 2, 0, 0, 1, -3, -4, -3, -1, -1, -1, -4, 3, 4, 0, 2, 4, 2, 4, -3, 0, 3, 1, 2, 0, 0, -2, 0, 0, 1, 0, 1, 3, -3, -2, -2, 4, 1, -5, -7, 0, -2, -4, 2, -2, 0, -2, 4, -3, 0, 0, -3, -4, 1, 0, 0, -1, 1, 1, 5, 0, 0, 0, -1, -5, 0, 0, 3, 3, 1, 0, -3, 0, -3, 3, -2, 3, 0, 1, -3, -3, 0, -4, 0, -1, 2, 3, 4, 0, 0, 3, 0, -4, 2, -2, 1, -5, -4, 3, 3, 5, 0, 3, 1, 3, 2, -3, -4, -2, 1, -2, -4, -1, -4, -1, -1, -8, 0, 0, -2, 1, -2, -3, -1, -3, -2, -2, -3, -3, 0, 3, 3, 5, 0, -1, 4, -1, 0, 0, 3, -4, -1, 3, 0, -2, -2, 4, -3, -5, -8, 0, -4, 1, 1, 0, 0, -1, -3, -1, -3, 2, -4, 0, 0, -1, 1, 0, -1, -2, -3, -2, 0, 0, -1, 0, 5, 3, -1, 6, -6, -1, -2, -4, -5, -3, -1, 1, 1, 0, 2, 0, 3, -3, 0, 2, 8, 6, 7, 7, 0, 2, 0, 0, -3, -1, 0, 2, 4, 5, 3, 2, -4, -5, -7, -1, -4, -1, -3, -4, 0, 1, 3, 2, 0, 2, 5, 8, 9, 13, 6, 5, 10, 11, 2, 9, 1, 0, 6, 0, 2, 3, 3, 1, 0, -6, -11, -1, 2, 0, 0, -4, 1, 3, 1, 3, 3, 11, 10, 9, 9, 15, 16, 11, 10, 12, 13, 13, 6, 4, 7, 9, 4, 7, 3, 0, 2, -3, -4, -7, -3, -1, 1, -1, 0, 6, 4, 3, 3, 8, 9, 18, 18, 16, 13, 12, 8, 10, 14, 11, 5, 5, 6, 5, 6, 8, 2, -2, -1, -6, -8, -2, -3, -3, 3, -2, -1, 4, 7, 9, 5, 9, 7, 16, 10, 15, 18, 17, 13, 12, 8, 5, 8, 5, 6, 6, 1, 0, 2, -3, 0, -6, -9, 0, -1, -3, -7, 0, 0, 4, 4, 8, 9, 3, 7, 4, 14, 11, 13, 6, 4, 8, 2, 6, 1, 3, 1, 1, 0, 0, -3, 0, -1, -10, -1, -2, -8, -2, -7, -1, -5, 0, 0, 3, 2, 0, 1, 2, 6, 7, 7, 1, 5, -2, -3, 5, 3, -4, -4, -4, -3, -7, -9, 0, -7, -1, -2, -6, -3, -9, -4, -8, -4, -9, -5, -2, -7, -1, -4, -6, 2, 1, -5, -5, -4, -4, -6, 0, 0, -8, -8, -7, -4, -6, -5, -4, 0, 2, 1, -7, -1, -9, -7, -10, -8, -8, -6, -7, -11, -5, -9, -5, -7, -8, -5, -7, -7, -7, -8, -4, -2, -9, -9, -11, -13, -8, -8, -1, 4, -3, 3, 1, 0, -5, -4, -9, -10, -14, -13, -8, -9, -9, -5, -3, -9, -9, -5, -7, -8, -7, -5, -4, -9, -7, -6, -5, -6, -4, -3, 0, 5, 6, 9, 6, 4, -3, -1, -5, -12, -6, -10, -5, -3, -8, -4, -8, -8, -3, -3, -2, -1, -8, -3, -8, -6, -6, -8, -10, -6, 2, 1, 3, 3, 3, 12, 4, 0, 0, -3, -5, -11, -8, -15, -12, -10, -10, -5, -11, -8, -3, -2, -5, -6, -7, -9, -10, -4, -7, -9, -6, -9, 0, -4, 3, 9, 6, 12, 3, 2, 7, 1, -2, -12, -11, -11, -7, -5, -8, -5, -5, -10, -4, -4, -7, -4, -8, -4, -3, -5, -5, -6, -11, -10, -6, 0, 2, 3, 4, 15, 6, 5, 0, -3, -5, -2, -9, -7, -3, -8, -2, -4, -1, -4, -7, 1, 0, -6, -5, -9, -5, -7, -2, -8, -7, -4, -3, -2, 7, 5, 8, 19, 14, 4, 1, 3, 0, -4, -8, -2, -4, -5, -2, -6, 0, -2, -7, -8, -2, -7, -6, -6, -4, -3, -5, -7, -3, -1, -2, 7, 6, 12, 11, 20, 17, 11, 10, 1, 3, 2, 2, -2, -2, 0, -2, -3, 0, 2, -3, 2, -3, 0, -2, 0, -4, -1, 1, -4, -1, 2, 6, 6, 11, 13, 16, 17, 16, 14, 8, 5, 11, 2, 3, -2, 3, 0, 4, 2, 2, -1, 3, 0, 0, 3, -1, 6, 4, -1, 0, 3, 1, 3, 7, 13, 16, 9, 13, 19, 16, 18, 19, 18, 12, 14, 9, 6, 5, 10, 12, 13, 12, 8, 13, 8, 11, 14, 7, 11, 7, 16, 9, 13, 12, 14, 14, 16, 20, 14, 17, 8, 6, 8, 12, 10, 14, 9, 10, 9, 9, 9, 9, 11, 7, 6, 11, 10, 12, 16, 9, 8, 15, 7, 14, 13, 6, 12, 11, 9, 12, 14, 10, 7, 6, 12, 6, 4, 10, 13, 7, 6, 4, 3, 6, 1, 3, 2, 0, 3, 9, 3, 5, 8, 1, 11, 11, 4, 11, 7, 5, 6, 13, 9, 9, 5, 4, 8, 4, 3, 11, 3, 2, 2, 1, -3, -4, -5, -4, -3, 2, -1, 2, 2, -4, -2, 1, 5, 5, 1, 6, 12, 5, 9, 7, 5, 4, 9, 3, 10, 9, 7, 10, 4, 4, 4, -3, -1, -3, 0, -2, -1, -7, -5, -2, -3, -2, -4, -2, 2, 1, 0, 8, 4, 6, 8, 9, 7, 4, 5, 7, 8, 6, 8, 6, 4, 5, 4, -4, -3, -7, -8, -4, -3, -4, -4, -3, -5, -4, 0, -2, 0, 0, 1, 3, 7, 2, 1, 7, 7, 1, 7, 0, 2, 6, 3, 1, 2, 5, 1, -4, 0, -8, -6, -3, -6, -2, -6, -4, -5, -7, -8, -2, -3, 0, -2, 5, 3, 3, 6, 1, 2, 8, 2, 4, 3, 4, 3, 6, 2, 0, 3, 1, -7, -1, -4, -7, -8, -9, -10, -5, -10, -10, -9, -3, 0, 2, 3, 1, 1, 5, 7, 6, 1, 2, 5, 6, 3, 3, 3, 6, 6, 0, -4, -2, -2, -7, -12, -11, -5, -7, -4, -11, -5, -5, -6, -3, -2, 4, 2, 6, 5, 0, 3, -1, 1, 0, 0, -1, 4, 5, -1, 5, 2, 2, -2, -5, -3, -7, -2, -8, -9, -8, -2, -6, -7, -2, -1, 2, 2, 1, 1, 0, 5, -1, 2, 5, 1, -4, 6, 2, -1, -1, 0, 5, 2, 2, 0, -1, -1, -5, -6, -4, 0, 0, -3, -9, -8, -4, 0, -2, 0, 3, 0, 3, -1, 0, 1, 0, 0, 1, 0, 0, -3, 0, 4, 0, -2, 2, 3, -2, -6, -8, -5, -4, -2, -4, 0, -3, -4, 0, -1, -4, 3, 0, -2, 2, 3, -3, -5, -5, 0, -3, -6, -6, -2, 0, 0, -2, 1, -4, -7, -6, -2, -8, -2, -6, -2, -4, -5, -6, -7, -3, -5, -1, -7, -4, -3, 0, -4, -1, -3, -1, 0, -4, -7, -4, 0, -7, -3, -1, -3, -3, -4, -3, -6, -6, -2, 0, -3, 0, -2, -4, 0, 0, -7, -3, -2, -2, -3, 1, -3, -2, -6, -3, -6, -11, -12, -7, -7, -6, 0, -4, -3, -8, -6, -4, -6, -6, -3, -6, -4, 2, -5, -1, -7, -7, -7, -8, -7, -2, -8, -6, -1, -7, -5, -3, -10, -10, -8, -6, -10, -8, -4, -8, -8, -5, -5, -8, -4, -2, -3, -4, -3, 0, -2, 0, -1, -2, -2, -7, -7, -3, -2, -4, -8, -7, -10, -6, -10, -10, -17, -12, -5, -9, -3, -10, -10, -6, 0, -3, -2, 0, -5, -2, -3, -1, 4, 6, 0, 1, 2, 0, -4, -1, -6, -7, -7, -7, -3, -7, -10, -15, -18, -10, -7, -8, -9, -4, -9, -1, -2, -6, 1, -2, -2, 1, 1, 6, 5, 2, -1, 3, -1, 3, 0, -6, -3, 0, -2, -1, -5, -10, -14, -16, -11, -7, -5, -8, -9, -5, -4, -7, 0, -8, -5, 5, 1, 3, 8, 6, 11, 10, 4, 5, 0, 4, 0, -4, -7, -5, -4, -8, -5, -11, -12, -11, -10, -16, -8, -11, -13, -7, -8, -6, -7, -8, 0, -4, 0, 1, 7, 1, 2, 0, -2, 0, -2, -1, -8, -4, -6, -10, -8, -5, -9, -12, -9, -14, -10, -8, -16, -16, -10, -10, -5, -4, -4, -4, -7, -9, -4, -2, 4, 1, -1, -1, -5, -5, -8, -2, -7, -10, -13, -12, -9, -10, -8, -8, -13, -13, -11, -10, -12, -12, -10, -8, -9, -9, -10, -8, -3, -5, -3, -2, -1, -2, -1, -1, -4, -11, -8, -10, -6, -11, -13, -10, -10, -11, -14, -13, -10, -11, -10, -10, -9, -10, -11, -16, -15, -15, -15, -9, -9, -15, -11, -4, -12, -10, -9, -9, -13, -9, -9, -5, -13, -16, -17, -13, -14, -21, -18, -12, -11, -8, -9, -9, -13, -12, -13, -16, -13, -15, -10, -12, -11, -8, -16, -10, -11, -13, -9, -7, -9, -10, -15, -9, -8, -17, -17, -17, -17, -18, -16, -13, -5, -11, -5, -6, -11, -13, -12, -17, -9, -16, -17, -11, -12, -15, -12, -8, -12, -10, -11, -12, -5, -13, -14, -12, -11, -10, -18, -14, -12, -11, -10, -11, -7, -9, 2, -3, -3, -11, -6, -10, -12, -12, -12, -17, -13, -6, -12, -12, -8, -13, -5, -8, -7, -8, -9, -14, -12, -10, -13, -16, -13, -9, -12, -3, -2, -7, 2, -5, -1, -4, -5, -9, -14, -14, -13, -14, -12, -14, -12, -14, -10, -12, -8, -10, -5, -7, -12, -14, -12, -14, -10, -12, -11, -3, -8, -6, 2, 1, 3, 0, 2, 0, -3, -5, -8, -15, -12, -14, -15, -14, -15, -12, -7, -13, -11, -7, -13, -7, -15, -9, -12, -11, -15, -13, -13, -12, -10, 0, 0, 0, 6, 4, 2, -6, -1, -10, -11, -9, -10, -12, -6, -7, -10, -8, -7, -12, -7, -8, -8, -14, -8, -9, -10, -7, -9, -10, -10, -5, -1, 2, 3, 8, 7, 4, 4, -3, -8, -8, -4, -10, -9, -8, -12, -9, -6, -8, -6, -4, -4, -2, -8, -11, -7, -10, -9, -13, -13, -11, -7, -5, 0, 5, 7, 5, 5, 7, 6, -1, 2, -4, -2, -4, -7, -11, -7, -5, -5, -7, -7, -10, -9, -10, -7, -2, -8, -5, -3, -5, -6, -1, -3, -6, -1, 2, 9, 3, 10, 8, 3, 2, 7, 0, 2, -1, -3, -3, 0, -6, -2, -5, 0, -6, 0, -5, 0, -5, 1, -7, -2, 0, 0, -4, -3, 2, 2, 2, 10, 10, 17, 8, 13, 8, 6, 9, 4, 1, 4, 2, 6, 2, 1, 10, 4, 1, 7, 5, 2, 10, 9, 8, 1, 10, 6, 9, 5, 12, 10, 10, 12, 9, 22, 20, 16, 14, 19, 17, 16, 15, 21, 22, 21, 15, 20, 18, 14, 23, 22, 15, 16, 17, 19, 18, 25, 20, 16, 15, 16, 20, 15, 19, 22, 20, 18, 20, 20, 15, 16, 18, 19, 17, 15, 12, 14, 13, 8, 8, 11, 8, 10, 13, 14, 15, 10, 13, 15, 17, 14, 13, 19, 17, 16, 15, 18, 12, 15, 17, 18, 15, 19, 17, 14, 11, 9, 7, 0, 7, 2, 8, 3, 8, 6, 8, 9, 6, 5, 10, 12, 12, 8, 16, 12, 17, 19, 11, 15, 10, 14, 18, 18, 12, 16, 10, 15, 14, 6, 1, 1, 0, 1, 4, 0, -1, 0, 2, 4, -1, 3, 5, 6, 11, 15, 12, 10, 8, 16, 10, 15, 15, 14, 16, 9, 9, 14, 16, 8, 7, 4, 5, -2, 1, -3, 1, -1, 1, -2, 3, 0, 4, 1, 0, 7, 3, 8, 15, 8, 11, 15, 9, 15, 12, 14, 13, 11, 6, 12, 12, 7, 8, 5, 8, 0, -2, -6, -4, -5, 0, -1, -4, -6, -2, -4, 5, 2, 1, 11, 11, 7, 8, 7, 14, 12, 6, 8, 9, 6, 10, 8, 13, 12, 5, 4, 6, -2, 0, -2, -4, -8, -1, -7, -5, -5, 0, 0, -1, 6, 2, 8, 6, 4, 12, 4, 4, 10, 5, 6, 10, 6, 8, 9, 5, 6, 8, 0, 6, -2, 0, -5, -8, -3, -4, 0, -7, -3, -6, 4, -1, 6, 5, 5, 6, 10, 3, 6, 7, 5, 4, 2, 1, 5, 3, 11, 11, 5, 8, 7, 0, 1, 1, 0, 0, 2, 1, 4, -1, -2, -3, -4, 2, 2, 2, 9, 8, 9, 3, 7, 8, 6, 6, 9, 0, 7, 2, 0, 1, 3, 3, 1, 4, -1, -2, 1, 1, 0, 0, -1, -1, -5, 0, -3, 2, 5, 1, 7, 6, 4, 0, 0, 3, 0, 4, 1, 5, 6, 8, 7, 3, 4, 0, 4, -1, 0, 3, 3, 0, -1, 4, -2, 0, -5, 0, -2, 6, 0, 1, 2, 6, 3, 4, 3, 5, 4, 1, 0, 5, 0, 4, 1, 2, 5, -3, 4, 3, -5, 1, -1, -1, 0, 4, 1, 1, -1, 2, 0, -2, 0, 0, -3, 1, -2, -1, 0, 2, -3, -3, -5, -4, 4, 2, 0, 0, -1, -2, 2, -1, -3, -2, -2, 4, -3, 0, 4, 1, -1, -4, -5, 0, -4, 1, 2, 3, -2, 2, 0, -3, -2, -4, -7, -4, 1, 1, -1, -3, 2, 0, -5, -5, -4, -3, -3, -1, 4, 2, 0, 0, 1, -1, 3, -4, 2, 0, 0, 0, 0, 2, -5, -5, -7, -9, -7, -8, -5, -5, 3, -3, 2, 0, 1, 0, 0, -4, 1, -2, 1, 6, 4, 0, 1, -3, 0, 0, 0, -3, -3, 0, 0, 0, -1, -5, -2, -12, -10, -7, -9, -7, -4, -5, -3, -6, 2, 0, -2, -2, 0, 5, 4, 2, 10, 3, 7, 5, 0, 0, 0, -1, -2, 0, 2, -1, -5, -2, -9, -12, -12, -7, -4, -5, -7, 1, 0, -2, -1, -1, 5, 3, 7, 9, 8, 11, 4, 9, 4, 3, 3, 6, 7, 4, -1, -3, -2, -4, -1, -3, -6, -14, -14, -8, -3, -3, 0, 0, 1, -2, -1, 3, 1, 7, 3, 12, 8, 13, 9, 11, 3, 7, 6, 5, 7, 0, -1, -2, -3, 0, -3, -10, -8, -16, -9, -9, -11, -3, -4, 2, -5, 3, 1, -2, 3, 1, 2, 13, 5, 14, 15, 8, 2, 6, 5, 0, 5, 3, 0, 0, 0, -7, -9, -9, -13, -15, -13, -13, -6, -6, -3, 0, 0, -2, -2, 1, 3, 1, -1, 3, 4, 8, 7, 7, 6, 3, 7, 6, 4, -6, 0, -2, -7, -8, -4, -4, -8, -12, -10, -11, -7, -8, -4, -3, 0, -7, -1, -4, 2, -3, -1, 2, 3, 0, 4, 0, 0, -2, -1, -1, 0, -7, -3, -8, -5, -10, -8, -7, -8, -9, -7, -10, -7, -11, -5, -7, -9, -8, -6, -6, -3, -6, -2, -1, 4, -1, -1, -2, 2, -2, 1, -3, -2, -6, -4, -6, -10, -15, -7, -4, -7, -9, -6, -6, -11, -5, -10, -9, -5, -6, -6, -1, -5, -6, -6, 1, -3, 0, -1, -5, 0, 0, -5, 0, -5, -2, -11, -2, -6, -10, -5, -8, -7, -5, -3, -10, -11, -10, -10, -9, -8, -9, -3, -2, -6, -7, -3, -1, 2, 0, 4, 2, -2, -5, -6, -2, 0, -1, -6, -7, -8, -6, -8, -7, -5, -2, -5, 0, -6, -3, -4, -9, -8, -3, -8, -8, -7, -6, 2, -5, -4, 0, 1, 1, 2, -1, -2, -2, -2, -6, -5, -9, -7, -1, -8, -5, -5, -1, 4, 3, 0, -3, -5, -1, -6, -5, -6, -10, 0, -2, -1, -6, -5, 1, -3, -4, -4, -5, -6, -2, -7, -2, -2, -5, -8, -3, -6, -5, -3, -2, 8, 5, -2, -2, -5, -3, -10, -10, -7, -10, -5, -1, -5, 0, -2, 2, 1, 1, 2, -5, 0, -3, -5, -4, -3, -4, -7, -5, -6, -3, 5, 1, 4, 1, 3, 4, 2, 0, -6, -6, -5, 0, -3, -7, 0, -6, 0, 3, -1, 2, -5, -4, -9, -7, -3, -8, -4, -8, -10, -4, -1, 2, 1, 6, 11, 3, 1, -1, 0, 2, -2, -2, -4, -6, -3, -5, -2, -2, -1, 0, 2, 0, -5, -7, -5, -5, -4, -6, -2, -4, -1, -7, -4, 4, 3, 7, 9, 7, 2, 0, -1, -3, -2, 0, 0, 0, 1, -5, -5, 0, -1, 2, 1, -1, 1, -4, -3, -2, 0, -4, -5, 0, -2, -2, 2, 4, 10, 7, 13, 6, 11, 7, 4, 1, 2, 2, 3, 2, 3, -1, 4, -1, 2, 0, 0, 2, 0, 3, 4, -2, 0, 0, 4, 2, 5, 4, 2, 6, 3, 12, 12, 8, 12, 14, 13, 9, 12, 6, 7, 10, 9, 4, 9, 9, 11, 9, 12, 9, 11, 8, 9, 7, 5, 4, 8, 10, 11, 13, 7, 13, 9, 15,

    others => 0);
end iwght_package;
