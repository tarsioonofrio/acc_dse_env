library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 40, 0, 50, 58, 8, 0, 0, 0, 0, 0, 136, 53, 28, 31, 27, 53, 9, 33, 32, 0, 41, 105, 114, 127, 100, 14, 129, 126, 141, 135, 169, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 96, 0, 0, 27, 0, 0, 0, 0, 4, 15, 0, 0, 28, 0, 0, 160, 59, 0, 27, 0, 100, 0, 39, 14, 0, 238, 125, 0, 0, 304, 0, 0, 0, 129, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 92, 0, 43, 0, 57, 34, 0, 0, 0, 0, 0, 0, 0, 85, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 107, 5, 78, 69, 57, 82, 184, 0, 43, 0, 9, 63, 0, 22, 57, 0, 35, 0, 0, 0, 84, 8, 120, 77, 0, 0, 0, 0, 0, 0, 0, 0, 48, 0, 72, 131, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 121, 9, 0, 0, 0, 0, 0, 0, 36, 0, 0, 19, 0, 0, 9, 0, 0, 0, 0, 9, 0, 118, 0, 0, 79, 0, 96, 0, 0, 160, 9, 0, 80, 0, 155, 14, 16, 0, 6, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 21, 0, 15, 62, 27, 44, 8, 50, 57, 4, 93, 175, 61, 0, 17, 12, 138, 15, 114, 86, 0, 0, 123, 66, 96, 38, 0, 13, 0, 264, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 11, 29, 44, 18, 0, 27, 28, 38, 45, 35, 80, 0, 37, 0, 136, 62, 94, 197, 50, 27, 0, 91, 119, 14, 87, 33, 0, 114, 0, 0, 0, 58, 34, 4, 0, 201, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 213, 192, 207, 256, 186, 163, 183, 211, 283, 147, 36, 66, 0, 0, 0, 62, 0, 0, 102, 0, 15, 0, 14, 0, 0, 0, 0, 2, 0, 67, 0, 0, 56, 0, 133, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 0, 6, 0, 0, 0, 25, 0, 4, 0, 0, 0, 0, 0, 116, 12, 0, 0, 0, 54, 0, 0, 0, 0, 0, 0, 26, 126, 0, 191, 0, 0, 0, 131, 0, 0, 0, 66, 0, 7, 0, 126, 108, 0, 0, 0, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 74, 0, 0, 0, 0, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 138, 0, 0, 21, 0, 76, 63, 124, 0, 0, 77, 54, 58, 0, 0, 0, 0, 52, 1, 103, 13, 45, 0, 25, 19, 0, 0, 63, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 101, 0, 72, 0, 0, 0, 0, 0, 50, 0, 0, 0, 95, 96, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 213, 0, 0, 0, 0, 0, 0, 186, 0, 53, 0, 0, 59, 0, 118, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 76, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 0, 0, 166, 0, 129, 0, 0, 0, 191, 0, 0, 222, 0, 0, 0, 245, 0, 0, 0, 0, 0, 0, 119, 0, 0, 0, 67, 0, 35, 0, 0, 181, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 9, 21, 40, 82, 65, 38, 62, 63, 66, 14, 110, 1, 32, 31, 0, 63, 26, 100, 63, 110, 78, 177, 43, 12, 41, 0, 35, 32, 127, 37, 26, 58, 107, 71, 0, 34, 76, 37, 36, 72, 20, 112, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 77, 82, 356, 0, 0, 0, 139, 197, 53, 0, 0, 0, 0, 132, 0, 0, 128, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 0, 96, 0, 173, 23, 0, 305, 0, 0, 192, 71, 0, 0, 0, 201, 0, 69, 0, 110, 105, 107, 93, 0, 55, 15, 111, 140, 144, 117, 0, 106, 0, 0, 0, 0, 0, 0, 70, 0, 0, 0, 0, 113, 0, 0, 0, 42, 0, 0, 7, 0, 0, 0, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 40, 0, 186, 62, 154, 46, 54, 33, 34, 0, 0, 13, 91, 185, 67, 100, 48, 180, 34, 0, 16, 0, 0, 0, 107, 181, 44, 13, 0, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 87, 69, 46, 111, 66, 130, 94, 0, 109, 26, 74, 0, 26, 42, 0, 23, 0, 56, 0, 58, 50, 48, 75, 0, 0, 0, 0, 27, 0, 0, 0, 0, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 10, 25, 71, 74, 29, 10, 0, 113, 52, 31, 81, 30, 33, 35, 168, 110, 47, 43, 44, 0, 33, 90, 63, 51, 54, 101, 21, 33, 152, 9, 20, 22, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 89, 0, 0, 0, 0, 114, 0, 43, 117, 0, 0, 0, 0, 0, 0, 0, 0, 0, 114, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 55, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 2, 0, 0, 0, 0, 80, 0, 181, 60, 64, 114, 75, 52, 23, 112, 83, 98, 101, 69, 3, 0, 0, 28, 0, 0, 36, 0, 17, 0, 0, 0, 0, 35, 0, 0, 0, 0, 0, 13, 0, 0, 3, 0, 29, 0, 0, 1, 0, 0, 1, 0, 112, 10, 0, 21, 0, 0, 11, 0, 0, 0, 10, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 9, 84, 45, 22, 0, 42, 194, 0, 127, 0, 26, 0, 0, 67, 91, 167, 0, 185, 0, 0, 0, 71, 0, 0, 0, 0, 136, 0, 0, 0, 0, 66, 0, 11, 0, 0, 0, 0, 0, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 58, 0, 91, 105, 33, 0, 0, 87, 81, 74, 40, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 87, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 0, 48, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 112, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 6, 0, 0, 0, 0, 67, 97, 0, 19, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 0, 0, 49, 0, 0, 0, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 0, 0, 0, 147, 0, 28, 0, 205, 0, 0, 203, 0, 0, 0, 0, 111, 0, 109, 0, 0, 0, 0, 0, 0, 0, 0, 74, 38, 0, 0, 0, 0, 0, 0, 75, 0, 0, 0, 0, 0, 0, 105, 100, 145, 92, 40, 34, 98, 69, 86, 0, 99, 23, 0, 113, 0, 159, 0, 0, 143, 27, 24, 0, 170, 48, 0, 70, 73, 60, 0, 0, 0, 61, 35, 0, 79, 0, 0, 0, 0, 6, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 52, 66, 53, 11, 0, 0, 0, 0, 0, 85, 0, 51, 0, 0, 9, 42, 112, 0, 107, 19, 0, 24, 49, 32, 0, 89, 0, 81, 0, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 41, 0, 0, 0, 0, 47, 101, 0, 0, 0, 38, 33, 55, 29, 52, 0, 0, 14, 0, 0, 0, 0, 49, 0, 83, 0, 60, 0, 0, 34, 0, 9, 0, 63, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 0, 0, 0, 0, 0, 63, 0, 0, 41, 0, 0, 26, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 40, 321, 0, 0, 65, 66, 106, 0, 0, 0, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 166, 0, 0, 0, 16, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 0, 113, 45, 106, 0, 0, 103, 0, 143, 136, 221, 0, 0, 199, 0, 226, 30, 222, 93, 0, 132, 0, 147, 0, 87, 0, 121, 0, 108, 29, 0, 0, 0, 145, 0, 10, 0, 0, 26, 0, 0, 0, 0, 0, 0, 5, 6, 0, 0, 92, 0, 0, 0, 0, 0, 0, 43, 0, 0, 0, 88, 0, 0, 84, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 5, 68, 0, 18, 0, 46, 0, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 152, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 169, 0, 0, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 106, 149, 0, 147, 32, 48, 119, 0, 82, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 0, 0, 0, 0, 0, 0, 0, 53, 64, 4, 75, 0, 0, 51, 101, 98, 104, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 68, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 70, 0, 0, 0, 0, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 195, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 240, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 0, 0, 0, 0, 0, 0, 30, 0, 133, 0, 42, 0, 0, 172, 0, 90, 7, 82, 0, 0, 195, 0, 65, 0, 199, 0, 0, 0, 126, 0, 0, 0, 0, 150, 130, 35, 0, 14, 0, 62, 32, 30, 0, 15, 0, 44, 42, 42, 7, 31, 38, 58, 30, 129, 0, 0, 28, 0, 33, 23, 0, 34, 0, 18, 52, 40, 71, 175, 0, 0, 0, 0, 23, 0, 86, 7, 62, 0, 0, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 50, 0, 0, 0, 0, 0, 0, 120, 0, 0, 0, 0, 36, 0, 99, 0, 28, 0, 0, 0, 10, 0, 0, 99, 14, 241, 0, 30, 42, 36, 39, 83, 0, 27, 22, 0, 27, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 3, 0, 0, 70, 0, 4, 93, 0, 129, 115, 78, 186, 0, 62, 58, 107, 81, 278, 377, 99, 50, 0, 48, 113, 52, 258, 0, 0, 0, 0, 38, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 83, 60, 22, 30, 33, 0, 62, 0, 7, 0, 35, 0, 0, 0, 0, 9, 0, 0, 0, 73, 99, 15, 68, 1, 0, 0, 0, 0, 0, 56, 76, 39, 74, 0, 6, 52, 0, 0, 0, 0, 274, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 48, 0, 30, 0, 0, 0, 0, 18, 0, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 0, 56, 0, 0, 0, 0, 0, 101, 0, 12, 0, 0, 87, 57, 42, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 101, 87, 0, 0, 0, 6, 92, 72, 66, 35, 0, 0, 11, 73, 90, 45, 25, 0, 80, 15, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 105, 15, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 33, 119, 36, 29, 111, 37, 0, 111, 0, 12, 0, 0, 87, 0, 0, 0, 27, 33, 0, 95, 0, 0, 0, 0, 69, 4, 39, 0, 49, 23, 0, 0, 0, 0, 0, 37, 103, 0, 0, 0, 0, 0, 0, 0, 49, 0, 0, 0, 0, 0, 19, 60, 36, 38, 36, 63, 3, 0, 76, 108, 43, 0, 94, 0, 0, 0, 0, 56, 0, 0, 0, 0, 0, 0, 27, 0, 0, 44, 33, 0, 63, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 94, 106, 15, 20, 0, 0, 39, 18, 54, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 8, 0, 0, 0, 3, 0, 0, 0, 2, 0, 58, 91, 0, 88, 0, 43, 74, 0, 3, 9, 0, 300, 0, 26, 22, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 80, 60, 98, 2, 14, 0, 32, 199, 157, 95, 0, 53, 12, 0, 0, 0, 0, 48, 192, 25, 0, 0, 23, 0, 0, 0, 0, 0, 0, 27, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 0, 0, 236, 0, 0, 0, 0, 42, 0, 0, 355, 0, 182, 0, 73, 0, 0, 0, 86, 0, 0, 0, 0, 34, 0, 0, 0, 0, 177, 0, 0, 0, 0, 0, 52, 0, 0, 0, 0, 376, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 49, 48, 0, 0, 0, 0, 0, 105, 232, 54, 83, 82, 70, 15, 51, 118, 73, 70, 67, 113, 0, 0, 0, 0, 0, 96, 0, 4, 0, 52, 151, 0, 75, 64, 0, 0, 0, 220, 0, 35, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 102, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51, 26, 28, 17, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 155, 105, 28, 0, 0, 0, 6, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 124, 0, 0, 0, 3, 0, 0, 0, 0, 69, 0, 117, 0, 0, 0, 0, 0, 0, 121, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 99, 117, 12, 0, 49, 164, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 67, 0, 0, 0, 71, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 56, 18, 18, 19, 80, 47, 63, 33, 45, 12, 34, 0, 0, 35, 0, 0, 162, 18, 8, 5, 0, 0, 79, 18, 0, 40, 3, 26, 2, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 163, 158, 0, 40, 0, 0, 73, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 93, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 106, 0, 0, 19, 0, 0, 0, 38, 0, 0, 0, 0, 449, 0, 0, 0, 0, 16, 39, 165, 0, 0, 0, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 83, 167, 126, 0, 0, 33, 107, 116, 79, 0, 15, 0, 0, 31, 44, 28, 36, 26, 47, 59, 62, 34, 50, 34, 0, 17, 9, 2, 21, 51, 0, 0, 27, 0, 0, 0, 52, 29, 0, 10, 82, 0, 32, 7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 129, 66, 152, 0, 0, 0, 0, 0, 151, 154, 0, 0, 0, 0, 0, 5, 100, 38, 0, 0, 0, 0, 0, 0, 0, 23, 76, 79, 8, 226, 202, 73, 80, 183, 200, 154, 218, 299, 239, 184, 121, 106, 131, 150, 0, 0, 0, 0, 0, 0, 0, 106, 0, 0, 37, 110, 0, 186, 0, 284, 0, 0, 315, 127, 0, 0, 61, 0, 0, 144, 125, 0, 0, 19, 78, 0, 0, 38, 0, 0, 0, 168, 0, 90, 48, 15, 172, 0, 104, 29, 25, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 191, 33, 0, 3, 0, 0, 0, 0, 64, 30, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 115, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 164, 75, 0, 0, 13, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 74, 0, 65, 54, 0, 0, 0, 70, 53, 67, 23, 0, 48, 0, 0, 0, 26, 0, 0, 30, 0, 42, 0, 93, 0, 61, 0, 0, 181, 0, 88, 99, 160, 34, 0, 63, 57, 42, 20, 183, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 12, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 159, 0, 27, 0, 0, 14, 0, 0, 37, 61, 7, 108, 3, 0, 121, 111, 125, 79, 117, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 0, 64, 38, 161, 4, 62, 490, 236, 130, 0, 451, 0, 0, 237, 0, 0, 11, 882, 0, 0, 84, 0, 130, 46, 373, 0, 5, 240, 843, 0, 0, 0, 0, 0, 0, 458, 0, 0, 0, 0, 0, 0, 0, 127, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 102, 0, 0, 0, 0, 0, 142, 157, 0, 0, 0, 0, 0, 66, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51, 65, 0, 0, 0, 61, 131, 160, 176, 365, 0, 127, 144, 138, 156, 126, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 178, 246, 0, 103, 0, 0, 127, 0, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 64, 53, 69, 0, 39, 0, 22, 47, 0, 0, 1, 91, 12, 51, 141, 0, 0, 74, 196, 102, 13, 172, 157, 51, 64, 166, 160, 20, 13, 123, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 82, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 50, 50, 0, 55, 6, 43, 7, 34, 89, 37, 128, 32, 13, 56, 53, 50, 102, 27, 15, 74, 0, 41, 0, 0, 129, 72, 35, 17, 66, 134, 2, 103, 77, 2, 31, 11, 61, 88, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 93, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 0, 0, 0, 0, 0, 0, 0, 83, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 61, 22, 93, 9, 63, 24, 96, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 104, 0, 42, 0, 0, 0, 0, 137, 120, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 35, 92, 71, 36, 0, 22, 120, 100, 21, 67, 34, 0, 0, 17, 24, 39, 34, 47, 67, 32, 60, 0, 9, 0, 6, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 40, 92, 0, 104, 0, 0, 0, 0, 49, 0, 26, 0, 42, 44, 29, 47, 0, 0, 0, 0, 36, 54, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 78, 153, 124, 0, 213, 226, 227, 218, 214, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 82, 0, 0, 0, 0, 0, 0, 125, 0, 0, 0, 0, 91, 0, 44, 0, 0, 207, 0, 0, 0, 0, 0, 0, 181, 190, 0, 78, 0, 0, 0, 0, 235, 0, 0, 0, 0, 46, 40, 59, 0, 0, 0, 0, 26, 116, 0, 0, 0, 120, 6, 61, 299, 14, 0, 0, 310, 111, 0, 144, 107, 44, 0, 286, 73, 104, 43, 207, 0, 55, 0, 0, 106, 48, 215, 0, 0, 48, 69, 51, 21, 55, 53, 68, 78, 96, 79, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 113, 173, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 72, 0, 0, 0, 156, 123, 79, 26, 100, 104, 99, 88, 23, 27, 70, 0, 62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 16, 0, 0, 0, 0, 0, 31, 63, 0, 26, 23, 3, 46, 0, 58, 0, 0, 0, 0, 111, 0, 79, 34, 11, 0, 0, 0, 5, 71, 0, 0, 0, 91, 7, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 34, 0, 0, 21, 117, 99, 80, 5, 189, 15, 66, 151, 74, 3, 0, 50, 32, 70, 78, 90, 39, 0, 194, 82, 0, 32, 9, 0, 15, 33, 108, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 178, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 22, 105, 0, 0, 0, 0, 0, 0, 0, 180, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 198, 102, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 63, 0, 0, 0, 79, 72, 117, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 90, 0, 0, 141, 0, 112, 21, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 310, 38, 0, 223, 0, 54, 71, 0, 0, 31, 0, 0, 0, 61, 0, 146, 0, 0, 0, 313, 343, 270, 177, 55, 84, 202, 96, 0, 0, 13, 0, 24, 0, 0, 0, 0, 0, 0, 151, 69, 0, 0, 0, 0, 0, 0, 19, 53, 182, 178, 180, 164, 0, 10, 203, 109, 38, 128, 49, 248, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 0, 0, 168, 0, 0, 0, 0, 80, 97, 135, 133, 132, 0, 70, 57, 108, 99, 129, 0, 0, 0, 0, 55, 0, 3, 185, 266, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 245, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 38, 0, 0, 0, 14, 0, 30, 80, 0, 33, 0, 17, 0, 23, 14, 0, 5, 32, 0, 12, 27, 29, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 56, 85, 32, 0, 0, 0, 74, 0, 0, 0, 0, 29, 0, 20, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end ifmap_package;
