LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
	PACKAGE gold_package is
		type padroes is array(0 to 4000000) of integer;
		constant gold: padroes := ( 1, 0, 224, 162, 1, 0, 202, 
		147, 0, 0, 0, 0, 133, 109, 
		73, 137, 135, 0, 198, 71, 111, 
		15, 79, 188, 172, 50, 243, 98, 
		6, 0, 0, 175, 105, 19, 2, 
		0, 89, 96, 0, 57, 165, 104, 
		187, 66, 39, 0, 0, 191, 106, 
		
		43, 45, 0, 93, 162, 26, 113, 
		0, 0, 59, 0, 242, 207, 141, 
		94, 29, 175, 0, 0, 147, 64, 
		115, 83, 100, 11, 208, 45, 90, 
		0, 80, 119, 0, 71, 179, 0, 
		225, 4, 14, 88, 0, 83, 97, 
		0, 153, 0, 125, 142, 109, 7, 
		
		0, 0, 0, 0, 159, 119, 0, 
		0, 42, 73, 0, 74, 0, 47, 
		0, 0, 0, 0, 0, 0, 0, 
		22, 85, 0, 0, 0, 0, 0, 
		0, 117, 173, 0, 36, 102, 17, 
		14, 0, 124, 81, 89, 0, 95, 
		166, 200, 112, 3, 144, 0, 0, 
		
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		
		0, 0, 86, 92, 0, 0, 0, 
		0, 0, 39, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 171, 192, 
		0, 0, 0, 116, 82, 147, 0, 
		0, 0, 0, 9, 0, 0, 0, 
		101, 20, 0, 0, 0, 0, 0, 
		
		77, 7, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		47, 0, 39, 225, 0, 186, 0, 
		31, 0, 0, 0, 0, 46, 2, 
		126, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		
		93, 23, 44, 77, 204, 119, 63, 
		92, 53, 188, 194, 249, 97, 144, 
		53, 87, 10, 237, 116, 28, 221, 
		108, 74, 225, 66, 73, 152, 158, 
		103, 139, 36, 99, 18, 90, 41, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 34, 0, 0, 0, 0, 0, 
		
		0, 24, 0, 0, 0, 31, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		56, 0, 148, 2, 0, 0, 133, 
		146, 0, 0, 0, 0, 0, 50, 
		0, 0, 0, 176, 50, 0, 22, 
		0, 0, 0, 111, 0, 0, 55, 
		72, 15, 0, 0, 0, 0, 0, 
		
		0, 3, 86, 51, 36, 44, 0, 
		45, 117, 66, 106, 0, 0, 0, 
		6, 0, 0, 113, 0, 57, 41, 
		12, 139, 0, 0, 0, 0, 0, 
		0, 0, 0, 15, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		
		15, 88, 59, 64, 54, 125, 136, 
		70, 103, 68, 65, 167, 242, 247, 
		82, 115, 251, 26, 86, 119, 120, 
		0, 42, 107, 143, 68, 76, 185, 
		0, 0, 17, 82, 117, 127, 189, 
		34, 8, 148, 0, 0, 24, 0, 
		42, 220, 147, 62, 14, 38, 0, 
		
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 32, 0, 29, 0, 
		0, 0, 0, 97, 0, 25, 0, 
		35, 0, 0, 0, 0, 127, 0, 
		162, 0, 0, 0, 0, 112, 0, 
		148, 3, 172, 93, 235, 102, 132, 
		54, 229, 169, 100, 17, 222, 202, 
		
		0, 33, 0, 0, 0, 76, 0, 
		149, 82, 0, 0, 81, 15, 164, 
		109, 243, 0, 0, 161, 46, 0, 
		0, 140, 0, 51, 92, 47, 0, 
		22, 57, 105, 0, 0, 0, 0, 
		0, 9, 214, 0, 161, 0, 0, 
		61, 0, 126, 0, 53, 68, 229, 
		
		0, 0, 0, 0, 0, 230, 0, 
		0, 0, 150, 0, 0, 0, 223, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 50, 0, 
		0, 0, 58, 104, 135, 0, 0, 
		0, 48, 0, 0, 55, 0, 0, 
		43, 0, 0, 0, 0, 69, 78, 
		
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		
		0, 0, 0, 0, 53, 0, 0, 
		0, 65, 0, 131, 0, 0, 0, 
		0, 0, 0, 0, 201, 0, 0, 
		0, 0, 0, 0, 0, 5, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 120, 0, 0, 
		0, 0, 0, 0, 0, 26, 50, 
		
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 46, 0, 0, 53, 0, 
		88, 0, 202, 0, 136, 175, 59, 
		206, 27, 22, 219, 48, 232, 207, 
		
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 78, 0, 0, 
		0, 0, 0, 16, 74, 0, 0, 
		0, 0, 124, 0, 70, 0, 0, 
		9, 156, 0, 0, 0, 0, 85, 
		179, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 51, 0, 0, 0, 
		
		38, 121, 60, 0, 0, 0, 105, 
		0, 32, 0, 0, 0, 7, 0, 
		0, 1, 0, 0, 135, 0, 0, 
		69, 0, 0, 0, 38, 0, 122, 
		21, 50, 9, 0, 0, 0, 0, 
		207, 41, 1, 188, 172, 179, 233, 
		204, 32, 139, 165, 76, 181, 224, 
		
		0, 0, 0, 12, 102, 197, 86, 
		194, 77, 202, 0, 115, 65, 26, 
		160, 0, 9, 55, 152, 0, 73, 
		0, 25, 0, 98, 0, 0, 30, 
		0, 121, 29, 0, 0, 131, 0, 
		54, 1, 0, 86, 69, 144, 165, 
		50, 0, 88, 0, 122, 124, 207, 
		
		73, 243, 106, 73, 203, 0, 93, 
		78, 87, 19, 44, 0, 0, 0, 
		0, 81, 0, 194, 0, 0, 0, 
		0, 35, 0, 0, 0, 0, 0, 
		61, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		
		176, 115, 45, 0, 90, 171, 163, 
		0, 88, 106, 103, 179, 101, 52, 
		0, 71, 223, 31, 29, 132, 0, 
		76, 26, 127, 192, 71, 181, 86, 
		0, 29, 134, 0, 145, 246, 26, 
		30, 0, 123, 110, 0, 0, 11, 
		22, 130, 61, 118, 113, 74, 0, 
		
		0, 0, 0, 0, 29, 0, 4, 
		116, 0, 0, 0, 65, 0, 0, 
		46, 0, 0, 0, 126, 0, 0, 
		0, 0, 70, 0, 126, 0, 0, 
		0, 109, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		
		46, 88, 13, 50, 122, 95, 27, 
		153, 137, 89, 20, 11, 122, 88, 
		0, 133, 0, 48, 0, 0, 24, 
		0, 54, 161, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		
		33, 12, 0, 34, 0, 96, 110, 
		0, 0, 29, 0, 0, 0, 97, 
		122, 0, 0, 0, 32, 24, 0, 
		0, 0, 114, 0, 0, 101, 157, 
		66, 93, 0, 98, 136, 145, 153, 
		132, 159, 222, 172, 236, 88, 83, 
		48, 26, 103, 243, 58, 197, 62, 
		
		0, 13, 0, 0, 40, 18, 54, 
		177, 174, 81, 34, 200, 50, 49, 
		0, 0, 0, 0, 102, 62, 0, 
		0, 14, 54, 0, 62, 0, 0, 
		0, 89, 182, 74, 0, 172, 77, 
		30, 84, 0, 26, 122, 96, 214, 
		0, 0, 52, 49, 0, 0, 26, 
		
		0, 2, 164, 143, 0, 0, 162, 
		64, 58, 0, 0, 0, 39, 15, 
		0, 106, 31, 0, 212, 0, 166, 
		0, 0, 0, 80, 99, 91, 0, 
		70, 0, 65, 35, 62, 147, 0, 
		48, 0, 0, 74, 170, 17, 197, 
		127, 69, 188, 98, 209, 222, 208, 
		
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 6, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		
		0, 0, 0, 101, 83, 25, 110, 
		0, 8, 0, 103, 0, 0, 0, 
		0, 0, 0, 0, 110, 0, 0, 
		0, 0, 215, 0, 62, 0, 0, 
		0, 0, 0, 0, 0, 20, 52, 
		33, 36, 0, 0, 33, 128, 53, 
		167, 0, 0, 19, 53, 4, 0, 
		
		150, 111, 8, 0, 0, 0, 42, 
		93, 0, 0, 118, 108, 161, 0, 
		0, 145, 93, 88, 0, 108, 111, 
		42, 0, 37, 0, 44, 53, 212, 
		220, 0, 0, 98, 0, 106, 76, 
		148, 81, 145, 101, 71, 145, 93, 
		82, 253, 107, 24, 127, 180, 81, 
		
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		131, 0, 0, 116, 0, 59, 0, 
		151, 0, 0, 0, 0, 0, 0, 
		31, 0, 0, 0, 0, 0, 0, 
		0, 0, 0, 0, 0, 0, 0, 
		0, 0, 26, 0, 0, 0, 0, 
		
		91, 184, 74, 100, 85, 85, 34, 
		101, 167, 0, 201, 151, 152, 0, 
		95, 49, 150, 254, 119, 20, 197, 
		158, 161, 50, 200, 152, 131, 111, 
		151, 141, 101, 116, 0, 0, 25, 
		47, 55, 51, 28, 78, 70, 15, 
		0, 0, 0, 59, 0, 148, 0, 
		
		others=>0 );
END gold_package;
