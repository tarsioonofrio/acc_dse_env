library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    127, 0, 106, 0, 0, 0, 0, 0, 0, 0, 482, 0, 187, 112, 0, 160, 0, 234, 0, 0, 102, 102, 66, 0, 34, 0, 0, 392, 477, 474, 482, 207, 252, 133, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 194, 49, 85, 0, 73, 61, 65, 412, 413, 237, 0, 0, 37, 0, 0, 27, 329, 16, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 85, 0, 0, 0, 0, 108, 0, 34, 15, 0, 0, 0, 0, 0, 49, 173, 256, 138, 259, 245, 62, 0, 360, 331, 0, 0, 0, 0, 0, 0, 0, 0, 0, 280, 0, 59, 0, 0, 54, 0, 0, 0, 222, 448, 433, 405, 101, 76, 195, 212, 46, 0, 0, 71, 0, 140, 250, 0, 0, 0, 0, 0, 0, 65, 0, 3, 245, 0, 80, 43, 105, 155, 0, 164, 247, 0, 264, 181, 0, 0, 0, 0, 66, 0, 0, 64, 174, 0, 0, 136, 7, 135, 25, 0, 43, 0, 0, 0, 21, 0, 5, 0, 0, 0, 0, 0, 199, 57, 256, 447, 278, 319, 260, 159, 0, 0, 13, 42, 0, 182, 226, 140, 393, 155, 3, 80, 150, 74, 0, 197, 83, 0, 96, 169, 258, 301, 164, 130, 358, 0, 106, 0, 17, 0, 0, 140, 0, 34, 103, 101, 53, 172, 78, 369, 316, 241, 387, 396, 280, 117, 0, 0, 0, 0, 0, 0, 147, 353, 0, 0, 0, 0, 200, 104, 129, 32, 124, 0, 0, 0, 0, 0, 10, 0, 35, 0, 278, 124, 281, 413, 239, 311, 457, 434, 436, 136, 247, 0, 2, 318, 0, 0, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 227, 227, 21, 118, 81, 262, 135, 208, 8, 0, 194, 84, 0, 310, 98, 0, 0, 0, 0, 0, 0, 0, 48, 0, 0, 0, 0, 162, 251, 83, 237, 69, 0, 238, 301, 254, 47, 175, 51, 138, 234, 52, 107, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 222, 291, 0, 0, 0, 0, 0, 0, 57, 8, 0, 76, 0, 0, 0, 91, 204, 0, 0, 0, 0, 0, 0, 0, 43, 151, 0, 130, 71, 439, 150, 288, 360, 217, 173, 0, 0, 59, 135, 323, 215, 317, 0, 0, 98, 274, 293, 278, 291, 403, 255, 216, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 197, 0, 148, 76, 0, 229, 0, 67, 41, 14, 0, 0, 0, 0, 0, 0, 112, 101, 0, 0, 0, 0, 0, 0, 0, 27, 148, 287, 308, 118, 0, 30, 45, 0, 0, 0, 0, 0, 0, 0, 0, 72, 175, 293, 191, 0, 0, 0, 0, 18, 0, 0, 0, 0, 139, 119, 39, 105, 176, 81, 15, 42, 34, 110, 251, 439, 156, 179, 88, 117, 50, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 158, 0, 44, 53, 0, 157, 125, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 0, 0, 0, 0, 245, 208, 0, 0, 0, 0, 0, 0, 167, 442, 354, 154, 232, 88, 13, 267, 206, 91, 0, 53, 0, 0, 43, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 187, 154, 232, 161, 321, 0, 126, 33, 370, 277, 408, 
    
    
    others => 0);
end ifmap_package;
