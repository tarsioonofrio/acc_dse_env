library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 4000000) of integer;

  constant input_wght : mem := (
    -- bias
    27969, 2595, -1981, -4314, -5392, -892, -20327, -10102, 19330, -2965,

    -- weights
    -- filter=0 channel=0
    25, 16, 10, 13, 14, 6, 0, 6, 6, 8, 7, 5, 6, 0, -4, -2, 0, 10, -5, 3, -5, -1, 9, 0, 7, 2, 15, 7, 16, 22, 22, 0, 5, -5, -7, 7, 1, 1, 4, -5, -2, 0, -3, -7, -8, 0, -3, 2, -1, -9, -3, -10, -10, -7, 4, 3, -4, -3, 14, 20, 7, 8, 2, 2, -6, -7, -9, -10, 4, 2, -1, 0, 6, 5, -9, 2, 3, -13, -6, -1, -8, -3, -10, 0, -11, -10, -10, -7, -3, 6, 12, -1, -4, -4, 1, -13, -12, -9, 0, 0, -6, 5, -1, -4, 2, 2, -8, -5, -9, -10, -4, -16, -4, -10, 0, -13, -8, -7, -6, 13, 11, -3, 1, -7, -7, -2, -12, -8, -2, 3, 0, 1, 7, -1, -4, 5, -3, -8, 1, 0, -11, -8, -16, -11, -13, -11, -2, 1, 0, 1, 9, 0, -13, -1, -15, -10, -3, -2, -11, 2, -1, 3, 5, -2, -2, 5, 9, 4, 4, -10, -11, -11, -9, -4, -13, -15, -4, 1, 0, 3, 8, -2, -10, -10, -8, 0, -3, -15, -7, -11, -3, 1, 4, 11, 12, 9, 5, -6, 0, -3, -1, -12, -9, -9, -3, -8, -15, -3, -3, -1, 12, -3, -12, -11, -8, -10, -6, 0, -12, -10, 3, 2, 2, 7, 9, 13, 1, 5, 5, 5, -10, 0, -2, -7, -12, -4, -2, -8, -1, 2, 8, -11, -11, 0, -10, -1, -12, -10, -15, 0, -1, 8, 4, 6, 13, 14, 12, 4, 4, 7, -5, -10, -4, -7, -12, -13, -17, -8, -4, 0, 6, -7, -7, -2, -6, -9, -3, -1, 0, -5, -1, 6, 7, 0, 15, 16, 6, 2, 0, 3, -3, -2, -11, -4, -18, -15, -9, -17, -6, 5, 4, -2, -14, 0, -6, -11, -12, -12, -3, 1, -5, -3, 6, 4, 11, 12, 15, 14, 3, 5, 4, 0, -10, -13, -4, -14, -3, -12, -14, 5, 4, -8, -2, -4, -1, -11, -6, -15, 0, -6, -7, 0, -1, 18, 10, 10, 20, 12, 14, 6, 7, -3, -8, -6, -17, -12, -8, -14, -11, 4, 2, 2, 0, -8, -6, -8, -15, -14, -5, -9, -2, -5, 0, 7, 18, 29, 24, 22, 25, 4, 8, 5, -10, -13, -6, -12, -15, -16, -3, 0, 8, -11, -4, -6, -1, -6, 0, -8, -13, -14, 1, 6, 13, 18, 24, 25, 32, 33, 16, 6, 13, 5, -4, -7, -9, -14, -18, -3, -9, 6, -4, 3, -14, -3, -16, -5, -7, -7, -4, -9, -7, -1, 8, 7, 30, 36, 25, 27, 19, 10, 6, 0, 1, -11, -16, -11, -6, -12, -6, 0, 5, -3, -8, -2, -12, -3, -8, -16, -12, -4, -5, 8, 5, 17, 26, 22, 34, 19, 30, 20, 15, 0, -9, -11, -4, -4, -11, -10, -8, 3, -4, -11, -7, -5, -2, -8, -7, -1, -9, -14, 3, -1, 8, 15, 12, 26, 33, 25, 15, 16, 0, -4, -10, -7, -8, -7, -16, -7, -3, 0, 3, -11, -4, -14, -9, -2, -13, -13, -5, 0, -12, 3, 13, 4, 18, 13, 21, 20, 21, 17, -1, 3, -7, -8, -7, -9, -5, -7, -9, -1, 2, -1, -11, -6, -3, -1, -8, -16, -12, -7, -9, 1, 10, 2, 8, 22, 22, 23, 12, 1, 1, -3, -12, -4, -11, -7, -5, -5, -4, 0, 9, -8, -11, -15, -14, -12, -2, -2, -17, -3, -5, 7, 5, 2, 11, 20, 7, 20, 13, 12, -4, 0, -5, -7, -17, -14, -6, -12, -11, 3, 0, -4, -3, -4, -10, -13, 0, -10, -6, -11, 3, -2, 2, 11, 8, 18, 7, 10, 7, 2, -3, -9, -14, -14, -7, -4, -11, -13, 0, 5, 6, -11, -14, -9, -12, -12, -9, -11, -10, -8, -9, -7, -2, 13, 15, 13, 6, 12, -1, 6, 5, -5, -13, -5, -6, -10, -3, -14, 2, 6, 11, 1, -9, 0, -6, -8, -5, -1, -5, -6, -3, 4, -3, 5, 7, 10, 3, 0, 5, -6, -10, -15, -15, -11, -13, -8, -5, -3, -5, 2, -1, 1, -7, -9, -13, -3, -5, -7, -6, -9, -8, 2, 1, 9, -2, 1, 0, 4, 0, 2, -11, -10, -15, -6, -4, -17, -4, -6, -7, 3, -1, 1, -6, -9, -14, -3, 0, 0, 3, 4, -5, -7, 2, 10, 7, -3, -4, -6, 3, -12, -10, -13, -6, -5, -4, -6, -1, -6, -1, 3, 2, -6, -5, -8, -13, -9, -11, -7, -12, 2, 0, 1, -6, -2, 7, 10, 0, 1, 1, -5, -15, -13, -8, -2, -2, -8, -15, -13, -2, 10, 15, -5, 3, -7, -10, -6, -12, -6, -11, -5, 5, 1, 6, -2, -2, -8, -1, 2, -5, -10, -17, -2, -4, -14, -15, -7, -4, 1, -7, 13, 15, 4, 5, -1, -7, -1, -6, 2, -8, -5, 4, 1, -7, -3, -3, 3, 2, 2, 0, -5, -9, -3, -13, -12, -4, -2, -8, 4, 10, 17, 12, 8, 0, 1, 5, -5, -8, -5, -8, 4, -11, 4, -6, -5, 2, -6, -3, 0, -12, -11, 0, -11, -7, -8, -9, -6, -5, 13, 16, 14, 23, 22, 19, 7, 4, 0, 10, 4, 5, 7, 2, 0, 0, 0, 0, 9, -5, -1, -4, 8, 4, 12, 1, 2, 7, 3, 10, 22, 16, 21,
    -- filter=0 channel=1
    9, 7, 11, 0, 5, 10, 8, 11, 0, 0, 0, 1, -8, -9, -11, -11, -1, -5, 1, -6, 1, 0, -7, 0, -7, -4, -10, 0, -5, -6, -1, -2, 13, 7, 14, 1, 10, 7, 0, -6, 2, -7, -7, -12, -10, -8, -11, -11, -12, -10, -1, -5, 0, -8, -1, -8, -11, -5, -13, 0, 2, 8, 0, 7, 14, 14, 10, 12, -3, 1, 1, -2, -1, -2, -5, -3, -1, -4, 0, 1, -3, 5, -3, 1, 2, -8, -11, 0, -15, 0, 7, 5, -1, 11, 12, 14, 8, 3, 2, 1, -10, -2, -5, -7, -19, -9, -8, 1, -7, 7, 0, -1, -5, 4, 2, 7, -5, 3, -8, 0, -1, 3, 10, 4, 7, 3, 15, 7, 12, -7, -3, -13, -4, -6, -13, -9, -10, -2, 6, 6, 9, 4, -1, 9, 13, 11, 0, 4, -10, -13, 0, -4, 12, 14, 16, 2, 13, 16, 10, 7, -5, -17, -15, -17, -17, -13, -14, 1, 0, 5, 0, 4, 15, 11, 10, 3, 4, 6, 0, -5, 6, 8, 0, 9, 6, 5, 3, 10, 5, -4, -11, -8, -12, -9, -18, -5, -16, 0, 0, 2, 13, 14, 9, 3, 5, 8, 12, 8, -7, 0, -7, 3, 7, 14, 6, 18, 8, 14, 1, 0, -3, -14, -19, -21, -20, -5, -16, 4, -5, 3, 11, 17, 16, 17, 17, 15, 13, -1, -8, 0, -1, 10, 1, 15, 5, 8, 17, 3, 10, 6, -1, -6, -7, -19, -20, -7, -15, -5, 0, 0, 2, 2, 4, 10, 16, 15, 5, 3, -4, -3, 4, 10, 4, 0, 3, 11, 3, 7, 11, 0, -12, -4, -20, -17, -19, -19, -11, -11, 5, 11, 11, 12, 8, 7, 12, 15, 4, 9, -5, 1, 0, -2, 0, 11, 12, 6, 13, 3, 0, -7, -5, -14, -17, -14, -25, -16, -5, -2, 7, 10, 10, 14, 17, 21, 11, 9, 9, 13, -5, 0, 0, 0, 10, 10, 1, 9, 2, 6, -2, -6, -14, -11, -16, -15, -24, -27, -8, -12, 0, -1, 8, 9, 16, 6, 10, 24, 8, 3, 5, 0, 4, 2, 4, 11, 11, 8, 2, 12, 0, 3, -3, -14, -13, -20, -27, -19, -6, -4, 0, 0, 10, 2, 12, 17, 9, 12, 13, 13, 9, 0, 7, 6, -1, 10, 14, 15, 5, 13, 2, -4, -1, -20, -15, -25, -19, -24, -17, -8, 0, -1, 1, 5, 2, 5, 10, 10, 18, 7, 4, -3, 1, 12, 6, 14, 10, 7, 1, 0, 7, 0, -13, -16, -20, -25, -32, -22, -18, -2, 0, 5, 14, 7, 8, 17, 11, 22, 17, 11, -2, -1, -2, 0, 8, 6, 11, 14, 9, 6, -4, 1, -1, -18, -13, -19, -32, -17, -16, 0, 4, 6, 6, 9, 11, 17, 20, 13, 13, 15, 2, 5, 4, -3, 7, 7, 7, 12, 8, 12, -2, 4, -3, -10, -20, -30, -24, -27, -11, -14, 5, 0, 11, 2, 13, 12, 17, 14, 16, 7, 13, 8, 6, -3, 11, 4, 10, 14, 9, 14, 8, -6, -6, -18, -13, -22, -25, -19, -16, -14, 2, 8, 8, 6, 16, 20, 7, 13, 5, 4, 13, 7, 9, 3, 13, 14, 11, 16, 5, 15, 1, 1, -5, -8, -12, -15, -26, -25, -17, -9, -6, 6, 1, 7, 6, 22, 21, 10, 17, 14, -3, 5, 5, -3, 1, 5, 10, 4, 6, 4, 7, 0, -13, -9, -19, -29, -14, -12, -8, 0, -8, 8, 0, 12, 10, 6, 10, 13, 19, 9, 5, 0, 2, 1, 0, 13, 6, 10, 8, 11, 6, 9, -10, -14, -23, -12, -25, -9, -4, -2, 0, 5, 10, 5, 4, 6, 11, 16, 17, 3, -5, 2, 2, 8, 7, 9, 2, 7, 12, 7, 0, -1, -6, -10, -12, -18, -13, -19, -8, -2, 4, 0, 2, 11, 7, 21, 10, 11, 7, -4, 8, -1, -6, 6, 6, -1, 12, 3, 5, 14, 1, -4, -6, -3, -7, -21, -9, -12, -12, -8, 2, 1, 11, 14, 14, 14, 5, 7, 8, 7, -9, -7, 0, 1, 0, 10, 13, 4, 5, 10, 0, -6, 4, -16, -17, -17, -18, -14, -15, -2, 3, 4, 13, 15, 8, 7, 3, 1, 9, -5, -1, 0, 5, 2, 8, 1, 12, 15, 4, 5, 10, 8, -2, -14, -17, -12, -20, -20, -1, 1, -1, 10, 4, 2, 2, 11, 1, 6, 7, -3, -10, 0, -2, 5, 5, 0, 14, 4, 2, 14, -2, -2, 2, -3, -3, -8, -14, -5, -13, 3, -4, -5, 9, 8, 2, 12, 9, 9, 9, -6, -5, -9, 2, 8, 5, 10, 7, 6, 7, 13, -5, -7, -10, -10, -6, -9, -4, -18, -8, 1, -1, -7, 1, 6, -4, 1, 0, 1, 0, -9, 0, -5, 4, 11, 1, 0, 1, 0, 5, 12, 5, -6, 0, -3, -7, -11, -9, -11, -6, -7, 2, 3, -4, -1, 5, -6, 0, 1, -5, -13, -4, -5, 3, 5, -3, -4, 13, -2, 12, -2, 7, -3, 2, 3, 2, -2, -15, -14, -9, -1, -9, 1, -10, -7, 0, 0, -8, -9, -12, -13, 1, -14, 4, 6, 8, -5, 7, 0, -5, 6, 1, 7, -5, 4, 3, -12, -6, -7, -7, -12, -12, 1, -11, -7, -7, -8, -9, -12, -8, -8, -11, -6,
    -- filter=0 channel=2
    -6, 0, 0, 7, 0, 5, 4, 3, 4, -8, 6, -5, 5, -3, -7, -10, -2, -6, 0, 1, 0, -1, -8, 3, -2, -9, 1, -2, 5, 4, 0, -2, -2, -1, 2, 0, -6, -4, -3, -9, 6, 1, -9, -1, -4, 1, -8, -1, 2, -4, -5, 3, 0, 1, -1, 0, 5, -3, -1, 3, -2, 3, -4, 0, 4, 5, 8, -3, -3, 6, -6, 5, -5, -9, -9, 0, -6, -11, -12, 0, -3, 2, 4, -2, 4, -2, -8, -2, 8, -5, 3, 9, 6, 8, 4, -5, 9, 1, 1, -2, 3, 1, 1, -8, -3, -11, 0, 0, 2, 1, -7, -5, -8, 0, 4, 0, 7, -3, 0, -6, -2, 7, 10, 8, 6, -5, 7, -5, -2, 2, -2, 2, -8, -10, -5, -7, -2, -8, -5, -6, -5, 3, -9, 3, 3, -2, 0, 6, 8, -5, -3, 11, 6, 5, 11, 5, 8, -6, 3, -8, -4, 0, -2, -7, 2, -10, -1, -4, 1, -13, 2, 2, -10, -7, -4, -5, 3, 1, 3, 0, 3, 2, 1, -2, 10, 11, 7, 7, 8, 2, -6, -6, -1, -5, 0, -12, -7, -2, -1, -9, 1, -11, 0, -3, 3, 4, 0, 4, 1, 4, 2, 12, 3, 4, 0, -3, 6, 2, 5, 5, -1, 4, 2, -12, -1, -6, 3, 1, -11, 3, 0, 3, 1, 5, 0, 3, -7, 6, 0, 0, -4, -3, -1, 0, -1, 7, -2, 1, 6, 1, 3, 6, -3, 4, 0, -6, -1, 0, 7, 4, -7, 5, -9, -9, -8, -3, 2, 3, 3, 0, 4, -2, 2, 13, -2, -3, 8, 7, -5, 0, -1, 2, -2, 5, 1, -4, -4, -4, 4, -7, -7, -2, -3, -7, -1, -6, -4, 9, 3, -6, -2, 3, 8, 10, 4, -1, 2, 1, 0, -1, 6, 4, -1, 9, 3, 10, 9, 0, 5, 0, 0, -3, -3, -2, 5, -2, 6, 3, 2, -2, -5, -3, 7, 9, 3, 8, -3, 7, -2, 8, -1, 7, 2, 5, 10, 13, 0, 0, -1, 0, -4, 3, 8, 6, -4, 1, 10, 11, 0, 9, 9, -2, 3, 4, 10, 11, 7, -1, 3, 4, 0, 8, 12, 10, 2, 16, 14, 4, 11, 7, 10, 11, -1, 2, -5, -1, -3, 11, 0, 8, 0, 6, 3, 2, 10, -4, 5, 2, 1, 6, 13, 12, 11, 18, 19, 10, 12, 16, 9, 14, 6, 8, 2, 8, -5, 10, 0, 4, -3, 2, 1, 7, 4, 11, 2, -4, 12, 4, 11, 4, 3, 13, 20, 19, 17, 15, 3, 10, 16, 1, 9, 9, 3, -3, 5, 0, 0, 8, 3, 4, -1, 5, 1, 3, 5, 5, 11, -3, 12, 6, 7, 18, 5, 17, 8, 4, 11, 7, 16, 2, 11, 2, 10, 0, -3, -2, -1, 0, 10, 6, 1, 9, 4, 1, -4, 4, 4, 4, 2, 0, 13, 11, 18, 4, 16, 1, 5, 0, 1, 2, 14, 3, 5, -4, 1, 9, 11, 12, -1, 6, -3, 2, 11, 5, 6, 3, -1, 7, 1, 13, -1, 7, 10, 8, 8, 3, 13, 10, 7, 10, 0, 0, -1, -3, 0, 3, 5, 6, 11, 8, -6, 9, -2, 10, -2, -4, -4, 0, 9, 0, -2, 2, 7, -2, 5, 3, 6, 1, 3, 10, 7, -1, -5, 0, 0, 7, 6, -3, 9, -2, 1, 9, 7, -4, 1, -3, 2, 2, 5, 6, 0, 10, 7, 3, 5, 9, 3, -2, -7, -2, -4, 4, 0, 1, -1, -1, 3, 5, 6, 6, 8, -2, 6, -3, -5, 0, 5, 0, -6, -7, 4, -3, -1, -8, 6, -6, -7, -6, 1, -4, -4, -7, -4, 0, 2, 4, -5, -4, -4, 4, 0, 11, 2, 0, -1, 5, -2, -5, 6, 1, -6, 0, 0, 1, 2, 4, -3, 2, 3, 4, 0, -4, -1, 4, -4, 7, 5, 9, 3, -3, 6, -2, 3, 7, 8, 6, 0, -1, -9, -6, 0, -3, 0, -5, -7, -8, -1, -4, -10, -9, 0, -5, -5, -6, 1, -7, 5, 8, -4, 5, 0, 6, 4, 7, 8, -2, 0, 0, 7, 0, -4, -4, -6, -7, -3, -5, -8, -14, -5, 1, -6, -12, -4, -4, -1, -6, 2, 3, -5, 5, 6, 4, 10, 0, 2, 1, -3, 7, -6, -1, -8, -2, 0, 1, 0, 0, -5, -7, -8, 0, 2, -6, -5, 0, 3, -2, -6, -3, -4, -1, 1, 5, -2, 9, 0, 10, 0, -4, -4, 5, 2, -2, -10, 0, -11, 0, -8, -13, 1, -11, -6, -11, -1, -2, -9, 5, 8, 3, -4, 6, 1, 6, 2, -5, 5, 3, 3, 2, 7, -9, -6, -6, -10, -1, -5, -4, -6, -9, -1, -10, 0, 0, -8, 5, -8, -7, -3, 0, 5, -7, 7, 7, 2, 0, -3, 0, 1, 3, -8, -7, 5, 6, -2, -2, 4, 4, 0, 4, -5, -5, 1, -8, -3, 0, -6, 7, -5, -3, -6, -8, 0, 7, 0, 0, 7, 6, -5, 8, 1, 2, 3, 5, 2, 0, -6, -1, -4, 1, 2, -7, 0, 3, -4, 0, -7, -3, 2, 5, 8, 0, 7, 2, -1, 0, -3, 0, -8, -6, -2, -1, 5, -8, -2, 5, -6, -5, -10, -1, -3, -11, 0, -2, -2, 1, -6, -7, -3, 8, 5, 8,
    -- filter=0 channel=3
    -1, 8, 7, 1, 1, 10, 7, 2, -2, -1, -1, 6, -4, 9, -6, -5, -5, -7, -4, -2, -5, 5, 5, 7, -2, -7, 3, 0, -4, -8, 0, 2, 5, -2, 6, 7, 4, 0, -2, 7, -4, 3, -1, 9, -2, -2, 9, -2, 0, 0, -2, 1, 8, -5, 2, 2, -5, -4, 0, -6, 0, 0, 6, 6, 11, -2, 5, -1, 8, 8, -3, -4, 2, 8, 5, -2, -5, 2, 6, -6, 0, 5, -2, -2, 4, -1, -4, 6, 6, -1, 10, 10, -2, 0, 6, 8, 5, -5, -3, 0, 1, 5, 3, 6, 10, -5, -3, -4, 7, 0, 0, 5, 2, -10, -9, -6, 6, -5, -1, 3, 3, 1, 11, 7, -3, 0, 0, -1, 5, 1, -5, -2, 2, 8, 9, 2, -6, 5, 4, 0, 0, -6, -1, -10, -1, 4, -7, 4, 0, -5, -3, -1, 1, 9, 1, -4, -4, 9, -6, 0, 0, 1, -1, 5, 2, 0, 2, 2, 2, -8, 0, 2, 2, -2, -9, -5, 4, -8, 0, 1, 8, 0, 9, 10, 8, 4, 10, 4, -1, 0, 3, -2, 8, -1, 4, 7, 2, -2, -4, -2, -6, -5, -9, 3, -5, -10, -2, -8, -5, -11, -1, 5, 7, 11, 13, -3, 4, 6, 8, -3, -3, 9, 10, -1, -3, 6, 0, -7, -9, -10, -2, -3, -3, 0, -3, -8, -11, -5, -5, -6, 0, 13, 7, 7, 4, 12, -1, 14, 13, 0, -2, 1, 0, 9, -3, -1, 6, 4, 5, -2, 0, -1, -9, -7, -10, 0, -9, -2, 0, -7, 3, 5, 12, 2, 6, 8, 8, 10, 14, 7, 0, 5, 6, 11, 7, -5, -5, -6, -3, -7, -9, 2, -8, -13, 0, -6, -12, -7, -2, -5, 11, 8, 18, 15, 8, 3, 10, 13, 11, 8, 1, 5, 4, 9, -1, -6, -3, 5, 3, -2, -7, 0, 0, -12, -9, -9, -10, -6, -1, -13, 13, 13, 11, 7, 13, 12, 7, 13, 18, 4, 5, 11, -1, 5, 0, -8, -8, -10, 0, -1, 2, -3, 0, -6, -9, -6, -10, -11, -15, -7, 11, 3, 12, 14, 11, 5, 4, 11, 15, 9, 3, 12, 2, -3, 0, -2, 3, -6, -9, -4, -9, -13, -4, -8, -3, -8, -8, -11, -12, -8, 8, 7, 15, 15, 18, 7, 11, 8, 7, 14, 1, -1, -3, 6, 0, -4, 0, -11, 2, 0, -9, -10, -2, -2, -11, -15, -18, -12, -12, -7, 10, 18, 20, 17, 10, 18, 6, 18, 12, 11, 3, 10, 9, 3, -6, -1, -7, -1, -10, -5, -2, -7, -13, -2, -13, -9, -8, -14, -9, -11, 16, 4, 21, 13, 14, 18, 17, 7, 2, 6, 10, 0, -2, 8, 5, -8, -11, -9, -4, 3, -5, -14, -15, -2, -6, -12, -10, -14, -5, -13, 7, 17, 12, 11, 18, 7, 9, 10, 6, 7, 8, 0, -1, -7, -4, 3, 2, 2, -10, -7, -5, -1, -11, -17, -16, -9, -11, -8, -17, -8, 13, 6, 5, 15, 5, 14, 20, 6, 15, 11, 8, 8, 9, 4, -4, -4, -9, 1, 0, -12, 0, -12, -3, -8, -2, -10, -5, -4, -10, 0, 2, 12, 7, 3, 3, 14, 3, 2, 3, 11, 14, -2, 4, 5, 1, 0, 5, 1, -5, 1, -8, -5, -14, -4, -15, -10, -13, -5, -4, -5, 6, 4, 3, 5, 5, 8, 8, 3, 2, 0, 9, 0, 9, -3, -2, -1, -3, -1, 3, -4, 1, -5, 1, -11, -3, -9, -5, -11, -11, -6, 4, 15, 12, 12, 0, 6, 0, 3, 0, 8, 9, -4, 4, 5, -1, 6, -1, -6, -2, -4, -4, 3, -12, 0, -7, -2, -6, -9, -7, -5, 11, 8, 2, 7, 10, 13, 7, 12, 3, 10, -2, 11, -5, -4, -3, -4, -3, -9, -3, 2, -2, -1, -2, -5, 0, -1, -8, 3, -8, 1, 0, 6, 3, 0, -1, 12, -2, 8, -1, -1, -2, 10, 0, -4, -4, 2, -1, 6, -1, -4, 0, -10, 0, -6, -8, 0, 0, 2, -8, -3, 2, 6, 10, 2, 1, -3, -3, -1, 9, 6, -4, 8, -1, 8, 5, 9, 4, -9, -1, -1, -10, -5, -3, 5, 2, 0, -6, -9, -2, -8, -2, 11, 0, 5, 1, 4, 9, 0, -1, 1, 0, 0, 4, 0, 2, 0, -7, 3, 0, 6, -3, -8, 0, -2, -1, 3, -7, -10, 3, -11, -2, 5, 12, -3, 6, 8, -1, 4, 9, 9, 5, -5, 10, 9, 0, -1, -4, 1, -3, 0, -4, -9, 1, 5, -1, -1, -6, -3, -8, 0, 9, 9, 8, -2, 8, 10, 4, 2, -5, 6, 2, 7, 1, 1, 11, -2, -5, -4, -4, -4, 5, 0, -5, 2, 2, 5, 5, -2, -9, 4, 7, 10, 9, 8, 8, -3, 2, 6, 7, 0, -3, 5, 7, 3, 8, 1, 0, 10, -2, 5, 2, 5, 0, 0, -4, 0, 6, 5, -3, -3, -5, 8, 7, 10, 1, -1, 6, -6, 9, 2, -6, 5, -6, 3, 8, 7, 2, 5, 0, 7, 7, -2, -1, -5, 0, -2, -2, 6, -3, -10, 4, -2, 6, 2, -3, 7, 1, -5, -3, -5, 7, 0, 2, -5, -5, -2, 9, 4, 0, -2, 0, 5, 4, 1, 0, -8, -7, 0, -8, -12,
    -- filter=0 channel=4
    4, -8, -6, -3, 0, -6, -5, 0, 5, -3, -6, 4, -6, -3, -9, 4, -8, -8, 0, -9, -5, -11, -11, -8, -10, 0, -2, -10, -12, -9, -4, 0, 4, 7, 4, 4, 2, 0, 0, -3, 0, 2, -7, -4, -5, -9, -8, -5, -8, -9, -1, 2, -8, 4, -3, -4, 0, 0, 0, -8, 0, -5, 0, -6, 1, -3, -5, -4, -1, -1, 4, 4, 0, 2, 7, 7, 1, -9, 3, -9, -1, -5, 0, 2, -6, 5, -7, 4, 0, -4, -8, -6, -5, -4, 0, 6, 6, -4, 7, -1, 0, 6, 2, 4, -5, -1, 0, -8, 6, 1, -6, -10, -3, 1, -4, -9, 5, 5, -9, -6, -7, -3, 8, -2, -4, 3, 8, 3, 7, 2, 1, -8, -3, 0, -3, -8, 2, 1, 6, -1, -8, 6, 2, -3, -8, -1, 0, -9, -7, -6, 5, -2, 9, 3, -1, 9, -3, 9, -2, 3, 0, -1, 2, 8, 0, -3, 0, -1, 2, 0, -1, 4, -10, 0, 4, -6, -4, -3, -3, 4, 0, 0, -1, 2, -3, 8, -2, -6, 7, 2, 3, 5, -7, 6, 3, 3, 0, 5, -1, -6, -9, -5, 4, -6, 0, -1, 2, -5, 5, -2, 4, 5, 1, 5, -5, 2, -5, -2, 0, 0, -4, -1, -8, 6, -8, -1, 2, 0, -7, -5, 3, 0, 2, -8, 0, -2, -5, -1, -6, -9, 7, -2, 0, 8, 8, -3, 0, -3, 0, 6, -1, 4, -2, -6, 0, 3, 0, -1, -7, -8, -5, -8, 4, 4, 4, -1, -5, 2, -6, -6, -5, 4, -2, 8, 6, 3, 2, 4, 7, 6, -1, -7, -1, 4, -6, 5, -4, -4, -6, 1, 0, -9, -8, 3, -8, -4, -6, -4, 5, -4, -7, -3, 3, -5, 2, 1, -3, -2, -4, 2, -5, -2, -6, 0, -8, 0, 4, -8, 0, -4, -7, -7, 0, -9, -7, 4, 2, 0, -2, 1, 6, 5, 10, -1, 0, 0, 3, -1, 8, -4, 7, 6, 5, 6, -6, 7, -8, 4, 0, -6, 0, -6, 0, 0, 0, -9, -7, 4, 1, 0, -7, -5, 5, 2, -2, 5, 5, 0, 2, -1, -4, -3, 0, 3, -1, 3, 5, -7, 2, 0, 1, -2, 1, -3, -3, -8, 6, -3, 5, -4, -1, 2, -2, -5, -1, -3, 6, 7, -3, -5, -6, 6, -3, 4, 0, -3, 7, -5, 3, -3, 0, -5, 2, 0, 2, 3, -3, -8, -7, -2, -1, -6, 6, -5, 9, 7, 6, 0, -2, 5, -5, -5, -5, -7, 8, 2, 2, -6, -3, 1, -7, -3, 1, 1, -3, 6, -6, -7, -7, -9, -4, 1, 4, -1, 1, 4, -3, -5, 2, -4, -5, -7, 1, 2, -3, 4, -7, -4, 2, -7, -6, -2, 3, 0, -5, -1, -9, 2, -7, -2, 5, -2, 3, -5, -6, 3, 0, 6, 2, -1, 3, 5, -4, 0, -7, 6, -6, -4, 0, 1, 5, -4, 5, 6, 0, 1, -7, -2, -5, -9, -4, 4, -4, 7, 8, -2, 1, 1, -3, 3, -2, 0, 5, 8, -6, 1, -5, 3, 3, 4, 5, -9, -2, 0, 5, 1, 2, -5, -1, 3, -5, 2, -5, 0, 9, -6, 3, 1, 4, 8, 1, -5, -7, 8, -5, 0, 2, 5, -3, -6, 5, 5, 4, 0, -1, -9, 0, -4, 0, 2, -4, 5, -3, -1, 9, 7, -2, 7, -1, -7, 1, 4, -4, -1, -6, 2, 2, 0, 0, 4, 0, -6, -5, 0, 4, 0, -5, 0, 2, 4, 7, -6, 5, -5, 0, 7, -5, 5, -2, 0, 2, -5, 1, -2, -6, -4, 6, 3, 6, -2, 3, 0, -1, -6, -8, 1, -5, -7, -2, 2, -2, 0, -5, -5, -3, 1, -5, -5, 6, 8, 6, 2, 7, -2, 1, -1, -4, -8, -6, -5, -8, 0, -3, -6, -10, 2, 0, 0, 0, -6, -4, 8, 0, 0, -3, -6, -5, 4, 3, -8, -6, 3, -3, 7, -4, -7, -1, 0, 2, 3, -6, -2, 3, -9, 0, -7, -9, -2, -10, 2, 1, -7, 0, 0, 9, 0, 2, -2, -6, -6, -7, 7, -6, 7, -2, 5, 6, 1, -4, 3, -5, 6, 2, -2, -3, -2, -8, -8, -1, 0, -4, -3, -3, -1, -5, 2, 0, 3, 6, -2, 7, 8, -1, 4, -4, 0, -2, -1, -8, -9, 3, -10, -9, 4, 0, -1, -7, 5, -8, -4, -5, 8, 8, 6, -2, 9, 0, -2, 0, 9, 7, 5, 7, -6, 0, 1, -7, -2, -7, -3, -3, -8, -7, 6, -5, 0, -4, -5, 1, -11, -9, 2, 1, 9, 9, 3, 2, 7, -3, 2, -6, -1, -2, 3, -4, 4, 2, -8, -4, -8, 0, -1, 0, -10, 0, -9, -2, -7, -1, 0, -7, 4, 3, -2, 1, -5, -1, 8, -2, -5, -5, 3, 8, 0, 1, 0, 1, 2, -2, -4, -3, -1, -8, -7, 0, 6, -6, -2, 4, -11, 4, 3, 0, 7, -5, -1, 4, -2, -7, -5, 2, 3, -8, -6, 2, -7, 1, -1, -7, 2, 0, 3, -8, 6, -1, -4, -9, 4, 0, -6, 1, 0, -7, -3, 0, -5, -4, -5, -3, -1, 2, 3, -1, 0, 4, -3, 4, -2, 2, 0, 2, -4, -1, -11, -5, -1, -3, -12, 0, -1,
    -- filter=0 channel=5
    1, 10, 0, 13, 3, 10, 2, -1, -5, 6, 8, -1, 6, 0, 9, 9, -4, 8, 0, 7, 6, 5, -1, -4, -1, 3, -2, -9, -2, 2, 10, 11, 4, 10, 4, 10, 13, 5, 0, 7, 5, 6, 3, 16, 13, 12, 5, 8, 9, 1, -3, 11, -3, 4, 6, 8, 9, 5, 3, -9, 0, 14, 10, 17, 17, 17, 19, 17, 13, 14, 14, 6, 19, 6, 5, 9, 4, 15, 18, 1, 5, 13, 13, -1, -2, 0, 4, -4, -9, -3, 10, 1, 15, 16, 8, 19, 10, 20, 6, 10, 13, 10, 20, 14, 20, 5, 4, 14, 4, 16, 9, 0, 5, 11, 0, 0, -2, 4, 4, -5, 0, 15, 9, 14, 15, 12, 13, 22, 6, 10, 20, 10, 13, 15, 13, 11, 12, 6, 7, -3, 0, 4, 5, -1, 7, 5, 0, 10, 1, -3, 3, 3, 11, 21, 21, 14, 16, 15, 18, 4, 14, 13, 12, 11, 1, 1, 8, 8, 7, -1, -4, -2, 5, 7, 7, -2, -5, 6, 2, -8, 6, 4, 19, 7, 6, 8, 9, 10, 13, 2, 2, 9, 7, 5, -2, 3, -6, -5, 2, 5, 0, -1, 4, 5, 3, 3, -1, -8, 2, -1, 5, 6, 12, 10, 2, 2, -2, 0, 11, 0, 13, 4, 10, 8, 4, -5, 6, 4, 1, -4, -10, -5, -9, -4, -8, 1, 1, 3, 0, -7, -5, 4, 10, 7, -2, 0, -6, 0, 8, 8, 7, 6, 4, -1, 7, 3, -4, -5, -11, -4, -10, -9, -8, -7, 0, -3, 2, -2, -13, -7, -2, 2, 12, 3, -4, 3, 2, 0, 5, -4, -2, 2, 6, -4, -1, -5, -9, -2, -15, -12, -7, -14, -12, -5, -16, -7, 3, 3, -4, -18, 5, 8, 0, -3, 0, -6, -10, -10, -11, 5, -1, 2, 0, 10, -3, 5, 0, -11, -17, -6, -20, -9, -9, -7, -16, -8, -4, -13, -13, -11, 0, -6, -2, -3, -6, -12, -4, -5, 0, 2, -1, 0, 8, -2, 5, -6, -6, -6, -10, -18, -20, -13, -5, -17, -9, -10, -6, -1, -10, -11, 3, 3, 2, 6, -11, -10, 0, -9, -7, -9, 0, -1, -4, -5, -4, -8, -1, -2, -5, -10, -9, -16, -6, -20, -13, -4, 0, 1, -7, -9, -6, 2, 2, -1, -1, -6, -2, -13, -1, -8, -7, -1, -4, 0, 0, -5, -13, -2, -18, -13, -18, -7, -20, -6, -11, -8, -14, -7, -14, -10, -8, -1, 0, -1, -6, -8, -14, -13, -3, -7, 5, 4, 2, 5, -1, 0, 0, -4, -7, -12, -13, -6, -8, -12, -8, -17, -2, -12, -2, -15, -1, -7, 5, -7, -12, -10, -5, -12, 2, -2, 2, -3, 7, 1, 2, -11, -1, -16, -6, -7, -21, -10, -18, -12, -15, -13, -11, -14, 0, -5, -8, 3, -4, -6, -9, -15, -2, -11, -9, -8, 6, -6, -2, 4, -1, -13, -3, -5, -5, -21, -7, -18, -14, -14, -18, -16, 0, -13, -16, -15, -10, 2, 4, -6, 2, -2, -2, 1, -7, -5, 0, 0, 6, -5, -2, 1, -16, -10, -17, -13, -14, -7, -18, -10, -9, -14, 0, -13, -2, -16, 2, 6, 4, 2, 0, 1, -10, -4, -5, 6, -5, 0, 4, 6, 4, -12, -12, -17, -19, -13, -9, -12, -18, -11, -12, -17, 1, -7, -10, -11, 5, 8, -3, 0, 4, -6, -8, -1, 5, 5, -3, -2, 4, -6, 6, 4, -1, -2, -11, -18, -20, -17, -8, -11, -6, -14, -11, 0, -4, -20, -7, -3, 11, 12, 7, -5, 0, 5, -8, 6, -5, 2, 0, -2, -2, -7, -1, -9, -9, -7, -3, -5, -9, -11, 0, 1, -1, -8, -12, -10, 2, 4, 4, 7, 10, 2, 0, 4, -4, 7, 9, 6, 3, 11, -3, 4, -4, 0, -8, -8, -13, -10, -8, -14, -8, 3, -9, -5, 1, -6, 4, -1, 13, 15, 16, 1, 9, 9, -4, 1, 7, 9, 8, 11, -2, 2, 2, 3, -9, -10, 3, -2, -8, 0, -1, -5, -5, 1, 0, -2, -3, 5, 13, 7, 16, 0, 11, 9, 1, 0, 12, 9, 0, 4, 8, -3, 2, 2, 4, -4, 5, -2, -3, -8, 6, -6, -4, -4, -2, -1, 10, 3, 20, 20, 12, 5, 10, 15, 7, 0, 14, 17, 2, 14, 10, 4, 9, 6, -3, 7, -2, -5, 0, 0, -1, 12, 7, -1, -3, -8, 0, 11, 7, 15, 20, 17, 8, 19, 19, 19, 20, 4, 5, 18, 2, 11, 9, 1, 4, 4, 9, 0, 12, -1, 5, 0, 4, 4, -4, 0, -5, 1, 11, 24, 19, 14, 7, 9, 10, 10, 18, 6, 14, 16, 17, 18, 12, 8, 6, 3, 6, 3, 1, 0, 7, -2, 10, 2, 0, -4, 7, 1, 15, 10, 17, 21, 5, 9, 11, 5, 6, 6, 11, 13, 8, 10, 12, 1, 12, 9, 12, 7, 1, 7, 11, 12, 3, -5, 0, -9, 3, 7, 9, 1, 9, 12, 3, 5, 9, 3, 6, 14, -1, 0, 2, 1, 13, 9, 4, 10, 1, 9, 7, 3, 5, 8, 6, -5, -1, 3, -2, 8, 11, 3, 7, 0, 6, 9, 0, -1, 2, -2, -1, -1, -4, 0, 0, -3, -2, 4, 0, -3, -6, -5, 4, -2, 4, 0, -5, -12,
    -- filter=0 channel=6
    -5, -6, -1, 1, 0, -14, -8, -7, -9, -4, -2, -3, -10, -7, -11, -9, -8, 1, 2, -2, -9, -12, -5, -2, -15, -3, -6, -5, -15, -23, 3, 6, -4, 8, -4, -3, 5, -9, -6, -6, 4, 4, -1, -7, 5, -3, 6, 0, 0, 5, -7, 0, -8, -7, -9, -2, -8, -3, 1, -5, 0, 10, 1, 10, 1, 0, -2, 6, 4, 0, -5, 7, 0, 8, 7, 4, 1, 3, 0, -8, 2, 6, 3, -2, 3, -5, -1, 2, -9, -1, -1, 7, 12, 9, 9, -1, 0, 5, -3, 6, 5, -1, 10, 7, 14, 5, 0, 10, -1, -2, -3, 5, -8, 0, 0, 2, 1, -1, 1, -9, 5, -1, -1, 2, 9, -4, 6, -6, -7, 2, -3, -1, 3, 4, 6, 9, 14, 5, -1, 7, 2, 5, 2, -4, -5, 3, -6, 0, -2, -4, 2, 0, 3, 8, -5, 5, 5, 1, 6, 8, 11, 2, 10, 18, 5, 7, 10, 9, 8, 6, 5, -4, 3, -7, -1, -7, 6, -1, 0, -3, 0, 9, 7, 4, 4, 5, 1, 8, 2, 3, 3, 1, 13, 3, 5, 7, 14, -1, 10, 3, 3, 6, 7, -3, -1, -6, -6, 5, -1, -9, 4, 10, 6, 6, 0, -4, 7, 0, -5, -5, 5, 3, 7, 5, 6, 2, 2, 14, 12, 10, 11, 0, 1, -2, -5, 5, -7, 1, 5, -1, 9, 11, 3, 8, 3, 9, 5, -3, -3, 5, 5, 11, 2, -1, 1, 3, -3, 9, 0, -2, 9, -3, 2, 7, -2, 4, -5, 4, -1, -1, -2, 0, 14, 6, 10, -4, 1, 11, 0, 11, -5, 9, -2, 3, 8, 4, 3, 0, 6, 2, 2, 9, 0, 8, 1, -1, 8, 5, 6, -7, 11, 7, 8, 1, -1, 2, 3, 7, 1, 10, 4, 7, 1, 0, -1, -4, 1, -1, 1, -6, 9, 4, 7, -2, 13, 7, -3, -1, 1, 2, 8, 5, 3, 7, 6, 13, 4, 7, -2, 12, 7, 1, -7, 0, -9, 0, -17, -17, -3, -3, 3, 8, 2, 11, 15, 12, 5, 5, -1, -7, 12, 0, -1, 13, 6, 10, 13, 2, 0, 9, 5, -6, 2, -4, -9, -2, -18, -4, -7, -8, 2, -1, 15, 9, 8, 10, 1, 0, 6, -3, 2, 10, 14, 2, 1, 11, 5, 10, 11, 5, 6, 9, -7, 0, -4, -3, -20, -6, -15, -3, -2, 4, 1, 14, 2, 5, 0, 3, 7, 7, 5, 8, 0, 0, 4, 7, 9, 3, 3, 14, 3, 8, -9, 1, -5, -8, -13, -11, -9, -9, -8, 11, 5, 8, 6, 4, 9, 3, 8, -1, 0, 10, 4, 2, 2, 7, 19, 7, 7, 4, -1, 0, 4, -2, -4, -5, -6, -14, -7, -6, -1, 9, 12, 4, 5, 6, 11, 1, 10, -1, 0, 5, 9, 10, 14, 10, 14, 10, 4, 13, -1, 10, 2, -8, -14, -11, -11, -18, -6, -7, 0, 3, 10, 15, 8, 0, 5, 8, 0, 0, -2, 0, 7, 3, 15, 12, 10, 9, 15, 13, 10, 8, 5, -7, -7, -6, -17, -10, -13, 1, -3, 7, 5, 4, 15, 0, -3, 6, 8, 5, 12, 3, 14, 11, 2, 6, 8, 14, 7, 7, 9, 7, 7, -5, -5, 0, -13, -10, 0, 1, 10, 0, 11, 14, 11, 7, -3, -1, 0, 1, 2, 3, 5, 7, 7, 10, -1, 6, 12, 2, 6, 0, 9, 4, -6, -9, 2, 3, 1, 8, 6, 0, 1, 5, -3, 6, -3, 5, 10, -1, 4, -1, 13, 13, 3, 0, -1, 3, 0, 3, -3, 8, 0, -4, -2, 1, 8, -2, 9, -3, 5, 8, 7, -1, 5, 8, 5, 0, 1, -7, 2, 2, 13, 3, 9, 11, 0, 1, 10, 0, 3, -2, 3, -2, 2, 4, 9, 2, 0, -2, 0, 0, 10, 0, 0, -6, 1, -7, 0, -4, 7, 3, 16, 5, -2, 2, 10, -4, -2, -1, -4, 1, -1, 3, 3, 11, 3, 12, 1, 6, -5, 0, -5, 0, -1, -6, 5, -6, 7, 2, 1, 3, 2, 10, 7, 2, -1, 5, -1, 2, 11, 10, 12, 1, 7, 4, 14, 7, -2, 3, 9, 0, -5, 0, -5, -3, -2, 4, 2, -2, -5, -1, 2, 0, -4, 3, 5, -7, 1, 4, 6, 9, 11, 14, 8, 14, 13, 14, 1, 6, 1, 4, -9, 0, -2, 2, -5, -4, -6, -7, 9, 10, 5, 5, 9, -1, -1, -4, 1, 8, -3, 4, 8, 5, 1, 6, 9, 2, 7, -5, -7, 3, -7, -9, 4, 4, 3, 4, 5, -13, 7, 1, 5, 8, 0, -2, 5, 5, 3, 6, 10, -3, 5, 6, 13, 9, -1, -1, -3, 4, 0, 7, 3, -1, -6, 1, 0, -6, -3, -8, 8, 9, 8, 9, 6, 2, -7, 6, 5, 4, 0, 4, 0, 9, 6, 4, -3, 7, 0, 1, 7, 6, -8, -3, 2, 0, -9, -6, -4, -14, -8, 5, 10, 0, -5, 0, -7, -1, -1, -9, -7, 2, 4, -1, 0, -3, 4, 0, -6, 4, 3, 3, 3, -2, -9, 0, 2, -7, -8, -17, -15, -5, -9, -2, 1, -1, -7, 3, 1, -2, 1, -7, -4, -10, 0, -5, -3, 4, -2, 0, -9, -9, -6, -8, -12, -10, -14, -18, -4, -17,
    -- filter=0 channel=7
    -12, -12, 0, -8, -12, -9, 3, 7, -3, 1, 0, -6, 3, -2, 3, 6, 0, 7, 0, -5, 5, -3, 1, 7, 0, 9, 6, 6, -1, -9, -6, -15, 2, -4, -6, 0, 0, 7, -4, 8, 0, -3, 1, -6, -6, 2, -3, -3, 5, 6, 5, 9, 4, -1, 5, 8, 7, 13, 7, 0, -17, -9, -3, 5, 2, 3, 4, 1, 4, 5, -3, 7, -5, 0, 1, 6, 7, -7, 4, 5, -4, -4, 0, 4, 1, 0, 0, 15, 3, 2, -3, -8, -9, -6, 3, -1, 6, 7, 12, 5, -1, 7, 4, -8, -2, -2, -5, -4, 2, -4, 0, -3, 0, 11, 6, -2, 5, 2, 13, 5, -15, -1, 1, -2, 5, 7, 0, 15, 2, 1, 0, 10, -4, -7, 4, -4, -4, 0, -4, 0, -4, 7, 3, -4, 5, 0, 8, 0, 4, 0, -12, -3, 1, 7, 3, 3, 5, 18, 10, 7, 0, 4, 3, 9, -4, 3, -5, -4, 4, -9, -7, 0, 0, 0, 5, -1, 3, 2, 1, -1, -9, -3, 3, -6, 2, -1, 8, 9, 12, 4, 2, 0, 6, 7, 1, 6, 3, 4, -7, 5, -3, 0, 1, -6, -3, -2, 0, -2, 8, -2, -11, -1, -6, 0, 4, 12, 12, 17, 19, 6, 18, 13, 16, 6, 11, -1, 6, -4, 0, 1, -10, 1, 1, 3, -7, -1, -4, 5, 13, 3, -7, -12, 0, 3, 0, -1, 3, 16, 14, 10, 7, 8, 17, 17, 6, 9, 6, 7, -1, -7, -3, -7, -5, -2, 2, -8, -4, 5, 0, 0, -2, -13, 1, -5, -3, 5, -2, 11, 14, 6, 17, 12, 13, 18, 7, 8, 14, -4, -10, -14, -15, -7, -10, -9, -6, -8, 2, 0, 4, 3, -6, -6, -9, -4, 3, -5, -4, 9, 9, 3, 18, 9, 6, 10, 7, 13, 17, 12, 0, -12, -6, -4, -1, 0, -3, 0, 5, 2, 8, -4, 0, -9, -4, -12, -13, -7, -2, 7, 2, 3, 3, 9, 9, 10, 13, 8, 16, 9, -4, -2, -8, -8, -11, -14, -9, -6, 5, -4, 11, 1, -9, 0, -12, -11, -7, -6, -9, -5, -3, 11, 14, 3, 9, 14, 6, 22, 17, 6, 6, -1, -10, -6, -4, -6, -6, -7, -3, 0, 1, -1, -10, -5, 0, -11, -9, 0, -12, -10, 4, 12, 11, 0, 10, 13, 20, 11, 9, 10, 8, -4, -9, -10, -4, -11, 1, -3, 5, -4, 8, 2, -13, -11, 0, -1, -4, -17, -12, -4, 1, -4, 12, 13, 14, 3, 19, 20, 13, 8, 0, -15, -13, -8, -7, -16, -7, -10, 3, -4, 11, 9, 2, -4, -11, -13, -3, -14, -8, -9, 0, -1, 6, -1, 16, 7, 8, 10, 10, 14, -8, -10, -16, -18, -14, -3, -4, -9, 1, 0, 1, 5, -13, 2, -12, -12, -5, -16, -8, -3, -4, 8, 9, 4, 9, 8, 11, 15, 12, 7, -4, 0, -15, -3, -15, -12, 3, 3, 0, 5, -2, 9, -3, -1, -5, -2, -15, -5, -6, 0, -6, -3, 4, 14, 14, 14, 12, 18, 10, 12, 6, -7, -7, -16, -15, -2, -1, 0, -6, 4, -3, -4, -3, 1, 0, -11, 0, -11, -3, 6, 3, 10, 11, 11, 7, 16, 9, 9, 18, 15, 3, 3, -8, -13, 0, -2, 0, 2, -6, 3, 11, 9, -2, -6, -7, 2, 1, 0, -2, 9, 6, 12, 9, 17, 14, 10, 17, 12, 12, 1, -2, -2, -4, -2, -7, -5, -6, 0, 6, 8, 9, 4, 0, -9, -9, 0, 3, 1, 11, 12, 10, 16, 15, 12, 14, 8, 4, 16, 7, -4, -2, -7, -15, -5, -2, -9, -9, 0, 0, -4, 11, 6, 2, -5, -11, 4, -2, 3, 8, 3, 15, 7, 17, 10, 17, 14, 7, 11, 2, -2, -2, 0, -2, -1, 0, -3, -2, -11, 0, -2, 12, -4, -6, -5, -8, 0, 5, -2, 2, 5, 6, 17, 6, 11, 13, -1, 12, 8, -5, 6, -6, 1, -12, -15, -9, -7, 0, 0, 1, 1, 3, 6, -10, -1, -2, 2, 1, -1, 3, 5, 10, 13, 3, 5, 8, 5, 3, 0, -4, -7, 2, 4, -12, -3, 2, -1, -2, 0, 5, 10, -1, 9, -5, -10, -7, 0, 5, 2, 1, 5, 7, 9, -2, 0, 0, 0, 3, -1, -8, -9, 0, 1, 3, 1, -2, -4, -7, -9, 8, 7, 5, 13, -5, 5, -9, 7, 1, 10, 6, 10, 6, 3, 1, 4, 4, -8, 4, -11, 0, -8, 2, -11, -3, -6, -9, 6, 6, 0, 9, 13, 0, 1, -2, -3, -5, 1, -7, 7, 2, 12, 5, 2, 4, 0, -12, -4, -9, -9, -7, -3, 3, -4, 2, 8, 7, 6, 0, 7, 3, 0, 0, -1, -11, 2, 2, 3, -5, 4, 7, 12, 3, 2, -2, -7, 5, 0, 0, -1, 0, 5, -1, 4, 8, 3, -3, 0, 13, 12, 0, 0, 11, -3, -10, -4, -3, 0, 5, 8, 2, 9, 2, 2, -4, 7, 6, 0, 2, 2, 3, -5, -4, 4, 7, -3, 10, 10, 11, 0, 2, 12, 7, -1, -12, -12, -12, -13, -11, 2, 3, -6, 7, -7, -1, 0, 6, 0, 4, 6, -5, 2, 1, -5, 3, -6, 9, 8, 7, 6, 4, 4, -3, -10,
    -- filter=0 channel=8
    3, 3, 3, 2, -10, -3, 1, -13, 1, 1, 1, -7, -2, 1, -13, -1, 2, -2, -2, 6, 8, 0, 1, 1, 15, 6, 8, 10, 21, 18, 2, -12, -5, -2, -10, -11, -18, -8, -15, -3, -16, -2, -10, -1, -8, -3, 0, -2, -3, -11, -5, -6, 5, 0, 8, 4, 10, 13, 13, 25, 2, -5, -5, -4, -11, -13, -5, -15, -5, -4, -10, -13, 0, -10, -9, 1, -10, -2, -7, -2, -7, 0, -2, 1, -2, -3, 9, -2, 5, 13, 0, -6, -16, -19, -5, -6, -19, -17, -5, -8, -11, -6, -10, -10, -9, -12, -10, -3, -1, -10, -4, -8, -5, 4, -6, 0, 6, 12, 12, 14, 0, -14, -13, -13, -17, -5, -21, -15, -17, -20, -8, 0, -6, -14, -11, 4, -8, 3, 3, 0, 0, 5, 2, 2, 3, -6, -4, 3, 5, 13, -2, -13, -10, -19, -13, -8, -20, -13, -9, -20, -15, -2, -5, 0, -4, -8, 8, 1, 0, -2, 6, -4, 10, -3, -4, -8, 9, 3, 9, 15, -1, -13, -2, -13, -18, -8, -7, -14, -18, -15, -3, -7, -12, -2, -2, -6, 0, 2, 11, 7, 14, 0, 6, 13, 10, -2, 11, 5, 14, 14, -9, -8, -10, -9, -18, -8, -15, -10, -13, -10, -6, -18, -5, -11, -3, -7, -6, -5, 0, 14, 1, 15, 4, 3, 0, 4, 9, 10, 11, 19, -4, -3, -4, -8, -10, -5, -16, -8, -6, -6, -13, -19, -14, -15, 0, -8, 7, 7, 9, 14, 10, 14, 14, 13, 3, 9, 6, 12, 7, 14, 0, 0, -7, -13, -12, -20, -8, -8, -15, -19, -7, -5, -6, -6, -4, 1, 8, -4, -2, 10, 2, 6, 0, 8, 13, 13, 7, 12, 17, 12, -3, -17, -17, -14, -19, -18, -9, -15, -10, -9, -14, -16, -11, -5, 0, -6, 2, 0, 9, 2, 15, 8, 14, 14, -1, 7, 3, 2, 15, 13, -2, -1, -11, -18, -19, -19, -17, -15, -14, -11, -23, -8, -9, -2, 2, 5, 9, 8, -2, 5, 5, 12, 11, 13, 10, 8, 0, 9, 17, 10, 0, -15, -11, -11, -19, -14, -16, -22, -16, -16, -16, -11, -15, 1, -6, 2, 3, 0, -4, 6, 6, 11, 11, 8, 15, 12, 11, 8, 9, 24, -1, -7, -7, -13, -12, -6, -6, -10, -21, -15, -6, -9, -4, -10, -3, -1, -4, 7, 4, 5, 9, 16, 8, 13, 1, 12, 1, 9, 18, 16, -8, -4, -5, -12, -12, -11, -14, -18, -24, -14, -12, -13, -11, -4, -2, -2, 4, -2, 10, 8, 0, 8, 5, 11, 8, 13, 7, 5, 12, 25, -11, -1, -4, -12, -6, -12, -12, -16, -9, -14, -9, -6, -7, -5, 2, 3, 1, 3, -1, 9, 7, 6, 17, 14, 3, 0, 10, 3, 8, 13, -9, -13, -7, -9, -15, -6, -12, -17, -24, -14, -22, -19, -2, -6, 0, 1, 3, 1, 1, 5, 3, 5, 1, 16, 11, 2, 13, 6, 11, 24, -1, -12, -15, -10, -6, -15, -15, -9, -21, -14, -13, -9, -12, -1, 0, 4, -7, 7, 11, -2, 11, 8, 12, 18, 16, 9, 11, 6, 14, 11, -10, -1, -4, -8, -18, -11, -9, -9, -17, -8, -21, -4, -9, 0, 1, -8, 2, -1, 10, 8, 12, 6, 3, 8, 15, 0, 0, 11, 14, 22, -6, -7, -9, -11, -9, -7, -8, -6, -18, -15, -21, -8, -17, -7, -6, 3, 0, 0, 9, 9, 9, 2, 15, 6, 14, 12, 11, 5, 20, 16, -10, -6, -8, -14, -5, -6, -5, -16, -15, -22, -16, -4, -16, -15, -8, 0, -2, 10, 11, 9, 12, 3, 1, 10, 13, 9, 2, 11, 16, 25, -4, -14, -14, -16, -19, -8, -12, -19, -8, -20, -17, -16, -5, -4, 0, -6, 7, 5, 0, 8, 7, 1, 9, 3, 5, 6, 0, 0, 15, 18, -2, -1, -17, -7, -13, -19, -6, -19, -5, -5, -13, -14, -14, -3, 3, 4, 9, 6, 8, 5, 14, 1, 2, 4, -2, 3, 11, 9, 16, 24, -5, -15, -15, -10, -8, -12, -5, -6, -21, -7, -15, -9, -4, 1, -10, -6, 1, -5, 8, 0, 1, 10, 14, 9, 5, 3, 7, 13, 15, 19, 1, -4, -7, -20, -15, -14, -14, -20, -9, -8, -4, -14, -12, -2, -3, -3, -4, -3, 0, 0, -1, 7, 11, 7, -3, 0, -1, 7, 5, 17, -1, -4, -6, -4, -17, -14, -16, -10, -17, -14, -4, -4, -12, -5, -8, 0, -3, 4, -6, 6, 9, 0, 8, -1, -4, 5, 8, -3, 9, 17, 5, -4, -9, -10, -7, -10, -7, -11, -8, -19, -2, -11, -9, 0, -8, 2, -8, -1, -3, -7, 2, -7, -5, -7, -9, -2, 3, 7, 0, 9, 2, -1, -8, -16, -11, -10, -8, -13, -13, -6, -6, -18, -17, -8, -11, -10, -14, 0, 2, 0, -4, 0, -8, 0, -3, 6, 2, 0, 10, 15, -1, -10, -6, -5, -4, -18, -8, -4, -15, -3, -18, -5, -15, -9, -5, -8, -1, 1, -11, -3, -1, -11, -4, 1, 1, -1, 2, 15, 3, 13, 5, 0, 1, -9, -1, 3, -5, -6, -4, 0, -3, -3, -4, -7, -13, -7, -1, 0, 4, 3, 4, 2, -1, 0, 0, -1, 8, 14, 10, 24,
    -- filter=0 channel=9
    -16, -1, -14, -6, -12, -3, -3, 6, 0, 4, 6, 16, 18, 8, 16, 13, 10, 19, 9, 17, 22, 17, 16, 7, 0, 0, 3, 2, 0, -17, -15, -11, -12, -13, -6, -6, 1, -13, -5, -9, 1, 2, 4, 1, 6, 13, 13, 8, 17, 21, 13, 5, 13, 5, 10, -1, -4, 3, -11, -3, 0, -15, -17, -18, -4, -17, -10, -1, 0, -9, -5, 3, 4, 2, -2, 14, 12, 15, 9, 4, 10, 15, 8, 7, 4, 1, -1, 5, -3, -1, -14, -6, -7, -16, -11, -11, -19, -17, -14, -3, -2, 3, 2, 3, 6, 8, 9, 8, 10, 16, 9, 8, 3, 9, 8, 7, 7, 1, -7, -9, -8, -3, -20, -14, -12, -10, -18, -13, -4, -5, -1, -12, 3, -3, -2, -2, 4, -1, -1, 5, 10, 7, 2, 0, 5, 5, 3, 0, 0, -2, -12, -8, -13, -21, -24, -16, -10, -9, -11, -1, 1, -1, 4, -3, -5, 8, -3, -1, 0, 7, 12, 14, 10, 9, 0, 6, 2, -3, -4, 4, -8, -5, -13, -20, -14, -10, -9, -19, -9, -1, -12, 0, 5, 2, 3, 3, 0, -3, 11, 15, 9, 5, 13, 8, 16, 8, 3, 4, 5, 4, -6, -6, -20, -9, -9, -3, -10, -12, -11, -4, 0, 1, 0, -4, 6, -2, -1, 6, 9, 6, 2, 0, 12, 12, 3, 15, 5, 11, 0, 4, -9, -15, -18, -13, -8, -15, -5, -7, -5, 1, 0, 0, 0, 7, 0, 0, -5, 3, 1, -3, 14, 11, 4, 4, 15, 3, -1, 0, -3, 6, 1, -9, -14, -2, -11, -1, -2, -13, -3, -9, 4, -6, 3, 7, -7, 4, -10, -5, 6, 0, 11, 9, 11, 12, 4, 16, 3, 11, 3, 4, -11, -5, -4, -12, -11, 0, 3, -7, 4, -7, 2, 6, 2, 0, -7, -4, -8, -6, -3, 10, 2, 13, 5, 11, 4, 12, 10, -2, 9, 5, 5, -4, 0, -14, 3, 5, 0, -6, -5, 8, -3, 9, 2, 1, -5, -3, 0, -3, -9, 7, 0, 13, 2, 9, 14, 2, 9, 5, 2, 0, -9, 0, -9, -10, 1, -3, 1, 5, -1, -1, -2, 0, 1, 3, 2, -15, -5, -12, 1, 5, 7, 13, 10, 3, 0, 11, 9, 4, 0, 2, -2, -5, -10, -10, 0, -1, 3, 1, -4, 0, -4, -5, -2, 2, -12, -4, -15, -7, -16, -1, -2, 11, 8, 2, 0, -1, 1, -5, 3, -2, 1, -14, -3, -5, -2, 9, 10, 3, -2, -5, 3, 0, 5, 0, -10, -11, -12, -10, -16, -11, 0, 13, 15, 13, 9, -2, -2, -4, 0, -8, -5, -6, -10, 0, -3, -4, -1, 3, 6, -2, 2, 0, -4, -2, -10, -14, -20, -20, -8, 3, 5, 9, 11, 9, 0, 4, 7, 5, -3, 2, -7, -5, -16, 0, 7, 9, 10, 8, 9, -2, -6, -3, 6, 2, -1, -7, -8, -8, -8, -5, 1, 11, 12, 15, 5, 2, 3, -3, -4, 3, 0, -8, -5, -4, 5, -2, 9, -6, 8, 7, 4, -1, -3, 5, -3, -13, -12, -7, -4, -2, 10, 9, 8, 2, 9, 13, 2, 0, -4, 7, -6, -11, -10, -12, -3, 5, 8, -7, 1, -5, 0, 0, 1, 9, -7, 3, -6, -6, -8, 1, 1, 11, 8, 10, 2, 9, 10, 8, -3, 1, -11, -4, -15, -15, -10, -1, -3, -4, 2, -7, 7, -2, -4, -2, 0, -5, -7, 0, -4, -2, 12, 9, 1, 12, 13, 14, 0, 2, -5, 5, -5, -7, -20, -17, -9, -5, 2, -12, 0, 1, -7, 5, 12, -2, 0, 0, -3, -3, -5, 10, 4, 9, 5, 10, 13, 15, 12, 0, 0, 0, -1, -1, -9, -21, -6, -4, -15, -14, -8, -5, 5, 0, 2, -1, -5, 1, 6, 2, 1, 13, 4, 4, 1, 16, 12, 7, 6, 7, -1, -4, 1, -15, -15, -15, -6, -7, -12, -11, 1, -1, 3, 5, 4, 5, 5, 0, 0, -4, 4, 4, 6, 14, 14, 17, 8, 14, -4, 0, -5, -7, -4, -12, -23, -9, -10, -18, -6, -11, -13, -12, 2, 7, 4, 11, 10, 8, -5, 3, -1, 7, 3, 3, 2, 1, 15, 3, 0, -2, 3, -1, -10, -9, -20, -13, -9, -11, -14, -6, -10, 3, 0, 0, -3, 11, 9, 10, -1, 5, 14, 16, 1, 1, 14, 9, 0, 2, 2, 0, -6, 0, -6, -5, -7, -20, -11, -14, -9, -11, -14, 2, -8, -5, 11, 2, 10, 8, -2, 12, 11, 14, 1, 8, 5, -1, 2, 1, -6, 2, 0, -3, -4, -12, -17, -11, -14, -16, -17, -3, 0, -2, -3, 7, 6, 3, 9, 8, 6, 8, 9, 15, 2, 1, 14, 7, 2, -3, 2, 5, 2, -4, -3, -2, -8, -8, -13, -10, -7, 2, -2, 6, -2, 3, 0, 12, 14, 15, 7, 8, 14, 5, 11, 16, 12, 12, 6, 3, -5, -8, 2, -13, -9, 0, -1, -14, -5, -13, 0, 0, -3, -1, 3, 16, 16, 12, 16, 19, 19, 21, 9, 15, 21, 15, 3, 15, 0, 9, 6, -3, -7, 0, -6, 0, -12, -5, -8, -10, 2, 1, 5, 12, 17, 8, 19, 15, 11, 19, 11, 24, 13, 20, 22, 16, 9, 6, 0, 1, 4, -13, -6, -15,

    others => 0);
end iwght_package;
