library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 4000000) of integer;

  constant input_wght : mem := (
    -- bias
    -- layer=3
    -6641, -4126, -2619, 3887, 8492, -5286, 12928, -7389, 3259, -4088,

    -- weights
    -- layer=3 filter=0 channel=0
    -35, -46, -27, 41, 4, 59, 1, -19, 1, -21, -3, -23, 17, 35, -10, -17, 11, -53, 6, 11, 19, 2, 0, 32, 60, -6, 6, 10, 31, 59, 30, 10, -28, 13, 0, -25, 1, -9, 20, 45, -20, -30, -3, -5, -48, -21, 46, 26, 4, -3, -5, -22, 24, -22, 17, -7, 13, -76, -13, -28, -33, 20, 37, -28, -21, 14, 0, -18, 15, 3, -4, 3, 12, 1, -3, -6, 38, 21, 21, -29, -29, 3, 13, -14, -35, -6, 16, 7, 5, 3, 20, -57, 31, -22, 15, 2, -6, 19, -51, 0, -24, -10, -52, -21, 20, -17, 13, 32, -1, 23, -38, -88, -24, 75, -21, -21, 3, -8, -57, 45, -17, -1, 2, 15, 44, 4, -1, -5, 4, -9, 45, 61, 12, 27, 8, 10, -28, -5, 1, -13, 26, 27, -34, 8, 8, -12, 32, 6, -19, 6, -10, -6, 40, -17, -7, -5, 0, -28, 14, 33, 2, -2, -27, -44, -6, -64, 30, 27, 32, 1, -3, 33, -46, -24, 35, -19, 10, 0, -13, -16, 12, 21, -2, 38, 6, -29, -17, 16, 24, -2, 24, -54, -21, 20, 16, -6, 13, -22, -1, -7, -26, -9, -27, 10, 15, 40, -4, -5, 20, 18, -1, 15, 9, 0, -27, -19, 14, 15, -11, 12, 0, -34, -26, -22, -14, 2, 23, -16, -43, -1, 13, -16, 4, -25, -1, -12, -5, -21, -4, 37, 4, 41, -36, 16, 3, -35, -6, 18, -10, 35, 11, -20, 1, -21, 0, 1, 24, 17, -13, 36, 19, 36, -17, -11, -4, 41, 29, -23, -12, -11, -14, -1, -2, -25, 12, -11, 3, -12, 5, -27, -19, 8, 5, 29, 35, -31, -26, 49, -25, 13, 27, -59, 2, 22, 13, -35, -1, 33, 4, 12, -18, 16, -55, -22, 3, -4, 31, -6, 28, 15, 5, -23, 39, -48, -17, -27, -16, 2, 0, 51, 0, 25, -4, 10, -21, -4, 10, -3, -85, 12, -33, -5, 27, 1, 12, 32, -13, 31, -16, -22, -8, 41, -46, 13, 10, -9, -51, -56, 21, -19, 14, -4, 28, -3, -114, -48, -46, -8, -40, -11, -12, -20, -20, -2, 8, -55, 15, -53, -22, -29, -17, 67, -3, -25, -71, -31, -13, 50, 15, -27, -26, 0, 1, -16, 17, -32, 85, 3, -8, 1, -15, 0, -31, -47, 9, -29, -27, -12, -40, -34, 0, -2, -5, 0, -19, -9, -11, 8, 59, -25, -18, 7, -23, 1, -37, -30, -35, -71, 4, -61, 11, -1, 55, 19, 30, -22, 4, -35, -18, -47, 10, 18, 31, 21, 15, -17, -2, 4, 11, 2, 20, -58, -21, -7, 23, -23, -7, -22, -18, -31, 38, -17, 31, -10, 13, 16, 9, -7, 42, 33, 10, 14, 19, 2, 20, -15, -13, -24, 15, 13, 12, 2, 2, -9, 7, -55, 2, -18, 32, 16, 22, 3, -11, 56, -5, -37, 0, -6, -9, -13, -18, -16, -14, 15, 37, -118, -5, 26, -28, -26, 9, 8, 1, 17, -17, 7, -6, 5, 17, 18, -19, -7, -10, 10, 25, -25, 24, -24, -15, 4, -43, -39, 34, 48, -51, -2, -31, 8, 8, -21, 2, 8, 24, -3, 15, 5, 0, -21, 2, -25, -7, -51, 8, 17, -33, -35, 17, -17, -17, -24, -14, 0, -8, 2, 2, 1, 47, 3, 32, -28, 0, -8, 26, -4, -7, 0, -10, -29, -56, 27, 26, -18, -7, 10, -3, -26, -2, -35, 0, -12, -4, -41, -9, -7, 30, 10, 9, 53, 11, -41, 2, -18, -25, 20, -13, -67, 22, -3, -26, 3, 0, 16, -55, 52, -2, 17, 1, -24, -6, 43, -38, 13, 9, -13, 25, -25, -12, -53, -5, -33, -10, 29, 4, 38, -17, -8, 0, -14, -20, 23, 43, -8, -15, 46, 24, 2, -10, -7, 4, -11, 24, -25, 44, -18, -11, -7, -1, 3, -46, -16, -6, 12, 16, 20, -36, -11, 4, -37, 36, 4, -24, -24, -15, -30, -13, -24, -4, 9, -9, 52, 11, 59, -22, -78, -2, -56, 6, 3, -6, -7, 38, 34, 18, 5, -11, -6, -24, 10, -60, -17, 15, 13, 3, -5, 12, -19, 21, -1, 0, -28, 0, -30, -10, -17, 13, 21, -6, -18, -15, -33, -6, -9, -6, 3, 0, -25, 3, -37, -42, 19, -11, 7, -10, -71, 32, 53, -16, -18, 14, 4, 3, -38, 2, 55, 12, 14, -6, -23, 1, -11, 12, -12, -4, -53, -4, -29, -13, -48, -11, 2, 41, -108, 0, 16, -18, 35, -41, 45, -56, -15, -16, 58, 18, 2, -16, -35, 9, -14, 20, 54, 29, 0, 39, -59, -19, -7, 3, -9, 16, 6, -38, -25, -38, 16, -8, -33, 44, 9, -32, -15, -16, 3, 30, 4, 19, 39, 25, -51, 12, -31, -5, 18, -17, -48, -16, 3, 35, -40, -1, 0, -11, -14, -19, 15, -2, -7, 9, 2, -39, -20, 18, -13, 13, 21, -18, -19, -24, 17, 64, 27, 27, -4, -11, -54, -4, -5, 38, -39, -13, 2, -17, 14, -49, -19, 30, 23, -33, 17, 27, 32, 13, -62, -5, -17, -10, -33, 0, 10, -42, 5, 48, -42, 21, 49, -7, -24, -25, -21, -22, -5, -50, 26, 12, 28, 10, 23, -8, -30, -16, -68, 12, 10, -14, 27, 55, 8, -74, 13, 2, -26, 31, 14, -9, 5, 55, 7, 4, 34, 19, 43, -26, -7, -4, -11, -7, -1, -31, 0, 12, -57, 34, 17, -6, 8, 3, 14, -11, 4, 3, -8, 4, 0, 18, -8, -35, -51, 15, -34, -16, 40, 22, -28, 1, -20, 12, 2, 15, 16, -16, 22, -16, 23, -12, -1, 11, -1, 20, 0, -2, -30, 11, 39, -10, 31, 19, -45, -4, 22, -16, 8, -14, -6, -33, -12, 31, -59, -11, 7, -23, -14, -22, 2, -38, -5, -28, 17, -14, 28, 1, -65, 13, 31, 9, -17, -17, 14, -51, 33, 21, -17, -24, 12, 9, 7, -12, -18, -54, -24, -18, 18, 44, -30, -6, -3, -7, 15, 27, 48, 9, 28, 37, 31, 20, -2, 30, 28, -1, 43, -38, 16, 12, 9, 34, 14, 35, -31, 20, 1, -12, -3, 2, -1, 1, -17, 61, 4, 21, 14, -49, 22, -9, 25, -29, -2, -15, -10, 9, 29, 2, 36, 12, 18, -9, 14, -6, -28, 11, 34, -25, -8, -19, -14, 4, 35, -81, -7, 13, -69, -60, -21, 4, 42, -20, -7, 17, -4, -13, 4, -2, 43, 19, 14, -23, 4, -2, 21, -5, -19, -3, 14, 38, 12, 22, 23, -3, -5, -13, 0, 10, -23, 2, -22, -3, 18, 6, -13, 7, -49, -37, 11, -13, -12, 2, -9, 14, -43, -7, -2, -3, -32, -70, 32, 44, 25, -10, -10, 27, 41, -7, -21, -6, 12, 8, 33, -1, -38, -5, 28, 78, -57, 25, 15, -42, 0, -3, 3, 18, 28, 30, -9, -13, -10,
    -- layer=3 filter=0 channel=1
    -24, -4, -54, 7, -32, -48, -1, 1, 0, 15, -9, -12, -5, -36, -7, 5, 12, 54, 16, 25, -17, -2, 7, 8, -40, 21, 18, 8, -41, -30, 0, -50, 3, 46, 13, 15, 4, 39, 22, 13, -10, -10, -14, -18, 25, 43, -23, -24, 41, 44, 13, -22, 4, -6, -18, -39, -5, -16, -5, 29, -6, -9, -2, 5, 4, 20, 18, -24, 11, -17, 16, -4, -42, 11, 18, -18, 5, -15, 19, 13, 6, 9, -4, 30, 26, -11, -53, -19, -8, -17, 4, -6, 36, 22, 6, 1, -31, -12, -46, 11, -7, 43, 2, 13, 31, 8, -37, -10, -6, -10, -28, -2, -1, -31, -42, 17, 0, 21, -26, -18, 8, -17, -28, -15, -27, 18, -38, 16, 12, 16, -18, -28, -64, -55, 5, 18, -13, 0, 12, -39, -29, -18, -10, -8, 3, 0, 3, 19, 29, 7, 8, -51, 7, -25, 0, 8, -10, 4, -28, -19, 11, 19, -1, -24, 15, -8, 39, 12, 4, -27, 9, 17, 17, -10, -6, 20, 6, -3, -19, -20, -49, 5, 17, -20, -11, 19, 5, 3, -6, 13, -1, 12, 9, -38, -11, -7, -49, 0, 0, -2, 22, -6, 34, -27, -15, -17, 29, -23, 14, -18, 3, -17, 15, 20, -51, -2, -1, -7, -43, 29, 39, -17, 9, -36, -4, 19, 52, 8, -16, 25, 12, -35, -7, 27, 13, 5, -1, 5, 14, -28, -13, -74, -14, -20, 0, -56, -9, 7, 4, -26, -6, 23, -15, 14, 18, 3, 16, -38, 46, -3, -22, 34, 3, -2, 6, 6, 14, 8, 6, -18, -5, 3, 5, -45, -18, 6, -8, 7, 5, 13, 12, 1, -9, 4, -37, 39, 35, -34, 20, 42, 1, 15, -6, -11, 3, -30, -1, 0, 14, 2, 3, 12, -21, 27, -28, -20, 3, 0, -12, 9, -9, -2, -34, -33, 32, 17, -18, 12, 22, -30, -13, 13, 7, -4, -33, 11, 14, -14, 23, 9, 21, -46, 30, -77, -25, -45, -13, -6, -8, 34, 20, 36, 34, -22, -2, -10, 33, 9, 18, 29, -5, -41, -28, 14, 35, 0, 1, -5, 12, 19, 26, 6, -18, -21, 1, 24, -37, -9, 15, -14, -26, -12, 38, -15, 20, -19, 7, 13, -34, -3, -13, -28, -3, 14, 4, -39, -44, 28, -27, 2, 6, 11, -23, -73, -23, -16, -44, 9, 16, 23, 9, -3, 32, 27, -38, -22, -13, -38, -19, 61, 18, 5, -7, -5, -9, -43, -14, -66, -3, 93, -11, -6, -17, 32, 24, 8, -7, 21, 24, -41, 0, 0, 19, 0, 16, -12, -29, -14, -1, 23, 8, 5, -4, -46, -22, 8, -23, -10, 8, -50, 5, -7, 51, -43, 0, 1, -36, -11, 29, -28, 8, -24, 13, 3, -11, -52, -15, 37, -10, 9, 38, -31, -3, -2, 26, -10, 25, -19, -32, -4, -47, 26, -2, 30, -22, -5, 28, -20, -35, 19, -12, 34, -6, -30, -57, 12, 8, -54, -15, -5, -5, 9, -9, 16, 14, -42, -14, 26, 0, -5, 39, -19, 27, -28, -21, -42, -39, -13, -3, -5, -13, -83, 11, -1, 31, 44, -4, -4, 16, -17, 36, 9, -26, 0, -18, -62, 48, 0, 16, 23, 61, 28, 28, 16, 0, -48, 11, -9, -10, 3, 3, 0, -3, 8, 8, 31, 34, -29, 22, 6, -37, -46, 35, -15, -8, 8, -7, -9, 27, 31, 15, -80, -5, -8, -15, -2, 2, -58, 11, 1, 45, -48, -12, -9, -38, 15, 43, 59, 26, -57, 9, -71, -28, -64, -12, -25, 17, -21, -37, -20, -1, 8, 15, -30, 32, 43, -5, 43, 6, 28, -28, 26, 10, -75, 12, -26, 8, -51, 31, -12, 9, -5, 10, 6, -6, -1, -59, 12, -27, -10, 2, 40, -15, 17, 17, 32, 44, -31, 43, 0, -51, 47, 14, 0, 0, 36, 3, -12, -46, -80, 7, 39, -4, 7, -47, -51, 5, -19, -13, 24, -75, 8, 3, -37, -19, 7, -12, -20, 39, -70, 5, 15, -30, 8, -8, 76, 2, 21, 11, -61, 19, 56, 7, 31, 17, 40, 7, -27, -52, -19, -9, 9, -18, 27, -17, -18, 25, 18, 22, -42, -55, 3, -21, -54, 10, -32, 12, -4, 31, -52, -6, -1, -29, -11, 18, -3, 16, -112, 18, -9, -37, -34, 1, -28, -1, 61, -71, -7, 0, 17, -8, -11, 59, 42, 27, -12, 7, 11, -54, -19, -39, -59, 34, -8, 1, -24, 20, 10, -14, 24, -52, 20, 3, 27, -38, -31, -17, -19, 2, -17, -1, -5, -6, -5, -26, 27, -24, 0, 1, -51, -22, -14, -23, 59, -7, -8, -27, -13, -51, 8, -36, -18, -23, -13, -8, 12, 4, 46, -30, -27, -2, 1, -20, 70, -1, -25, -42, -38, -38, 9, -6, 13, 1, 13, 3, 13, -4, 30, -31, -8, -11, 31, -38, -19, -4, 2, -4, -14, -26, -12, -107, -77, -14, -6, -6, -3, 64, -25, -55, -49, -10, -80, -16, 44, 41, -18, 6, 6, 12, -18, 22, -17, -1, 35, -68, 11, -72, -65, -18, -16, -4, -30, 8, -44, -41, -3, -3, -15, -32, -23, 32, 24, 7, -41, -4, 6, -80, 18, -33, 25, 57, 19, 17, -2, -24, 16, -18, 30, 26, -31, 15, -11, -7, 15, -37, 7, 50, 34, -16, -16, -15, -18, 25, 3, -52, 7, 1, -9, 81, -16, 10, 23, 2, -6, -31, 34, -10, 26, -37, -5, 13, 33, 9, -49, 27, 17, 38, -21, -16, -48, 17, 10, 1, 4, 43, 0, 32, 26, -29, 8, 61, 24, -11, 11, -26, 18, 49, -25, 8, 8, 3, -29, -25, -31, -38, -14, -22, -5, -14, -11, -16, -53, -45, 3, 58, 38, 33, -33, -8, -2, -13, 37, -10, -5, 24, -38, 15, 8, 43, -4, 13, 36, 50, 34, -43, -20, -5, -35, -9, 24, -2, 3, -54, 10, 7, -7, -15, -54, 48, -11, 6, -60, -21, 0, -5, 65, 2, -76, 37, -17, -54, 1, 38, -11, 3, 22, -9, -1, 9, -52, 36, 25, -39, 36, 7, -4, 7, 55, 9, -1, 25, -21, -14, -6, -24, 0, 28, 0, 26, -9, -8, 15, -9, 9, -61, -9, -10, 12, 67, -16, -19, -33, -10, 25, 38, 21, -10, -32, -43, 22, -19, 10, 100, -8, 0, 12, -83, 31, 64, 5, 17, 61, -12, -47, 11, -37, -17, 55, 18, 6, -88, 17, -8, -25, -50, -12, -22, 12, -4, 18, -13, -15, 35, -17, 7, -24, -35, -10, -5, -30, -67, -1, 17, -58, 6, -2, -26, -15, 34, -10, 37, -3, 0, 62, -84, 21, 5, 0, 22, -17, -48, 11, -15, -16, -53, -57, -9, -16, 48, -5, 15, 29, -94, -31, -42, -34, 9, -17, 9, 7, -25, 15, 9, 0, 26, -38, -2, -32, -44, 68, -60, 18, 52, 20, -16, 19, 7, -22, -17, 19, -20, -15,
    -- layer=3 filter=0 channel=2
    19, 16, 75, -6, 19, -41, -11, 11, 10, 0, 19, -44, -7, 6, -2, -33, -4, -10, -8, -31, -34, 6, -4, -5, -27, -11, 4, -55, -5, 9, -31, -2, -20, 49, -17, -31, 10, -27, -25, -24, 12, 21, 5, -9, -22, -7, 0, -7, 19, 2, 12, 8, -7, -7, 0, 5, 0, 4, -5, -3, 15, 24, 13, -17, -2, -2, -1, 1, -1, 34, -4, -3, 3, 7, -37, -22, -11, 23, -1, 18, 35, 8, 13, -10, -46, 15, -20, -34, 0, -14, -7, 56, -4, -39, 11, -6, 28, 10, 33, -20, 16, -49, 34, 0, -18, 29, -46, -1, 3, 11, -4, -28, 5, -40, -2, 0, -2, -7, -33, 21, -6, 16, 34, -21, 2, -16, -23, 21, 36, 58, 34, 38, -7, 1, 9, -1, 10, 38, -21, 32, -22, -38, 20, -28, -8, 17, -27, 7, 25, -14, -6, -21, 9, -23, -10, 6, -42, 28, -5, 1, -40, 13, -38, -16, -17, -33, 25, 5, -1, -25, 13, 29, 23, 8, -6, -12, 27, -47, -23, -8, -6, -8, 16, 0, -34, -34, -5, -8, 9, -28, 4, 18, -1, 31, 7, -3, -43, -7, -13, 5, 6, 9, -55, -29, 12, -17, -9, 24, -5, -8, 7, -46, -28, 30, 6, -5, -8, -13, -6, -32, -16, -8, -40, 13, 40, 44, 3, -8, 7, 5, 12, 22, -8, -11, 1, 30, -9, -23, -8, -21, -7, -17, -12, -22, 1, -8, -18, -29, 1, -38, 15, -7, 5, -14, -17, -28, 6, -22, -21, -3, -42, 4, 3, -15, 12, 12, 9, 11, 0, -9, 27, 12, -15, 12, -16, -34, 0, 11, 5, -12, 31, -64, -8, 37, -12, -16, -33, -37, -10, 12, 1, 3, -19, 13, 16, -13, -7, 18, -6, -29, 10, -26, 2, -12, -1, -15, 21, -21, -27, -9, 18, -6, 0, 3, -5, -25, 2, -33, 5, 16, 0, -6, 27, -20, 10, 26, 10, 4, 22, -10, 6, 10, -14, 13, 27, 10, -11, 7, 3, -77, -12, -36, 19, -8, 8, 4, -23, 21, 19, -20, -9, -11, 4, 6, 18, -4, 40, 19, 11, 10, -1, 28, -7, -28, 7, 12, -17, -6, -6, -10, -27, -45, 25, -10, -6, 34, -6, -33, 6, -12, 0, 46, 9, -6, -36, 1, -13, 0, -6, 33, -10, -9, -2, 4, 10, 28, 12, 34, 1, 9, 4, -21, 12, 3, 22, -12, 8, 24, 16, -64, 3, -22, 8, -56, -19, 2, -5, -25, -34, 31, -2, -37, 19, 33, 11, 8, 10, 2, -32, -13, 7, 13, 42, 6, -19, -9, 16, 24, 8, 13, 25, 2, -24, 13, 43, 21, 45, -25, -3, 12, 14, 2, 16, -7, 1, 16, 12, -9, 8, 17, -8, -17, -16, 18, 40, 0, 7, -42, 3, 3, 7, -12, 17, 9, 8, 16, 62, -9, 17, -17, -8, -24, 21, -27, -9, -3, 1, 0, 56, -4, -1, -48, 8, -40, -9, -32, -14, 6, -29, -34, 42, -20, -33, 32, 17, 39, -5, 0, -5, -25, 11, 0, 40, 40, -32, 7, -19, 10, 10, -7, -10, 32, -55, 20, -20, -38, 14, -6, 0, 7, 31, -24, -7, -12, -14, 1, 33, -25, -25, -2, -1, -11, -31, 15, -14, -39, -42, -55, 0, 17, 26, 28, 35, 24, -3, -17, 24, -44, -48, -10, 29, 40, 23, 10, -15, -19, 1, -13, -11, 3, -5, -1, -16, -2, -17, 82, 2, 8, -3, -9, -47, 35, 11, 18, -1, -14, -9, 15, 21, -28, 9, 8, -5, -24, -7, -17, 25, 8, -14, 9, -12, 7, -28, 0, 19, 28, -15, -14, -19, -47, 27, -15, -15, -51, 3, 25, 5, 6, -30, -21, -3, -3, -44, -47, -4, 8, 44, 24, -25, -19, 3, -3, 24, -1, -92, 12, 22, 24, 7, 7, 28, 54, -10, 25, -2, 55, -15, 0, 13, 22, 9, -30, 26, -27, 19, -12, 11, 0, 38, 3, 5, 6, 13, -1, 19, -83, 5, 17, -2, -4, -36, 27, -24, 6, -8, -44, -9, 19, -1, 54, -22, -47, -1, -20, 14, 0, 6, 31, 32, 23, 28, -13, -9, 9, -7, -3, -25, -11, -3, 8, -5, 9, -13, 10, 0, 18, -23, -20, 24, 48, 11, -12, 33, 3, 6, -9, -31, 9, 6, 42, -9, 50, 6, -28, 6, -64, 4, 17, 17, 18, 1, -13, -34, 11, -2, -45, -19, 66, 26, 48, 10, 2, -23, 14, -10, -20, 28, -43, 0, 28, 49, -31, 7, 6, -41, -1, 7, -24, -37, -5, -10, 20, 3, -14, -19, 13, 39, -15, 55, 15, 20, -19, 15, -76, 4, 4, 3, -36, 50, -5, 9, 2, 34, 2, -27, -22, 4, -23, 21, -21, 9, -13, 41, -57, -10, -1, 50, -30, 39, 28, 30, -39, 2, -22, 3, -20, 42, -17, -34, -2, -12, 3, -17, 11, 14, -7, 20, -10, 30, -6, 42, 25, 14, 1, 37, 16, 3, -3, 43, -10, -17, 23, -1, 4, -3, 6, 21, 31, 12, 11, -38, 10, 4, 38, -29, -22, 16, -11, 4, 23, -5, 26, -51, -10, 61, -14, -13, 5, -19, 9, -28, -17, -36, 14, 59, -5, 28, -12, 17, -8, -1, 1, 20, 34, -18, -43, 11, -21, -18, -27, 8, 30, 18, -24, 43, -27, -34, 11, 5, 27, 29, 30, -13, -62, 35, -1, -9, 53, -11, 28, 30, 1, 2, -13, 4, -30, 9, -31, -4, 11, 7, -29, -1, 4, 46, -19, -17, 0, 5, 21, 18, 47, -6, 32, 20, -11, -6, 3, 14, -18, -40, 10, 7, -34, -34, 24, -5, 28, -19, -4, -4, -24, -18, 1, 37, 23, -41, 13, 50, -12, 7, -5, 14, 15, -21, -33, -96, -9, -68, 38, -15, -10, 23, -4, -31, 34, 9, -13, -26, -6, -15, -7, -23, 0, -6, -23, 8, 70, -12, 9, -27, 6, 5, -14, 5, 11, 23, -3, -42, 5, -68, 33, 15, -42, -28, 29, 17, -19, -29, 7, 35, 5, 3, -41, 5, -26, -7, -21, -13, 28, 45, -17, 7, -12, -17, -13, -2, -15, 8, -18, 36, -32, -8, -31, -3, 80, 16, 7, -5, -17, -17, 11, 3, -18, 29, 0, 50, 18, 19, -51, -6, 25, 40, -18, -35, -6, -1, 34, 34, -19, -8, -3, -31, -51, 3, -24, -29, 18, -45, -15, 7, -14, -19, 63, 51, 32, 11, 0, -18, 12, 19, 12, 20, -2, -7, 18, 48, -3, -7, -8, -26, 14, -39, 19, -11, 7, 12, 8, -5, 6, 11, 16, 24, 5, 2, 16, -31, 15, 11, -15, -79, -8, -20, -25, 47, 52, -4, -24, -30, 3, -2, -18, -10, 1, 2, 16, -32, 31, 2, -25, 5, 4, 24, 23, 23, 28, -40, -21, 31, 28, -8, -27, -13, 14, 0, -12, 5, 28, -1, -54, -10, -3, -26, 33, 6, -8, -17, -1, 46, -69, -17, -19,
    -- layer=3 filter=0 channel=3
    -1, 6, -33, -5, 21, -5, -4, 0, 7, 22, 0, 33, -41, -17, 24, 20, -14, 42, 5, 12, -15, -1, -11, -14, -22, -33, -2, 38, -18, -10, -41, 15, 13, -32, 21, -10, -12, -14, -23, 32, -25, 0, 5, -6, 7, 0, 1, -17, -5, -3, -43, -2, 20, -26, 15, 14, -16, -28, -14, 0, 14, -27, -5, 36, 0, 5, 22, 15, 3, 30, -10, 7, 29, 8, 16, 1, -1, 35, -23, -23, -42, -47, -6, 20, 33, -46, 14, 7, 17, 6, -1, 3, -58, 16, -18, 1, 18, -30, -28, -19, -32, 26, -8, -38, -1, -15, 15, -12, -14, 20, 19, 20, 5, 0, 56, -27, -23, 23, 22, -53, 9, -16, -13, -21, 24, -8, -8, -5, 29, 35, -3, -11, 23, -9, -12, -8, 16, 51, -11, 2, 14, -16, 1, -12, 5, -5, -15, 21, -21, -4, -5, 24, -22, -7, 2, -39, -14, 39, 29, -28, 19, -10, 19, 49, -27, -13, -10, -24, -22, -5, 8, 0, 30, 17, -8, 10, 14, 19, -33, -15, -4, -28, 17, -5, 47, 3, -3, 4, 0, -10, 8, 27, 0, 15, -16, 1, 5, -19, -8, -2, 22, 19, 0, 17, 0, -14, -9, -18, 29, -30, -12, 21, 26, -13, 0, -6, 2, 2, 4, 13, -37, 24, -18, 9, -6, -29, -43, -2, -12, 9, -11, 27, -1, 19, 8, 0, -10, -19, -24, -15, 2, -23, 83, 17, -4, 26, 24, 12, 0, -28, 6, 5, -5, 33, 23, -9, -8, 53, -15, -11, 8, 43, 9, 9, 20, 50, -34, -13, 4, -17, 2, -11, -23, -29, 0, 21, 5, -15, 2, 5, -27, 34, 16, 4, 15, -22, -1, -36, -8, 11, -12, -8, 19, -11, -50, 14, 20, 10, -5, 16, 8, -30, -2, -27, 18, 26, -66, -1, -16, 26, -9, -23, -3, -2, -12, 35, 5, -16, 29, -12, -17, -17, -12, 4, 0, -11, -2, -14, 0, -15, -24, 10, -24, 0, 7, -22, 32, 0, 12, 75, 9, -8, -36, -35, 8, 5, 28, 2, -14, 37, -23, 0, 27, 15, -7, 39, -26, -11, 24, -36, -19, -36, -23, -38, 14, -11, 23, -31, -8, -35, 22, -3, -1, 15, -2, -6, 6, -2, -34, -19, -12, -25, -22, -4, -5, 28, -10, 30, 3, 6, 0, -10, 22, -7, -19, -7, 12, 0, -9, -30, 17, 19, 0, 3, 3, -5, 11, -15, -18, -17, -10, 48, -13, 10, -40, -27, -3, 4, 9, 8, -8, -17, -24, 16, -34, -20, -5, -18, -13, 4, 17, 0, 6, -3, 9, -3, 7, -8, 15, 17, -13, 0, -54, -3, -11, -16, -7, 9, -11, 2, -31, -16, 1, -3, -6, -3, -20, 5, -57, 6, -26, -39, -9, 1, -6, 51, -8, -17, -7, -44, -11, 4, 17, 3, -32, -9, -19, 26, 17, -15, -5, 29, -7, -16, 25, 12, -45, 9, -9, -18, 28, -25, 6, -39, 13, 3, 9, -17, -12, 30, 25, -2, 6, -43, -22, -13, -6, -22, -3, -3, 5, 16, 10, 15, 44, 31, 8, -45, -11, 1, 11, -28, -7, -4, -3, 22, -2, 0, -8, 28, 8, -37, -13, -17, 6, 34, -43, -8, 14, -50, -44, 8, -10, -10, 10, 53, -40, -17, -16, -62, 11, -9, 16, -7, -5, -31, -56, 16, -11, 7, -36, -7, 32, -10, 2, -5, -17, 0, 5, 6, 0, 33, -2, 11, -27, 11, -5, 0, -25, 9, -44, 8, -15, 14, -21, 7, -29, -21, -19, 23, 6, -17, -26, 7, 15, -3, -36, 53, 42, -4, -16, -12, 9, -6, -27, -18, 14, -6, 10, -10, -48, -48, 32, 31, 1, 33, 33, 62, 22, 55, 4, -34, -13, 58, -17, -70, -51, -12, 25, -13, 5, -12, -3, 13, -8, -15, 5, -15, 5, -9, 22, 7, 0, -9, 0, -2, -11, -15, 22, 45, -6, 9, -23, -9, 3, 12, 1, 6, -45, -20, 16, 2, -13, 18, -21, -9, 14, -1, 0, -10, -70, -69, 18, 6, -10, -6, 2, -53, 6, 15, -16, 2, -2, -15, 4, -5, 11, 35, -14, 19, -22, 13, -9, 18, 0, 9, 24, 0, 12, 27, 10, 35, -1, -10, -12, -16, -32, -8, 2, 38, -13, 9, 15, 4, -10, 5, -23, -8, -17, 9, 3, 10, -4, 30, 16, 4, 5, 9, 6, -5, 0, 35, -19, -17, -22, -4, 25, -28, 18, -27, -2, -5, 29, 38, 0, -8, 19, 27, -2, 7, 10, 0, 11, -38, 29, 12, 56, -10, -25, -4, 5, -38, -28, 19, 16, -30, 6, -4, -5, 13, 4, 43, -8, 19, -4, 5, -21, 1, -8, 21, -1, -8, 13, 1, 3, -6, -21, 0, 22, -5, -3, -42, 19, -17, -9, -1, -2, -4, -14, 14, -15, -49, -22, -30, -10, 3, -22, 29, 33, -22, 15, -13, -19, -39, -15, 38, -3, -3, -11, 8, 0, 21, -11, 20, -11, -17, -28, 13, 9, 10, -13, 11, 2, 29, -12, 10, -27, 14, 3, 3, 32, -7, -2, -15, 18, -31, 17, -16, 9, -25, 10, 1, -36, -13, -22, 4, 12, 8, 8, 10, -15, 21, 4, 12, -42, 35, 34, 12, 3, -9, -36, -22, 38, 14, -3, -8, 8, -49, 18, 13, -9, 16, 13, -33, -30, 0, 13, 42, -10, 18, -18, -38, -25, -10, -20, 0, 27, -14, 11, 19, -21, -17, -12, 16, -31, 13, 20, 20, 21, -29, -18, -15, 3, 13, 11, -57, 41, -18, -16, -20, -14, 32, -9, 7, -18, 30, 4, -39, 16, 12, -54, -6, -1, -11, -14, 11, -25, 10, -6, -64, -5, -14, 4, -7, -21, 22, 16, 12, -17, 25, -12, 29, 1, 0, -62, 11, 18, 11, 10, -23, -21, -23, 20, -6, -22, -27, -2, -18, -6, -17, -8, -1, -52, 4, 27, 5, 0, -32, 0, 2, 11, 10, -19, 21, -4, -13, -23, 13, 20, 7, 30, 6, 25, -6, 10, 9, 31, 19, -14, 6, -17, 39, 13, -6, 6, -30, -48, -1, -7, 0, -25, -24, 13, -25, 38, -6, 8, 24, -14, -20, -14, -18, 47, -13, -19, 11, -3, -19, -27, 19, -5, -8, -7, -2, -11, -19, -18, -4, 21, -19, -23, 19, 16, -20, 8, 15, -13, -30, -24, 0, 9, 0, -6, 13, 6, -27, 14, -28, 0, 3, 10, -32, -31, -17, 1, -21, 13, -9, -15, -17, 17, -4, 44, -3, 23, 13, -5, -6, -13, 0, -19, -25, -39, -5, -18, 20, 0, 34, 0, 12, 29, 11, -46, 38, 12, -15, -25, -13, 20, 20, -9, 4, -12, -24, 25, 3, -8, 39, 22, -25, -9, -3, 2, -3, 1, 9, -10, 5, -3, -3, 32, -22, 3, 17, -36, -19, 20, 18, 9, -38, 6, 20, 9, -14, -8, -10, 7, -32, -33, -26, 52, -16, -25, -22, 17, 38, 2, -11, -29, -30, 22, -4,
    -- layer=3 filter=0 channel=4
    -43, -37, 28, 13, -42, 33, -17, 7, 4, 6, -29, 21, -16, 12, 7, -19, -16, 32, 23, -15, 43, 5, -7, 15, -32, 24, -13, 23, 25, 25, -10, 6, 6, 16, -24, 14, -2, 15, 41, -23, -85, 1, 10, 15, -34, -37, 6, -1, -56, -2, -9, 9, -24, 8, -4, -14, 15, 5, 2, 6, 30, -11, -26, -57, 13, -11, 31, -9, 15, -49, 16, 15, 24, 17, -19, 19, 25, -13, -1, -9, -14, -21, 8, -13, -15, -10, -65, -6, 2, -9, 6, 17, 12, -67, 14, -33, -19, 12, 17, -5, 13, 41, -40, 6, 12, 15, -11, 2, -7, -11, 2, 27, -21, 9, -26, -12, -29, 13, 36, 43, -1, -15, -32, 0, 35, -62, -32, -10, -5, -11, 12, -23, -43, -18, -6, -8, 16, -3, -11, -21, 23, 60, 8, -5, 7, -41, -11, 0, 18, 14, -7, 47, -72, -18, -22, -36, 52, 27, 7, -14, -9, 34, 25, 25, -14, -42, -2, -28, -31, 14, 9, -27, -38, 31, 7, 0, -15, 58, -21, -2, 11, -42, 13, 23, -8, 18, -25, -19, 44, -1, 7, -15, -22, -22, 40, 0, 53, -7, -8, -16, 15, -8, 30, 22, 9, 10, -10, 30, -25, 39, -9, 15, -33, -23, -82, -18, -8, 4, -17, -27, -24, -33, 58, -26, 0, -12, -63, -4, 25, 12, -36, -24, -8, 12, -15, -27, 15, -14, -10, 33, -1, -28, -44, -7, -7, 20, 24, -10, 2, -12, 38, 2, -37, -101, -22, -14, 5, -22, 39, -37, 38, -46, -11, -15, 7, -19, 13, -31, 28, 29, 24, 31, -9, -21, 6, -2, -14, -12, 13, -18, -34, -57, 3, -38, 17, 23, 14, 12, 15, 34, -2, -4, -11, 8, 24, -64, 3, -4, -9, 0, -20, 43, 29, -9, 0, -1, -22, -9, 20, -32, 5, 5, 23, 10, -17, 14, 48, 30, -36, -42, 8, 11, -8, 9, 24, -27, -2, 0, -17, -13, 32, -9, -24, -26, -36, -38, 9, -6, 7, -50, -2, -16, -24, -12, -6, -20, 2, 24, -37, -61, 65, 5, 40, 5, -69, -12, 20, -6, -96, -6, 8, -26, -19, -17, 5, -77, 11, 42, 14, -32, -15, 34, -12, 18, 23, 15, -6, 29, 14, -56, -41, -17, 26, 5, -3, -55, 6, -24, -8, -10, 3, 0, -6, 5, -16, -10, -6, 33, -9, 19, -20, -12, 6, -24, -22, 8, 15, 21, 4, -28, -12, -16, 18, 38, 13, 9, 8, 24, -48, 8, -19, 19, -8, -40, 18, -16, 9, -47, 24, 0, 4, 0, -45, -17, 22, -24, 2, 2, -13, 42, 7, 24, 15, 10, -13, 14, -11, -105, -20, 19, -4, -7, 4, 17, 16, 4, 28, -8, -23, 14, 19, -30, 24, 19, -23, -28, 9, 0, 11, -21, -39, -16, 15, 0, 4, -20, -28, 17, -4, 21, -17, 16, 25, -1, -6, -24, -2, -12, 8, 8, -45, 46, -8, -11, -19, 20, 5, 48, 56, -30, 33, -24, 31, -16, 6, 58, 42, 29, -14, -14, -32, 4, -12, 4, -119, -41, 0, 37, -8, 9, -3, -33, -47, -31, 0, 16, -3, 2, -15, 13, -22, -35, -10, -27, -1, 2, -25, 8, -45, -51, -2, 55, 35, -58, 0, 6, -9, 21, -10, 33, -50, -34, 26, -23, 11, -40, 15, -8, -23, -5, 9, -56, -32, -25, 51, -43, -14, -37, -10, -3, -20, 0, -58, 7, 21, 46, 0, 16, 20, -2, -22, 21, -15, -5, 2, 5, -29, -27, 52, 1, -35, 44, 14, -39, -5, -9, -15, -46, -5, -24, 12, -6, 25, -33, -55, -2, -34, 14, 5, -33, -23, -7, 18, 6, 1, 11, -17, -1, 1, 38, -5, 0, 2, -59, 0, 34, 54, 45, 13, -12, -7, -26, 12, 0, 15, 11, -7, -6, -46, 9, 3, 0, -61, 11, 19, 10, -12, -14, -5, -23, 10, 4, 1, 21, 4, -6, 11, 47, 4, -7, -8, -18, -7, -8, -45, 14, -3, 18, -11, -13, 54, -21, -3, 10, -5, 12, -5, 26, -24, -8, -30, -35, 10, -35, 3, 30, -18, -45, -31, -39, 5, -20, 39, -22, 8, -7, -23, -2, 3, 16, 16, -15, 9, 22, -12, -10, -30, -3, -2, -7, 10, 10, -2, -7, -29, -1, 31, 45, 2, 23, 11, 8, -17, -13, 0, -26, -13, -6, 9, -4, -14, 4, -9, -67, -61, 33, 30, -10, -6, 29, 0, 18, -49, 5, 13, 14, -31, 27, 5, -10, -45, -9, -9, 0, 25, 19, -12, 0, 20, 9, -20, 22, 9, -7, 15, -10, 22, -10, 19, 1, -67, -8, 29, -46, -20, 12, 9, 35, 34, 4, -4, -19, 38, 14, -1, -14, 25, 24, 22, -21, -5, 26, -71, -17, -3, -27, -7, -30, -3, -35, 14, 42, -5, 59, 8, 11, -33, -12, 8, 7, 7, -68, 54, 25, 4, -86, -4, 48, -79, 8, 20, 19, -15, -10, 12, 0, -2, -15, -8, 41, 21, -15, -5, -5, -58, -11, 9, 17, -8, -1, -24, -3, -49, 27, 33, -26, 51, 25, 3, 8, -5, 3, -9, 7, 1, -28, -4, -12, 22, 0, -44, -23, 11, 37, 3, 31, -7, 23, 0, -33, 2, 27, -18, 6, -23, 45, -5, 17, 29, 69, -3, 26, -12, -23, -5, -18, 20, -9, -2, 39, 5, -3, -58, -22, -1, -1, -51, 33, -25, 15, 7, -8, -3, 9, 5, 37, 11, 0, 25, -87, 61, 25, -5, -7, -36, 3, 9, -10, 0, -2, -77, -59, -29, -72, -24, -7, 29, -88, 14, -1, -75, 35, -23, 5, -27, 9, 29, 11, -7, -52, 46, -5, 3, -43, 25, 52, 26, 5, 22, -3, -17, -21, 31, -25, 2, -4, -37, 14, 10, -16, 10, 5, -45, -20, -3, 21, -4, -14, 7, 5, -54, 19, 21, 20, -35, 33, 5, 32, -4, -3, 17, 31, -16, -28, -1, 17, 31, 12, -24, 14, -23, 43, -24, -44, -19, -38, 10, 19, 17, -5, 10, 8, -43, -91, 0, 21, -6, -9, -3, 8, 35, -70, -56, 0, 4, -31, -11, -13, 8, -68, -16, 18, 21, -23, -14, 5, -44, 3, 25, 43, 16, 0, 50, 0, 45, 16, 22, -31, 34, -10, -15, -5, -27, 1, 28, -24, -6, 43, 0, -17, -7, 25, 18, -22, 7, -86, -19, -27, -56, 26, 2, 3, -6, 10, 31, 22, 10, -41, -4, 20, 9, -7, -14, 17, -10, 3, 41, 0, 7, 9, 3, 19, -23, -16, -17, -9, 13, -23, -24, -41, -24, 8, 15, 21, 2, 3, 10, 4, -33, 26, 34, 29, -32, -34, -7, -32, -17, -10, -18, 25, -15, -7, -19, -9, 18, 36, 1, -18, -23, 2, -6, -25, 6, -7, 8, -21, -19, -3, -17, -6, 29, 35, 0, 5, 25, 46, 0, -8, 23, -67, -10, 23, 3, 4, 9, 0, -4, 11, 10, 30, -33, -20,
    -- layer=3 filter=0 channel=5
    10, -1, -3, -12, 43, 41, 14, -16, 9, -8, 14, -31, 37, 10, -14, 7, -2, -11, -65, -25, -51, -10, -10, -10, -53, -30, -20, -58, 17, -85, 16, 25, -14, -37, 5, 40, 4, -27, -50, -2, 41, 49, -8, 3, 21, -10, -8, -9, -27, -33, 57, 16, -37, 6, -6, -21, -15, 3, 33, 4, -1, -39, 6, 50, 4, -10, -27, -8, -10, 16, -16, 15, -8, 0, -35, -15, -9, -10, -20, 39, 36, 2, 12, 18, 32, -13, 24, -2, -12, -12, -26, -11, -28, 32, -35, 0, 20, -6, 32, -9, 12, -15, 36, -23, -29, 31, -3, -26, 9, 4, 31, -52, 12, -25, 30, -1, -21, 16, 32, -74, 0, 11, -25, -54, -12, 19, 67, 10, -23, 1, -33, -10, 24, 65, -7, 4, 30, -54, 24, 46, -5, -8, -23, 4, -17, 18, 48, -2, 10, 0, -15, -9, -16, -4, -4, -34, -46, -25, 20, -42, 14, -33, 12, -20, 20, 39, -31, -7, 24, -11, 11, 7, 59, -30, -16, 22, -4, -28, 13, 15, -15, -3, 13, -60, 40, -18, 62, 11, -59, 34, -14, 40, -4, 7, -29, -7, -4, 44, -16, -7, -11, 8, -32, 34, -13, 2, 21, 68, 12, -36, -14, -15, 8, -28, 34, 0, 2, -6, 10, 7, 46, -1, -41, 8, 19, -44, 28, 26, 9, 21, 30, -29, -49, 31, -2, -27, -9, -9, 23, -48, -5, 13, 34, -22, 31, 20, -18, 0, -7, 29, 5, 22, 0, 10, 32, -9, -14, 14, -9, -11, -6, -2, 6, 6, -21, -83, -38, 30, -45, -1, -14, -2, -8, 46, -16, -29, 12, -13, -2, 34, -3, 11, -16, -2, -21, -30, 43, 0, 44, 5, -5, -15, -15, 21, -49, 45, -5, -21, -7, 6, 20, 7, 29, 2, 6, 26, -89, 4, 6, -29, -12, 7, 50, 0, 17, 17, -37, 14, -15, 13, 0, 19, 17, -10, 4, 32, -16, 9, 55, 10, 30, -18, 9, -5, 32, 74, -20, -8, -2, 9, 14, -48, -12, 5, 12, -21, 0, 13, -18, 56, -24, 28, -9, -21, -17, 43, 17, -15, 36, -6, -1, 5, -10, 5, 5, 12, -10, -15, -17, 32, 62, -20, 1, -30, -19, -9, -13, 0, -59, 10, 22, 39, 0, -17, 37, -18, -26, 20, -13, -21, -13, -11, 23, 18, 5, -18, 9, 38, 27, 22, 10, -14, -73, 0, -5, 17, 0, -14, -35, -43, -12, -22, -23, -123, -19, -10, -8, -8, 14, -1, -14, -3, -32, -36, 2, 9, -6, 15, 27, 9, -10, 27, 7, 0, 5, -5, -19, -7, 2, 17, 8, 14, -20, -5, 7, 17, -18, 4, -10, 10, -35, 2, -13, -8, -8, 7, 6, -14, 4, -11, 32, 7, -4, 11, 3, 29, 0, 26, 17, -54, 56, 4, -15, -1, -6, -24, -3, 1, -3, 18, 19, 8, -62, 0, -17, 9, 32, -15, 6, -8, -5, 12, 3, -28, 0, -6, 1, 35, 40, -32, -23, 15, 11, -40, -3, -11, -3, -36, -15, -13, 3, -7, 8, -33, 57, -27, -2, 7, -13, -16, 15, 6, -62, -9, -20, 21, -28, 30, 0, 16, -23, -28, 8, 10, 0, 10, -4, -5, 0, -21, 1, -2, 27, -39, 11, 14, 18, 12, -19, -24, -40, 16, -19, -12, 9, 6, -19, 6, -12, 23, 0, -1, -8, -12, -14, -1, 11, 23, -32, -6, 12, 27, 17, -55, -17, -7, 6, -27, -26, -8, -71, -5, -12, -9, -14, 3, -38, 14, -18, -21, -73, -7, -5, -11, -17, 41, 41, -50, -12, -25, 11, 9, -23, -2, 15, 1, 33, -13, 20, -23, 3, -33, 8, 56, 33, -17, 14, -4, -7, -20, -18, 3, 22, 17, -17, -21, -9, -52, 10, 13, 12, -60, -3, -2, 4, 0, -12, 5, -6, -18, -17, 16, 5, -4, 16, -8, 4, -7, -33, 17, -63, 26, -10, -3, 0, -7, 5, -25, -39, 6, -1, -9, -11, -6, 10, 27, 0, -27, 11, -109, 29, -67, 13, 27, 7, 22, 0, -31, -86, 16, -56, -23, -17, -25, -10, -28, 25, 4, 21, 16, 3, 0, -16, 25, 2, 0, -2, -27, -30, 35, 8, 11, 46, 19, -15, 6, 18, -8, 7, -15, -12, -1, 1, -11, -32, 16, 1, 49, 0, -27, -12, -15, 17, 38, 7, -15, -37, -12, 0, 0, 29, 31, -37, 16, -33, 17, -26, -39, -26, -12, 1, -16, 10, 35, 2, 31, -10, 46, 12, -6, 5, -8, -11, -8, -27, -18, -20, -17, 19, -7, 0, 21, 25, -3, 17, -25, -20, -18, -21, -2, 1, 40, -5, 21, 0, -5, 7, 20, -14, -17, 2, 22, -12, -21, -9, -16, -33, -53, -7, -14, 6, -25, -18, -9, 8, 36, -8, -61, -41, -50, -18, -12, -60, 4, 3, -38, -46, -27, 0, 18, 0, -34, -4, 14, -17, 22, 0, -29, 4, -8, 11, 53, -19, 10, 6, -26, -99, 11, 10, 3, 51, 17, 8, 10, -22, -5, 5, -8, -14, 12, 29, 16, -13, -11, 5, -41, 8, 4, -3, 38, -17, -19, -10, -20, 0, -9, 9, 13, 7, -35, 18, 4, -1, -27, -13, 37, 1, -19, -13, -31, 19, 22, 5, -47, 26, 8, 3, 10, 9, 16, -10, -8, 32, 17, -28, 1, 15, -36, 6, 1, 5, 26, 12, -3, 17, -11, -2, -39, -22, -25, -7, 11, 4, 0, 27, 12, -10, 0, 13, -1, -24, -15, -11, 19, 2, -35, 36, -9, 7, -14, 13, -10, -7, 20, 0, -17, 4, -59, 10, -52, 14, 19, -14, 24, -43, 10, 28, 16, 0, -31, 4, -22, -7, -19, 14, 12, -14, -5, -36, -11, 0, -7, -17, -10, -30, -4, -13, 3, 28, -20, -26, 3, -50, -17, -18, 33, -4, 2, 2, 1, -13, -37, 14, -20, -17, -4, 16, -21, 17, 23, 9, -49, -28, -29, -20, -8, 1, 25, -7, -7, -9, 23, -4, 38, 19, -59, -7, 23, -11, 0, -1, -38, 47, -8, -19, -41, 9, 36, -13, 12, -36, -11, 15, -16, 12, -27, -14, -32, 0, 23, 2, -10, -28, 8, -12, 13, -51, 18, -34, 7, -2, 11, -8, 53, -3, 23, 0, -10, -48, -14, -4, 11, 2, -44, 13, 4, -8, -38, 6, -2, -8, -45, -36, -30, -60, -16, 30, -31, -34, -2, -11, -40, -45, 20, -27, -31, -11, -63, 23, 1, 12, 36, 20, 0, -7, 8, -24, 15, 12, 31, 13, -4, -24, 5, -25, 0, 48, 13, 2, 18, 2, 3, -9, 21, 6, 12, -3, 3, -19, 9, -18, -3, 17, -10, 19, -42, 0, 18, -34, -37, -40, -11, 3, 17, 5, -7, -40, 4, -57, 0, -15, 0, -22, -30, 12, -17, -26, 2, 7, -26, 21, 21, -9, -3, -10, 4, 7, 9, 17, -17, 24, -44, -12, 18, 3, 6, 0, -16, -8, -11, -11, -7,
    -- layer=3 filter=0 channel=6
    -35, 36, 26, -6, -29, -49, 7, 13, -11, -11, -46, -14, 52, -8, -10, -8, -1, -17, 14, 9, -6, -5, 5, 29, -37, 26, -34, -1, -24, -18, -19, 24, -20, -5, 10, -63, -7, -2, -72, -8, 6, 4, -18, 6, 8, 49, -31, -21, 14, -15, 29, 0, 16, -23, 16, 3, 2, 26, -10, 37, -77, 24, -12, 5, 3, -25, 21, -18, -8, -39, 3, 5, 1, -19, 0, -16, -106, 15, -5, -17, 3, 40, -13, 18, -32, 66, -13, -54, 6, 3, 12, -8, -80, 9, -23, 12, -3, 4, -52, 11, 33, -2, 12, -9, -6, 9, -8, -43, 1, -23, -52, -24, -20, -63, -30, 3, 27, -32, -37, -1, 0, -27, -12, 18, -41, 11, 2, 13, -6, -4, -56, 1, 10, -52, -1, -7, 26, -30, 7, -21, 28, -6, 33, -15, 4, 19, -2, 14, 4, 3, 12, 25, -10, 31, -15, 8, -11, -96, 2, 27, 5, 47, -24, -6, -10, 43, -39, -32, -8, -1, 12, -50, 28, -27, 5, -87, 13, -9, 13, -9, 5, -35, 17, -6, 1, 12, 2, 1, 40, 10, 3, -42, -19, -56, 17, 9, 5, 23, 8, -14, -35, 8, -16, -30, -18, -28, 28, -36, -20, -25, -2, 26, -47, 23, -22, -13, -15, -17, 47, 23, 0, 11, -42, -14, 0, -18, -63, -8, 18, -40, -55, 4, -7, 16, -45, -11, -16, 24, -13, 26, -16, 44, 13, 15, -10, 41, 37, -34, -10, -59, -39, 21, -49, -33, -44, 0, 46, -14, -3, -25, -26, -7, 6, 14, 20, -14, 3, 16, -50, -28, 13, -60, 1, 7, -45, 14, -2, -29, 5, 19, -29, -5, 0, -30, -19, -74, -16, -7, 30, -8, -9, 26, -12, -10, -34, 0, -54, -31, 1, -3, -4, -33, 25, -19, 16, 19, -15, -12, -11, -46, 9, -23, -54, 15, 6, 5, -45, 12, 26, -24, 2, -11, 49, 6, 17, -8, -2, 15, -2, 6, -32, 6, -36, -3, 11, 12, -4, -33, -1, 21, -47, -31, 7, 5, 4, -4, 21, -10, 8, -84, -51, -39, 5, 46, -25, -31, 10, -14, 22, 19, 26, -8, -51, -56, -13, 30, -55, 6, 3, 57, -50, 7, -7, 72, -18, -44, 8, -37, -38, 7, -17, 4, 19, -7, -67, 97, -11, -13, -2, -31, 0, -1, 7, 0, -7, -21, 18, -11, 19, -11, -7, -7, -36, -55, 0, -10, 3, 0, -46, 27, -20, 24, 23, 29, -51, -22, 12, 2, 19, -69, 11, -5, -37, 25, 31, 49, 16, -8, -31, 8, 36, -2, -20, 34, 32, -3, -9, -39, 6, -23, -19, -42, -32, -19, -53, 2, -1, 11, 7, -20, 14, -11, -31, 39, -2, -13, 7, 9, 22, 29, -64, 68, 19, 16, -26, -18, 2, -17, -35, 40, -27, 5, -18, 1, -18, -6, -91, 56, 8, -32, -3, 19, -24, 15, 22, 61, 24, 12, 6, 0, 27, 34, 7, 12, -65, -5, 2, -72, -1, -25, -25, -18, -47, 31, -13, -80, 1, -20, 0, 33, 4, 11, -9, 17, 9, 30, 6, 14, -10, 5, 11, 29, 42, 48, 10, -63, 26, -29, -11, 12, -55, -39, -38, -13, 8, 55, -63, -9, 10, 31, -18, -66, -40, -4, 10, 26, 40, -114, -17, -36, -12, -61, 14, 38, 0, 33, -60, 0, 72, 6, 79, 11, -3, 5, -5, 61, 5, -20, 47, 75, -10, -2, -4, 4, 24, 2, -34, 8, 33, 1, 67, 52, 9, -13, -19, -4, 4, -70, -97, -35, 25, 14, 34, 8, -14, -29, -38, -13, 36, -12, 16, -14, -11, 18, -3, 10, -30, -36, 60, -28, 6, 50, 13, -24, 1, 70, 61, 26, -51, 18, 0, -10, -97, -26, 6, -3, -15, -16, 26, -1, 27, 3, -19, -108, -47, -29, -15, -43, 60, -22, 45, -11, -64, 53, -1, -111, 0, -18, 4, -5, -39, -3, 14, -50, 32, -8, -5, -5, -30, -59, 38, 4, -6, 35, -58, 1, 9, -5, -15, 13, -71, -48, -11, -15, 19, -17, -11, 20, -55, 29, -4, 4, 13, 58, -24, 30, -43, -15, 21, -18, 33, 1, -13, 49, -16, -13, -2, -25, -35, 29, -24, -10, -16, 18, -11, 0, 25, -1, -7, 38, 6, -15, 27, 7, -5, -43, -73, -46, -19, 4, 37, 15, 7, 10, 22, -6, 11, -36, -17, 17, 6, 21, 16, 28, -11, -14, 47, -9, -41, -32, 22, 13, -24, 44, 12, 45, -7, -1, 12, 14, -99, -27, 2, -34, -60, 7, -4, 30, -21, -48, 3, -40, -28, 4, -19, -13, 28, -5, -51, -49, 31, -3, -30, 18, -7, 7, 31, -11, -9, 11, 49, -12, 15, -23, 9, -2, -18, -64, 34, -12, 12, 26, 21, -25, -15, -4, 8, 0, 8, 23, 31, -21, 0, -15, 16, -29, -35, 18, 41, 57, -4, -27, -38, 10, 37, 47, -19, -15, 66, 7, -31, -11, -6, 48, -4, -2, -45, 11, -39, -12, -19, -19, 0, -21, 37, -18, -4, -40, -4, -16, 22, 4, 26, 47, -42, 2, -13, 14, 12, -50, -7, -33, 12, -22, -21, 5, -16, -13, 15, 22, -33, 3, 6, -4, -17, 11, -48, -8, 17, 36, 10, -21, 3, 10, -36, -36, 1, -16, -41, -59, -14, -9, -51, -14, 19, 19, -28, 10, 15, -12, 46, -26, 27, 6, 9, 5, -52, -22, -92, -38, -35, 6, 12, -17, -1, -7, -17, -2, -54, 8, -36, -15, 4, 28, 3, -15, -19, -3, -7, 17, -20, -39, -20, -26, 17, -48, -48, 5, 20, -19, 13, -32, -20, -9, -67, 2, -14, -48, 5, 15, 3, 29, 4, 9, -14, -17, -7, 0, -14, -6, -8, 23, -16, -14, -31, 16, -16, -70, -33, 20, 7, -39, -1, 12, -13, -29, 5, -5, 9, -11, 64, 22, -30, -9, 12, -44, 14, -86, -4, 6, 35, 0, 11, 1, 15, -18, -17, 22, -68, -3, 39, 14, -14, -13, 0, -5, 3, 38, -19, 0, 2, -3, -10, 44, -3, 10, -9, -14, 0, -17, 42, -45, -8, 6, 2, -22, 3, 23, 0, 14, -12, -5, 0, -19, 13, -24, 30, -17, -28, -27, 0, -2, 1, 31, -14, -4, 7, -21, 36, 2, 4, 28, 25, -16, 8, -13, -10, -2, -33, -69, -22, -23, -16, -8, -9, 4, 7, 9, 46, -46, -23, -2, -42, -34, -35, -6, -1, 3, 9, 34, -4, 7, -6, -45, 26, -3, 5, 30, 13, 54, 18, 6, -44, 25, -32, -7, 10, 23, -19, -39, -43, 4, 7, 0, 6, 14, -14, 15, -31, -72, -33, 9, 11, -12, 19, -34, -8, 24, 69, -43, -28, -38, 14, -13, -1, 66, -16, 8, -16, 47, 5, -20, -36, -11, 20, 26, 4, 8, -23, 41, 0, -87, 11, 5, -25, -18, 0, -31, -7, 9, -21, 53, -8, -37, -24, -16, 16, 35, 6, 0, 18, 9,
    -- layer=3 filter=0 channel=7
    9, 15, 0, -39, -5, -15, 17, 14, -37, -57, 3, 13, 2, -9, 12, -20, 12, 27, -8, 17, 11, -1, -8, 29, 23, -56, 4, -39, 8, 3, 13, -7, 37, -24, 17, 14, 6, -6, 18, -14, -19, -20, 9, -18, -14, -7, -4, 40, -31, -10, -18, -9, 20, -19, 10, -23, 3, 34, 11, -28, 22, 10, -16, 2, 17, 4, -29, 1, 9, -2, -15, 13, -25, 3, 29, 15, 3, -77, -17, -20, -27, -37, 15, -15, -28, -27, 7, -24, -12, 11, 33, -22, 23, 4, 25, -18, 0, -7, -20, 15, -36, -24, 0, 28, -44, -31, 16, 11, -14, 26, 27, 24, -2, -8, 1, -36, 37, -27, -21, -25, 12, -2, 40, 29, 0, 0, 80, -9, -33, -7, -6, -11, -22, -2, -19, 7, -15, -66, -66, -12, -13, 39, -5, -18, 10, 30, -2, -63, -67, 11, -18, 8, -15, -2, -13, 35, 27, -64, 1, 2, -22, -69, 28, -1, 3, -3, -56, 9, 33, -21, 0, -15, -29, -22, 3, 13, -45, -2, 22, -7, -7, 12, -16, -10, -64, 1, -25, 12, 1, -13, -41, -39, 11, 12, -3, -3, -6, 9, -14, -4, -4, 11, 53, -47, 17, 2, -53, -8, -16, -32, 13, 0, 47, -53, 37, 17, -10, 11, -2, 17, 81, 19, 29, 13, -25, -31, -64, -15, -38, -11, 21, -9, 17, -42, 23, 5, -14, -31, -22, -14, 13, 45, -28, 30, -50, -42, -10, -47, 0, 28, -4, -30, 50, -6, 16, -10, 9, 13, -30, 20, 4, 5, 15, -7, -64, -51, 16, -16, 34, 5, 11, -21, 20, 9, -6, 19, 8, -8, 1, 0, 20, 5, -30, -35, 21, -31, -3, -23, 1, -66, -3, -7, 12, -8, 7, 28, 25, 40, -8, 7, 38, 38, 11, 4, -42, -45, 19, 20, 28, -3, -16, -17, 0, -26, 7, -15, 9, -30, -53, 20, 19, -33, -15, 0, 22, -19, -16, 5, -6, 23, -21, 25, -1, 13, -27, -45, -23, -5, -14, -58, 1, 0, -22, -10, 8, -7, -38, 4, -20, 34, 33, -5, -29, -18, 24, 13, -17, 8, 2, 36, 15, -6, 0, 59, -3, -27, 29, 32, -6, -23, 16, 26, 1, -28, -25, -7, -1, 5, 29, 41, 32, 27, -7, 0, 34, 28, -39, 9, 21, 8, 2, 3, -18, 43, -16, -12, 17, -39, -22, 14, 10, 27, 20, -54, -1, 17, -3, -4, -42, -6, -20, 34, 32, -60, 21, 2, -7, 79, 7, -3, -17, -14, -9, -56, 57, -20, -2, -29, 39, 18, -69, -53, 14, 13, 15, -8, -37, 44, 0, -7, -17, 46, 18, 21, -41, 0, -44, 26, -15, 24, -26, 14, -30, 19, 7, 11, 32, -5, -77, -23, 1, -7, -37, 18, 9, -29, 8, 17, 1, 10, -50, -38, 11, 14, 1, 23, 27, -27, -30, 13, 76, -53, 5, -34, 9, -4, -34, 28, -56, 0, 7, -16, 13, 31, 15, 37, -18, 15, -23, 15, -21, -13, -17, -73, 3, 7, -11, -14, -3, -6, -22, -28, -29, -9, -28, 12, 27, -2, 7, 9, 13, -1, -7, 12, -14, -6, -55, 1, -10, -63, 34, 25, -25, -30, 15, -26, 21, -34, -23, 18, -26, -104, 33, -74, -9, 29, -57, 43, -21, 12, -16, 24, -12, -6, -12, -15, 50, -36, -68, -29, -90, -31, 2, 12, -49, -3, -13, 32, 14, -124, 9, 25, 27, 41, 7, -34, 2, 27, -7, -8, 9, -44, 3, 5, -16, 0, 11, 30, -19, 28, -44, 0, 9, -9, 1, 84, 0, -10, -27, -7, -1, 17, 29, -34, 32, -27, 47, 19, -81, -12, 5, -109, -60, 33, 22, -43, -70, 0, 38, -3, 6, 44, 21, -1, -2, 54, -12, 20, 2, 11, -97, -67, -12, 22, 65, 3, 6, 10, -4, -5, -74, 0, -35, 21, -20, 0, 14, 6, 20, -13, 31, -27, -6, 38, -32, 35, 15, 18, -63, -45, 26, 10, 15, -25, 12, -30, 11, -94, -42, -37, 15, -87, 23, 17, -47, 43, -14, 6, 15, 12, 9, 36, -2, -93, 27, -15, 12, 20, -55, 23, -9, 19, 6, -51, -2, 8, -50, -17, -12, -11, -48, 5, 24, 32, 15, 8, 29, 16, 0, -9, -7, -5, 22, 11, 24, 56, 20, -20, -76, 39, 2, -43, -1, -10, -70, -14, -15, -2, 0, 9, -5, -22, 16, 12, 5, -24, -75, -18, -17, 35, -14, 5, 34, -29, -1, 24, -7, 17, -5, -14, 12, 16, -12, -11, -54, -34, 41, -13, 36, -10, 6, 15, 35, 5, 15, 20, -3, -21, 20, 34, -14, -1, 85, -66, 14, 16, 42, -4, -15, -17, -30, 9, 8, 37, 2, 30, 25, 22, -2, -3, -1, -10, -32, -22, 13, -5, 14, -4, 1, -56, 41, 29, 2, -29, -20, 55, 49, 0, -8, 7, 6, -50, 29, 68, -9, -33, 31, 18, -36, 8, 62, -7, 0, -16, 21, 23, 14, 18, 46, 26, 14, -4, -26, 56, -68, 9, -3, -3, -19, 13, -4, 2, -22, -73, 73, 67, -20, 25, 18, 30, 5, 9, 16, 50, -112, -39, 9, 16, 1, -11, -20, -14, -20, 22, 41, -8, -68, 27, 45, 3, -31, 0, -24, -6, 13, -5, -4, -18, 48, 36, -4, 22, 37, 8, -12, 17, 0, -56, -12, -25, -12, 0, -45, -5, -87, -2, -9, -42, -22, 4, 27, -23, -14, 0, 33, -4, -12, -60, 43, 15, -21, 21, -7, -22, -63, -37, 9, -19, -5, 45, 1, -14, 18, 2, 4, -47, -19, -75, -4, 5, -28, -27, -15, -7, 50, -6, 42, 12, 2, -50, -4, 27, 24, 8, 9, 20, 18, 5, 74, -16, 1, -4, 4, 37, -2, -4, -61, 28, 29, 35, 2, 49, -59, -23, 60, 25, -3, 12, 8, -1, -11, -5, 18, -1, 22, -5, 28, -3, 9, -8, -18, -6, -34, -11, 1, 2, 23, 7, -17, 16, -24, -9, 13, 35, -48, 42, 26, 3, -45, 6, -16, 19, -29, -6, 9, 6, 58, -2, -12, -58, 16, -28, -29, -3, -67, -21, 0, -19, 8, 50, 5, -28, -28, -12, -39, -65, -51, 44, 49, 41, -17, 0, 41, -13, -1, -9, -11, -9, -16, 33, -10, -10, -39, -40, 30, -28, -10, -1, 37, 2, 0, -59, -17, -27, 23, -97, -23, 2, -60, 10, 0, -36, -3, 14, -7, -7, 5, -34, 17, -13, 22, 12, -3, 47, -4, 4, 1, -4, 0, -40, 10, 17, 20, -21, 14, 6, 21, -26, 2, 1, 4, -15, 7, 8, 11, -10, 60, 0, -81, 11, 7, -8, -33, 54, -2, 16, 3, 28, 0, 7, -13, 0, 10, -8, -7, -17, 16, -41, -2, 3, -52, -15, -8, 34, 41, -9, 29, 23, 25, 30, -28, 59, 0, 20, 29, 18, -13, 21, -20, -86, -23, 22, 32, -35, -9, 1, 20, -21, 4, -11, -5, -13,
    -- layer=3 filter=0 channel=8
    32, 13, -60, -3, -72, -15, -18, 7, -7, -25, 5, 2, 22, -53, -61, 48, 10, 0, 5, -8, 17, 6, 12, -52, 15, 21, -24, 25, 19, -31, 25, 13, 21, 17, 12, -46, -10, 3, 25, -2, 1, -7, 5, -23, -14, -20, -14, 0, -9, 13, 1, -18, 40, 32, 1, 24, 29, 15, -5, -8, 66, 25, 36, -63, 16, -11, -36, -5, 0, -77, 0, 18, -67, 7, -21, 32, -1, -12, 0, -28, -40, 14, 11, -43, -3, -28, -5, 0, -11, -9, -42, -27, 19, -17, -2, -3, -36, 23, -60, -51, -78, 22, -10, 24, 4, 4, 14, 25, -3, 13, -32, 7, 3, 21, 21, 30, 0, -25, 1, -20, -16, 10, 17, 3, -18, -35, -2, 0, 6, -39, 3, -16, 14, -11, -11, -14, 4, 33, 25, -20, 13, -17, -10, 34, 0, 19, -20, -8, 26, -16, 7, -6, 7, 14, -7, 8, 13, -4, -19, -5, -8, 2, 4, -23, 1, 13, -20, 27, -13, 6, -16, 31, -43, 0, -20, 25, 0, 34, 24, -24, 26, 19, 15, 0, 25, -1, -35, -47, -33, 6, 34, -26, 13, 7, -50, 10, -31, -91, -9, 0, -61, -6, -33, -4, -7, 14, -22, -46, -42, 59, -15, -23, -37, 47, -6, -13, -5, -10, -5, 16, -1, -22, 22, -1, -20, -14, 10, 9, -31, -24, -22, -1, 30, -20, 16, -14, 3, 19, 23, -21, -26, 16, -37, 9, -11, -32, -28, 25, -12, 17, -18, -14, -16, -46, -22, -22, -11, 5, -39, -7, 12, -9, 9, -9, 67, -4, 23, -10, 40, 0, -5, -18, 14, 1, 43, -1, 17, -17, -17, -14, 25, 15, -13, -6, -4, 2, 42, 41, 3, 61, 23, 25, 1, 14, 35, 16, 39, 9, -2, 12, -42, -7, -18, 5, 9, 16, -8, -3, -6, -35, 9, 18, -13, -4, -14, 32, 9, 24, 22, -41, 9, -6, -64, -9, -15, -59, 11, 11, -58, -5, -3, -16, 14, 21, -55, 2, 31, -9, -7, -21, 14, 55, 42, 0, 17, 1, -16, -31, -10, -48, 8, 19, -51, -5, -24, -13, -30, -17, -27, -1, 4, 10, 3, 11, -18, 11, 26, -2, -6, 25, 34, 0, 33, -42, -12, 4, -2, -7, 23, 17, -42, 0, 4, -25, -43, -31, -37, -36, -36, -14, -15, -12, -31, -51, 9, 8, -6, -48, -22, 49, -27, 30, 33, 16, 37, -1, -13, -5, 16, 29, -15, -26, 27, -7, 46, 12, 13, -23, 1, -2, 3, 58, 6, -49, -53, -17, 10, 35, 1, 14, -19, -2, -49, 0, -4, -15, 21, 9, 8, -56, 37, 31, -17, -31, -48, -33, 38, -18, -12, 42, -7, -15, -71, -4, -2, -10, -28, 14, 4, -26, -24, -62, 6, -10, -27, 41, -8, -22, -21, 32, 16, 5, 13, 0, -15, -4, -24, -8, 10, -4, -73, 17, 25, -3, -26, -19, -9, -44, 30, -8, 12, -3, -13, -15, 0, 16, -6, 5, 14, 25, 6, -75, 20, 8, -14, 10, 10, 8, -1, -25, -23, 1, 9, -49, 0, -12, 6, -41, -14, 0, -36, 6, -12, -36, -7, -7, 3, 36, 6, 20, -19, 17, 49, -30, -6, -1, -22, 73, -13, 31, 0, 26, -9, 50, -10, -61, 12, -14, -21, -1, 35, 2, -25, 32, -9, -1, -16, 67, 17, 21, -10, 26, -19, 7, 7, 32, 0, -16, -11, -10, 2, 24, 53, -18, 28, -63, -5, 61, 32, 6, -6, -2, 0, 2, -16, -20, -29, -34, -11, -45, 54, -25, 22, 64, -9, -37, -18, 49, 24, -19, 15, 8, 18, 36, -26, -13, -4, -27, -17, 2, 50, 40, -19, 28, -15, -32, 35, -48, -3, -28, -18, 17, 15, -5, -1, 17, -37, -9, 53, -47, 29, 30, -2, -6, -32, -25, -23, 10, -20, 3, -15, -18, -1, -4, 16, 0, -10, -4, 27, -7, -18, -7, 0, -28, -29, -30, 7, 33, 26, 6, 38, -23, 0, -32, 38, 23, -13, 35, -43, 6, -12, 19, 27, -39, 21, 1, -16, -14, 28, -31, 28, -1, 0, 28, -44, 0, 13, -16, 14, 30, -21, -4, -37, -21, -7, -49, 4, 28, -30, -47, 35, 27, 12, -16, -4, -40, 11, -14, -75, -37, -6, 8, -10, 0, -4, 24, -15, 20, 30, -96, 19, 9, 7, -39, -16, -5, 34, -29, 11, -7, -14, -3, 1, -52, 15, 0, -2, -6, -12, -32, -17, 5, -42, -18, -48, -70, 26, 36, 12, -39, 4, 45, 9, 92, -11, 24, 22, -61, 15, 36, -23, -34, -41, 0, -29, 7, -12, 11, -56, -47, -5, -38, -55, 54, 3, 8, -30, 41, 10, 30, 19, 7, -13, -87, -24, 39, 13, -12, -32, 5, 9, 16, 12, 21, 2, 29, 11, -7, -12, 7, -6, -18, -18, -21, -8, 13, -19, -51, -23, -44, 13, 31, -31, -89, -9, 53, -76, -5, 18, 8, -39, -14, -18, -42, -26, -44, 9, -8, -65, -2, -16, 35, -15, 24, 20, 11, -70, 70, -8, -15, 19, -15, 14, -2, 0, 45, 44, -18, -27, -27, -6, -45, -20, 46, 65, 11, 13, -5, -12, 0, -89, 20, 17, -13, -13, -2, 36, 33, -42, -39, -47, -54, -2, -36, 41, 6, 11, 0, -20, -36, 4, -49, -52, -9, -31, -75, -23, 0, -3, -15, -29, -19, 72, 23, 27, 13, 56, -14, -21, -20, -59, -13, -20, 9, -26, 4, 41, 35, -45, 53, 8, -88, -2, -53, 23, 35, -24, -6, 11, 3, -3, 28, 14, 5, -27, 32, 8, 61, 21, 11, -8, -8, 2, 15, 32, -23, -11, -22, -12, -1, -61, 6, 37, 1, 43, -32, 10, 1, -13, 27, 18, -29, -2, -19, 1, -5, 69, 14, -23, -14, 17, -11, 44, 13, 0, 5, -11, 8, -24, 3, 13, -20, 38, -8, 67, 28, -57, 16, 8, 33, -51, 1, 67, -1, -5, 0, -8, -47, 7, 0, 15, -10, 34, 40, 50, -7, 27, -6, -8, -52, 11, 17, 26, -4, 12, -55, -63, -27, 2, 0, -49, 20, -31, 36, -47, 26, 12, -30, 44, -10, -8, 8, 2, -10, 25, 22, -54, -2, -11, -55, 6, 12, 3, 34, -38, 2, -51, 20, -21, -8, -24, -54, -45, 57, -63, -14, -4, -59, 1, 30, 3, 12, -32, 4, 21, 40, 81, -9, 7, 10, -24, -47, -6, -26, 48, 51, 0, 34, -49, -54, 7, -42, 56, -32, -14, -10, 21, 23, 13, -41, 19, -45, 2, 30, 14, 26, -16, 3, -3, 16, 18, 13, -111, 0, -1, -4, -35, -5, 30, 12, 40, -74, 97, 1, -1, 27, -5, -20, -4, 2, 47, -5, 12, -8, -63, 1, -26, -4, 60, 2, 103, 19, -58, -22, -22, -21, -1, -32, -58, -54, 12, -43, 13, -56, -78, 13, 8, -45, -41, 10, 12, -15, -7, 7, 19, 0, -12, 10, -33, 9, 0, 4,
    -- layer=3 filter=0 channel=9
    33, 6, -37, -28, 36, 46, -5, -4, -68, 24, 10, -1, -30, 15, 14, 27, 0, -37, 28, 7, 17, -5, 0, -44, -7, 43, 17, -4, -16, 19, -25, -76, 35, -35, 39, 11, 18, 28, 2, 12, 30, 25, -7, 17, 9, 10, -14, -10, 2, -22, 5, 8, 0, -1, 11, -10, 7, -23, 19, 23, -28, 0, -46, 8, -6, 18, -39, 8, -11, 56, 10, -1, 11, 2, 29, -4, 14, -20, 1, -20, 15, -10, -6, -58, -5, 12, -25, -11, -10, 15, -18, -18, -12, 31, 18, 2, -61, -5, 26, 4, -41, -82, -18, 19, -21, 15, 29, 18, -12, -35, 11, -2, -10, -2, -12, 23, 11, -59, 40, 14, -5, -10, -2, 6, -6, -14, 0, 12, -36, -5, -30, -32, 31, -4, -2, -12, -7, 8, 0, 2, -41, 39, -59, 31, 3, -27, 2, 30, -2, -6, 14, -35, -3, 23, -21, 41, 40, 1, 34, -27, -2, -57, 17, -2, 6, -8, -11, -19, 21, 36, 15, -21, -14, 15, -31, 2, 8, -1, 20, 11, 44, 46, -14, -12, -9, 5, 32, -15, -7, 22, -31, -20, 9, -18, 21, -9, -15, 33, 17, 4, -6, 4, 0, 9, 16, -30, 23, -60, 22, -21, 9, -70, -19, 3, -28, -17, 14, 1, 8, -22, 6, 66, 7, 29, 2, 17, -17, 32, 40, -41, 10, -24, 9, 56, 29, -11, 12, 42, -7, -36, 1, -26, 17, -31, 7, -25, -65, 24, 9, -17, 5, 3, 37, 20, -23, 6, -33, -37, -31, 16, 2, -50, -1, -15, -29, 20, -8, 37, -25, 0, -41, 11, 1, -11, 17, 23, 2, 5, -2, -30, 23, 2, -11, -3, -33, 4, -18, -20, 0, -92, -21, -10, -1, -21, -10, -11, 39, 6, 17, -19, -21, -51, -13, 10, 44, 27, 41, -9, 36, 21, 15, 8, -29, -27, 19, -11, 9, -11, -7, -6, -21, -21, -52, -14, -9, 27, -8, 0, 48, -15, 5, 16, 30, -23, 62, -35, 0, -4, -6, -36, -12, -23, -43, -19, 11, 10, 16, 29, 8, -15, -14, -16, 5, 17, 21, -3, 46, -29, -8, 4, -36, -10, 52, 23, 8, 27, 4, -45, -22, 4, 29, -43, -18, -72, 24, 7, 20, -9, 10, 28, 45, -24, 0, -10, 31, -39, 20, -67, 14, 13, -14, -15, 3, 63, 0, 0, 1, 14, -15, -13, -2, 21, -26, 13, -7, 17, -5, -9, 8, -30, -25, 3, -31, 14, 14, -18, 16, 0, 5, -10, -15, -24, 11, -9, -43, -1, -1, 16, -20, 42, -53, 20, -33, 12, -53, 0, -12, -49, -17, -15, -31, 1, 29, -8, -15, 38, 41, 1, -16, 5, 25, -4, -23, -9, 12, 8, -62, 0, 31, -2, 24, 21, 5, 11, -36, -12, 20, -36, -35, -6, -53, 3, 9, 4, -34, 31, 2, -22, 2, 1, 9, -52, 3, 14, -20, 2, 0, -76, -28, -3, -7, -26, 0, 29, 42, 12, 16, -1, 61, 22, -8, 33, 0, -17, -10, 13, 38, 6, -37, -24, 3, 5, -14, -96, -57, 10, -13, -12, -11, -10, 11, 86, 7, -33, 11, -9, 11, 43, -20, -49, -3, 58, 29, -19, -7, -1, 21, -28, 18, 46, 18, -28, -23, -23, 28, -21, 12, 34, 5, 32, 3, 12, -45, 30, -5, 1, 1, 15, -15, 9, -23, 42, 18, 4, 28, -11, 8, 43, -14, -24, -15, 9, -15, 8, 48, 20, -10, 37, -26, 0, 61, -5, -16, -3, 16, 17, 22, -36, 3, 91, 28, -1, 1, 29, -8, -49, -72, 10, -48, -27, 13, 6, -26, -18, -7, -9, 3, 4, -7, -15, -46, 33, -9, -20, -10, -22, -49, 18, 22, 27, -19, -18, 10, -74, -3, -47, 56, -11, 15, 39, -34, 15, 4, -2, 35, -34, -7, -31, -3, -31, -19, -77, 13, 2, -31, 2, 4, -1, 35, -11, 7, 6, -20, -15, 25, 44, 16, -14, 14, 26, 43, -19, 0, -2, 0, 34, 20, 24, -5, 4, 38, -18, 28, -35, 15, -8, -5, 58, 5, 19, 23, 3, -5, 0, 4, -9, 15, 0, -1, -32, -23, -3, 0, -31, 2, 12, -6, -16, -11, -39, -16, -30, -34, -48, -3, 12, -27, 2, 22, 7, -12, -12, 11, 15, 22, 0, 26, -8, 10, -3, -26, 44, -6, -9, 23, -9, -12, -42, 8, 5, -5, -9, -19, 1, -14, 7, -33, 36, 1, 0, 0, 26, -4, -8, -33, -44, -1, 30, -15, -15, 1, -31, -9, -39, 68, 29, 42, 6, 28, 17, -7, -38, 1, -37, 20, 0, -14, 4, 13, 7, 7, -91, -40, 28, -17, 0, -21, 25, -64, -26, 14, -9, -92, -20, -13, -18, -17, 45, -52, 18, 11, 23, 21, 20, -5, -59, -78, 13, -1, -4, -26, 30, 31, 15, -17, -2, 14, 36, -4, -91, 8, 50, 6, -15, -44, -24, 6, 14, 5, 2, -56, -76, 3, -31, -20, 30, 52, -7, 8, -72, -20, -45, -14, -34, 29, -3, -11, -51, -16, 0, -15, -2, 51, -1, 3, 7, -53, -12, -2, -64, -8, 42, 15, 4, -2, -12, -14, -11, 35, 6, 49, -26, 7, -31, -25, -41, 17, 4, -28, 18, 35, 26, -42, -14, -25, -23, -11, 6, -30, -6, -18, -14, 34, 27, 24, -14, 67, -11, 14, 17, -89, -31, -13, 37, -27, -17, -10, 33, 4, -39, 40, 18, -6, 16, 8, 1, 2, 20, 22, -32, -52, 48, -4, -3, -33, 17, 17, 11, -11, -20, 41, 0, -5, 4, 6, -17, -1, 11, -19, 23, 13, -1, 9, 14, 24, -24, -49, -49, 0, 23, -18, 28, -19, 15, -43, -60, -37, 16, -14, -15, 8, 4, 33, -2, 4, 1, -10, -57, 61, 14, 1, -23, 39, 19, -3, 13, -5, -1, -9, -3, 10, -11, -15, 47, -70, -6, -29, 25, 12, -21, -3, -6, -14, -14, 12, 13, -2, 9, 11, 8, -9, -50, 0, 5, -7, -37, -46, -6, 47, 0, -36, -12, -71, 33, -14, -15, 23, -44, -19, -1, -14, 53, 42, -41, 28, 10, -21, 6, -32, 5, -47, 0, 27, -21, -18, -8, 36, -65, -27, -13, 7, -6, -3, -46, -17, 21, -7, -14, 0, 34, -1, -28, -31, -7, 15, -15, 9, 14, 20, -8, -35, 24, -1, 21, 33, -2, -14, -37, 64, 11, 12, 19, 29, -35, -4, 0, -3, 50, 21, 6, -46, -25, -78, -42, -53, -15, -50, -17, 2, -68, -5, 16, 55, -22, -14, -103, -45, -26, -8, -36, -10, -8, -4, -24, 0, 15, 15, -8, 22, 12, -27, -21, -76, 9, -21, 19, -7, 10, 17, 17, 7, -3, 4, 7, 18, -50, 23, 41, 2, -58, -17, 11, 20, -3, -56, 31, 4, -4, 18, -21, -10, -21, -1, -26, 20, 5, -4, 0, -1, 70, -40, -27, 43, -15, 11, 12, -49, 0, -27, 26, 19, 0,

    others => 0);
end iwght_package;
