LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
	PACKAGE inmem_package is
		type padroes is array(0 to 4000000) of integer;

		constant input_mem: padroes := ( 
					-- bias

					-- weights

			0, 11, 0, 0, 32, 0, 4, 
			213, 44, 0, 8, 97, 7, 42, 
			66, 42, 0, 0, 340, 30, 0, 
			0, 78, 0, 40, 66, 0, 0, 
			0, 320, 30, 0, 0, 76, 0, 
			0, 0, 50, 0, 66, 15, 0, 
			24, 0, 60, 12, 4, 4, 0, 
			

			0, 0, 0, 123, 122, 0, 2, 
			59, 0, 0, 41, 0, 16, 118, 
			0, 122, 0, 0, 116, 132, 0, 
			0, 48, 0, 103, 0, 199, 0, 
			0, 162, 15, 0, 95, 175, 0, 
			0, 0, 365, 33, 73, 0, 0, 
			139, 0, 120, 25, 0, 4, 0, 
			

			71, 62, 74, 60, 68, 93, 117, 
			104, 91, 103, 90, 45, 103, 112, 
			66, 60, 77, 93, 0, 76, 86, 
			0, 40, 18, 92, 53, 115, 146, 
			0, 16, 60, 50, 38, 40, 112, 
			2, 0, 0, 0, 0, 0, 0, 
			0, 27, 0, 0, 0, 0, 0, 
			

			54, 113, 69, 0, 0, 0, 0, 
			0, 0, 18, 31, 0, 42, 0, 
			0, 0, 0, 14, 0, 0, 27, 
			0, 0, 1, 26, 0, 54, 77, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 38, 0, 176, 0, 
			259, 0, 119, 66, 14, 71, 309, 
			181, 336, 0, 60, 100, 93, 0, 
			41, 57, 0, 0, 314, 39, 0, 
			0, 0, 271, 0, 83, 16, 24, 
			0, 325, 98, 0, 0, 0, 0, 
			468, 0, 0, 1, 0, 0, 28, 
			

			60, 134, 70, 8, 0, 0, 0, 
			0, 0, 0, 29, 0, 50, 0, 
			7, 0, 14, 64, 0, 78, 0, 
			27, 0, 0, 105, 0, 52, 0, 
			49, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 22, 0, 
			0, 0, 0, 85, 0, 68, 0, 
			85, 0, 0, 39, 0, 46, 0, 
			84, 0, 54, 0, 0, 0, 0, 
			0, 0, 192, 0, 57, 0, 0, 
			93, 0, 98, 56, 43, 3, 69, 
			

			0, 0, 37, 1, 68, 70, 0, 
			3, 117, 115, 48, 0, 16, 0, 
			0, 0, 77, 134, 0, 4, 68, 
			132, 0, 0, 0, 0, 0, 0, 
			88, 116, 12, 146, 0, 0, 0, 
			0, 0, 0, 0, 16, 105, 83, 
			0, 0, 0, 9, 21, 0, 0, 
			

			0, 5, 0, 141, 0, 0, 0, 
			0, 0, 41, 32, 0, 73, 0, 
			1, 0, 0, 97, 0, 105, 0, 
			72, 0, 79, 103, 0, 20, 0, 
			92, 0, 0, 0, 106, 0, 0, 
			0, 0, 35, 0, 0, 0, 0, 
			0, 141, 0, 0, 0, 0, 0, 
			

			0, 5, 0, 0, 0, 0, 0, 
			0, 0, 0, 28, 0, 0, 32, 
			0, 0, 0, 35, 0, 57, 72, 
			0, 0, 0, 0, 0, 65, 0, 
			0, 0, 0, 23, 20, 46, 0, 
			0, 0, 0, 26, 0, 0, 0, 
			0, 202, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 52, 166, 3, 0, 
			69, 0, 0, 0, 0, 0, 0, 
			12, 263, 79, 0, 0, 0, 0, 
			0, 3, 0, 0, 34, 46, 39, 
			0, 0, 0, 30, 40, 75, 30, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 151, 0, 0, 
			0, 78, 0, 0, 262, 0, 0, 
			0, 0, 46, 0, 216, 0, 0, 
			0, 101, 40, 0, 0, 0, 0, 
			184, 113, 0, 0, 0, 31, 42, 
			330, 0, 0, 16, 14, 127, 15, 
			

			0, 0, 9, 0, 0, 0, 0, 
			0, 0, 0, 44, 0, 32, 0, 
			0, 0, 0, 81, 0, 0, 0, 
			0, 0, 0, 0, 0, 18, 9, 
			0, 0, 6, 90, 0, 0, 0, 
			0, 79, 0, 0, 18, 34, 3, 
			0, 0, 60, 35, 41, 2, 73, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 24, 0, 0, 92, 
			0, 97, 0, 0, 0, 0, 0, 
			0, 7, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			149, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 23, 0, 10, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 149, 131, 56, 0, 28, 
			27, 99, 131, 77, 67, 70, 21, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			1, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 1, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 3, 
			0, 0, 0, 0, 0, 107, 10, 
			0, 0, 0, 0, 20, 0, 0, 
			

			0, 137, 0, 0, 0, 49, 0, 
			0, 20, 52, 114, 0, 161, 0, 
			0, 0, 0, 200, 0, 144, 95, 
			128, 0, 0, 59, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 86, 19, 15, 
			0, 0, 43, 105, 101, 31, 0, 
			

			32, 0, 0, 40, 32, 93, 108, 
			0, 0, 0, 0, 0, 0, 115, 
			10, 0, 0, 0, 0, 0, 15, 
			0, 9, 0, 0, 0, 0, 1, 
			0, 0, 0, 0, 30, 54, 149, 
			216, 0, 57, 133, 101, 145, 163, 
			270, 112, 90, 96, 106, 123, 75, 
			

			0, 0, 0, 0, 9, 35, 0, 
			53, 0, 93, 26, 0, 24, 0, 
			0, 0, 0, 23, 0, 0, 11, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 35, 0, 16, 117, 0, 
			0, 0, 39, 82, 54, 46, 37, 
			39, 0, 0, 0, 32, 0, 38, 
			

			78, 89, 167, 82, 75, 89, 69, 
			241, 109, 119, 128, 216, 145, 85, 
			188, 156, 62, 157, 410, 120, 36, 
			55, 78, 218, 130, 307, 100, 110, 
			74, 274, 123, 83, 46, 0, 83, 
			0, 320, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			54, 44, 57, 43, 31, 0, 8, 
			106, 11, 0, 0, 38, 0, 39, 
			145, 20, 52, 0, 82, 25, 12, 
			53, 0, 0, 39, 90, 52, 77, 
			24, 119, 0, 20, 44, 50, 8, 
			0, 133, 125, 46, 53, 80, 77, 
			49, 63, 23, 76, 62, 72, 101, 
			

			132, 145, 147, 46, 81, 67, 90, 
			120, 202, 116, 96, 138, 89, 94, 
			137, 108, 111, 93, 156, 85, 96, 
			55, 120, 32, 34, 107, 89, 139, 
			34, 207, 93, 117, 0, 0, 110, 
			0, 9, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 89, 0, 87, 0, 0, 
			144, 64, 7, 0, 229, 0, 0, 
			37, 8, 47, 0, 488, 0, 0, 
			0, 0, 189, 0, 266, 0, 43, 
			0, 236, 0, 0, 0, 0, 155, 
			87, 394, 0, 0, 0, 107, 51, 
			138, 0, 14, 23, 80, 87, 147, 
			

			0, 25, 0, 83, 0, 77, 0, 
			0, 0, 13, 165, 0, 189, 59, 
			158, 0, 0, 305, 0, 243, 72, 
			292, 13, 0, 137, 0, 182, 0, 
			203, 0, 27, 51, 103, 0, 0, 
			0, 0, 229, 0, 47, 0, 0, 
			0, 0, 53, 49, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 42, 0, 11, 46, 
			0, 0, 0, 0, 0, 114, 0, 
			116, 0, 0, 0, 0, 0, 0, 
			0, 0, 7, 0, 0, 0, 0, 
			

			38, 0, 14, 157, 117, 66, 89, 
			0, 0, 35, 26, 0, 0, 24, 
			0, 107, 121, 0, 0, 2, 0, 
			0, 30, 83, 53, 0, 67, 0, 
			0, 0, 12, 33, 154, 98, 63, 
			192, 35, 228, 132, 24, 0, 16, 
			0, 258, 55, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 24, 23, 0, 
			0, 0, 0, 30, 61, 9, 64, 
			122, 0, 0, 0, 0, 36, 0, 
			157, 137, 22, 90, 16, 72, 0, 
			254, 167, 185, 248, 245, 278, 316, 
			290, 316, 279, 270, 286, 295, 339, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 67, 50, 60, 
			135, 0, 0, 27, 161, 31, 65, 
			87, 11, 0, 0, 190, 0, 46, 
			89, 95, 0, 26, 0, 0, 72, 
			0, 185, 0, 0, 124, 172, 84, 
			242, 0, 93, 171, 201, 178, 192, 
			

			131, 170, 185, 115, 98, 96, 98, 
			169, 184, 163, 88, 97, 30, 97, 
			0, 136, 0, 14, 126, 4, 57, 
			0, 108, 101, 0, 98, 0, 61, 
			0, 17, 43, 0, 11, 31, 108, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			252, 227, 107, 240, 141, 92, 199, 
			75, 201, 118, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 11, 
			0, 0, 0, 0, 56, 32, 36, 
			0, 0, 0, 30, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			29, 19, 0, 0, 0, 0, 0, 
			279, 30, 122, 189, 101, 140, 153, 
			199, 274, 141, 136, 155, 206, 205, 
			
