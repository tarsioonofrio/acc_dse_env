-- https://docs.xilinx.com/r/en-US/ug953-vivado-7series-libraries/BRAM_SINGLE_MACRO

library UNISIM;
use UNISIM.vcomponents.all;
library UNIMACRO;
use unimacro.Vcomponents.all;


-- BRAM_SINGLE_MACRO: Single Port RAM
--                    7 Series
-- Xilinx HDL Language Template, version 2021.2

-- Note -  This Unimacro model assumes the port directions to be "downto".
--         Simulation of this model with "to" in the port directions could lead to erroneous results.

---------------------------------------------------------------------
--  READ_WIDTH | BRAM_SIZE | READ Depth  | ADDR Width |            --
-- WRITE_WIDTH |           | WRITE Depth |            |  WE Width  --
-- ============|===========|=============|============|============--
--    37-72    |  "36Kb"   |      512    |    9-bit   |    8-bit   --
--    19-36    |  "36Kb"   |     1024    |   10-bit   |    4-bit   --
--    19-36    |  "18Kb"   |      512    |    9-bit   |    4-bit   --
--    10-18    |  "36Kb"   |     2048    |   11-bit   |    2-bit   --
--    10-18    |  "18Kb"   |     1024    |   10-bit   |    2-bit   --
--     5-9     |  "36Kb"   |     4096    |   12-bit   |    1-bit   --
--     5-9     |  "18Kb"   |     2048    |   11-bit   |    1-bit   --
--     3-4     |  "36Kb"   |     8192    |   13-bit   |    1-bit   --
--     3-4     |  "18Kb"   |     4096    |   12-bit   |    1-bit   --
--       2     |  "36Kb"   |    16384    |   14-bit   |    1-bit   --
--       2     |  "18Kb"   |     8192    |   13-bit   |    1-bit   --
--       1     |  "36Kb"   |    32768    |   15-bit   |    1-bit   --
--       1     |  "18Kb"   |    16384    |   14-bit   |    1-bit   --
---------------------------------------------------------------------

entity ifmap_18k_layer1_entity2 is
    generic (
        DEVICE: string := "7SERIES"
        );
  
    port (
        RST  : in std_logic;
        CLK  : in std_logic;
        EN   : in std_logic;
        WE   : in std_logic_vector(2-1 downto 0);;
        DI   : in std_logic_vector(INPUT_SIZE-1 downto 0);
        ADDR : in std_logic_vector(10-1 downto 0);
        DO   : out std_logic_vector(INPUT_SIZE-1 downto 0)
    );
  end ifmap_18k_layer1_entity2;

  architecture a1 of bram is

    begin

    BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
    generic map (
       BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
       DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
       DO_REG => 0,                     -- Optional output register (0 or 1)
       INIT => X"000000000000000000",   -- Initial values on output port
       INIT_FILE => "NONE",
       WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       SRVAL => X"000000000000000000",  -- Set/Reset value for port output
       WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
       -- The following INIT_xx declarations specify the initial contents of the RAM
       INIT_00 => X"001f0034003500240021001a000a00260024000b000a00080051003300280020",
       INIT_01 => X"0053005e004b002b0019001a00330014000e00120019002e0045002f0036005b",
       INIT_02 => X"005d0042003b0015001b0071005e00150035007e00440064003b0033003b0067",
       INIT_03 => X"0038003900250001007f009e0028001300bd007e007d004b002e005b007f0050",
       INIT_04 => X"0047003c0015007a009400430017005a007500a80065004e007800810046003b",
       INIT_05 => X"004c0033008e00a500400039003900a50085006a0050005f0078004c0048004b",
       INIT_06 => X"002600b000b800660073003800660059004e0051003300650041002c002b000e",
       INIT_07 => X"00c000b300860075006f0033005f00790042005a00400025002f0027002700c7",
       INIT_08 => X"00ab008b00a2009e0065009100b90079003c00400047005a0071006800c100cb",
       INIT_09 => X"009d00c900e700a5008a0085007c006f007800800088008a008e008c00a100b1",
       INIT_0A => X"00e500af007a00750070007100760084008c0095009a00a3009d008500a600ef",
       INIT_0B => X"008800800079007300770082008c009b009300a300ab0097008f007f00a70074",
       INIT_0C => X"007f0089007e007c008800860085009a00af008d000000000000000000000000",
       INIT_0D => X"0000000000000013001c000b000000000000000000000000000000000000000b",
       INIT_0E => X"00140033000000000014001e00000000003f0000000000000000003e001c0028",
       INIT_0F => X"00000000000000000007001e00000019000000000000000c0000000000000000",
       INIT_10 => X"00000000001a0006000e0000000000000009000000000000000f0004001d0000",
       INIT_11 => X"00000008000000000025002f00000002004f0003000000000000000600000026",
       INIT_12 => X"001c00000000000000000018000d000d00000000000500000009000000180008",
       INIT_13 => X"000000000000000200000007000000000000003d001e000000000000001c0000",
       INIT_14 => X"0010000000000000002e00000022003200030000000000360026003a000d0000",
       INIT_15 => X"000000000000000a00000012001500000000002e001f00310001000000000008",
       INIT_16 => X"00000000002200000000000000000019000f000d000000000000001600210041",
       INIT_17 => X"00000000000000a20052003f0037000c000600000002000000000000000d0036",
       INIT_18 => X"0000004100560000000200000000000000000000000300000000000200000025",
       INIT_19 => X"003e0006000000000001000000000007000a000000000042000c000000180036",
       INIT_1A => X"0024001300090000000000000005000000000000000400000000000000000000",
       INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_1D => X"00000004001f000000000000000000000000000b000000000000000000000000",
       INIT_1E => X"0005002d00000007000000020001000000020000000000000000000000000002",
       INIT_1F => X"003b000000000003000000100001000600000000002c0000000000000000005d",
       INIT_20 => X"00000000000e000000000000000000000000001c000f00000000000000520000",
       INIT_21 => X"00000012001300000004000000000000000c0017000000050000002d00000000",
       INIT_22 => X"001d00030000000000160000001100000012000000000008000000110000001b",
       INIT_23 => X"00000000000900190000003b0000000300100000000500000000001200120000",
       INIT_24 => X"00000033000d0000005800000000002d00040000000200280033003e002c001d",
       INIT_25 => X"007000360000003b0000002e004e004e00440049004f00560058005a0053005a",
       INIT_26 => X"006f00480008000000490048004a004c0054005b005b0057005d005e005a0060",
       INIT_27 => X"008a0000003100500045004d005300570061006400610074005e005000670067",
       INIT_28 => X"00410049005f00550049005200520052005e006b00530045002f002e0033002e",
       INIT_29 => X"002f002f0031002f002b0023001c0027002600270024003200320035002d0034",
       INIT_2A => X"00550013002500040021001300150024002d0028001a003b0034002e0038002c",
       INIT_2B => X"00000000001a004f000a000b00040027003900000079002c003600250023001a",
       INIT_2C => X"000800180053000000120000000e005300000063000a0049002c001a00000000",
       INIT_2D => X"0008005f000b0000001e00000039000000380000002e00490000000000000000",
       INIT_2E => X"00bf0000000000230004000d00000015000c000000610050000a0000000000a4",
       INIT_2F => X"00000000001e0027000d000000000001000000450068000000080000007c0000",
       INIT_30 => X"0000002a00220012000000170000003c001100030000001c0031000600220000",
       INIT_31 => X"0026003a0044000a00180000004a00000019002a000e0017000a000000050048",
       INIT_32 => X"0056001c00510011000000a30000000b005600000000000000140028002d001e",
       INIT_33 => X"0000004000280000009800000000000000000000000900100010000e00110000",
       INIT_34 => X"000300410048001f000000090005000a00080010001400170010000800170000",
       INIT_35 => X"0010007400000000001100000009000d0010000d00090000002600000000000d",
       INIT_36 => X"0019000000000016000c0009001800100000000b003100030000000000000000",
       INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_38 => X"0000000400000000000000000001000000000000000000000000000000000000",
       INIT_39 => X"0000000000000000000000000000000000000000000400120000000000000000",
       INIT_3A => X"0005000000000000000000000000000000000001002700000000003800080000",
       INIT_3B => X"0000000000000000000000000004000000000000000000000000000000000000",
       INIT_3C => X"000000140000000000000000000f000000000000000000000000000000000000",
       INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_3F => X"0000000000000000000000000000000000000000000000120000000000000000",

       -- The next set of INITP_xx are for the parity bits
       INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

    port map (
       DO => DO,      -- Output data, width defined by READ_WIDTH parameter
       ADDR => ADDR,  -- Input address, width defined by read/write port depth
       CLK => CLK,    -- 1-bit input clock
       DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
       EN => EN,      -- 1-bit input RAM enable
       REGCE => REGCE, -- 1-bit input output register enable
       RST => RST,    -- 1-bit input reset
       WE => WE       -- Input write enable, width defined by write port depth
    );


-- End of BRAM_SINGLE_MACRO_inst instantiation
