library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    234, 234, 239, 238, 237, 225, 247, 258, 240, 209, 183, 193, 199, 202, 201, 
    236, 241, 247, 244, 249, 228, 206, 211, 169, 130, 76, 82, 128, 190, 202, 
    164, 236, 247, 248, 255, 246, 143, 100, 86, 124, 74, 72, 51, 114, 191, 
    33, 157, 235, 251, 204, 182, 120, 68, 69, 156, 82, 88, 54, 40, 179, 
    41, 137, 193, 260, 170, 123, 88, 55, 50, 137, 105, 52, 75, 36, 91, 
    48, 135, 181, 178, 199, 139, 106, 78, 25, 196, 93, 51, 92, 58, 34, 
    48, 84, 170, 172, 182, 171, 152, 95, 47, 191, 73, 47, 69, 86, 67, 
    65, 87, 74, 148, 168, 210, 90, 109, 79, 187, 99, 48, 86, 103, 132, 
    72, 110, 11, 130, 106, 124, 98, 86, 119, 116, 128, 51, 79, 138, 195, 
    127, 117, 24, 107, 70, 85, 126, 94, 69, 121, 52, 40, 92, 196, 201, 
    151, 117, 34, 188, 50, 49, 120, 101, 30, 18, 4, 3, 12, 63, 48, 
    74, 117, 91, 219, 63, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 54, 139, 141, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 102, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=1
    47, 65, 51, 50, 40, 60, 57, 51, 43, 53, 67, 69, 64, 54, 45, 
    39, 64, 51, 53, 43, 50, 49, 73, 83, 44, 35, 43, 55, 55, 48, 
    82, 62, 48, 52, 41, 88, 78, 51, 35, 35, 68, 52, 43, 35, 61, 
    68, 0, 49, 45, 60, 32, 58, 43, 40, 46, 88, 67, 66, 40, 38, 
    65, 27, 50, 3, 84, 48, 106, 74, 65, 1, 64, 62, 46, 46, 17, 
    62, 86, 75, 56, 156, 118, 112, 63, 62, 0, 98, 83, 50, 45, 30, 
    53, 107, 78, 93, 64, 57, 123, 74, 88, 22, 100, 60, 33, 38, 48, 
    73, 110, 15, 67, 11, 101, 120, 90, 86, 42, 89, 71, 47, 70, 53, 
    93, 96, 76, 70, 42, 85, 76, 56, 32, 40, 93, 95, 51, 44, 35, 
    108, 84, 109, 32, 100, 44, 37, 78, 41, 106, 86, 47, 34, 39, 55, 
    92, 88, 110, 11, 64, 32, 66, 136, 102, 38, 12, 9, 10, 18, 21, 
    65, 97, 80, 43, 170, 103, 68, 69, 52, 28, 25, 27, 28, 22, 35, 
    9, 48, 41, 136, 120, 39, 42, 35, 24, 16, 12, 17, 34, 33, 14, 
    26, 22, 32, 177, 49, 27, 30, 35, 35, 31, 24, 36, 24, 12, 59, 
    36, 32, 27, 78, 27, 35, 45, 37, 25, 23, 29, 16, 0, 29, 36, 
    
    -- channel=2
    132, 151, 150, 146, 139, 154, 149, 142, 135, 114, 106, 120, 140, 133, 117, 
    134, 163, 156, 147, 153, 241, 155, 139, 103, 132, 140, 112, 96, 104, 120, 
    95, 99, 145, 146, 141, 142, 110, 80, 101, 198, 166, 149, 111, 61, 127, 
    112, 140, 138, 151, 152, 152, 185, 126, 110, 156, 171, 124, 97, 52, 104, 
    182, 234, 152, 197, 335, 292, 210, 142, 88, 168, 212, 146, 129, 91, 69, 
    178, 224, 167, 161, 213, 237, 255, 167, 113, 246, 212, 116, 124, 120, 108, 
    206, 219, 116, 137, 180, 258, 237, 204, 124, 251, 181, 131, 123, 147, 123, 
    247, 259, 147, 154, 167, 267, 193, 146, 119, 216, 178, 116, 122, 137, 121, 
    273, 275, 159, 190, 164, 139, 138, 153, 145, 159, 106, 69, 90, 133, 157, 
    257, 261, 178, 227, 150, 148, 201, 245, 146, 107, 70, 59, 119, 171, 135, 
    250, 265, 176, 327, 341, 224, 251, 215, 138, 112, 95, 131, 129, 104, 85, 
    119, 228, 232, 381, 197, 68, 96, 95, 80, 90, 96, 109, 121, 121, 113, 
    92, 119, 245, 302, 86, 119, 112, 105, 95, 99, 114, 128, 122, 121, 155, 
    92, 103, 174, 177, 95, 123, 118, 106, 111, 119, 111, 98, 103, 132, 96, 
    110, 111, 109, 66, 60, 73, 84, 111, 140, 145, 110, 107, 175, 168, 81, 
    
    -- channel=3
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 67, 0, 0, 96, 40, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 89, 0, 0, 111, 29, 42, 0, 0, 89, 19, 0, 0, 0, 0, 
    0, 77, 0, 0, 17, 73, 78, 0, 0, 112, 0, 0, 0, 0, 0, 
    45, 60, 0, 0, 0, 136, 0, 0, 0, 69, 0, 0, 0, 0, 0, 
    82, 109, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    97, 107, 0, 50, 0, 0, 0, 38, 0, 0, 0, 0, 0, 0, 0, 
    125, 97, 0, 167, 91, 10, 92, 55, 0, 0, 0, 0, 0, 0, 0, 
    49, 91, 34, 259, 76, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 30, 92, 194, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 87, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 20, 0, 
    
    -- channel=4
    123, 115, 120, 123, 123, 114, 126, 126, 119, 111, 97, 96, 100, 106, 103, 
    120, 117, 120, 126, 122, 137, 130, 113, 85, 73, 84, 79, 76, 95, 108, 
    101, 97, 130, 124, 131, 112, 98, 59, 63, 84, 101, 75, 79, 72, 94, 
    85, 93, 135, 122, 122, 93, 107, 82, 77, 82, 104, 82, 64, 60, 67, 
    100, 131, 142, 98, 145, 132, 108, 82, 65, 64, 108, 94, 70, 60, 61, 
    122, 134, 145, 132, 93, 109, 128, 88, 75, 93, 141, 82, 69, 68, 59, 
    117, 140, 110, 106, 79, 129, 139, 119, 78, 105, 121, 87, 72, 79, 89, 
    137, 115, 107, 111, 97, 138, 127, 95, 84, 111, 114, 84, 65, 94, 88, 
    146, 132, 128, 96, 132, 78, 89, 95, 82, 112, 91, 60, 54, 80, 118, 
    141, 140, 118, 86, 104, 84, 82, 121, 109, 84, 58, 28, 59, 114, 115, 
    126, 143, 115, 117, 171, 126, 129, 117, 90, 57, 48, 59, 71, 89, 92, 
    88, 118, 121, 185, 173, 74, 60, 56, 56, 58, 63, 61, 65, 72, 68, 
    82, 85, 114, 198, 77, 60, 59, 57, 58, 60, 60, 71, 74, 66, 75, 
    69, 64, 97, 136, 76, 63, 66, 58, 53, 59, 66, 67, 62, 74, 91, 
    76, 56, 76, 54, 64, 57, 59, 60, 65, 71, 70, 58, 75, 97, 63, 
    
    -- channel=5
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 12, 0, 2, 0, 29, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 27, 14, 0, 0, 41, 24, 44, 0, 0, 
    122, 0, 0, 0, 0, 0, 27, 35, 9, 0, 63, 7, 35, 16, 0, 
    147, 0, 20, 0, 51, 41, 72, 50, 18, 0, 43, 77, 1, 47, 0, 
    111, 0, 40, 0, 0, 34, 73, 59, 71, 0, 92, 82, 0, 34, 28, 
    112, 56, 0, 32, 0, 0, 50, 63, 90, 0, 112, 62, 0, 0, 34, 
    96, 76, 58, 34, 0, 0, 96, 10, 46, 0, 61, 65, 0, 0, 0, 
    106, 33, 135, 0, 27, 0, 36, 16, 0, 19, 0, 54, 0, 0, 0, 
    43, 31, 148, 0, 86, 2, 0, 63, 23, 5, 53, 7, 0, 0, 0, 
    0, 40, 137, 0, 179, 94, 0, 55, 113, 57, 25, 20, 13, 3, 41, 
    0, 0, 86, 0, 172, 97, 21, 22, 50, 30, 31, 29, 36, 38, 56, 
    69, 0, 0, 52, 179, 39, 43, 33, 38, 34, 35, 39, 46, 45, 43, 
    84, 38, 0, 114, 78, 31, 57, 39, 31, 35, 40, 40, 53, 25, 61, 
    90, 42, 23, 31, 45, 9, 25, 37, 31, 45, 61, 35, 11, 84, 112, 
    
    -- channel=6
    134, 134, 137, 136, 137, 139, 138, 139, 135, 123, 114, 119, 126, 124, 118, 
    133, 143, 141, 138, 143, 162, 138, 130, 109, 114, 108, 104, 108, 117, 122, 
    103, 131, 142, 139, 142, 136, 98, 98, 95, 129, 91, 88, 79, 96, 119, 
    77, 142, 139, 144, 131, 140, 119, 86, 82, 121, 90, 88, 66, 59, 119, 
    90, 149, 131, 171, 172, 161, 108, 79, 66, 132, 122, 85, 88, 63, 94, 
    99, 126, 124, 130, 125, 122, 115, 96, 67, 168, 109, 70, 91, 79, 78, 
    106, 108, 114, 104, 135, 150, 124, 112, 67, 168, 93, 80, 92, 98, 83, 
    119, 115, 113, 124, 137, 151, 97, 92, 76, 143, 93, 74, 89, 95, 90, 
    123, 136, 77, 114, 118, 106, 93, 96, 111, 130, 88, 52, 83, 102, 128, 
    122, 130, 70, 141, 83, 103, 131, 121, 103, 72, 57, 61, 98, 135, 124, 
    143, 137, 81, 184, 128, 116, 136, 100, 66, 81, 76, 82, 90, 112, 101, 
    97, 124, 114, 206, 85, 43, 70, 66, 50, 62, 58, 64, 63, 61, 53, 
    50, 93, 146, 145, 34, 59, 56, 56, 53, 55, 61, 64, 59, 61, 74, 
    38, 58, 128, 67, 51, 66, 58, 55, 56, 58, 57, 49, 50, 63, 45, 
    40, 47, 64, 54, 48, 49, 47, 55, 67, 68, 51, 55, 84, 66, 28, 
    
    -- channel=7
    0, 0, 0, 0, 0, 0, 0, 0, 3, 10, 5, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 30, 5, 22, 0, 7, 0, 0, 0, 0, 
    19, 0, 0, 0, 0, 0, 31, 15, 5, 0, 22, 3, 27, 0, 0, 
    89, 0, 0, 0, 6, 0, 10, 33, 0, 0, 29, 9, 23, 21, 0, 
    93, 0, 32, 0, 0, 19, 38, 33, 9, 0, 9, 60, 0, 30, 0, 
    89, 0, 42, 18, 0, 26, 19, 35, 39, 0, 56, 61, 0, 17, 18, 
    87, 0, 1, 44, 0, 0, 9, 26, 60, 0, 69, 41, 0, 0, 23, 
    65, 0, 42, 11, 0, 0, 58, 0, 30, 0, 32, 45, 0, 0, 0, 
    52, 0, 101, 0, 34, 0, 16, 0, 0, 0, 0, 43, 0, 0, 0, 
    0, 0, 89, 0, 67, 4, 0, 5, 19, 16, 35, 5, 0, 0, 6, 
    0, 0, 75, 0, 75, 62, 0, 6, 66, 19, 0, 0, 0, 0, 12, 
    0, 0, 34, 0, 113, 53, 0, 0, 14, 0, 0, 0, 0, 0, 4, 
    10, 0, 0, 0, 123, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 0, 0, 20, 37, 0, 7, 1, 0, 0, 0, 0, 0, 0, 8, 
    25, 0, 0, 0, 11, 0, 0, 0, 0, 0, 11, 0, 0, 9, 44, 
    
    -- channel=8
    293, 295, 297, 305, 299, 293, 309, 307, 294, 276, 246, 244, 255, 259, 242, 
    291, 298, 304, 313, 307, 386, 331, 291, 219, 209, 231, 197, 187, 233, 258, 
    250, 246, 309, 306, 306, 314, 249, 162, 155, 250, 286, 234, 201, 158, 236, 
    242, 216, 319, 310, 307, 257, 305, 210, 189, 239, 299, 211, 167, 119, 175, 
    339, 378, 348, 319, 510, 393, 338, 221, 155, 178, 342, 251, 193, 157, 111, 
    342, 414, 370, 247, 341, 358, 402, 274, 195, 268, 402, 233, 202, 194, 147, 
    349, 403, 299, 267, 248, 371, 456, 341, 245, 311, 363, 231, 185, 222, 226, 
    401, 413, 299, 312, 261, 445, 379, 273, 236, 296, 332, 226, 185, 239, 226, 
    453, 442, 318, 309, 294, 234, 260, 253, 255, 272, 240, 158, 119, 214, 287, 
    441, 436, 358, 282, 327, 210, 271, 385, 263, 239, 160, 80, 174, 291, 302, 
    406, 438, 352, 398, 547, 380, 381, 399, 292, 164, 134, 165, 198, 253, 245, 
    272, 386, 413, 560, 495, 210, 169, 164, 166, 159, 171, 172, 190, 202, 196, 
    204, 232, 369, 569, 265, 178, 171, 159, 156, 161, 178, 206, 216, 204, 241, 
    198, 175, 270, 439, 211, 187, 186, 164, 159, 177, 182, 190, 179, 214, 229, 
    209, 166, 178, 200, 149, 143, 170, 178, 194, 211, 191, 169, 238, 289, 186, 
    
    -- channel=9
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 20, 136, 181, 156, 94, 0, 0, 
    17, 0, 0, 0, 0, 0, 0, 93, 134, 123, 71, 84, 118, 90, 0, 
    182, 106, 0, 0, 0, 0, 49, 94, 128, 100, 75, 75, 119, 114, 0, 
    261, 192, 0, 0, 99, 19, 45, 60, 107, 180, 114, 102, 135, 142, 109, 
    249, 212, 0, 0, 0, 33, 94, 80, 110, 202, 128, 130, 142, 160, 96, 
    249, 239, 76, 0, 0, 148, 126, 105, 75, 76, 105, 122, 165, 106, 0, 
    298, 311, 231, 133, 0, 57, 33, 100, 95, 0, 63, 85, 113, 0, 0, 
    249, 294, 241, 253, 159, 82, 91, 146, 139, 58, 98, 147, 105, 0, 0, 
    311, 240, 221, 318, 260, 270, 336, 313, 269, 207, 338, 412, 437, 334, 303, 
    612, 405, 257, 269, 331, 463, 488, 496, 537, 556, 613, 641, 678, 678, 683, 
    765, 580, 360, 298, 440, 593, 593, 578, 594, 636, 689, 713, 705, 717, 762, 
    811, 712, 571, 422, 525, 614, 607, 600, 624, 670, 725, 750, 749, 827, 793, 
    789, 774, 666, 544, 577, 629, 635, 614, 627, 666, 692, 700, 742, 806, 757, 
    
    -- channel=10
    242, 243, 248, 246, 248, 237, 252, 268, 262, 233, 210, 212, 216, 224, 231, 
    247, 253, 255, 251, 252, 193, 220, 235, 216, 149, 93, 110, 153, 203, 220, 
    201, 230, 254, 259, 264, 221, 183, 150, 129, 84, 53, 60, 73, 142, 190, 
    71, 130, 231, 259, 225, 191, 109, 93, 81, 114, 71, 102, 85, 94, 171, 
    30, 47, 188, 237, 75, 89, 69, 79, 79, 123, 68, 75, 80, 71, 135, 
    45, 34, 171, 241, 120, 118, 60, 74, 52, 116, 57, 77, 84, 71, 73, 
    42, 12, 159, 210, 143, 120, 67, 71, 56, 88, 51, 67, 78, 78, 73, 
    42, 0, 73, 134, 157, 95, 52, 90, 83, 114, 78, 67, 86, 87, 130, 
    14, 9, 30, 73, 125, 114, 97, 85, 86, 115, 130, 92, 104, 122, 188, 
    42, 23, 6, 45, 54, 107, 94, 33, 71, 126, 87, 92, 84, 168, 209, 
    33, 36, 10, 51, 0, 16, 41, 22, 23, 47, 28, 11, 3, 30, 45, 
    0, 12, 16, 37, 8, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 41, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=11
    168, 178, 169, 175, 174, 163, 181, 185, 174, 165, 149, 142, 143, 150, 146, 
    164, 171, 177, 183, 171, 173, 185, 173, 161, 87, 89, 86, 93, 124, 144, 
    164, 139, 173, 180, 176, 230, 162, 91, 47, 91, 137, 109, 115, 73, 126, 
    134, 43, 172, 177, 178, 112, 136, 95, 89, 104, 168, 117, 96, 60, 83, 
    155, 133, 193, 132, 203, 171, 184, 110, 96, 34, 151, 127, 83, 81, 52, 
    153, 181, 196, 164, 191, 190, 203, 137, 110, 36, 218, 134, 91, 94, 52, 
    131, 229, 146, 181, 142, 139, 249, 162, 145, 108, 198, 108, 76, 79, 100, 
    159, 203, 123, 147, 118, 201, 238, 169, 118, 142, 185, 122, 79, 120, 123, 
    204, 198, 152, 131, 121, 154, 134, 118, 88, 170, 119, 129, 54, 98, 147, 
    212, 201, 192, 107, 152, 96, 100, 172, 113, 150, 132, 40, 51, 141, 175, 
    162, 194, 198, 76, 229, 124, 159, 224, 155, 81, 11, 22, 57, 91, 85, 
    117, 165, 175, 226, 336, 114, 79, 73, 54, 44, 46, 47, 44, 58, 53, 
    56, 88, 104, 305, 162, 51, 57, 49, 42, 33, 36, 42, 71, 62, 44, 
    55, 41, 70, 283, 79, 53, 54, 47, 44, 45, 51, 58, 51, 27, 106, 
    69, 39, 55, 111, 53, 41, 62, 54, 51, 56, 57, 38, 34, 96, 66, 
    
    -- channel=12
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=13
    77, 71, 70, 67, 66, 68, 70, 65, 58, 76, 89, 90, 73, 59, 51, 
    65, 58, 68, 67, 72, 82, 49, 70, 79, 84, 66, 66, 93, 92, 63, 
    83, 140, 70, 62, 71, 137, 75, 61, 65, 142, 114, 109, 70, 96, 95, 
    10, 117, 70, 70, 58, 86, 72, 78, 99, 182, 107, 108, 83, 60, 128, 
    77, 147, 69, 117, 108, 97, 97, 74, 88, 152, 102, 59, 93, 52, 90, 
    136, 208, 80, 80, 250, 163, 111, 76, 41, 213, 141, 89, 120, 84, 50, 
    123, 165, 125, 27, 170, 166, 179, 119, 64, 236, 120, 75, 102, 107, 84, 
    146, 153, 99, 68, 118, 235, 168, 158, 96, 195, 135, 77, 124, 135, 96, 
    170, 210, 93, 167, 88, 164, 99, 91, 136, 87, 127, 99, 110, 107, 79, 
    213, 212, 98, 175, 101, 124, 148, 101, 113, 145, 105, 72, 115, 116, 87, 
    250, 195, 111, 243, 102, 86, 224, 227, 135, 80, 78, 101, 142, 168, 134, 
    290, 272, 164, 284, 209, 172, 170, 164, 146, 146, 160, 166, 168, 173, 164, 
    175, 256, 266, 247, 144, 152, 148, 149, 145, 150, 164, 171, 188, 192, 191, 
    176, 172, 299, 243, 151, 165, 142, 143, 157, 165, 180, 192, 179, 198, 222, 
    171, 176, 182, 193, 150, 178, 188, 166, 161, 160, 155, 169, 191, 183, 147, 
    
    -- channel=14
    0, 0, 0, 0, 0, 0, 0, 0, 8, 10, 6, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 23, 8, 24, 0, 6, 0, 0, 0, 0, 
    28, 0, 0, 0, 0, 0, 51, 12, 0, 0, 8, 3, 26, 0, 0, 
    84, 0, 0, 0, 21, 0, 5, 20, 0, 0, 42, 0, 29, 14, 0, 
    84, 0, 26, 0, 0, 0, 34, 34, 13, 0, 0, 47, 0, 31, 0, 
    57, 0, 37, 4, 0, 10, 37, 26, 48, 0, 53, 62, 0, 16, 10, 
    52, 8, 0, 53, 0, 0, 6, 31, 57, 0, 68, 35, 0, 0, 11, 
    38, 13, 17, 16, 0, 0, 73, 1, 29, 0, 42, 40, 0, 0, 0, 
    43, 0, 92, 0, 17, 0, 12, 2, 0, 3, 0, 55, 0, 0, 0, 
    2, 0, 98, 0, 35, 0, 0, 4, 0, 14, 52, 0, 0, 0, 11, 
    0, 0, 82, 0, 94, 20, 0, 12, 72, 31, 0, 0, 0, 0, 15, 
    0, 0, 18, 0, 114, 60, 0, 0, 8, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 133, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 72, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 
    
    -- channel=15
    205, 218, 219, 220, 213, 218, 218, 217, 211, 187, 164, 178, 193, 179, 171, 
    215, 220, 224, 221, 235, 365, 195, 196, 131, 207, 192, 135, 135, 183, 185, 
    144, 205, 224, 220, 223, 232, 164, 101, 137, 288, 222, 200, 132, 107, 208, 
    118, 246, 218, 235, 215, 230, 254, 152, 159, 255, 218, 160, 132, 74, 185, 
    236, 358, 197, 307, 454, 281, 229, 157, 110, 256, 283, 153, 180, 115, 71, 
    203, 379, 212, 160, 383, 277, 333, 201, 124, 413, 255, 135, 189, 157, 111, 
    230, 316, 202, 164, 277, 387, 362, 259, 154, 406, 235, 161, 171, 228, 161, 
    292, 355, 178, 226, 249, 434, 211, 209, 179, 328, 261, 146, 188, 193, 177, 
    347, 391, 169, 327, 193, 185, 207, 227, 249, 172, 213, 70, 123, 218, 227, 
    395, 382, 230, 323, 209, 143, 282, 340, 161, 176, 80, 79, 196, 259, 208, 
    452, 369, 222, 529, 444, 280, 356, 312, 184, 117, 149, 189, 193, 217, 188, 
    270, 385, 336, 586, 273, 145, 160, 155, 162, 165, 183, 188, 214, 214, 201, 
    185, 237, 411, 449, 124, 190, 170, 169, 171, 185, 210, 227, 216, 218, 277, 
    192, 186, 302, 332, 189, 201, 186, 168, 180, 197, 196, 204, 197, 263, 186, 
    186, 197, 183, 182, 137, 167, 183, 191, 220, 230, 186, 196, 309, 271, 154, 
    
    -- channel=16
    216, 226, 225, 224, 214, 228, 229, 212, 203, 199, 187, 192, 201, 188, 160, 
    205, 220, 229, 228, 234, 345, 251, 217, 177, 209, 232, 179, 158, 180, 177, 
    180, 194, 221, 219, 221, 282, 223, 136, 152, 317, 339, 278, 202, 131, 195, 
    195, 199, 235, 228, 229, 232, 305, 224, 209, 319, 336, 248, 190, 106, 165, 
    387, 420, 281, 320, 544, 453, 387, 247, 166, 265, 393, 264, 214, 150, 95, 
    438, 507, 324, 248, 490, 479, 468, 299, 179, 391, 464, 261, 237, 215, 149, 
    458, 485, 287, 191, 303, 467, 533, 392, 253, 438, 425, 257, 219, 270, 234, 
    531, 520, 324, 265, 291, 559, 441, 339, 255, 383, 402, 249, 237, 278, 223, 
    594, 591, 377, 389, 306, 315, 299, 281, 293, 267, 276, 169, 150, 230, 250, 
    582, 585, 420, 407, 370, 250, 351, 443, 297, 273, 165, 95, 192, 268, 241, 
    552, 570, 417, 578, 648, 433, 510, 524, 349, 185, 170, 228, 273, 299, 272, 
    425, 555, 524, 742, 621, 328, 291, 286, 269, 253, 276, 293, 321, 336, 326, 
    326, 381, 553, 710, 359, 296, 284, 268, 260, 271, 304, 337, 352, 351, 394, 
    337, 306, 463, 549, 307, 309, 298, 275, 283, 307, 320, 334, 322, 373, 376, 
    348, 318, 320, 301, 236, 260, 292, 296, 324, 344, 316, 304, 406, 442, 305, 
    
    -- channel=17
    186, 201, 194, 205, 197, 191, 201, 204, 203, 194, 170, 158, 167, 169, 165, 
    189, 196, 199, 211, 200, 262, 221, 208, 160, 122, 141, 106, 93, 139, 171, 
    196, 137, 199, 204, 197, 202, 182, 85, 81, 127, 193, 153, 139, 68, 141, 
    195, 67, 195, 203, 222, 146, 208, 144, 121, 107, 221, 132, 119, 77, 63, 
    253, 207, 228, 173, 362, 245, 237, 160, 108, 39, 214, 182, 119, 120, 29, 
    223, 253, 248, 163, 198, 232, 293, 185, 153, 87, 290, 173, 115, 134, 88, 
    219, 279, 169, 218, 127, 219, 324, 234, 194, 126, 260, 157, 96, 126, 147, 
    261, 279, 170, 203, 136, 285, 289, 178, 167, 145, 238, 155, 99, 143, 139, 
    311, 272, 235, 181, 187, 118, 157, 170, 133, 150, 146, 129, 47, 112, 178, 
    297, 269, 283, 119, 231, 126, 137, 263, 150, 186, 134, 42, 80, 170, 207, 
    229, 269, 261, 174, 415, 258, 246, 290, 236, 105, 62, 93, 105, 128, 137, 
    114, 225, 270, 311, 384, 135, 68, 67, 93, 85, 92, 87, 95, 102, 111, 
    113, 85, 172, 393, 217, 99, 96, 83, 82, 82, 89, 108, 125, 115, 125, 
    119, 83, 82, 352, 148, 96, 106, 87, 85, 94, 95, 102, 94, 110, 141, 
    131, 87, 77, 100, 80, 68, 99, 104, 107, 114, 107, 79, 112, 180, 123, 
    
    -- channel=18
    84, 67, 76, 80, 82, 67, 75, 75, 78, 83, 76, 72, 70, 82, 88, 
    85, 64, 78, 77, 79, 65, 76, 60, 55, 68, 89, 88, 82, 82, 88, 
    78, 76, 75, 73, 83, 71, 48, 70, 94, 102, 104, 105, 115, 111, 79, 
    95, 127, 78, 73, 63, 66, 85, 111, 116, 111, 74, 96, 92, 121, 103, 
    80, 129, 81, 75, 57, 75, 57, 86, 109, 96, 79, 95, 111, 118, 125, 
    75, 86, 63, 57, 21, 22, 48, 92, 111, 119, 69, 76, 113, 111, 115, 
    66, 81, 62, 56, 97, 56, 63, 68, 96, 114, 57, 91, 108, 105, 120, 
    50, 56, 107, 68, 114, 88, 65, 76, 87, 113, 64, 88, 109, 107, 101, 
    49, 61, 75, 78, 82, 62, 67, 93, 109, 80, 80, 83, 106, 103, 102, 
    50, 72, 66, 87, 81, 97, 74, 81, 116, 82, 93, 107, 131, 108, 85, 
    63, 56, 63, 99, 69, 120, 105, 61, 86, 100, 126, 134, 133, 103, 90, 
    131, 59, 76, 96, 36, 53, 86, 86, 111, 132, 142, 139, 138, 147, 140, 
    168, 128, 67, 57, 56, 129, 134, 136, 145, 151, 153, 154, 151, 140, 147, 
    157, 145, 125, 53, 118, 141, 137, 139, 138, 143, 151, 148, 144, 158, 153, 
    153, 147, 136, 117, 145, 145, 144, 139, 143, 143, 151, 152, 153, 158, 154, 
    
    -- channel=19
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 35, 21, 70, 51, 3, 0, 0, 
    29, 0, 0, 0, 0, 3, 50, 51, 26, 25, 114, 93, 109, 0, 0, 
    174, 0, 0, 0, 0, 0, 75, 85, 74, 0, 132, 76, 108, 67, 0, 
    184, 20, 0, 0, 95, 87, 148, 115, 103, 0, 98, 128, 71, 110, 0, 
    148, 67, 19, 0, 30, 82, 142, 116, 150, 0, 154, 138, 58, 101, 79, 
    130, 165, 0, 58, 0, 0, 133, 113, 166, 0, 168, 118, 61, 55, 80, 
    130, 179, 64, 54, 0, 26, 181, 91, 100, 0, 123, 131, 49, 61, 23, 
    170, 128, 178, 40, 50, 68, 85, 87, 14, 82, 42, 136, 36, 0, 0, 
    126, 115, 223, 47, 135, 51, 26, 144, 72, 76, 139, 79, 11, 0, 0, 
    59, 112, 218, 0, 223, 130, 75, 169, 182, 137, 93, 99, 101, 76, 96, 
    85, 90, 136, 14, 295, 186, 143, 143, 148, 139, 143, 153, 158, 159, 174, 
    183, 72, 0, 178, 268, 155, 165, 151, 151, 147, 153, 157, 172, 172, 159, 
    209, 159, 0, 269, 167, 148, 169, 157, 155, 161, 171, 172, 182, 151, 214, 
    222, 180, 144, 173, 153, 130, 147, 153, 150, 167, 184, 156, 127, 224, 234, 
    
    -- channel=20
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 66, 0, 0, 0, 8, 0, 
    0, 73, 0, 0, 0, 0, 0, 0, 5, 89, 0, 0, 0, 0, 24, 
    0, 44, 0, 0, 0, 0, 0, 0, 0, 106, 0, 0, 5, 0, 52, 
    0, 0, 0, 0, 19, 0, 0, 0, 0, 218, 0, 0, 21, 0, 0, 
    0, 0, 0, 0, 54, 23, 0, 0, 0, 182, 0, 0, 21, 24, 0, 
    0, 0, 0, 0, 32, 69, 0, 0, 0, 97, 0, 0, 42, 9, 0, 
    0, 5, 0, 10, 0, 0, 0, 0, 14, 0, 5, 0, 40, 0, 0, 
    0, 3, 0, 88, 0, 17, 16, 0, 17, 0, 0, 13, 53, 0, 0, 
    68, 0, 0, 185, 0, 6, 109, 0, 0, 0, 65, 97, 101, 64, 27, 
    170, 51, 0, 133, 0, 0, 69, 66, 55, 95, 107, 116, 116, 116, 101, 
    114, 172, 98, 0, 0, 90, 90, 94, 96, 114, 126, 131, 116, 119, 130, 
    97, 127, 249, 0, 29, 106, 80, 99, 110, 119, 128, 124, 111, 173, 114, 
    88, 131, 132, 42, 83, 125, 104, 91, 113, 107, 100, 120, 161, 106, 52, 
    
    -- channel=21
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 26, 29, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 16, 17, 14, 16, 6, 11, 
    19, 0, 0, 0, 0, 14, 13, 14, 18, 21, 19, 14, 3, 7, 11, 
    21, 18, 0, 0, 10, 7, 17, 14, 16, 14, 13, 7, 19, 14, 0, 
    19, 21, 7, 0, 15, 9, 5, 14, 13, 13, 14, 17, 9, 0, 28, 
    
    -- channel=22
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 7, 0, 0, 10, 10, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 11, 2, 0, 0, 0, 12, 0, 0, 0, 8, 0, 0, 0, 0, 
    0, 4, 0, 0, 0, 12, 14, 7, 0, 0, 5, 0, 0, 5, 0, 
    4, 11, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 12, 5, 0, 5, 0, 0, 0, 0, 7, 6, 0, 0, 0, 0, 
    10, 6, 8, 0, 0, 0, 15, 27, 16, 0, 0, 0, 0, 0, 0, 
    33, 25, 17, 4, 43, 18, 8, 9, 9, 7, 11, 11, 11, 13, 14, 
    20, 23, 9, 21, 14, 8, 12, 9, 8, 7, 9, 8, 20, 20, 8, 
    22, 15, 20, 36, 12, 9, 8, 9, 12, 11, 16, 21, 18, 9, 40, 
    22, 17, 21, 20, 12, 15, 22, 14, 11, 7, 15, 13, 7, 16, 25, 
    
    -- channel=23
    295, 309, 307, 309, 306, 294, 317, 338, 315, 267, 241, 249, 262, 276, 277, 
    304, 320, 315, 318, 306, 279, 273, 285, 234, 143, 93, 106, 156, 230, 269, 
    241, 257, 319, 326, 321, 262, 210, 129, 103, 77, 70, 69, 84, 127, 233, 
    107, 135, 290, 314, 284, 194, 140, 94, 82, 84, 114, 99, 86, 91, 168, 
    49, 87, 250, 215, 160, 119, 111, 97, 86, 71, 88, 94, 83, 82, 111, 
    25, 80, 246, 255, 132, 126, 128, 92, 87, 71, 100, 88, 76, 71, 72, 
    21, 72, 184, 274, 146, 131, 116, 105, 86, 64, 81, 74, 66, 66, 93, 
    39, 43, 63, 176, 136, 116, 106, 98, 111, 119, 107, 76, 66, 103, 170, 
    32, 19, 49, 87, 131, 95, 105, 97, 81, 132, 120, 103, 88, 146, 235, 
    69, 35, 52, 16, 67, 97, 77, 78, 72, 135, 97, 56, 84, 209, 252, 
    35, 47, 48, 18, 45, 18, 37, 41, 42, 25, 0, 0, 0, 0, 0, 
    0, 0, 31, 54, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=24
    159, 158, 156, 162, 163, 151, 165, 169, 168, 162, 146, 135, 134, 141, 139, 
    158, 151, 157, 169, 155, 159, 187, 167, 152, 105, 117, 118, 115, 120, 138, 
    176, 118, 163, 167, 169, 209, 188, 128, 74, 83, 154, 113, 126, 94, 110, 
    165, 61, 168, 161, 183, 119, 147, 113, 106, 91, 184, 134, 120, 91, 64, 
    176, 129, 194, 101, 168, 164, 199, 140, 118, 39, 166, 151, 96, 93, 72, 
    214, 194, 206, 194, 190, 194, 213, 148, 135, 20, 244, 167, 98, 104, 72, 
    191, 246, 170, 174, 112, 154, 239, 183, 158, 83, 233, 149, 103, 99, 121, 
    217, 208, 160, 160, 100, 169, 251, 178, 141, 123, 207, 165, 90, 131, 123, 
    246, 212, 225, 127, 178, 165, 168, 149, 94, 192, 156, 150, 78, 91, 132, 
    239, 222, 236, 112, 184, 114, 106, 175, 161, 151, 137, 53, 44, 123, 174, 
    175, 223, 243, 75, 240, 151, 145, 215, 172, 109, 56, 48, 87, 134, 145, 
    148, 177, 185, 207, 394, 208, 147, 140, 115, 90, 90, 94, 95, 112, 114, 
    126, 130, 131, 335, 244, 95, 96, 92, 92, 85, 86, 95, 115, 108, 99, 
    124, 96, 109, 306, 136, 96, 106, 92, 84, 90, 108, 114, 108, 94, 163, 
    133, 91, 117, 156, 117, 94, 101, 90, 86, 104, 115, 90, 77, 154, 126, 
    
    -- channel=25
    132, 159, 154, 146, 135, 161, 157, 148, 135, 119, 116, 132, 145, 133, 112, 
    137, 172, 164, 149, 156, 222, 146, 152, 113, 118, 103, 82, 88, 118, 118, 
    97, 127, 146, 150, 139, 131, 90, 55, 86, 158, 112, 100, 61, 60, 137, 
    58, 122, 137, 158, 140, 136, 150, 85, 65, 149, 108, 92, 51, 28, 124, 
    117, 196, 124, 215, 310, 229, 155, 91, 44, 149, 161, 93, 87, 52, 53, 
    93, 180, 139, 114, 225, 211, 194, 117, 48, 241, 133, 63, 94, 73, 70, 
    123, 142, 125, 118, 173, 223, 201, 136, 79, 220, 109, 73, 73, 108, 77, 
    168, 182, 101, 127, 152, 264, 99, 101, 84, 171, 118, 56, 97, 100, 91, 
    179, 205, 65, 174, 102, 104, 99, 98, 129, 76, 106, 21, 59, 117, 148, 
    179, 182, 93, 170, 129, 98, 161, 181, 83, 100, 27, 45, 120, 159, 124, 
    207, 189, 86, 285, 222, 166, 208, 165, 94, 40, 47, 79, 65, 50, 30, 
    68, 171, 176, 301, 82, 0, 20, 20, 15, 15, 15, 19, 26, 19, 16, 
    0, 57, 196, 196, 0, 37, 32, 22, 7, 9, 17, 28, 26, 26, 46, 
    0, 11, 131, 76, 12, 32, 21, 25, 31, 28, 4, 1, 0, 27, 0, 
    0, 12, 12, 0, 0, 0, 10, 27, 50, 38, 6, 6, 72, 30, 0, 
    
    -- channel=26
    14, 15, 18, 7, 9, 20, 17, 12, 10, 13, 12, 26, 15, 4, 0, 
    17, 21, 26, 6, 25, 28, 0, 13, 4, 32, 0, 0, 34, 35, 1, 
    0, 71, 14, 8, 23, 66, 0, 0, 16, 86, 0, 0, 0, 41, 42, 
    0, 117, 9, 30, 0, 35, 0, 0, 0, 131, 0, 4, 0, 0, 119, 
    0, 71, 0, 121, 0, 0, 0, 0, 0, 143, 0, 0, 0, 0, 57, 
    0, 30, 0, 16, 146, 0, 0, 0, 0, 258, 0, 0, 28, 0, 0, 
    0, 0, 6, 0, 146, 76, 0, 0, 0, 231, 0, 0, 10, 24, 0, 
    0, 0, 0, 0, 91, 132, 0, 0, 0, 147, 0, 0, 45, 9, 0, 
    0, 18, 0, 63, 0, 39, 0, 0, 47, 0, 49, 0, 34, 36, 28, 
    0, 9, 0, 113, 0, 0, 54, 0, 0, 0, 0, 7, 73, 72, 1, 
    114, 1, 0, 214, 0, 0, 82, 0, 0, 0, 4, 15, 30, 40, 0, 
    135, 58, 0, 179, 0, 0, 17, 10, 0, 0, 0, 2, 0, 0, 0, 
    0, 113, 110, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 200, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 
    0, 0, 11, 7, 0, 18, 1, 0, 1, 0, 0, 0, 39, 0, 0, 
    
    -- channel=27
    324, 349, 346, 348, 336, 339, 358, 365, 338, 295, 265, 276, 300, 298, 281, 
    329, 363, 359, 358, 355, 419, 341, 324, 256, 200, 175, 141, 163, 251, 287, 
    243, 290, 354, 359, 348, 328, 244, 133, 124, 216, 201, 176, 134, 111, 267, 
    174, 170, 337, 360, 326, 273, 270, 156, 128, 195, 244, 158, 120, 54, 188, 
    255, 288, 331, 356, 498, 356, 283, 168, 97, 158, 274, 186, 144, 108, 64, 
    206, 307, 351, 257, 320, 339, 357, 220, 129, 236, 304, 167, 148, 141, 97, 
    226, 283, 261, 315, 252, 334, 380, 280, 181, 260, 267, 152, 119, 161, 156, 
    280, 324, 183, 293, 244, 385, 295, 210, 188, 253, 263, 142, 130, 181, 211, 
    324, 325, 181, 255, 217, 194, 200, 184, 196, 218, 172, 114, 82, 197, 290, 
    342, 312, 239, 208, 222, 164, 238, 314, 148, 202, 123, 49, 141, 292, 311, 
    310, 323, 236, 320, 431, 245, 287, 305, 199, 94, 31, 63, 57, 99, 92, 
    74, 273, 312, 446, 307, 46, 17, 12, 8, 6, 3, 2, 10, 7, 6, 
    0, 45, 261, 402, 104, 25, 17, 6, 0, 0, 0, 9, 22, 19, 36, 
    0, 0, 93, 286, 58, 22, 18, 1, 6, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 23, 0, 0, 4, 24, 38, 32, 0, 0, 50, 50, 0, 
    
    -- channel=28
    43, 53, 46, 53, 48, 54, 44, 32, 41, 62, 69, 59, 64, 50, 43, 
    45, 41, 43, 53, 50, 147, 87, 67, 69, 109, 165, 112, 64, 56, 57, 
    79, 44, 40, 43, 30, 65, 110, 74, 86, 164, 216, 201, 170, 54, 69, 
    208, 66, 58, 44, 84, 92, 187, 156, 154, 114, 232, 135, 155, 98, 37, 
    316, 231, 122, 76, 343, 236, 240, 176, 136, 82, 232, 196, 154, 161, 26, 
    259, 280, 153, 15, 170, 211, 294, 205, 192, 104, 284, 197, 147, 178, 139, 
    268, 306, 117, 99, 99, 194, 304, 250, 223, 154, 283, 187, 140, 165, 168, 
    291, 348, 192, 177, 100, 242, 292, 183, 183, 123, 245, 181, 134, 153, 117, 
    351, 331, 267, 215, 147, 132, 167, 177, 165, 144, 104, 149, 79, 106, 81, 
    318, 310, 333, 203, 242, 132, 178, 300, 156, 153, 167, 101, 127, 100, 96, 
    285, 299, 316, 228, 490, 300, 276, 333, 296, 194, 170, 211, 217, 222, 217, 
    235, 310, 334, 323, 392, 243, 196, 198, 231, 230, 251, 256, 279, 277, 285, 
    310, 204, 254, 381, 319, 257, 253, 241, 241, 250, 276, 291, 298, 298, 330, 
    329, 275, 172, 425, 270, 260, 272, 244, 250, 268, 280, 286, 296, 306, 321, 
    335, 290, 248, 250, 224, 217, 251, 266, 273, 294, 284, 269, 309, 376, 334, 
    
    -- channel=29
    175, 188, 182, 181, 169, 194, 181, 160, 153, 168, 165, 171, 174, 146, 121, 
    161, 180, 187, 183, 200, 344, 187, 177, 150, 220, 240, 171, 150, 166, 149, 
    146, 197, 178, 169, 178, 290, 163, 111, 160, 403, 364, 303, 205, 136, 194, 
    164, 247, 191, 190, 181, 237, 321, 232, 236, 407, 328, 263, 191, 94, 204, 
    380, 499, 218, 346, 602, 467, 376, 233, 177, 335, 412, 246, 247, 154, 104, 
    421, 564, 250, 206, 562, 462, 463, 300, 173, 544, 453, 231, 283, 237, 150, 
    431, 518, 247, 137, 388, 508, 576, 393, 246, 598, 400, 245, 248, 315, 238, 
    517, 561, 298, 257, 345, 676, 426, 353, 252, 481, 396, 232, 285, 314, 205, 
    603, 659, 326, 445, 286, 334, 285, 300, 337, 262, 298, 146, 182, 246, 234, 
    627, 642, 392, 502, 362, 256, 395, 492, 298, 283, 164, 119, 257, 293, 210, 
    675, 616, 398, 738, 654, 467, 625, 586, 352, 205, 223, 308, 346, 367, 311, 
    575, 656, 559, 905, 611, 321, 347, 338, 320, 338, 372, 395, 429, 439, 421, 
    421, 506, 645, 780, 326, 380, 369, 352, 347, 370, 416, 451, 463, 465, 520, 
    433, 407, 609, 602, 362, 407, 377, 360, 380, 411, 429, 446, 426, 509, 488, 
    440, 429, 408, 392, 312, 358, 392, 390, 429, 447, 409, 410, 550, 562, 379, 
    
    -- channel=30
    0, 4, 0, 2, 0, 0, 0, 3, 13, 24, 21, 0, 0, 13, 29, 
    0, 0, 0, 13, 0, 0, 78, 31, 89, 0, 36, 19, 0, 0, 10, 
    91, 0, 0, 8, 0, 3, 135, 65, 0, 0, 57, 27, 123, 0, 0, 
    343, 0, 0, 0, 64, 0, 54, 45, 8, 0, 166, 5, 103, 48, 0, 
    265, 0, 99, 0, 43, 0, 174, 115, 81, 0, 43, 166, 0, 126, 0, 
    116, 0, 127, 0, 0, 0, 168, 119, 226, 0, 187, 194, 0, 66, 40, 
    72, 147, 0, 213, 0, 0, 96, 106, 249, 0, 241, 121, 0, 0, 58, 
    38, 140, 20, 121, 0, 0, 262, 32, 118, 0, 130, 162, 0, 0, 12, 
    105, 0, 245, 0, 5, 0, 71, 31, 0, 109, 0, 201, 0, 0, 0, 
    10, 0, 340, 0, 141, 0, 0, 109, 0, 28, 200, 5, 0, 0, 37, 
    0, 0, 325, 0, 291, 46, 0, 79, 218, 120, 0, 0, 0, 0, 19, 
    0, 0, 64, 0, 426, 160, 0, 0, 14, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 81, 387, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    42, 0, 0, 345, 74, 0, 12, 0, 0, 0, 0, 0, 0, 0, 41, 
    74, 0, 0, 49, 16, 0, 0, 0, 0, 0, 7, 0, 0, 36, 146, 
    
    -- channel=31
    28, 22, 24, 22, 24, 19, 29, 30, 21, 22, 24, 26, 23, 28, 29, 
    27, 25, 26, 23, 21, 0, 14, 18, 22, 0, 0, 9, 26, 34, 28, 
    17, 47, 26, 24, 26, 8, 0, 10, 9, 0, 0, 0, 0, 37, 31, 
    0, 30, 29, 21, 5, 0, 0, 0, 0, 0, 0, 0, 0, 18, 51, 
    0, 0, 11, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 42, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 11, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 12, 21, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 19, 27, 19, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=32
    187, 199, 195, 196, 195, 189, 204, 220, 206, 171, 152, 156, 167, 176, 178, 
    186, 211, 204, 203, 197, 144, 193, 187, 168, 85, 40, 63, 95, 133, 165, 
    148, 147, 204, 211, 204, 190, 150, 113, 59, 12, 23, 21, 27, 59, 125, 
    77, 17, 181, 205, 184, 134, 75, 41, 13, 18, 62, 49, 42, 19, 73, 
    36, 0, 165, 151, 75, 86, 88, 55, 31, 10, 54, 56, 24, 22, 44, 
    36, 0, 163, 179, 65, 112, 73, 65, 35, 0, 68, 67, 21, 25, 18, 
    39, 2, 111, 205, 65, 51, 61, 60, 52, 0, 66, 41, 16, 8, 27, 
    31, 24, 30, 115, 71, 21, 88, 56, 57, 28, 55, 51, 11, 33, 88, 
    21, 0, 32, 1, 79, 80, 72, 36, 12, 102, 61, 76, 29, 53, 120, 
    28, 1, 29, 0, 40, 57, 42, 26, 27, 70, 57, 23, 0, 93, 162, 
    0, 23, 42, 0, 0, 0, 0, 12, 7, 15, 0, 0, 0, 0, 0, 
    0, 0, 10, 0, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=33
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=34
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 0, 0, 0, 33, 0, 0, 0, 4, 0, 0, 0, 3, 0, 
    0, 12, 0, 0, 0, 31, 0, 0, 0, 37, 0, 0, 0, 0, 20, 
    0, 35, 0, 0, 1, 0, 8, 0, 0, 31, 0, 0, 0, 0, 33, 
    0, 51, 0, 0, 25, 0, 0, 0, 0, 16, 0, 0, 4, 0, 0, 
    0, 30, 0, 0, 62, 0, 1, 0, 0, 79, 0, 0, 7, 0, 0, 
    0, 41, 0, 0, 65, 17, 22, 0, 0, 96, 0, 0, 0, 7, 0, 
    0, 11, 0, 0, 14, 61, 0, 0, 0, 63, 0, 0, 7, 5, 0, 
    0, 10, 0, 39, 0, 0, 0, 12, 1, 3, 15, 0, 2, 13, 5, 
    0, 1, 0, 43, 0, 0, 0, 28, 0, 0, 0, 0, 30, 36, 0, 
    72, 0, 0, 61, 0, 0, 33, 2, 0, 0, 0, 5, 9, 6, 0, 
    43, 19, 0, 94, 0, 0, 0, 0, 0, 0, 1, 2, 2, 5, 0, 
    0, 28, 0, 46, 0, 0, 0, 0, 0, 1, 5, 3, 5, 0, 1, 
    0, 1, 25, 23, 0, 0, 0, 0, 1, 2, 1, 4, 0, 8, 5, 
    0, 5, 6, 17, 0, 5, 2, 0, 6, 3, 0, 0, 17, 4, 0, 
    
    -- channel=35
    395, 419, 419, 418, 411, 404, 436, 456, 421, 346, 299, 325, 353, 369, 364, 
    409, 449, 436, 429, 423, 445, 378, 382, 275, 206, 136, 152, 210, 304, 356, 
    288, 335, 434, 442, 433, 368, 245, 166, 137, 157, 91, 87, 83, 148, 321, 
    125, 231, 402, 437, 387, 285, 222, 97, 77, 138, 133, 111, 75, 65, 246, 
    48, 197, 330, 348, 330, 212, 166, 112, 75, 134, 166, 104, 113, 75, 123, 
    0, 145, 316, 296, 228, 174, 211, 138, 95, 203, 117, 69, 103, 74, 76, 
    1, 114, 239, 360, 243, 234, 191, 136, 96, 185, 86, 80, 81, 101, 103, 
    41, 118, 72, 267, 205, 232, 91, 111, 119, 218, 116, 77, 85, 121, 203, 
    51, 90, 0, 155, 155, 114, 141, 141, 129, 187, 162, 61, 92, 207, 331, 
    111, 81, 36, 94, 88, 97, 144, 169, 78, 134, 53, 43, 123, 313, 331, 
    126, 104, 41, 179, 100, 60, 75, 52, 0, 13, 0, 0, 0, 0, 0, 
    0, 23, 62, 212, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 39, 133, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=36
    37, 37, 37, 37, 37, 34, 38, 42, 42, 41, 38, 38, 33, 39, 44, 
    37, 38, 37, 37, 34, 1, 32, 42, 35, 14, 2, 19, 30, 35, 42, 
    47, 28, 37, 38, 37, 12, 18, 23, 29, 0, 0, 0, 9, 34, 30, 
    16, 11, 34, 36, 36, 14, 2, 16, 7, 0, 0, 7, 9, 34, 26, 
    0, 0, 20, 12, 0, 0, 0, 9, 17, 0, 0, 5, 9, 22, 40, 
    0, 0, 11, 23, 0, 0, 0, 0, 13, 0, 0, 0, 5, 6, 19, 
    0, 0, 8, 42, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 6, 1, 0, 0, 0, 1, 0, 0, 0, 6, 0, 15, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 17, 18, 13, 8, 25, 
    0, 0, 0, 0, 0, 8, 0, 0, 0, 22, 13, 29, 13, 12, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=37
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 67, 40, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 8, 0, 0, 30, 63, 11, 8, 0, 0, 
    93, 61, 0, 0, 108, 26, 81, 16, 6, 0, 62, 12, 5, 0, 0, 
    88, 148, 0, 0, 154, 80, 106, 33, 13, 0, 111, 39, 21, 13, 0, 
    76, 161, 0, 0, 21, 38, 166, 64, 59, 62, 110, 21, 0, 16, 4, 
    103, 183, 3, 0, 0, 147, 138, 69, 38, 33, 82, 32, 16, 34, 0, 
    165, 188, 71, 79, 0, 48, 31, 20, 22, 0, 31, 27, 0, 0, 0, 
    178, 169, 138, 74, 95, 0, 28, 109, 13, 48, 32, 0, 0, 0, 0, 
    183, 151, 143, 102, 175, 76, 135, 213, 127, 17, 11, 33, 61, 75, 54, 
    202, 201, 155, 181, 262, 144, 115, 111, 109, 94, 114, 125, 140, 142, 146, 
    153, 149, 130, 251, 181, 120, 119, 107, 103, 108, 130, 145, 165, 163, 175, 
    181, 138, 134, 307, 120, 124, 118, 111, 119, 134, 147, 168, 156, 170, 212, 
    182, 160, 121, 182, 99, 115, 139, 128, 124, 140, 142, 134, 153, 212, 173, 
    
    -- channel=38
    315, 331, 324, 326, 316, 321, 341, 344, 314, 281, 256, 271, 280, 277, 258, 
    307, 339, 336, 335, 332, 372, 316, 306, 243, 200, 161, 161, 199, 250, 266, 
    252, 297, 334, 336, 335, 412, 243, 168, 118, 236, 223, 180, 129, 148, 264, 
    146, 198, 332, 337, 309, 261, 251, 140, 132, 263, 246, 190, 129, 60, 223, 
    203, 308, 315, 333, 415, 319, 300, 168, 124, 186, 289, 166, 154, 83, 105, 
    231, 372, 331, 270, 454, 355, 345, 218, 120, 281, 324, 175, 180, 132, 72, 
    228, 347, 295, 276, 315, 346, 422, 270, 180, 343, 287, 161, 146, 173, 156, 
    285, 363, 190, 277, 244, 448, 331, 269, 194, 342, 277, 174, 164, 222, 219, 
    343, 391, 182, 285, 218, 279, 242, 207, 213, 261, 255, 144, 129, 215, 277, 
    400, 384, 239, 272, 246, 170, 254, 308, 198, 233, 132, 54, 139, 294, 300, 
    399, 384, 265, 384, 324, 207, 307, 358, 184, 92, 41, 43, 90, 164, 133, 
    258, 355, 315, 530, 418, 151, 144, 135, 74, 58, 59, 69, 74, 86, 74, 
    36, 204, 330, 519, 173, 76, 69, 64, 51, 44, 54, 73, 93, 85, 100, 
    40, 46, 261, 390, 91, 86, 65, 60, 60, 67, 64, 77, 52, 72, 105, 
    54, 45, 67, 180, 48, 62, 79, 72, 80, 88, 63, 55, 108, 126, 20, 
    
    -- channel=39
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=40
    40, 47, 50, 51, 51, 48, 50, 55, 59, 46, 31, 30, 37, 39, 38, 
    51, 55, 55, 54, 53, 83, 60, 57, 23, 12, 12, 3, 1, 17, 37, 
    39, 11, 51, 53, 53, 23, 19, 0, 0, 6, 0, 0, 0, 0, 15, 
    13, 11, 39, 59, 65, 30, 34, 6, 0, 0, 10, 0, 0, 0, 0, 
    12, 27, 41, 54, 92, 66, 20, 5, 0, 0, 19, 12, 0, 0, 0, 
    2, 4, 38, 46, 0, 15, 36, 11, 0, 18, 27, 0, 0, 0, 0, 
    7, 7, 0, 44, 7, 41, 27, 21, 0, 10, 3, 0, 0, 0, 0, 
    26, 7, 12, 29, 17, 32, 11, 0, 0, 5, 4, 0, 0, 0, 0, 
    27, 11, 7, 0, 33, 0, 0, 10, 0, 14, 0, 0, 0, 0, 32, 
    11, 6, 3, 0, 0, 14, 8, 28, 6, 0, 0, 0, 0, 39, 48, 
    0, 17, 0, 25, 69, 42, 30, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=41
    286, 306, 310, 311, 301, 303, 316, 313, 302, 269, 229, 241, 263, 251, 233, 
    294, 316, 319, 318, 325, 476, 313, 299, 202, 221, 217, 153, 147, 220, 251, 
    226, 243, 315, 313, 314, 307, 219, 97, 128, 299, 264, 214, 154, 93, 246, 
    169, 231, 309, 329, 322, 274, 323, 181, 160, 257, 281, 180, 123, 47, 173, 
    300, 418, 310, 380, 624, 432, 323, 193, 104, 218, 345, 207, 180, 111, 52, 
    274, 438, 329, 259, 405, 372, 439, 245, 143, 407, 376, 166, 184, 164, 102, 
    296, 408, 244, 264, 295, 460, 484, 341, 191, 425, 314, 183, 156, 223, 180, 
    390, 434, 231, 297, 285, 545, 330, 248, 190, 361, 319, 160, 172, 214, 190, 
    463, 477, 244, 349, 274, 193, 219, 255, 247, 230, 216, 76, 79, 207, 296, 
    480, 461, 307, 325, 275, 188, 300, 424, 205, 221, 92, 29, 171, 325, 294, 
    489, 463, 290, 551, 612, 379, 459, 414, 246, 117, 97, 165, 179, 211, 188, 
    231, 424, 408, 718, 422, 100, 96, 90, 97, 108, 123, 127, 147, 154, 143, 
    123, 189, 424, 619, 130, 138, 121, 109, 102, 113, 137, 169, 172, 164, 218, 
    118, 116, 279, 415, 155, 146, 135, 109, 120, 138, 130, 131, 120, 191, 145, 
    133, 118, 121, 103, 65, 84, 117, 136, 173, 179, 127, 114, 245, 249, 87, 
    
    -- channel=42
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=43
    25, 26, 0, 0, 0, 5, 8, 12, 0, 46, 83, 65, 9, 0, 1, 
    0, 0, 0, 2, 0, 0, 0, 39, 150, 0, 0, 0, 67, 46, 0, 
    114, 130, 1, 1, 16, 227, 82, 78, 0, 0, 0, 0, 0, 75, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 97, 0, 64, 23, 1, 67, 
    0, 0, 0, 0, 0, 0, 0, 0, 44, 0, 0, 0, 0, 0, 59, 
    19, 0, 0, 146, 288, 97, 0, 0, 0, 0, 0, 35, 8, 0, 0, 
    0, 0, 80, 5, 104, 0, 28, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 46, 105, 131, 9, 46, 19, 5, 23, 51, 0, 
    0, 0, 0, 0, 0, 214, 29, 0, 0, 2, 164, 153, 85, 0, 0, 
    24, 0, 0, 0, 0, 18, 0, 0, 0, 171, 122, 35, 0, 0, 6, 
    10, 0, 0, 0, 0, 0, 0, 116, 0, 0, 0, 0, 0, 11, 11, 
    241, 85, 0, 0, 266, 232, 162, 154, 45, 0, 0, 0, 0, 0, 0, 
    0, 185, 0, 69, 182, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 189, 179, 11, 0, 0, 0, 0, 0, 0, 25, 0, 0, 105, 
    0, 0, 16, 184, 48, 72, 65, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=44
    99, 107, 105, 110, 109, 105, 110, 119, 115, 93, 84, 78, 91, 106, 99, 
    104, 115, 108, 115, 100, 80, 149, 110, 86, 31, 52, 58, 45, 56, 89, 
    90, 28, 108, 116, 101, 41, 107, 66, 40, 0, 46, 42, 62, 28, 43, 
    123, 0, 102, 107, 115, 58, 61, 65, 25, 0, 85, 37, 45, 51, 0, 
    121, 0, 145, 53, 81, 126, 104, 81, 35, 0, 61, 106, 19, 59, 30, 
    119, 0, 163, 105, 0, 101, 91, 83, 76, 0, 113, 102, 0, 46, 65, 
    139, 29, 81, 132, 0, 16, 37, 90, 83, 0, 110, 78, 17, 2, 62, 
    123, 41, 113, 78, 15, 0, 120, 33, 61, 0, 70, 76, 0, 16, 73, 
    99, 5, 147, 0, 97, 21, 58, 28, 7, 72, 0, 78, 0, 15, 73, 
    24, 15, 118, 0, 82, 77, 21, 38, 73, 34, 62, 15, 0, 35, 102, 
    0, 37, 103, 0, 144, 84, 0, 17, 87, 49, 0, 0, 0, 0, 0, 
    0, 0, 63, 0, 90, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 100, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=45
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=46
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 7, 35, 0, 0, 0, 12, 0, 0, 0, 5, 0, 
    0, 34, 0, 0, 3, 18, 0, 0, 0, 89, 0, 0, 0, 10, 22, 
    0, 121, 0, 6, 0, 18, 0, 0, 0, 113, 0, 0, 0, 0, 89, 
    0, 83, 0, 99, 0, 0, 0, 0, 0, 141, 0, 0, 0, 0, 38, 
    0, 30, 0, 0, 96, 0, 0, 0, 0, 268, 0, 0, 19, 0, 0, 
    0, 0, 0, 0, 121, 75, 0, 0, 0, 228, 0, 0, 7, 22, 0, 
    0, 0, 0, 0, 83, 113, 0, 0, 0, 147, 0, 0, 35, 2, 0, 
    0, 9, 0, 53, 0, 3, 0, 0, 43, 0, 8, 0, 23, 39, 23, 
    0, 11, 0, 108, 0, 0, 52, 0, 0, 0, 0, 0, 68, 59, 0, 
    96, 0, 0, 239, 0, 0, 83, 0, 0, 0, 0, 25, 34, 12, 0, 
    95, 47, 0, 193, 0, 0, 0, 0, 0, 0, 4, 10, 9, 13, 0, 
    0, 91, 115, 0, 0, 0, 0, 0, 0, 8, 19, 17, 4, 6, 25, 
    0, 8, 180, 0, 0, 12, 0, 0, 9, 10, 6, 3, 0, 42, 0, 
    0, 9, 17, 0, 0, 18, 4, 0, 20, 6, 0, 11, 72, 0, 0, 
    
    -- channel=47
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=48
    15, 15, 16, 12, 8, 22, 11, 3, 0, 7, 16, 27, 25, 8, 0, 
    14, 13, 14, 7, 21, 82, 1, 7, 0, 70, 63, 46, 49, 40, 10, 
    0, 61, 13, 7, 7, 42, 11, 29, 54, 138, 81, 89, 30, 48, 52, 
    0, 124, 18, 19, 4, 67, 64, 42, 58, 140, 61, 56, 42, 20, 90, 
    72, 158, 11, 109, 145, 88, 66, 43, 35, 159, 106, 29, 73, 28, 41, 
    85, 179, 26, 0, 195, 115, 100, 64, 16, 237, 74, 39, 90, 58, 43, 
    108, 109, 77, 0, 122, 161, 124, 86, 32, 222, 72, 51, 80, 101, 54, 
    125, 150, 78, 49, 87, 187, 64, 85, 60, 152, 83, 43, 96, 80, 56, 
    143, 190, 43, 155, 42, 94, 76, 70, 130, 34, 79, 15, 70, 91, 42, 
    168, 178, 61, 183, 74, 67, 149, 111, 68, 56, 17, 46, 106, 75, 22, 
    231, 167, 68, 303, 133, 102, 167, 144, 73, 53, 94, 109, 123, 132, 96, 
    214, 224, 154, 269, 64, 102, 128, 127, 119, 118, 133, 141, 155, 152, 142, 
    140, 192, 261, 159, 66, 135, 123, 125, 123, 134, 155, 163, 153, 161, 199, 
    148, 152, 244, 130, 108, 147, 127, 125, 134, 146, 148, 157, 152, 193, 138, 
    136, 158, 142, 144, 102, 135, 138, 139, 148, 155, 132, 154, 211, 167, 119, 
    
    -- channel=49
    255, 266, 273, 278, 275, 255, 279, 294, 278, 223, 182, 195, 228, 244, 248, 
    278, 283, 284, 282, 284, 317, 256, 227, 155, 149, 134, 104, 110, 196, 241, 
    153, 195, 280, 287, 280, 171, 156, 94, 116, 133, 105, 118, 111, 94, 210, 
    140, 173, 264, 284, 244, 198, 187, 118, 99, 89, 126, 84, 88, 83, 151, 
    148, 187, 243, 258, 295, 182, 121, 106, 67, 114, 155, 125, 115, 120, 73, 
    39, 119, 234, 140, 58, 111, 182, 145, 118, 151, 102, 81, 97, 111, 116, 
    74, 89, 149, 239, 126, 171, 140, 137, 118, 112, 98, 97, 88, 118, 126, 
    78, 126, 110, 203, 174, 143, 66, 68, 118, 125, 117, 81, 83, 90, 175, 
    83, 82, 55, 137, 116, 43, 112, 123, 137, 117, 76, 44, 59, 173, 244, 
    94, 83, 95, 83, 96, 76, 128, 180, 63, 84, 54, 64, 128, 221, 226, 
    80, 87, 73, 158, 247, 148, 77, 41, 62, 59, 55, 64, 20, 9, 14, 
    0, 24, 128, 156, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 58, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    
    -- channel=50
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 13, 0, 0, 2, 11, 
    0, 0, 0, 0, 0, 0, 32, 0, 63, 0, 0, 0, 0, 0, 0, 
    35, 0, 0, 0, 0, 30, 80, 54, 0, 0, 28, 11, 43, 0, 0, 
    132, 0, 0, 0, 0, 0, 0, 28, 0, 0, 73, 24, 62, 28, 0, 
    125, 0, 51, 0, 0, 0, 80, 54, 43, 0, 0, 77, 0, 42, 0, 
    135, 0, 72, 28, 0, 60, 26, 53, 70, 0, 106, 130, 0, 26, 0, 
    110, 19, 14, 86, 0, 0, 26, 41, 114, 0, 141, 61, 0, 0, 24, 
    58, 29, 31, 8, 0, 0, 177, 49, 69, 0, 77, 95, 0, 0, 32, 
    62, 0, 150, 0, 8, 58, 54, 0, 0, 45, 0, 151, 0, 0, 0, 
    13, 0, 158, 0, 80, 5, 0, 0, 17, 52, 127, 16, 0, 0, 11, 
    0, 0, 167, 0, 29, 0, 0, 48, 113, 42, 0, 0, 0, 0, 0, 
    0, 0, 41, 0, 272, 166, 32, 34, 27, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 295, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    33, 0, 0, 152, 61, 0, 2, 0, 0, 0, 0, 0, 3, 0, 49, 
    49, 0, 0, 62, 37, 0, 0, 0, 0, 0, 13, 0, 0, 0, 84, 
    
    -- channel=51
    269, 260, 270, 273, 275, 250, 277, 296, 283, 246, 222, 228, 235, 247, 259, 
    276, 269, 273, 276, 275, 218, 241, 240, 210, 162, 110, 129, 173, 228, 251, 
    208, 259, 282, 284, 288, 230, 200, 169, 140, 93, 71, 89, 95, 161, 218, 
    107, 164, 265, 279, 242, 209, 125, 107, 104, 105, 100, 105, 112, 116, 188, 
    59, 69, 226, 226, 86, 73, 81, 100, 103, 118, 85, 92, 107, 103, 142, 
    45, 60, 212, 204, 95, 94, 80, 99, 93, 91, 71, 103, 104, 97, 97, 
    47, 27, 187, 238, 129, 110, 72, 94, 88, 69, 75, 92, 99, 95, 106, 
    28, 31, 85, 179, 145, 70, 84, 102, 121, 111, 93, 96, 95, 105, 176, 
    10, 12, 48, 85, 130, 112, 121, 103, 112, 138, 128, 124, 120, 155, 207, 
    51, 25, 40, 39, 66, 110, 106, 56, 80, 132, 116, 107, 101, 189, 233, 
    39, 36, 45, 42, 0, 18, 12, 25, 44, 77, 53, 21, 8, 53, 68, 
    0, 19, 38, 14, 0, 31, 9, 11, 4, 3, 0, 0, 0, 0, 0, 
    0, 0, 41, 3, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 17, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=52
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=53
    51, 60, 52, 63, 60, 48, 58, 74, 68, 49, 48, 34, 53, 65, 71, 
    53, 56, 48, 68, 44, 0, 97, 47, 86, 2, 21, 6, 0, 20, 53, 
    44, 3, 53, 75, 41, 0, 145, 79, 0, 0, 16, 36, 54, 0, 1, 
    184, 0, 52, 42, 60, 20, 14, 36, 0, 0, 115, 0, 84, 37, 0, 
    208, 0, 119, 0, 0, 0, 104, 83, 30, 0, 27, 106, 0, 77, 0, 
    121, 0, 165, 0, 0, 90, 108, 84, 102, 0, 109, 164, 0, 45, 42, 
    143, 0, 73, 162, 0, 0, 14, 95, 139, 0, 177, 87, 0, 0, 44, 
    82, 70, 50, 91, 0, 0, 173, 24, 113, 0, 110, 106, 0, 0, 83, 
    82, 0, 177, 0, 12, 18, 87, 0, 0, 38, 0, 153, 0, 0, 0, 
    18, 0, 210, 0, 84, 0, 0, 16, 0, 30, 130, 21, 0, 0, 64, 
    0, 0, 199, 0, 180, 0, 0, 14, 146, 63, 0, 0, 0, 0, 0, 
    0, 0, 84, 0, 176, 146, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 298, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 130, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 
    
    -- channel=54
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 83, 63, 40, 0, 0, 
    36, 0, 0, 0, 0, 0, 0, 12, 40, 0, 31, 0, 32, 0, 0, 
    145, 48, 0, 0, 20, 0, 19, 27, 35, 0, 24, 30, 30, 52, 0, 
    122, 101, 0, 0, 0, 0, 44, 11, 75, 0, 66, 34, 22, 57, 32, 
    109, 159, 0, 0, 0, 0, 61, 35, 73, 24, 80, 53, 29, 47, 20, 
    125, 180, 5, 0, 0, 34, 69, 4, 9, 0, 39, 44, 29, 0, 0, 
    190, 190, 144, 47, 0, 0, 0, 32, 0, 0, 0, 3, 0, 0, 0, 
    131, 153, 197, 100, 90, 0, 0, 122, 21, 0, 34, 31, 8, 0, 0, 
    171, 123, 169, 101, 285, 196, 189, 206, 195, 126, 192, 257, 267, 211, 197, 
    327, 225, 161, 126, 251, 260, 260, 268, 322, 340, 383, 397, 429, 422, 433, 
    506, 293, 139, 215, 287, 368, 369, 353, 363, 393, 435, 455, 451, 455, 497, 
    540, 454, 234, 347, 327, 375, 388, 368, 382, 418, 455, 470, 479, 526, 519, 
    529, 493, 404, 328, 343, 361, 380, 380, 392, 428, 441, 429, 463, 554, 521, 
    
    -- channel=55
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=56
    3, 0, 0, 0, 0, 0, 2, 0, 0, 0, 3, 2, 0, 1, 0, 
    3, 0, 0, 0, 0, 0, 14, 2, 0, 0, 0, 8, 8, 0, 0, 
    10, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 2, 17, 0, 
    0, 12, 4, 0, 0, 0, 0, 9, 5, 0, 3, 2, 0, 23, 0, 
    0, 0, 25, 0, 0, 17, 0, 10, 3, 0, 0, 11, 0, 0, 31, 
    44, 0, 37, 33, 0, 14, 0, 0, 0, 0, 21, 15, 0, 0, 14, 
    48, 0, 27, 0, 0, 0, 0, 10, 0, 0, 6, 9, 0, 0, 12, 
    49, 0, 49, 0, 0, 0, 24, 0, 0, 0, 0, 2, 0, 3, 9, 
    20, 0, 58, 0, 45, 0, 0, 0, 0, 0, 0, 12, 0, 0, 3, 
    0, 0, 7, 0, 5, 44, 0, 0, 43, 4, 4, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 11, 7, 0, 21, 0, 0, 0, 9, 0, 3, 
    0, 0, 0, 0, 4, 22, 0, 0, 2, 0, 0, 0, 0, 0, 1, 
    22, 9, 18, 0, 15, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    7, 11, 27, 0, 5, 0, 2, 0, 0, 0, 1, 0, 0, 0, 13, 
    12, 0, 23, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    
    -- channel=57
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=58
    36, 36, 37, 34, 37, 38, 29, 30, 37, 41, 50, 52, 50, 43, 50, 
    37, 34, 36, 31, 40, 26, 16, 32, 59, 78, 63, 57, 60, 57, 47, 
    32, 65, 32, 32, 32, 27, 40, 68, 83, 81, 41, 70, 64, 72, 60, 
    37, 78, 23, 37, 26, 70, 39, 68, 75, 79, 33, 58, 72, 78, 86, 
    41, 33, 11, 81, 10, 28, 16, 50, 68, 111, 30, 42, 74, 78, 86, 
    25, 15, 1, 37, 33, 28, 4, 45, 52, 104, 0, 46, 75, 77, 84, 
    32, 0, 24, 30, 73, 39, 0, 32, 42, 80, 10, 47, 76, 74, 54, 
    12, 15, 39, 29, 82, 23, 7, 42, 50, 60, 29, 41, 82, 53, 60, 
    1, 11, 11, 56, 27, 58, 41, 47, 73, 34, 40, 63, 89, 73, 43, 
    11, 13, 5, 74, 13, 70, 77, 23, 33, 52, 73, 106, 92, 48, 34, 
    34, 8, 5, 72, 0, 25, 47, 20, 42, 82, 98, 102, 91, 70, 68, 
    59, 43, 28, 8, 0, 48, 69, 70, 81, 94, 93, 93, 89, 83, 81, 
    77, 67, 66, 0, 31, 88, 87, 90, 93, 96, 97, 86, 79, 90, 85, 
    82, 89, 72, 0, 77, 89, 83, 87, 97, 92, 89, 84, 93, 88, 60, 
    74, 95, 81, 63, 87, 93, 92, 93, 92, 83, 79, 97, 97, 57, 79, 
    
    -- channel=59
    193, 207, 207, 204, 193, 209, 212, 206, 187, 160, 140, 159, 171, 159, 133, 
    189, 214, 214, 207, 217, 323, 199, 188, 106, 142, 121, 95, 111, 146, 148, 
    127, 180, 211, 206, 208, 240, 133, 64, 77, 228, 178, 141, 57, 68, 164, 
    40, 186, 205, 219, 193, 191, 196, 93, 83, 228, 179, 122, 55, 0, 143, 
    168, 308, 201, 298, 419, 315, 229, 113, 44, 209, 250, 108, 106, 17, 40, 
    220, 354, 230, 185, 395, 327, 303, 156, 36, 364, 270, 100, 127, 80, 35, 
    250, 282, 207, 128, 245, 372, 350, 234, 85, 370, 219, 109, 106, 150, 102, 
    322, 319, 171, 177, 201, 434, 245, 196, 120, 311, 224, 97, 126, 159, 133, 
    365, 394, 158, 265, 190, 188, 165, 157, 191, 154, 172, 31, 68, 157, 200, 
    387, 384, 183, 281, 189, 148, 253, 269, 165, 147, 21, 0, 109, 223, 185, 
    404, 382, 189, 499, 371, 236, 344, 313, 139, 41, 37, 73, 106, 148, 108, 
    241, 373, 309, 591, 302, 99, 107, 101, 66, 59, 70, 83, 101, 106, 92, 
    65, 208, 409, 475, 95, 90, 72, 66, 53, 61, 84, 112, 113, 111, 161, 
    62, 78, 322, 281, 84, 102, 78, 67, 73, 89, 85, 92, 74, 141, 97, 
    72, 77, 93, 94, 26, 61, 76, 85, 111, 120, 75, 79, 185, 161, 21, 
    
    -- channel=60
    392, 402, 402, 403, 393, 387, 416, 414, 383, 354, 324, 339, 346, 332, 311, 
    388, 395, 409, 413, 415, 521, 372, 374, 291, 280, 242, 201, 241, 328, 336, 
    316, 404, 415, 409, 416, 461, 314, 170, 165, 359, 320, 272, 194, 194, 352, 
    169, 319, 409, 415, 385, 339, 346, 213, 224, 370, 350, 254, 191, 107, 295, 
    309, 473, 395, 436, 602, 416, 369, 231, 176, 297, 382, 226, 231, 140, 130, 
    330, 567, 422, 331, 604, 462, 483, 276, 166, 478, 447, 234, 259, 206, 121, 
    329, 503, 384, 314, 409, 526, 578, 397, 230, 531, 391, 225, 220, 275, 234, 
    425, 498, 273, 357, 340, 648, 446, 368, 276, 479, 411, 221, 246, 315, 295, 
    511, 562, 284, 446, 316, 336, 308, 301, 331, 306, 327, 180, 180, 312, 373, 
    594, 561, 355, 399, 327, 245, 369, 440, 266, 332, 188, 79, 237, 404, 379, 
    621, 545, 360, 612, 566, 334, 518, 528, 307, 144, 107, 159, 212, 307, 265, 
    412, 573, 474, 808, 561, 247, 213, 200, 180, 170, 190, 194, 212, 223, 205, 
    194, 343, 553, 738, 242, 195, 176, 172, 162, 168, 191, 218, 242, 235, 273, 
    190, 182, 428, 593, 230, 208, 183, 162, 177, 194, 202, 221, 195, 248, 266, 
    197, 183, 208, 256, 154, 182, 216, 205, 218, 226, 185, 184, 289, 294, 147, 
    
    -- channel=61
    338, 348, 340, 351, 345, 333, 357, 368, 351, 325, 288, 279, 286, 294, 288, 
    333, 346, 350, 365, 349, 366, 355, 339, 285, 199, 180, 168, 192, 260, 292, 
    305, 294, 357, 363, 362, 399, 301, 188, 123, 169, 223, 170, 161, 151, 254, 
    226, 140, 354, 357, 348, 256, 262, 159, 143, 185, 266, 188, 152, 95, 170, 
    264, 252, 357, 298, 395, 278, 298, 181, 137, 94, 273, 202, 142, 117, 83, 
    263, 329, 370, 291, 360, 325, 347, 225, 159, 127, 349, 215, 156, 144, 82, 
    243, 345, 308, 328, 235, 292, 416, 279, 221, 198, 328, 186, 132, 156, 170, 
    290, 331, 212, 303, 216, 368, 354, 260, 218, 236, 307, 203, 135, 200, 213, 
    347, 335, 249, 243, 244, 242, 248, 215, 183, 265, 252, 178, 99, 187, 281, 
    374, 339, 304, 179, 277, 148, 193, 298, 190, 248, 171, 57, 101, 262, 332, 
    317, 342, 312, 211, 376, 228, 251, 337, 231, 107, 38, 35, 77, 181, 190, 
    179, 289, 308, 394, 501, 195, 117, 110, 87, 59, 53, 50, 53, 64, 65, 
    51, 129, 230, 499, 253, 58, 55, 46, 42, 32, 34, 48, 75, 68, 63, 
    53, 32, 130, 427, 127, 58, 59, 45, 38, 42, 46, 63, 45, 40, 110, 
    61, 22, 50, 159, 64, 45, 69, 56, 52, 62, 58, 31, 51, 114, 53, 
    
    -- channel=62
    52, 66, 56, 62, 52, 63, 67, 59, 45, 42, 38, 38, 47, 44, 26, 
    48, 65, 58, 68, 56, 120, 91, 62, 32, 19, 51, 31, 13, 25, 37, 
    48, 22, 61, 62, 52, 89, 63, 4, 0, 57, 117, 75, 50, 0, 36, 
    94, 0, 77, 55, 70, 33, 105, 44, 33, 44, 138, 56, 37, 0, 0, 
    168, 145, 116, 34, 248, 171, 173, 76, 28, 0, 149, 96, 36, 25, 0, 
    162, 200, 152, 36, 156, 173, 216, 108, 67, 12, 211, 94, 39, 45, 10, 
    165, 223, 100, 79, 48, 131, 238, 156, 109, 70, 195, 82, 29, 50, 68, 
    204, 236, 99, 113, 30, 189, 211, 110, 89, 76, 156, 87, 26, 77, 57, 
    251, 236, 163, 113, 91, 81, 99, 78, 60, 93, 64, 47, 0, 37, 60, 
    231, 225, 212, 93, 161, 39, 75, 191, 87, 73, 42, 0, 12, 65, 73, 
    185, 225, 209, 125, 318, 164, 154, 220, 145, 32, 0, 12, 28, 56, 51, 
    101, 190, 215, 256, 324, 104, 59, 55, 47, 28, 42, 47, 64, 72, 74, 
    76, 74, 139, 331, 160, 57, 56, 44, 36, 36, 48, 69, 84, 73, 94, 
    84, 57, 67, 286, 73, 58, 66, 49, 43, 55, 59, 69, 63, 69, 116, 
    100, 60, 57, 88, 30, 24, 47, 57, 62, 80, 73, 49, 79, 148, 90, 
    
    -- channel=63
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end ifmap_package;
