library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    0, 0, 0, 
    0, 76, 58, 
    135, 292, 0, 
    
    -- channel=1
    193, 0, 0, 
    0, 0, 136, 
    171, 555, 457, 
    
    -- channel=2
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=3
    180, 277, 241, 
    0, 0, 0, 
    222, 0, 182, 
    
    -- channel=4
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=5
    94, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=6
    549, 859, 586, 
    1015, 424, 401, 
    734, 430, 487, 
    
    -- channel=7
    168, 0, 0, 
    0, 0, 0, 
    289, 103, 0, 
    
    -- channel=8
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=9
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=10
    107, 0, 0, 
    0, 0, 24, 
    151, 0, 0, 
    
    -- channel=11
    563, 481, 428, 
    279, 396, 178, 
    764, 593, 729, 
    
    -- channel=12
    0, 0, 304, 
    0, 0, 0, 
    307, 0, 0, 
    
    -- channel=13
    328, 84, 216, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=14
    0, 0, 0, 
    0, 40, 0, 
    315, 0, 0, 
    
    -- channel=15
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=16
    0, 79, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=17
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 157, 
    
    -- channel=18
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=19
    0, 0, 0, 
    0, 0, 0, 
    267, 76, 0, 
    
    -- channel=20
    143, 45, 257, 
    0, 29, 303, 
    0, 0, 0, 
    
    -- channel=21
    0, 38, 185, 
    0, 0, 0, 
    0, 0, 64, 
    
    -- channel=22
    68, 0, 61, 
    0, 172, 8, 
    13, 24, 31, 
    
    -- channel=23
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=24
    0, 0, 0, 
    0, 0, 0, 
    0, 190, 358, 
    
    -- channel=25
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=26
    29, 217, 519, 
    0, 305, 319, 
    0, 0, 0, 
    
    -- channel=27
    0, 0, 0, 
    0, 0, 164, 
    0, 0, 0, 
    
    -- channel=28
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 200, 
    
    -- channel=29
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=30
    0, 53, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=31
    0, 159, 207, 
    0, 10, 0, 
    0, 0, 0, 
    
    -- channel=32
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=33
    130, 128, 11, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=34
    0, 40, 66, 
    0, 0, 0, 
    0, 375, 668, 
    
    -- channel=35
    0, 65, 0, 
    0, 0, 37, 
    0, 0, 0, 
    
    -- channel=36
    332, 421, 406, 
    36, 391, 188, 
    0, 0, 0, 
    
    -- channel=37
    804, 589, 385, 
    712, 697, 736, 
    518, 0, 0, 
    
    -- channel=38
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=39
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=40
    0, 0, 0, 
    0, 0, 0, 
    384, 157, 283, 
    
    -- channel=41
    0, 0, 90, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=42
    0, 0, 0, 
    0, 83, 30, 
    0, 0, 0, 
    
    -- channel=43
    0, 0, 0, 
    0, 0, 93, 
    0, 164, 0, 
    
    -- channel=44
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=45
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=46
    0, 0, 0, 
    0, 0, 0, 
    81, 315, 292, 
    
    -- channel=47
    0, 0, 0, 
    79, 242, 276, 
    0, 81, 61, 
    
    -- channel=48
    15, 136, 124, 
    383, 320, 97, 
    357, 94, 0, 
    
    -- channel=49
    0, 0, 0, 
    0, 0, 0, 
    13, 0, 0, 
    
    -- channel=50
    34, 165, 268, 
    562, 307, 233, 
    0, 0, 0, 
    
    -- channel=51
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=52
    0, 0, 0, 
    285, 143, 0, 
    436, 187, 221, 
    
    -- channel=53
    0, 0, 186, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=54
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=55
    302, 386, 347, 
    442, 521, 360, 
    18, 166, 19, 
    
    -- channel=56
    234, 238, 448, 
    183, 317, 0, 
    30, 0, 0, 
    
    -- channel=57
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=58
    285, 213, 143, 
    243, 387, 417, 
    256, 80, 0, 
    
    -- channel=59
    0, 0, 0, 
    0, 0, 0, 
    0, 16, 0, 
    
    -- channel=60
    0, 0, 0, 
    0, 0, 52, 
    0, 279, 0, 
    
    -- channel=61
    0, 0, 0, 
    359, 0, 0, 
    172, 0, 0, 
    
    -- channel=62
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=63
    0, 164, 0, 
    0, 31, 0, 
    0, 0, 0, 
    
    
    others => 0);
end ifmap_package;
