library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 5, 0, 0, 2, 84, 0, 0, 0, 27, 2, 0, 2, 5, 0, 
    0, 4, 0, 0, 0, 0, 0, 0, 7, 74, 0, 0, 0, 0, 28, 
    0, 117, 0, 9, 1, 12, 13, 0, 0, 49, 0, 0, 0, 0, 54, 
    0, 84, 0, 40, 52, 0, 0, 0, 0, 88, 0, 0, 10, 0, 6, 
    0, 31, 0, 0, 66, 0, 0, 0, 0, 217, 0, 0, 7, 0, 0, 
    0, 0, 0, 0, 68, 77, 0, 0, 0, 168, 0, 0, 4, 27, 0, 
    0, 0, 0, 0, 22, 81, 0, 0, 0, 98, 0, 0, 17, 0, 0, 
    0, 0, 0, 56, 0, 0, 0, 18, 23, 0, 18, 0, 6, 29, 18, 
    0, 0, 0, 71, 0, 0, 26, 14, 0, 0, 0, 0, 52, 55, 0, 
    97, 0, 0, 203, 0, 0, 43, 0, 0, 0, 23, 36, 16, 5, 0, 
    29, 14, 0, 146, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    0, 31, 56, 0, 0, 0, 0, 0, 0, 4, 9, 13, 0, 0, 21, 
    0, 0, 79, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 5, 0, 0, 56, 0, 0, 
    
    -- channel=1
    164, 171, 171, 172, 168, 172, 174, 171, 163, 149, 131, 139, 147, 138, 122, 
    164, 171, 176, 175, 183, 273, 179, 158, 112, 149, 148, 116, 111, 132, 134, 
    120, 154, 173, 172, 174, 238, 142, 94, 84, 228, 205, 174, 116, 83, 147, 
    107, 170, 180, 185, 174, 181, 204, 122, 124, 223, 209, 146, 103, 40, 133, 
    224, 305, 191, 252, 381, 291, 242, 136, 92, 191, 264, 143, 137, 76, 57, 
    244, 351, 208, 149, 348, 287, 302, 188, 102, 299, 285, 140, 155, 128, 72, 
    256, 324, 187, 128, 238, 321, 359, 247, 145, 342, 256, 146, 140, 174, 133, 
    308, 353, 196, 190, 205, 387, 271, 216, 146, 291, 248, 144, 150, 173, 147, 
    365, 394, 193, 267, 180, 210, 191, 184, 201, 199, 173, 86, 89, 158, 173, 
    386, 388, 239, 296, 207, 145, 249, 299, 177, 156, 87, 41, 125, 206, 179, 
    399, 378, 250, 432, 405, 253, 327, 332, 186, 112, 97, 126, 167, 205, 169, 
    293, 373, 328, 549, 375, 174, 178, 169, 141, 139, 156, 171, 187, 201, 185, 
    182, 252, 377, 481, 186, 166, 155, 150, 147, 154, 181, 201, 206, 205, 246, 
    185, 173, 308, 363, 165, 185, 168, 151, 157, 175, 185, 193, 185, 224, 210, 
    189, 177, 178, 206, 129, 146, 163, 168, 188, 207, 176, 178, 259, 270, 156, 
    
    -- channel=2
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 0, 0, 0, 51, 0, 0, 0, 35, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 71, 0, 9, 0, 0, 19, 
    0, 30, 0, 18, 5, 0, 6, 0, 0, 39, 11, 0, 0, 0, 0, 
    17, 71, 0, 4, 156, 58, 10, 0, 0, 98, 18, 0, 12, 0, 0, 
    8, 44, 12, 0, 72, 56, 63, 0, 0, 115, 5, 0, 0, 4, 0, 
    31, 42, 0, 0, 16, 122, 24, 38, 0, 87, 15, 0, 17, 23, 0, 
    48, 89, 0, 43, 0, 57, 7, 0, 14, 0, 52, 0, 12, 4, 0, 
    82, 86, 0, 66, 9, 0, 28, 6, 8, 25, 0, 0, 0, 0, 0, 
    117, 77, 0, 128, 0, 0, 80, 78, 0, 0, 0, 0, 9, 26, 1, 
    141, 114, 34, 148, 80, 41, 59, 56, 21, 16, 19, 29, 30, 32, 26, 
    14, 115, 109, 122, 9, 20, 18, 16, 11, 14, 22, 30, 38, 41, 40, 
    20, 27, 158, 77, 7, 28, 9, 18, 23, 28, 34, 47, 28, 52, 59, 
    17, 35, 39, 67, 13, 41, 40, 21, 24, 24, 21, 27, 48, 37, 0, 
    
    -- channel=3
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 6, 13, 23, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 11, 11, 3, 6, 3, 17, 10, 0, 
    36, 0, 0, 0, 0, 0, 5, 14, 8, 21, 6, 10, 10, 15, 0, 
    45, 5, 0, 0, 0, 15, 0, 8, 6, 4, 6, 23, 11, 20, 21, 
    58, 0, 0, 0, 0, 0, 0, 14, 11, 0, 20, 19, 15, 17, 8, 
    45, 28, 17, 0, 0, 0, 12, 4, 13, 0, 6, 16, 17, 3, 0, 
    38, 29, 37, 9, 0, 7, 8, 0, 14, 0, 0, 17, 11, 0, 0, 
    21, 24, 31, 24, 20, 17, 24, 5, 8, 1, 13, 28, 5, 0, 0, 
    19, 24, 28, 29, 30, 27, 16, 31, 40, 35, 51, 53, 48, 36, 38, 
    52, 49, 42, 0, 11, 77, 63, 67, 72, 69, 73, 77, 83, 78, 83, 
    87, 57, 59, 0, 80, 76, 73, 72, 73, 77, 83, 84, 79, 87, 96, 
    100, 88, 56, 29, 70, 75, 76, 74, 78, 81, 84, 87, 93, 95, 80, 
    97, 94, 75, 62, 68, 72, 74, 78, 74, 79, 81, 88, 90, 85, 97, 
    
    -- channel=4
    129, 134, 133, 134, 132, 128, 139, 146, 134, 114, 100, 105, 108, 117, 114, 
    128, 139, 141, 136, 136, 120, 120, 120, 89, 54, 28, 44, 70, 95, 110, 
    98, 113, 136, 138, 140, 148, 65, 53, 39, 54, 32, 30, 25, 57, 97, 
    21, 73, 124, 140, 114, 87, 57, 31, 24, 72, 32, 41, 14, 17, 92, 
    0, 63, 102, 133, 81, 73, 47, 26, 25, 51, 46, 25, 33, 15, 57, 
    3, 45, 89, 99, 84, 60, 42, 40, 16, 81, 39, 16, 41, 23, 16, 
    0, 31, 72, 101, 103, 64, 65, 32, 23, 85, 17, 15, 25, 27, 30, 
    6, 24, 32, 64, 85, 97, 46, 48, 26, 98, 27, 17, 35, 46, 65, 
    11, 31, 0, 40, 43, 55, 34, 33, 46, 62, 53, 26, 34, 65, 108, 
    32, 33, 0, 36, 25, 48, 49, 32, 39, 54, 24, 15, 41, 105, 107, 
    34, 34, 0, 68, 0, 14, 45, 32, 0, 0, 0, 0, 0, 0, 0, 
    9, 15, 16, 89, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 22, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=5
    42, 36, 37, 37, 39, 35, 42, 42, 35, 33, 32, 38, 31, 37, 33, 
    42, 39, 38, 37, 35, 32, 27, 34, 9, 15, 10, 33, 49, 43, 38, 
    39, 49, 44, 37, 44, 58, 1, 17, 18, 33, 11, 7, 14, 54, 45, 
    0, 87, 48, 39, 32, 16, 10, 6, 21, 53, 0, 22, 2, 30, 67, 
    0, 61, 27, 17, 0, 0, 0, 1, 26, 40, 4, 0, 24, 7, 67, 
    0, 39, 16, 25, 39, 0, 0, 0, 9, 79, 0, 0, 31, 5, 14, 
    0, 25, 35, 2, 59, 18, 4, 0, 0, 81, 0, 2, 28, 19, 21, 
    0, 0, 14, 12, 28, 44, 0, 17, 1, 74, 0, 4, 30, 36, 28, 
    0, 2, 0, 27, 15, 19, 7, 19, 32, 28, 41, 2, 40, 39, 43, 
    0, 6, 0, 33, 0, 19, 12, 0, 40, 14, 0, 14, 49, 63, 33, 
    35, 4, 0, 55, 0, 0, 25, 0, 0, 0, 17, 9, 29, 29, 6, 
    72, 12, 0, 57, 0, 0, 23, 17, 4, 9, 15, 15, 10, 19, 8, 
    17, 68, 19, 23, 0, 8, 9, 14, 15, 16, 14, 17, 16, 4, 9, 
    2, 19, 82, 0, 0, 16, 5, 15, 10, 13, 15, 17, 5, 21, 22, 
    0, 12, 25, 32, 17, 29, 17, 8, 9, 9, 10, 13, 13, 6, 0, 
    
    -- channel=6
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 18, 18, 5, 0, 0, 
    0, 0, 0, 0, 0, 12, 0, 1, 5, 59, 63, 46, 28, 11, 0, 
    6, 21, 0, 0, 0, 0, 16, 20, 38, 66, 43, 41, 33, 19, 4, 
    33, 68, 0, 0, 20, 18, 44, 30, 43, 41, 49, 21, 39, 19, 15, 
    70, 104, 0, 0, 110, 38, 49, 31, 32, 78, 65, 33, 49, 34, 13, 
    57, 111, 2, 0, 51, 51, 81, 42, 35, 108, 59, 40, 47, 49, 31, 
    72, 98, 30, 0, 11, 97, 72, 68, 32, 86, 56, 48, 53, 54, 4, 
    99, 124, 59, 66, 21, 61, 41, 49, 41, 32, 57, 34, 42, 21, 0, 
    111, 122, 72, 99, 54, 27, 45, 64, 58, 38, 31, 22, 30, 0, 0, 
    137, 107, 79, 122, 64, 56, 104, 114, 58, 43, 60, 69, 94, 99, 78, 
    197, 143, 78, 153, 147, 124, 139, 135, 119, 118, 133, 142, 150, 157, 150, 
    167, 177, 119, 165, 108, 128, 127, 127, 127, 135, 147, 156, 160, 157, 169, 
    172, 156, 177, 166, 110, 138, 130, 130, 132, 145, 161, 172, 163, 183, 194, 
    170, 167, 155, 165, 130, 145, 143, 131, 134, 149, 151, 153, 164, 189, 153, 
    
    -- channel=7
    120, 123, 123, 127, 126, 118, 124, 139, 130, 101, 83, 86, 97, 110, 115, 
    122, 129, 126, 129, 127, 97, 111, 99, 80, 50, 29, 32, 47, 80, 105, 
    71, 80, 129, 133, 131, 103, 78, 57, 42, 19, 29, 30, 29, 41, 77, 
    49, 33, 115, 127, 103, 83, 50, 41, 26, 26, 41, 35, 34, 31, 49, 
    40, 12, 103, 105, 43, 49, 41, 37, 24, 29, 40, 42, 28, 32, 34, 
    34, 6, 102, 104, 21, 54, 39, 47, 30, 4, 36, 41, 25, 30, 29, 
    43, 0, 62, 109, 40, 39, 28, 40, 37, 0, 39, 34, 25, 26, 38, 
    29, 12, 34, 59, 67, 14, 38, 30, 45, 34, 43, 38, 22, 30, 79, 
    18, 0, 28, 12, 49, 41, 50, 31, 29, 52, 41, 40, 28, 59, 92, 
    22, 12, 22, 0, 24, 35, 33, 24, 29, 37, 27, 20, 12, 64, 94, 
    0, 15, 22, 0, 20, 10, 0, 0, 1, 4, 0, 0, 0, 0, 0, 
    0, 0, 22, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=8
    5, 0, 4, 0, 0, 1, 3, 0, 0, 0, 2, 17, 4, 0, 0, 
    2, 0, 5, 0, 8, 0, 0, 0, 0, 21, 0, 0, 22, 28, 0, 
    0, 68, 4, 0, 8, 28, 0, 0, 9, 61, 0, 0, 0, 36, 34, 
    0, 95, 0, 8, 0, 22, 0, 0, 0, 109, 0, 2, 0, 0, 95, 
    0, 28, 0, 82, 0, 0, 0, 0, 0, 134, 0, 0, 0, 0, 51, 
    0, 24, 0, 25, 118, 9, 0, 0, 0, 210, 0, 0, 19, 0, 0, 
    0, 0, 15, 0, 95, 64, 0, 0, 0, 177, 0, 0, 11, 16, 0, 
    0, 0, 0, 0, 61, 84, 0, 5, 0, 116, 0, 0, 37, 15, 0, 
    0, 7, 0, 49, 0, 46, 0, 0, 39, 0, 32, 0, 43, 37, 11, 
    0, 13, 0, 85, 0, 12, 52, 0, 0, 3, 0, 4, 47, 41, 0, 
    90, 5, 0, 170, 0, 0, 62, 0, 0, 0, 0, 6, 22, 31, 0, 
    117, 76, 0, 122, 0, 0, 31, 26, 0, 8, 12, 16, 12, 13, 0, 
    0, 113, 132, 0, 0, 2, 0, 6, 2, 9, 13, 8, 6, 15, 14, 
    0, 17, 189, 0, 0, 12, 0, 1, 14, 11, 11, 16, 4, 32, 0, 
    0, 12, 35, 7, 0, 37, 24, 6, 11, 0, 0, 15, 45, 0, 0, 
    
    -- channel=9
    4, 0, 0, 0, 0, 0, 0, 0, 0, 22, 37, 28, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 14, 69, 12, 0, 0, 29, 24, 0, 
    39, 67, 0, 0, 0, 78, 37, 43, 1, 0, 0, 0, 0, 30, 6, 
    0, 0, 0, 0, 0, 12, 0, 0, 0, 39, 0, 16, 10, 0, 31, 
    0, 0, 0, 14, 0, 0, 0, 0, 9, 7, 0, 0, 0, 0, 20, 
    10, 0, 0, 41, 100, 34, 0, 0, 0, 0, 0, 13, 5, 0, 0, 
    0, 0, 26, 0, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 6, 32, 43, 0, 5, 1, 0, 11, 7, 0, 
    0, 0, 0, 0, 0, 84, 6, 0, 0, 0, 49, 58, 31, 0, 0, 
    8, 0, 0, 0, 0, 14, 0, 0, 0, 63, 55, 26, 0, 0, 5, 
    16, 0, 0, 0, 0, 0, 0, 47, 8, 0, 0, 0, 0, 39, 43, 
    101, 50, 0, 0, 80, 104, 70, 67, 30, 19, 5, 9, 0, 0, 0, 
    0, 73, 25, 0, 86, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 
    0, 0, 81, 65, 23, 0, 0, 0, 2, 0, 6, 19, 8, 0, 38, 
    0, 0, 11, 78, 31, 36, 36, 1, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=10
    168, 166, 175, 173, 173, 164, 184, 183, 170, 145, 123, 134, 143, 150, 138, 
    171, 179, 181, 178, 180, 196, 179, 160, 100, 87, 79, 82, 93, 128, 146, 
    114, 141, 182, 177, 182, 139, 84, 53, 65, 101, 70, 59, 53, 81, 133, 
    42, 148, 185, 183, 162, 127, 113, 63, 52, 105, 67, 61, 20, 30, 118, 
    47, 163, 173, 191, 198, 172, 90, 54, 28, 99, 105, 64, 59, 31, 79, 
    57, 119, 164, 132, 87, 103, 104, 73, 33, 172, 98, 31, 62, 44, 47, 
    68, 90, 124, 119, 110, 149, 123, 93, 36, 158, 61, 46, 53, 67, 66, 
    92, 84, 105, 124, 128, 174, 71, 65, 42, 143, 62, 34, 56, 75, 88, 
    90, 109, 43, 101, 116, 54, 59, 72, 95, 100, 68, 4, 34, 94, 163, 
    90, 105, 34, 94, 75, 83, 99, 106, 89, 64, 8, 8, 76, 167, 148, 
    109, 116, 31, 179, 124, 119, 133, 77, 31, 21, 17, 32, 41, 60, 45, 
    36, 79, 89, 222, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 33, 111, 141, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 90, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 
    
    -- channel=11
    12, 17, 11, 17, 14, 9, 13, 17, 13, 13, 14, 3, 9, 15, 19, 
    6, 9, 8, 20, 7, 0, 33, 9, 39, 0, 6, 0, 0, 0, 11, 
    19, 0, 9, 18, 7, 14, 58, 16, 0, 0, 49, 38, 46, 0, 0, 
    94, 0, 10, 1, 15, 0, 20, 39, 21, 0, 84, 26, 53, 19, 0, 
    125, 0, 55, 0, 24, 40, 82, 57, 34, 0, 35, 73, 7, 45, 0, 
    108, 9, 78, 27, 0, 76, 81, 59, 64, 0, 107, 95, 0, 39, 20, 
    104, 63, 19, 71, 0, 0, 65, 74, 89, 0, 121, 57, 2, 0, 40, 
    87, 78, 35, 33, 0, 0, 144, 50, 66, 0, 90, 69, 0, 19, 44, 
    101, 36, 125, 0, 29, 38, 49, 15, 0, 40, 0, 91, 0, 0, 0, 
    70, 48, 143, 0, 68, 21, 0, 47, 21, 45, 84, 7, 0, 0, 23, 
    0, 44, 137, 0, 141, 35, 0, 78, 105, 40, 0, 0, 0, 0, 0, 
    0, 12, 84, 0, 194, 100, 16, 17, 28, 9, 8, 8, 12, 15, 27, 
    33, 0, 0, 65, 182, 20, 26, 17, 17, 8, 4, 3, 21, 23, 3, 
    49, 6, 0, 145, 65, 11, 32, 16, 14, 12, 18, 20, 31, 0, 55, 
    64, 17, 7, 29, 31, 0, 21, 26, 11, 17, 34, 16, 0, 47, 80, 
    
    -- channel=12
    77, 83, 75, 83, 79, 74, 84, 85, 78, 74, 71, 64, 72, 75, 73, 
    74, 79, 74, 88, 73, 76, 104, 79, 84, 44, 65, 52, 38, 58, 72, 
    79, 50, 82, 87, 75, 73, 124, 64, 31, 9, 98, 80, 83, 23, 54, 
    142, 0, 91, 71, 89, 47, 86, 69, 58, 0, 142, 67, 92, 54, 0, 
    178, 37, 130, 4, 122, 83, 143, 101, 69, 0, 106, 117, 50, 80, 0, 
    148, 104, 161, 59, 68, 137, 170, 109, 108, 0, 169, 139, 41, 74, 54, 
    149, 149, 111, 134, 0, 56, 151, 137, 138, 0, 190, 107, 43, 47, 86, 
    149, 164, 86, 119, 9, 42, 190, 103, 123, 0, 153, 119, 28, 65, 90, 
    173, 121, 178, 66, 86, 80, 116, 77, 41, 92, 62, 119, 22, 50, 59, 
    151, 122, 214, 14, 141, 44, 43, 128, 63, 93, 109, 33, 3, 38, 95, 
    66, 127, 206, 0, 236, 96, 35, 146, 157, 74, 21, 13, 15, 40, 67, 
    6, 96, 157, 22, 273, 158, 63, 67, 74, 42, 41, 39, 48, 48, 64, 
    67, 1, 39, 172, 225, 54, 54, 47, 46, 37, 35, 40, 55, 54, 48, 
    84, 42, 0, 243, 102, 43, 66, 47, 40, 41, 45, 55, 62, 24, 87, 
    94, 47, 43, 85, 58, 30, 50, 56, 41, 54, 65, 43, 20, 87, 111, 
    
    -- channel=13
    58, 52, 59, 56, 57, 52, 66, 70, 57, 47, 47, 52, 50, 50, 44, 
    64, 59, 58, 59, 55, 31, 57, 55, 39, 12, 0, 8, 35, 55, 48, 
    36, 79, 65, 64, 60, 17, 37, 19, 1, 0, 0, 0, 0, 26, 46, 
    0, 28, 68, 61, 46, 31, 0, 0, 0, 0, 0, 0, 0, 0, 37, 
    0, 0, 56, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 61, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 71, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 26, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 49, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=14
    36, 36, 32, 30, 31, 28, 39, 41, 32, 36, 45, 41, 30, 33, 30, 
    31, 29, 33, 33, 23, 0, 29, 40, 61, 0, 0, 7, 35, 29, 25, 
    59, 49, 31, 35, 36, 66, 51, 34, 0, 0, 0, 0, 0, 30, 20, 
    0, 0, 25, 26, 27, 0, 0, 0, 0, 0, 10, 21, 13, 17, 20, 
    0, 0, 26, 0, 0, 0, 9, 6, 24, 0, 0, 0, 0, 0, 34, 
    8, 0, 30, 68, 43, 31, 0, 0, 0, 0, 16, 27, 0, 0, 0, 
    0, 2, 43, 32, 15, 0, 0, 0, 1, 0, 12, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 50, 37, 10, 0, 13, 13, 0, 16, 19, 
    0, 0, 12, 0, 8, 56, 13, 0, 0, 30, 21, 61, 24, 0, 4, 
    0, 0, 0, 0, 0, 22, 0, 0, 14, 40, 51, 7, 0, 0, 30, 
    0, 0, 10, 0, 0, 0, 0, 10, 7, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 71, 46, 18, 13, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 23, 18, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 14, 28, 0, 0, 0, 13, 12, 0, 
    34, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 21, 9, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 18, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 29, 20, 6, 0, 0, 0, 0, 0, 5, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 5, 12, 0, 0, 0, 
    0, 0, 0, 0, 4, 20, 0, 0, 0, 39, 22, 0, 7, 0, 0, 
    9, 0, 0, 0, 0, 0, 47, 46, 35, 0, 0, 0, 5, 25, 27, 
    45, 33, 0, 0, 21, 14, 0, 0, 0, 2, 1, 0, 0, 0, 0, 
    0, 28, 11, 11, 3, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 49, 31, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 
    0, 0, 0, 0, 0, 3, 10, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end ifmap_package;
