library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=1
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 14, 7, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 11, 8, 25, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 11, 11, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 16, 13, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 13, 11, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 7, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 15, 12, 29, 6, 0, 0, 0, 0, 0, 0, 0, 17, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 20, 22, 34, 21, 0, 0, 0, 0, 0, 0, 0, 7, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 30, 29, 35, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 37, 36, 39, 43, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 30, 36, 38, 40, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 20, 28, 27, 30, 24, 7, 12, 13, 0, 0, 0, 0, 0, 0, 11, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 16, 25, 18, 19, 17, 3, 20, 57, 52, 11, 0, 6, 3, 20, 33, 27, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 31, 37, 21, 23, 26, 11, 15, 46, 69, 55, 17, 13, 17, 26, 22, 20, 15, 4, 0, 0, 4, 10, 20, 31, 26, 24, 24, 19, 16, 21, 34, 
    0, 42, 49, 37, 38, 38, 19, 25, 46, 35, 32, 32, 12, 13, 15, 11, 22, 28, 18, 15, 31, 39, 39, 43, 51, 58, 61, 59, 58, 57, 61, 60, 
    3, 47, 37, 42, 39, 28, 19, 33, 39, 36, 44, 31, 29, 31, 31, 30, 32, 37, 37, 39, 48, 51, 54, 58, 63, 70, 71, 67, 66, 66, 70, 69, 
    29, 74, 45, 31, 41, 30, 15, 31, 35, 41, 41, 42, 44, 45, 45, 43, 43, 44, 46, 50, 53, 59, 63, 67, 71, 73, 70, 68, 73, 80, 86, 80, 
    35, 89, 64, 39, 34, 30, 32, 42, 45, 36, 37, 51, 51, 50, 49, 47, 46, 47, 50, 53, 59, 67, 73, 74, 72, 71, 67, 71, 85, 93, 89, 85, 
    35, 92, 77, 59, 38, 25, 46, 61, 51, 34, 43, 51, 56, 52, 47, 47, 49, 52, 55, 60, 64, 68, 73, 77, 79, 73, 73, 82, 91, 90, 85, 78, 
    34, 92, 83, 73, 58, 31, 35, 61, 45, 37, 49, 55, 57, 59, 53, 47, 47, 51, 58, 62, 67, 74, 74, 73, 75, 78, 84, 88, 92, 91, 75, 61, 
    39, 92, 83, 80, 73, 51, 29, 38, 43, 32, 41, 48, 55, 59, 59, 57, 55, 57, 60, 64, 69, 70, 71, 71, 74, 81, 89, 100, 107, 91, 63, 51, 
    35, 94, 80, 79, 78, 67, 50, 41, 35, 41, 40, 41, 43, 45, 51, 52, 52, 57, 66, 72, 71, 69, 68, 67, 70, 81, 96, 105, 97, 87, 67, 51, 
    33, 88, 74, 72, 74, 68, 57, 49, 43, 45, 43, 45, 46, 43, 38, 35, 38, 47, 57, 65, 70, 68, 61, 58, 63, 74, 86, 93, 90, 80, 67, 57, 
    0, 5, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 11, 4, 2, 0, 
    
    -- channel=2
    293, 198, 206, 190, 181, 196, 201, 193, 194, 201, 203, 195, 194, 204, 212, 211, 208, 206, 204, 194, 180, 177, 179, 184, 181, 174, 176, 181, 183, 177, 170, 55, 
    354, 289, 306, 290, 279, 292, 295, 290, 288, 286, 290, 283, 282, 299, 311, 312, 306, 293, 279, 268, 253, 249, 255, 262, 266, 260, 251, 255, 264, 257, 247, 108, 
    355, 292, 313, 295, 282, 297, 296, 291, 291, 293, 290, 258, 243, 282, 306, 301, 292, 260, 243, 228, 202, 180, 192, 222, 235, 261, 266, 260, 265, 262, 250, 104, 
    357, 291, 304, 298, 287, 303, 302, 294, 297, 307, 338, 253, 166, 233, 285, 262, 247, 238, 220, 199, 150, 114, 101, 124, 160, 192, 242, 267, 268, 259, 254, 107, 
    346, 276, 288, 295, 293, 304, 308, 296, 301, 315, 381, 333, 173, 200, 243, 234, 193, 194, 222, 188, 132, 101, 77, 85, 99, 119, 167, 250, 275, 253, 242, 104, 
    323, 211, 256, 327, 315, 303, 307, 300, 299, 311, 336, 311, 226, 182, 152, 160, 157, 160, 213, 189, 125, 105, 104, 109, 104, 78, 96, 194, 276, 264, 234, 98, 
    283, 115, 146, 312, 331, 301, 308, 311, 298, 291, 284, 265, 237, 173, 103, 117, 131, 123, 200, 229, 136, 82, 116, 147, 121, 80, 85, 130, 239, 278, 241, 93, 
    253, 39, 97, 229, 267, 284, 307, 308, 293, 238, 229, 248, 230, 153, 87, 113, 138, 118, 163, 257, 206, 91, 96, 145, 139, 103, 80, 97, 185, 280, 260, 88, 
    278, 0, 94, 199, 173, 241, 300, 317, 283, 160, 89, 189, 199, 125, 77, 96, 129, 120, 139, 228, 241, 133, 78, 95, 131, 124, 91, 68, 114, 251, 294, 96, 
    301, 47, 114, 169, 135, 209, 273, 352, 347, 171, 47, 116, 159, 91, 86, 79, 107, 95, 130, 237, 216, 130, 80, 69, 120, 126, 104, 77, 67, 164, 278, 125, 
    286, 70, 181, 152, 117, 191, 245, 307, 411, 243, 83, 120, 163, 72, 78, 98, 85, 73, 140, 281, 195, 101, 85, 66, 135, 148, 103, 84, 59, 97, 194, 119, 
    271, 57, 209, 163, 118, 191, 246, 220, 331, 296, 125, 177, 218, 97, 45, 105, 106, 36, 147, 314, 188, 77, 83, 75, 134, 159, 132, 100, 75, 77, 125, 76, 
    263, 45, 210, 130, 111, 223, 267, 196, 262, 282, 152, 198, 263, 142, 36, 90, 128, 53, 148, 303, 162, 70, 74, 91, 123, 148, 155, 128, 94, 89, 110, 44, 
    264, 56, 216, 73, 46, 230, 287, 204, 234, 271, 212, 220, 218, 174, 95, 101, 106, 69, 174, 282, 143, 72, 71, 73, 104, 122, 148, 149, 103, 103, 143, 48, 
    282, 64, 205, 62, 0, 168, 272, 201, 204, 245, 267, 243, 100, 98, 133, 145, 120, 77, 182, 277, 156, 78, 94, 91, 118, 145, 145, 155, 125, 131, 185, 72, 
    304, 65, 178, 87, 0, 88, 226, 181, 175, 254, 296, 281, 130, 63, 140, 148, 143, 126, 200, 255, 188, 117, 73, 74, 115, 162, 160, 158, 160, 182, 225, 80, 
    325, 52, 146, 117, 0, 30, 203, 166, 121, 203, 287, 225, 176, 133, 145, 147, 142, 159, 188, 227, 241, 207, 98, 78, 116, 163, 177, 162, 179, 222, 239, 78, 
    358, 53, 114, 125, 20, 0, 161, 192, 96, 126, 188, 191, 179, 145, 158, 121, 106, 189, 175, 123, 180, 222, 132, 87, 131, 158, 194, 205, 207, 241, 248, 87, 
    390, 91, 106, 124, 58, 0, 106, 193, 136, 108, 62, 159, 207, 157, 197, 98, 31, 180, 205, 134, 124, 107, 112, 114, 133, 158, 191, 242, 235, 246, 256, 95, 
    412, 143, 113, 133, 89, 2, 69, 164, 93, 103, 81, 120, 208, 183, 215, 106, 0, 91, 201, 186, 150, 90, 94, 125, 147, 179, 206, 254, 240, 250, 257, 96, 
    411, 193, 114, 141, 105, 22, 98, 216, 78, 0, 21, 91, 135, 166, 173, 91, 6, 17, 77, 119, 121, 106, 81, 77, 99, 121, 168, 200, 183, 182, 191, 60, 
    379, 215, 100, 133, 100, 18, 130, 272, 168, 0, 0, 55, 138, 161, 155, 122, 61, 44, 51, 44, 62, 69, 72, 59, 47, 55, 88, 108, 101, 92, 94, 0, 
    322, 225, 125, 125, 94, 36, 161, 269, 176, 62, 0, 38, 128, 142, 131, 126, 83, 52, 57, 53, 49, 41, 46, 45, 33, 25, 33, 45, 36, 25, 24, 0, 
    224, 158, 183, 166, 105, 113, 225, 244, 116, 26, 0, 35, 64, 62, 58, 59, 53, 37, 36, 43, 43, 33, 29, 26, 25, 18, 11, 16, 12, 9, 9, 0, 
    151, 25, 130, 199, 128, 155, 274, 198, 38, 0, 10, 27, 31, 23, 22, 30, 33, 26, 25, 29, 29, 20, 16, 20, 18, 15, 6, 6, 1, 2, 4, 0, 
    151, 0, 35, 132, 159, 209, 268, 116, 0, 0, 41, 24, 20, 18, 20, 26, 28, 26, 24, 25, 21, 17, 9, 10, 14, 13, 14, 21, 17, 8, 11, 0, 
    162, 0, 0, 41, 119, 264, 267, 43, 0, 1, 32, 33, 15, 6, 23, 29, 26, 23, 22, 21, 14, 16, 23, 14, 0, 0, 10, 26, 25, 9, 15, 0, 
    162, 0, 0, 0, 41, 201, 291, 48, 0, 37, 30, 30, 23, 0, 6, 20, 27, 29, 23, 17, 12, 3, 13, 16, 3, 0, 3, 13, 5, 0, 15, 0, 
    154, 0, 0, 0, 0, 76, 206, 115, 0, 55, 54, 52, 43, 21, 6, 5, 16, 17, 16, 10, 6, 2, 1, 10, 17, 13, 7, 0, 0, 0, 1, 0, 
    171, 0, 0, 0, 0, 7, 64, 81, 28, 29, 47, 56, 56, 54, 41, 30, 34, 28, 18, 2, 0, 0, 0, 15, 40, 46, 11, 0, 0, 0, 0, 0, 
    180, 0, 0, 0, 0, 0, 12, 30, 26, 13, 32, 35, 33, 39, 46, 64, 73, 65, 56, 29, 0, 0, 4, 33, 67, 75, 36, 0, 0, 0, 0, 0, 
    218, 87, 85, 94, 95, 97, 95, 101, 98, 87, 97, 100, 96, 95, 88, 107, 133, 146, 153, 140, 109, 102, 105, 122, 161, 176, 159, 104, 60, 72, 79, 19, 
    
    -- channel=3
    0, 2, 6, 5, 4, 4, 6, 6, 3, 4, 5, 4, 3, 6, 6, 7, 8, 7, 6, 5, 3, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=4
    0, 137, 137, 154, 161, 147, 148, 154, 151, 147, 140, 145, 148, 151, 156, 159, 160, 155, 145, 145, 146, 138, 132, 131, 137, 142, 137, 133, 133, 134, 128, 188, 
    0, 90, 82, 108, 122, 103, 109, 116, 120, 113, 102, 103, 106, 108, 117, 124, 131, 126, 104, 90, 75, 61, 51, 52, 72, 86, 102, 105, 106, 112, 107, 235, 
    0, 95, 85, 112, 124, 108, 113, 119, 123, 118, 112, 125, 146, 127, 119, 124, 127, 118, 97, 59, 64, 58, 40, 22, 17, 29, 52, 85, 101, 111, 109, 244, 
    0, 107, 99, 122, 126, 108, 108, 121, 116, 102, 82, 145, 235, 154, 104, 101, 86, 77, 45, 44, 69, 85, 77, 51, 42, 9, 18, 39, 69, 95, 106, 246, 
    0, 95, 81, 95, 118, 106, 108, 121, 115, 87, 0, 62, 190, 126, 55, 49, 49, 45, 0, 0, 34, 64, 79, 76, 55, 46, 4, 0, 14, 77, 107, 254, 
    0, 69, 26, 0, 64, 109, 116, 127, 122, 100, 0, 29, 143, 127, 102, 71, 70, 22, 0, 0, 26, 45, 45, 43, 45, 79, 38, 0, 0, 37, 102, 259, 
    0, 136, 35, 0, 6, 101, 116, 121, 125, 116, 78, 75, 83, 127, 162, 78, 37, 6, 0, 0, 31, 83, 50, 2, 34, 75, 67, 0, 0, 0, 82, 265, 
    0, 219, 86, 0, 22, 106, 114, 111, 127, 135, 132, 66, 44, 110, 142, 49, 2, 11, 0, 0, 0, 114, 74, 5, 22, 60, 67, 27, 0, 0, 40, 267, 
    0, 239, 69, 0, 85, 127, 105, 96, 111, 237, 240, 96, 27, 105, 132, 61, 2, 14, 0, 0, 0, 106, 119, 69, 34, 47, 67, 72, 0, 0, 0, 232, 
    0, 201, 0, 0, 141, 144, 90, 5, 0, 182, 255, 92, 46, 128, 144, 88, 42, 25, 9, 0, 0, 100, 145, 123, 36, 23, 60, 88, 63, 0, 0, 174, 
    0, 103, 0, 0, 166, 165, 126, 0, 0, 0, 187, 103, 75, 160, 145, 106, 67, 83, 0, 0, 0, 106, 126, 120, 12, 6, 43, 83, 103, 18, 0, 132, 
    0, 62, 0, 0, 168, 156, 157, 29, 0, 0, 111, 51, 13, 177, 181, 118, 87, 138, 0, 0, 0, 108, 126, 106, 0, 0, 26, 55, 84, 61, 7, 132, 
    0, 83, 0, 1, 142, 95, 129, 177, 0, 0, 77, 11, 0, 148, 232, 124, 69, 159, 0, 0, 14, 139, 127, 83, 1, 0, 0, 21, 65, 62, 69, 167, 
    0, 85, 0, 76, 150, 42, 70, 196, 3, 0, 25, 0, 0, 72, 162, 106, 67, 143, 0, 0, 35, 146, 126, 92, 42, 0, 0, 4, 53, 57, 74, 191, 
    0, 68, 0, 140, 197, 27, 13, 181, 69, 0, 0, 0, 68, 107, 72, 55, 68, 111, 0, 0, 32, 119, 102, 67, 14, 0, 0, 0, 44, 62, 49, 217, 
    0, 71, 0, 119, 236, 61, 0, 144, 89, 0, 0, 0, 93, 97, 29, 3, 46, 83, 0, 0, 29, 97, 102, 96, 17, 0, 0, 0, 37, 57, 49, 245, 
    0, 91, 0, 57, 235, 85, 0, 63, 135, 0, 0, 0, 27, 79, 25, 16, 29, 38, 0, 0, 0, 0, 98, 97, 0, 0, 0, 0, 52, 55, 76, 275, 
    0, 97, 0, 7, 202, 135, 0, 0, 160, 47, 0, 0, 0, 81, 45, 60, 50, 0, 6, 93, 2, 0, 57, 59, 4, 0, 0, 10, 56, 63, 94, 288, 
    0, 76, 3, 0, 143, 183, 0, 0, 75, 93, 103, 20, 0, 51, 0, 108, 114, 0, 0, 134, 60, 22, 56, 51, 0, 0, 0, 14, 71, 90, 104, 290, 
    0, 32, 26, 0, 87, 190, 22, 0, 29, 87, 129, 0, 0, 0, 0, 136, 200, 0, 0, 0, 22, 57, 25, 1, 0, 0, 0, 13, 89, 104, 96, 277, 
    0, 0, 50, 5, 61, 168, 21, 0, 102, 204, 213, 77, 22, 0, 0, 118, 233, 129, 25, 15, 11, 33, 29, 0, 0, 0, 0, 0, 53, 53, 43, 216, 
    0, 0, 58, 16, 69, 172, 0, 0, 79, 295, 234, 96, 0, 0, 0, 0, 89, 89, 67, 67, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 158, 
    0, 0, 0, 0, 81, 181, 0, 0, 0, 159, 173, 0, 0, 0, 0, 0, 0, 0, 8, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 121, 
    0, 0, 0, 0, 20, 82, 0, 0, 19, 118, 115, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 120, 
    0, 0, 0, 0, 0, 0, 0, 0, 115, 160, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 162, 
    0, 0, 0, 0, 0, 0, 0, 16, 216, 119, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 180, 
    0, 0, 0, 0, 0, 0, 0, 110, 250, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 145, 
    0, 0, 0, 0, 0, 0, 0, 79, 182, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 102, 
    0, 0, 0, 0, 0, 0, 0, 0, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 73, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 61, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 70, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    
    -- channel=5
    93, 90, 98, 95, 89, 93, 93, 92, 89, 88, 94, 94, 93, 95, 95, 95, 94, 92, 93, 89, 83, 81, 79, 83, 82, 80, 77, 75, 74, 71, 67, 7, 
    69, 18, 27, 21, 20, 28, 27, 24, 23, 24, 23, 22, 21, 22, 23, 23, 23, 21, 14, 6, 1, 0, 3, 8, 12, 18, 15, 13, 15, 13, 10, 0, 
    69, 18, 28, 25, 22, 28, 27, 23, 23, 29, 46, 38, 9, 11, 23, 23, 24, 9, 0, 4, 0, 0, 0, 0, 0, 0, 13, 16, 16, 16, 14, 0, 
    73, 24, 27, 25, 25, 30, 28, 22, 24, 34, 88, 72, 0, 5, 20, 8, 0, 0, 13, 17, 15, 4, 0, 0, 0, 0, 0, 7, 17, 14, 12, 0, 
    73, 16, 18, 23, 21, 26, 24, 20, 21, 30, 69, 51, 3, 0, 0, 0, 0, 0, 17, 39, 30, 19, 5, 5, 11, 0, 0, 0, 18, 14, 8, 0, 
    68, 0, 0, 20, 28, 23, 25, 23, 23, 26, 34, 0, 0, 0, 0, 0, 0, 0, 50, 56, 19, 0, 0, 10, 1, 0, 0, 0, 15, 21, 11, 0, 
    69, 0, 0, 3, 21, 21, 26, 29, 28, 22, 11, 8, 14, 5, 0, 10, 18, 10, 39, 60, 25, 0, 0, 0, 0, 0, 0, 0, 8, 19, 10, 0, 
    88, 0, 0, 54, 16, 11, 26, 31, 36, 13, 0, 34, 49, 18, 0, 0, 12, 0, 8, 35, 29, 0, 0, 0, 0, 0, 0, 0, 0, 25, 18, 0, 
    112, 0, 27, 69, 22, 4, 24, 62, 95, 49, 7, 31, 51, 8, 0, 0, 0, 0, 0, 33, 27, 0, 0, 0, 0, 0, 0, 0, 0, 6, 24, 0, 
    104, 0, 66, 54, 0, 0, 16, 80, 139, 84, 27, 55, 41, 0, 0, 0, 0, 0, 0, 65, 64, 11, 0, 0, 9, 8, 0, 0, 0, 0, 7, 0, 
    94, 0, 52, 46, 0, 0, 9, 41, 92, 59, 0, 14, 38, 0, 0, 0, 0, 0, 11, 115, 75, 10, 0, 0, 3, 15, 1, 0, 0, 0, 2, 0, 
    85, 0, 57, 21, 0, 0, 16, 10, 55, 12, 0, 8, 68, 12, 0, 0, 6, 0, 27, 128, 54, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 
    80, 0, 72, 0, 0, 0, 18, 0, 53, 39, 0, 28, 68, 28, 0, 0, 11, 0, 49, 116, 24, 0, 0, 0, 0, 0, 1, 6, 0, 0, 0, 0, 
    85, 0, 83, 0, 0, 0, 16, 0, 29, 43, 33, 65, 59, 4, 0, 10, 1, 0, 42, 102, 6, 0, 0, 0, 0, 2, 10, 17, 4, 0, 0, 0, 
    100, 2, 72, 0, 0, 0, 20, 0, 20, 45, 75, 105, 19, 0, 0, 0, 0, 0, 30, 75, 13, 0, 0, 0, 4, 22, 29, 23, 0, 0, 11, 0, 
    117, 2, 59, 7, 0, 0, 29, 0, 0, 48, 97, 62, 0, 0, 0, 0, 0, 0, 40, 65, 8, 0, 0, 0, 0, 7, 9, 0, 0, 4, 21, 0, 
    135, 0, 44, 22, 0, 0, 36, 25, 0, 20, 31, 0, 0, 0, 0, 0, 0, 4, 17, 0, 5, 19, 0, 0, 0, 3, 4, 0, 0, 14, 22, 0, 
    149, 6, 33, 23, 0, 0, 23, 31, 0, 0, 0, 0, 0, 0, 13, 1, 0, 24, 24, 0, 0, 0, 0, 0, 0, 0, 7, 21, 28, 32, 27, 0, 
    149, 9, 25, 24, 0, 0, 10, 27, 0, 11, 0, 0, 18, 21, 68, 29, 0, 11, 26, 16, 16, 0, 0, 0, 3, 17, 29, 42, 30, 25, 16, 0, 
    143, 19, 13, 21, 0, 0, 2, 50, 0, 0, 0, 15, 26, 46, 72, 23, 0, 0, 0, 0, 0, 0, 0, 0, 16, 25, 40, 41, 12, 5, 6, 0, 
    138, 33, 5, 21, 0, 0, 7, 114, 73, 0, 0, 9, 55, 62, 70, 25, 0, 0, 0, 0, 0, 0, 0, 2, 4, 7, 0, 1, 0, 0, 0, 0, 
    137, 44, 1, 17, 0, 0, 34, 134, 96, 50, 28, 18, 61, 62, 33, 0, 0, 0, 0, 0, 0, 0, 10, 23, 21, 8, 1, 0, 0, 0, 0, 0, 
    110, 36, 10, 22, 7, 0, 83, 142, 72, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 12, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    70, 0, 0, 27, 0, 11, 118, 120, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    65, 0, 0, 0, 0, 26, 101, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 9, 0, 
    71, 0, 0, 0, 0, 64, 110, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 12, 10, 0, 
    69, 0, 0, 0, 0, 65, 102, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    67, 0, 0, 0, 0, 30, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    73, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 18, 3, 0, 0, 0, 0, 
    76, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 8, 10, 1, 0, 0, 0, 0, 13, 36, 30, 0, 0, 0, 0, 0, 
    71, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 9, 3, 0, 0, 0, 0, 28, 38, 18, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=6
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=7
    0, 23, 24, 22, 23, 26, 25, 26, 26, 27, 26, 23, 21, 25, 28, 28, 31, 32, 30, 27, 24, 21, 19, 20, 19, 21, 20, 20, 21, 23, 23, 12, 
    0, 8, 7, 5, 8, 8, 8, 10, 10, 11, 6, 4, 5, 7, 11, 13, 15, 15, 9, 4, 0, 0, 0, 0, 0, 0, 2, 7, 8, 10, 11, 4, 
    0, 10, 8, 7, 11, 8, 8, 9, 10, 11, 8, 5, 5, 7, 12, 11, 6, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 8, 9, 3, 
    0, 11, 7, 6, 10, 9, 8, 8, 9, 9, 15, 2, 3, 7, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 6, 2, 
    0, 4, 0, 0, 7, 9, 8, 10, 11, 8, 3, 0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 3, 9, 9, 11, 12, 8, 0, 0, 9, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 5, 11, 12, 12, 11, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 0, 0, 1, 12, 12, 10, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 0, 0, 1, 10, 11, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 3, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 2, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 7, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=8
    0, 30, 32, 41, 37, 30, 34, 35, 35, 31, 31, 35, 31, 28, 29, 27, 29, 29, 30, 37, 41, 38, 35, 30, 33, 32, 30, 24, 23, 26, 27, 74, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 9, 12, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 76, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 17, 0, 0, 0, 0, 19, 15, 16, 29, 31, 17, 0, 0, 0, 0, 0, 0, 0, 1, 79, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 72, 80, 20, 0, 11, 13, 6, 6, 44, 73, 86, 68, 46, 22, 0, 0, 0, 0, 0, 0, 80, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 91, 48, 15, 4, 3, 0, 25, 64, 106, 122, 124, 95, 69, 61, 10, 0, 0, 0, 1, 82, 
    0, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 66, 62, 42, 19, 37, 36, 23, 70, 128, 135, 119, 102, 110, 88, 53, 0, 0, 0, 6, 83, 
    0, 76, 3, 0, 0, 0, 0, 0, 0, 0, 5, 3, 35, 81, 95, 69, 63, 65, 33, 63, 133, 138, 102, 93, 95, 98, 76, 15, 0, 0, 1, 86, 
    14, 129, 50, 0, 0, 0, 0, 0, 1, 35, 24, 17, 59, 109, 123, 90, 70, 78, 50, 27, 94, 140, 110, 73, 69, 88, 76, 49, 0, 0, 0, 92, 
    38, 177, 96, 55, 46, 12, 0, 0, 35, 113, 123, 82, 98, 126, 130, 92, 72, 78, 48, 0, 58, 132, 127, 87, 69, 77, 83, 66, 17, 0, 0, 88, 
    45, 190, 133, 100, 102, 34, 13, 0, 76, 186, 215, 121, 119, 145, 129, 114, 79, 75, 36, 4, 69, 133, 155, 120, 71, 77, 89, 84, 53, 0, 0, 68, 
    52, 177, 142, 128, 126, 54, 25, 15, 29, 147, 208, 152, 128, 172, 138, 116, 93, 94, 24, 8, 120, 163, 160, 123, 75, 74, 91, 91, 80, 26, 0, 41, 
    65, 178, 106, 152, 138, 58, 23, 39, 0, 97, 172, 122, 109, 192, 169, 115, 113, 117, 36, 26, 142, 184, 149, 120, 75, 63, 92, 92, 91, 62, 18, 41, 
    66, 176, 106, 176, 128, 37, 9, 54, 8, 44, 115, 100, 109, 197, 209, 137, 116, 136, 56, 38, 150, 194, 143, 112, 75, 57, 63, 88, 99, 81, 46, 70, 
    63, 180, 118, 196, 141, 22, 0, 51, 28, 18, 80, 122, 133, 181, 190, 147, 131, 132, 65, 50, 167, 180, 145, 120, 84, 69, 67, 90, 106, 88, 44, 92, 
    58, 190, 125, 207, 195, 38, 1, 51, 39, 28, 66, 133, 214, 177, 159, 140, 125, 114, 65, 57, 152, 181, 149, 116, 78, 72, 77, 83, 101, 69, 29, 103, 
    53, 207, 135, 204, 240, 94, 36, 66, 75, 28, 64, 133, 206, 174, 124, 102, 101, 100, 47, 52, 130, 162, 137, 119, 83, 62, 76, 71, 59, 37, 22, 99, 
    54, 229, 161, 202, 252, 152, 53, 94, 110, 38, 62, 80, 123, 148, 87, 97, 90, 69, 64, 61, 49, 98, 151, 113, 65, 39, 43, 50, 31, 23, 16, 100, 
    47, 247, 191, 200, 245, 202, 72, 103, 133, 105, 54, 48, 79, 97, 86, 120, 104, 57, 76, 61, 56, 77, 98, 79, 43, 21, 10, 29, 33, 20, 14, 111, 
    23, 244, 209, 202, 234, 231, 105, 88, 135, 129, 108, 49, 69, 79, 84, 154, 154, 55, 67, 111, 113, 69, 59, 62, 26, 26, 7, 13, 31, 17, 16, 106, 
    0, 214, 212, 197, 219, 233, 137, 92, 164, 153, 125, 61, 37, 72, 107, 182, 200, 94, 52, 86, 87, 75, 57, 32, 35, 23, 10, 8, 25, 17, 16, 95, 
    0, 182, 207, 186, 211, 224, 136, 94, 210, 227, 161, 125, 86, 137, 155, 200, 233, 158, 83, 69, 55, 68, 69, 62, 73, 56, 60, 48, 61, 59, 55, 101, 
    0, 159, 211, 187, 205, 209, 120, 120, 244, 326, 272, 194, 150, 157, 161, 192, 212, 170, 122, 94, 91, 93, 105, 120, 120, 116, 107, 105, 122, 123, 113, 141, 
    0, 127, 198, 191, 206, 214, 148, 155, 241, 338, 307, 181, 131, 128, 131, 140, 157, 148, 133, 140, 132, 130, 134, 144, 154, 160, 159, 165, 169, 173, 174, 169, 
    42, 116, 148, 167, 209, 187, 152, 188, 288, 295, 232, 178, 132, 126, 129, 128, 145, 154, 142, 143, 147, 155, 155, 158, 165, 178, 182, 180, 183, 187, 181, 179, 
    86, 153, 120, 129, 175, 144, 151, 232, 310, 252, 208, 167, 150, 152, 146, 145, 145, 149, 150, 151, 156, 163, 168, 170, 179, 187, 191, 191, 194, 189, 192, 215, 
    110, 203, 147, 108, 123, 127, 158, 273, 292, 230, 179, 162, 162, 158, 151, 148, 150, 152, 154, 160, 164, 172, 181, 188, 193, 188, 190, 187, 193, 208, 225, 232, 
    105, 220, 178, 135, 108, 95, 159, 296, 284, 217, 163, 160, 165, 163, 152, 149, 152, 157, 161, 163, 176, 182, 184, 192, 194, 191, 183, 183, 209, 230, 211, 203, 
    101, 220, 196, 170, 139, 84, 120, 278, 269, 186, 163, 158, 171, 174, 163, 155, 152, 155, 161, 170, 180, 182, 182, 188, 192, 192, 189, 212, 222, 211, 171, 175, 
    108, 226, 199, 186, 168, 123, 90, 201, 224, 162, 150, 152, 161, 177, 176, 162, 156, 163, 172, 177, 181, 189, 184, 174, 176, 192, 217, 233, 229, 217, 164, 150, 
    106, 225, 194, 189, 181, 161, 120, 137, 192, 147, 134, 140, 146, 155, 159, 160, 161, 170, 176, 190, 199, 190, 179, 169, 172, 194, 236, 258, 258, 216, 173, 130, 
    89, 222, 194, 182, 183, 175, 162, 142, 160, 150, 133, 133, 134, 139, 139, 133, 134, 151, 172, 196, 204, 188, 178, 164, 165, 190, 235, 266, 246, 200, 181, 133, 
    24, 118, 105, 94, 98, 96, 90, 83, 79, 82, 73, 72, 76, 74, 68, 59, 60, 71, 83, 96, 107, 103, 93, 84, 81, 91, 110, 135, 133, 112, 96, 82, 
    
    -- channel=9
    19, 4, 5, 10, 8, 2, 3, 4, 1, 0, 0, 11, 5, 0, 0, 0, 0, 0, 0, 11, 23, 26, 23, 19, 18, 18, 15, 8, 3, 6, 16, 58, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 58, 81, 74, 36, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 72, 103, 115, 108, 101, 82, 46, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 74, 96, 99, 82, 69, 72, 82, 73, 26, 0, 0, 0, 0, 0, 
    21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 72, 93, 86, 71, 71, 77, 60, 37, 41, 52, 47, 52, 25, 0, 0, 0, 0, 
    98, 67, 63, 35, 0, 0, 0, 0, 0, 0, 0, 0, 7, 46, 51, 64, 73, 71, 50, 17, 14, 35, 38, 28, 22, 47, 68, 50, 0, 0, 0, 0, 
    136, 122, 128, 108, 0, 0, 0, 0, 0, 43, 52, 45, 54, 46, 38, 53, 58, 47, 36, 19, 11, 27, 56, 55, 42, 59, 84, 83, 29, 0, 0, 0, 
    120, 105, 157, 116, 0, 0, 0, 0, 6, 81, 89, 76, 59, 34, 39, 60, 72, 55, 38, 60, 88, 69, 63, 67, 70, 76, 78, 79, 66, 8, 0, 0, 
    136, 81, 125, 93, 0, 0, 0, 0, 0, 0, 0, 9, 46, 49, 44, 58, 72, 67, 61, 104, 128, 79, 51, 38, 48, 72, 78, 82, 82, 68, 0, 0, 
    139, 88, 114, 65, 0, 0, 0, 0, 0, 0, 0, 0, 23, 58, 61, 53, 79, 97, 87, 118, 102, 41, 26, 25, 53, 54, 57, 79, 95, 94, 48, 8, 
    139, 93, 136, 75, 0, 0, 0, 0, 0, 0, 0, 0, 36, 56, 60, 64, 69, 84, 98, 124, 67, 22, 24, 34, 59, 52, 49, 73, 98, 88, 47, 25, 
    141, 97, 148, 101, 0, 0, 0, 0, 0, 0, 0, 47, 59, 14, 8, 54, 69, 55, 74, 108, 59, 36, 58, 76, 85, 82, 79, 92, 95, 61, 10, 12, 
    145, 104, 137, 98, 42, 0, 0, 0, 0, 12, 32, 106, 105, 32, 0, 7, 34, 43, 59, 72, 41, 31, 42, 51, 63, 81, 91, 79, 47, 4, 0, 0, 
    149, 111, 131, 105, 98, 60, 0, 0, 0, 5, 19, 30, 11, 0, 0, 0, 1, 15, 37, 32, 0, 26, 58, 55, 56, 64, 58, 28, 0, 0, 0, 0, 
    163, 126, 133, 112, 114, 87, 58, 19, 12, 0, 2, 0, 0, 0, 0, 16, 33, 34, 10, 0, 0, 0, 25, 35, 38, 42, 30, 5, 0, 0, 0, 0, 
    160, 129, 144, 119, 110, 108, 89, 53, 40, 38, 17, 0, 0, 3, 37, 80, 71, 43, 32, 9, 0, 0, 0, 0, 20, 35, 15, 0, 0, 0, 0, 0, 
    131, 99, 130, 118, 103, 109, 109, 69, 37, 68, 63, 11, 21, 33, 72, 127, 103, 49, 11, 19, 68, 50, 0, 11, 67, 74, 30, 0, 0, 0, 0, 0, 
    99, 70, 103, 101, 95, 102, 122, 137, 98, 47, 34, 39, 50, 53, 101, 125, 119, 74, 0, 0, 0, 6, 28, 62, 90, 73, 5, 0, 0, 0, 0, 0, 
    88, 69, 89, 86, 83, 74, 98, 165, 228, 200, 128, 138, 168, 163, 168, 132, 123, 132, 74, 14, 10, 52, 125, 165, 180, 136, 58, 12, 0, 0, 0, 6, 
    125, 114, 100, 93, 92, 85, 115, 176, 194, 222, 230, 193, 164, 147, 98, 60, 69, 84, 103, 126, 161, 192, 209, 234, 244, 216, 178, 141, 123, 132, 145, 104, 
    167, 135, 100, 112, 116, 122, 162, 200, 137, 76, 89, 97, 80, 63, 35, 34, 67, 101, 128, 174, 229, 250, 247, 243, 247, 257, 255, 239, 233, 239, 255, 177, 
    226, 157, 86, 103, 102, 91, 134, 158, 88, 49, 42, 96, 152, 159, 154, 158, 173, 193, 208, 224, 240, 247, 254, 261, 269, 280, 285, 277, 268, 273, 286, 196, 
    294, 261, 159, 108, 94, 79, 114, 113, 54, 41, 108, 201, 234, 241, 235, 233, 237, 238, 241, 253, 265, 270, 275, 287, 297, 295, 287, 287, 292, 303, 320, 230, 
    310, 316, 258, 169, 104, 109, 148, 106, 55, 84, 188, 243, 247, 241, 236, 235, 238, 245, 255, 268, 283, 293, 304, 305, 296, 278, 265, 277, 306, 326, 332, 225, 
    302, 314, 293, 246, 166, 133, 144, 107, 83, 163, 238, 247, 250, 243, 236, 239, 246, 256, 266, 277, 287, 290, 292, 296, 289, 273, 277, 303, 328, 318, 282, 159, 
    299, 315, 309, 291, 247, 165, 105, 78, 103, 191, 246, 253, 256, 262, 258, 247, 242, 251, 265, 274, 286, 291, 286, 277, 277, 294, 321, 344, 332, 274, 227, 138, 
    310, 322, 315, 307, 285, 226, 116, 58, 106, 186, 214, 233, 246, 254, 264, 264, 264, 271, 276, 279, 282, 285, 286, 279, 285, 316, 353, 368, 334, 280, 247, 170, 
    299, 313, 308, 308, 294, 269, 213, 141, 152, 216, 221, 223, 218, 216, 224, 238, 255, 272, 286, 295, 294, 284, 276, 280, 297, 329, 358, 349, 317, 297, 282, 184, 
    282, 291, 295, 296, 288, 271, 253, 228, 220, 236, 245, 246, 236, 223, 205, 196, 207, 227, 251, 271, 275, 270, 266, 272, 285, 296, 300, 294, 285, 276, 285, 189, 
    120, 65, 79, 88, 84, 78, 68, 68, 74, 81, 91, 91, 87, 91, 85, 71, 58, 50, 44, 39, 38, 50, 66, 66, 55, 31, 11, 18, 50, 82, 98, 68, 
    
    -- channel=10
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 17, 10, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    59, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    88, 11, 19, 11, 0, 0, 0, 0, 0, 7, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    111, 14, 43, 45, 0, 0, 0, 0, 0, 65, 38, 0, 15, 15, 0, 0, 0, 0, 0, 0, 41, 3, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    124, 9, 61, 56, 0, 0, 0, 0, 0, 38, 22, 0, 16, 31, 0, 0, 0, 0, 0, 0, 59, 19, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    130, 4, 65, 70, 0, 0, 0, 0, 0, 5, 0, 0, 0, 45, 0, 0, 0, 0, 0, 26, 67, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    130, 0, 68, 91, 0, 0, 0, 0, 0, 0, 0, 0, 11, 39, 11, 0, 0, 0, 0, 42, 61, 15, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    127, 9, 71, 92, 0, 0, 0, 0, 0, 0, 0, 37, 60, 23, 10, 0, 0, 0, 0, 22, 49, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    130, 28, 74, 89, 41, 0, 0, 0, 0, 0, 0, 35, 58, 29, 0, 0, 0, 0, 0, 0, 5, 10, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    138, 56, 80, 91, 77, 0, 0, 0, 0, 0, 0, 25, 21, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    138, 81, 92, 98, 95, 20, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    121, 85, 92, 99, 96, 45, 0, 36, 10, 0, 0, 0, 0, 0, 0, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    86, 82, 78, 82, 89, 60, 10, 52, 58, 0, 0, 0, 0, 0, 9, 48, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    52, 86, 65, 67, 81, 58, 5, 59, 114, 68, 1, 0, 16, 18, 53, 78, 48, 5, 0, 0, 0, 0, 0, 1, 11, 10, 0, 0, 0, 0, 0, 0, 
    45, 110, 77, 64, 79, 57, 3, 72, 120, 110, 76, 26, 50, 79, 92, 95, 79, 39, 25, 10, 9, 21, 36, 52, 73, 67, 62, 48, 36, 27, 35, 31, 
    61, 129, 109, 86, 88, 60, 14, 94, 132, 131, 87, 84, 82, 96, 95, 93, 96, 76, 61, 50, 65, 82, 92, 103, 115, 122, 124, 120, 119, 115, 120, 89, 
    98, 139, 113, 114, 104, 45, 49, 119, 136, 126, 105, 82, 88, 95, 90, 92, 95, 92, 94, 96, 108, 117, 120, 131, 136, 144, 145, 145, 146, 143, 148, 113, 
    130, 153, 118, 107, 116, 50, 72, 130, 129, 99, 92, 93, 101, 105, 100, 100, 105, 110, 111, 116, 125, 134, 136, 140, 151, 152, 152, 152, 157, 156, 166, 130, 
    145, 165, 135, 115, 100, 63, 108, 147, 114, 84, 95, 118, 118, 116, 113, 110, 108, 109, 114, 120, 132, 143, 150, 153, 155, 156, 156, 157, 173, 178, 178, 142, 
    153, 176, 151, 131, 103, 70, 151, 167, 92, 80, 109, 119, 129, 119, 110, 112, 112, 116, 121, 129, 143, 147, 158, 167, 169, 161, 158, 170, 188, 186, 180, 141, 
    153, 180, 166, 149, 127, 95, 140, 183, 74, 94, 116, 124, 129, 123, 118, 113, 115, 121, 132, 139, 148, 157, 160, 164, 163, 165, 168, 186, 194, 192, 159, 122, 
    159, 178, 171, 168, 148, 123, 122, 147, 91, 95, 109, 121, 132, 129, 127, 121, 122, 128, 134, 141, 150, 152, 155, 155, 157, 166, 181, 203, 208, 181, 129, 105, 
    155, 181, 165, 171, 159, 139, 123, 123, 90, 99, 104, 115, 119, 122, 125, 121, 122, 131, 141, 151, 149, 145, 145, 141, 148, 167, 197, 209, 192, 164, 137, 92, 
    148, 174, 156, 161, 157, 145, 123, 115, 104, 101, 101, 114, 113, 116, 108, 103, 113, 126, 137, 150, 149, 140, 135, 127, 144, 166, 194, 200, 181, 156, 144, 89, 
    51, 85, 75, 77, 74, 69, 57, 46, 46, 41, 39, 44, 42, 45, 44, 37, 37, 45, 56, 70, 70, 61, 59, 55, 64, 79, 97, 101, 90, 70, 70, 33, 
    
    -- channel=11
    155, 255, 251, 258, 263, 258, 260, 262, 262, 262, 252, 250, 259, 267, 270, 270, 267, 261, 256, 255, 252, 244, 241, 238, 239, 240, 235, 233, 230, 227, 219, 197, 
    51, 148, 138, 144, 153, 152, 159, 162, 163, 160, 149, 145, 151, 157, 159, 161, 163, 163, 155, 142, 124, 111, 103, 106, 118, 127, 141, 145, 143, 147, 148, 173, 
    58, 155, 143, 142, 149, 153, 163, 164, 167, 164, 153, 165, 186, 169, 155, 160, 160, 157, 132, 101, 102, 101, 96, 77, 74, 84, 100, 131, 148, 155, 155, 180, 
    60, 160, 157, 156, 154, 154, 159, 164, 161, 157, 153, 205, 260, 192, 149, 142, 124, 83, 67, 97, 135, 143, 134, 116, 91, 78, 95, 107, 130, 148, 153, 178, 
    53, 150, 142, 143, 150, 152, 153, 158, 156, 151, 130, 146, 184, 153, 110, 67, 39, 53, 64, 104, 135, 153, 164, 147, 133, 127, 99, 72, 93, 132, 152, 180, 
    31, 118, 93, 67, 124, 159, 160, 161, 165, 157, 88, 83, 109, 116, 104, 82, 91, 99, 71, 91, 138, 147, 125, 124, 135, 136, 102, 73, 63, 107, 147, 180, 
    28, 123, 81, 54, 115, 163, 162, 160, 164, 167, 135, 110, 111, 154, 179, 145, 131, 119, 78, 78, 134, 153, 122, 101, 110, 123, 109, 76, 53, 76, 128, 180, 
    50, 204, 130, 101, 166, 172, 159, 158, 158, 167, 153, 118, 139, 180, 183, 134, 109, 107, 73, 44, 80, 149, 140, 92, 84, 99, 116, 100, 55, 48, 108, 187, 
    53, 229, 178, 157, 211, 195, 161, 146, 166, 239, 261, 199, 153, 168, 153, 118, 93, 98, 58, 11, 57, 144, 152, 128, 103, 110, 125, 126, 86, 43, 64, 165, 
    39, 213, 145, 183, 223, 197, 151, 121, 131, 267, 284, 190, 134, 159, 150, 136, 115, 89, 78, 33, 93, 174, 186, 169, 113, 114, 137, 137, 111, 53, 40, 124, 
    13, 175, 101, 157, 222, 208, 157, 84, 4, 66, 175, 141, 131, 173, 179, 138, 129, 126, 85, 47, 150, 204, 173, 150, 100, 101, 125, 138, 134, 94, 57, 109, 
    27, 146, 57, 137, 221, 201, 177, 86, 0, 0, 120, 92, 103, 197, 210, 164, 141, 164, 109, 46, 153, 174, 149, 125, 87, 92, 111, 124, 132, 127, 102, 127, 
    27, 146, 59, 146, 189, 141, 161, 157, 42, 15, 92, 91, 118, 205, 245, 189, 155, 175, 106, 36, 139, 166, 147, 121, 90, 76, 81, 104, 136, 139, 139, 158, 
    34, 164, 78, 158, 172, 115, 133, 174, 84, 37, 99, 125, 148, 167, 180, 163, 154, 166, 73, 39, 141, 168, 151, 145, 116, 95, 105, 116, 144, 149, 149, 171, 
    34, 164, 89, 177, 196, 132, 119, 178, 119, 82, 98, 137, 195, 169, 118, 132, 124, 133, 74, 46, 120, 167, 162, 128, 102, 96, 107, 118, 136, 137, 138, 184, 
    27, 166, 99, 175, 225, 163, 111, 184, 172, 107, 54, 117, 146, 134, 97, 78, 100, 128, 83, 62, 124, 136, 143, 135, 99, 75, 82, 94, 107, 122, 143, 196, 
    16, 175, 116, 159, 228, 175, 89, 148, 189, 122, 23, 9, 52, 83, 86, 88, 103, 113, 122, 103, 48, 66, 152, 142, 73, 44, 45, 74, 119, 140, 160, 200, 
    3, 178, 130, 138, 210, 180, 95, 105, 199, 155, 77, 25, 48, 119, 121, 141, 140, 112, 117, 123, 84, 83, 84, 71, 51, 38, 63, 101, 149, 158, 158, 196, 
    0, 163, 139, 132, 195, 203, 104, 70, 145, 147, 149, 103, 77, 132, 122, 182, 187, 98, 104, 179, 153, 109, 75, 62, 64, 84, 120, 139, 162, 160, 157, 198, 
    0, 132, 151, 135, 171, 202, 123, 68, 138, 175, 139, 82, 63, 89, 126, 211, 212, 129, 84, 80, 76, 72, 65, 60, 53, 91, 115, 140, 161, 156, 148, 192, 
    0, 105, 164, 138, 157, 190, 117, 84, 186, 253, 230, 144, 150, 162, 166, 208, 236, 182, 119, 63, 35, 57, 76, 92, 78, 83, 90, 106, 117, 120, 114, 165, 
    0, 84, 167, 144, 151, 176, 114, 102, 258, 332, 325, 248, 154, 108, 92, 104, 137, 142, 116, 107, 104, 111, 123, 118, 109, 94, 74, 81, 102, 101, 93, 156, 
    0, 35, 106, 130, 161, 207, 165, 132, 203, 261, 216, 90, 9, 0, 0, 0, 8, 43, 83, 106, 112, 106, 94, 83, 79, 76, 78, 81, 90, 92, 92, 158, 
    0, 0, 15, 59, 143, 178, 118, 146, 188, 150, 84, 39, 20, 18, 19, 23, 48, 67, 75, 72, 73, 79, 74, 68, 72, 82, 90, 87, 91, 92, 89, 159, 
    0, 35, 2, 6, 65, 105, 89, 161, 177, 123, 73, 85, 87, 88, 88, 81, 78, 78, 75, 74, 74, 76, 80, 82, 88, 101, 104, 98, 96, 92, 101, 197, 
    9, 105, 44, 2, 33, 56, 97, 173, 178, 104, 74, 81, 87, 80, 73, 75, 80, 83, 85, 87, 85, 87, 95, 102, 97, 88, 80, 72, 77, 107, 131, 212, 
    0, 110, 79, 33, 28, 3, 50, 180, 202, 116, 91, 80, 80, 86, 76, 74, 80, 86, 87, 86, 86, 87, 82, 79, 80, 73, 59, 58, 91, 113, 86, 154, 
    0, 102, 90, 73, 36, 0, 0, 128, 184, 101, 87, 81, 93, 102, 94, 83, 72, 69, 71, 78, 78, 71, 67, 67, 72, 74, 80, 91, 93, 63, 31, 113, 
    0, 114, 86, 76, 64, 0, 0, 40, 98, 75, 64, 58, 77, 98, 103, 94, 80, 81, 86, 82, 83, 83, 75, 65, 67, 90, 111, 109, 95, 88, 60, 116, 
    0, 108, 83, 69, 78, 52, 2, 42, 73, 69, 50, 43, 50, 54, 67, 79, 87, 92, 95, 104, 111, 99, 82, 76, 83, 105, 126, 146, 138, 118, 71, 124, 
    0, 102, 87, 71, 74, 87, 76, 75, 83, 83, 64, 53, 48, 43, 48, 40, 37, 55, 80, 106, 117, 104, 95, 85, 76, 90, 115, 132, 117, 96, 74, 130, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 
    
    -- channel=12
    117, 162, 171, 173, 165, 160, 164, 163, 160, 158, 161, 166, 166, 169, 169, 168, 163, 157, 156, 158, 156, 151, 150, 148, 148, 141, 136, 133, 129, 121, 110, 63, 
    122, 128, 137, 144, 139, 138, 144, 142, 141, 136, 133, 141, 145, 145, 143, 140, 136, 131, 129, 125, 119, 111, 111, 113, 120, 121, 120, 113, 108, 99, 89, 47, 
    121, 123, 131, 140, 135, 139, 147, 145, 143, 142, 151, 163, 154, 142, 143, 145, 145, 135, 116, 102, 92, 81, 75, 77, 86, 95, 112, 115, 113, 107, 98, 52, 
    124, 130, 136, 146, 140, 144, 150, 148, 143, 147, 185, 234, 207, 154, 145, 144, 126, 102, 87, 99, 117, 116, 99, 76, 62, 63, 78, 101, 116, 114, 105, 57, 
    128, 136, 141, 149, 142, 140, 143, 142, 137, 140, 181, 259, 226, 146, 115, 96, 62, 41, 65, 131, 155, 158, 144, 121, 102, 82, 69, 75, 103, 116, 108, 57, 
    120, 109, 91, 114, 140, 142, 142, 141, 138, 135, 132, 157, 128, 105, 67, 34, 33, 47, 95, 157, 171, 160, 142, 130, 120, 100, 49, 40, 80, 119, 117, 64, 
    110, 83, 24, 53, 127, 149, 144, 147, 148, 142, 125, 122, 120, 129, 107, 78, 86, 80, 102, 169, 197, 160, 121, 116, 120, 89, 46, 30, 52, 101, 116, 65, 
    138, 112, 51, 95, 148, 150, 141, 148, 160, 152, 121, 123, 155, 176, 140, 99, 102, 92, 86, 138, 192, 172, 120, 100, 95, 70, 45, 23, 29, 77, 113, 70, 
    192, 163, 113, 181, 205, 161, 144, 168, 215, 231, 182, 167, 207, 203, 144, 92, 81, 75, 61, 87, 154, 175, 139, 98, 77, 78, 67, 44, 12, 39, 99, 75, 
    214, 201, 187, 246, 231, 170, 140, 174, 292, 371, 315, 250, 235, 198, 147, 106, 83, 61, 42, 88, 182, 200, 174, 126, 98, 97, 88, 71, 28, 11, 55, 55, 
    209, 189, 213, 274, 242, 170, 135, 128, 240, 336, 306, 237, 246, 214, 163, 128, 97, 61, 45, 136, 250, 239, 196, 128, 96, 111, 105, 82, 51, 21, 33, 26, 
    216, 169, 210, 266, 252, 185, 153, 96, 125, 217, 242, 209, 258, 259, 192, 146, 120, 93, 60, 184, 292, 236, 175, 104, 82, 102, 109, 99, 79, 57, 46, 16, 
    216, 160, 209, 261, 224, 172, 163, 115, 89, 180, 195, 186, 258, 306, 238, 175, 154, 131, 96, 210, 279, 208, 150, 94, 82, 84, 95, 98, 100, 86, 77, 26, 
    221, 174, 237, 266, 172, 132, 158, 130, 78, 150, 190, 231, 286, 305, 251, 202, 168, 131, 103, 221, 262, 203, 150, 105, 85, 80, 95, 118, 127, 106, 97, 47, 
    235, 199, 256, 272, 165, 127, 156, 141, 85, 133, 197, 300, 304, 245, 193, 188, 171, 125, 100, 203, 244, 197, 157, 123, 100, 106, 124, 141, 138, 108, 100, 62, 
    250, 227, 268, 280, 198, 140, 170, 167, 116, 143, 210, 315, 315, 221, 158, 149, 130, 112, 114, 184, 212, 190, 151, 96, 68, 91, 116, 124, 117, 101, 109, 77, 
    267, 256, 275, 294, 241, 149, 174, 196, 147, 118, 155, 200, 176, 130, 125, 117, 111, 120, 130, 150, 151, 171, 159, 111, 67, 68, 89, 100, 102, 112, 135, 85, 
    280, 282, 281, 294, 263, 153, 152, 204, 203, 133, 128, 111, 117, 120, 125, 135, 112, 138, 165, 130, 69, 105, 110, 54, 18, 27, 61, 103, 128, 144, 147, 85, 
    271, 289, 283, 288, 274, 186, 143, 190, 208, 178, 132, 82, 130, 156, 181, 203, 133, 123, 178, 172, 137, 110, 48, 14, 24, 54, 89, 132, 152, 151, 137, 81, 
    241, 283, 278, 280, 275, 210, 146, 182, 196, 177, 150, 95, 129, 157, 218, 260, 177, 113, 129, 130, 117, 73, 18, 13, 36, 95, 136, 167, 165, 148, 135, 81, 
    199, 279, 281, 276, 268, 212, 156, 234, 292, 226, 148, 115, 170, 212, 287, 304, 231, 155, 108, 48, 22, 12, 19, 31, 48, 94, 126, 158, 153, 134, 127, 73, 
    158, 283, 291, 277, 263, 199, 158, 278, 413, 393, 299, 234, 249, 277, 295, 280, 233, 179, 134, 77, 40, 52, 79, 99, 113, 115, 127, 135, 131, 117, 111, 66, 
    114, 260, 286, 286, 275, 233, 231, 356, 434, 398, 294, 203, 152, 148, 141, 135, 118, 94, 92, 84, 94, 102, 104, 106, 110, 108, 111, 119, 125, 114, 108, 74, 
    60, 161, 210, 265, 278, 263, 302, 410, 404, 301, 161, 75, 67, 66, 60, 61, 65, 72, 81, 78, 86, 94, 95, 95, 100, 109, 113, 116, 116, 109, 111, 77, 
    52, 95, 118, 190, 235, 236, 314, 406, 340, 200, 94, 86, 95, 96, 93, 88, 84, 81, 77, 75, 81, 89, 93, 101, 114, 128, 132, 130, 128, 125, 134, 103, 
    76, 110, 97, 128, 179, 233, 356, 386, 258, 110, 80, 100, 101, 96, 89, 85, 81, 79, 80, 85, 93, 103, 112, 122, 130, 134, 128, 126, 136, 152, 174, 143, 
    80, 112, 96, 95, 125, 211, 362, 355, 198, 92, 97, 103, 104, 89, 83, 87, 89, 91, 93, 100, 104, 109, 124, 131, 125, 108, 99, 110, 143, 167, 170, 121, 
    76, 110, 101, 99, 102, 154, 285, 303, 161, 107, 106, 106, 110, 102, 91, 87, 87, 92, 98, 104, 106, 102, 102, 107, 108, 101, 106, 129, 153, 136, 102, 69, 
    82, 111, 101, 103, 101, 100, 161, 188, 109, 80, 89, 100, 117, 119, 112, 100, 91, 93, 100, 105, 105, 99, 97, 94, 99, 117, 141, 159, 139, 89, 56, 57, 
    96, 121, 99, 101, 102, 93, 87, 98, 58, 57, 53, 65, 83, 95, 104, 105, 112, 121, 128, 128, 118, 103, 92, 90, 114, 158, 191, 187, 144, 102, 67, 53, 
    89, 118, 98, 99, 99, 101, 91, 85, 68, 56, 51, 56, 54, 53, 56, 68, 89, 111, 132, 150, 141, 114, 98, 101, 137, 184, 216, 193, 134, 89, 69, 43, 
    21, 42, 29, 26, 23, 26, 24, 16, 12, 0, 0, 2, 0, 0, 0, 0, 0, 16, 39, 56, 51, 36, 31, 31, 51, 79, 94, 74, 36, 10, 14, 2, 
    
    -- channel=13
    162, 129, 139, 135, 125, 127, 127, 125, 121, 117, 125, 133, 136, 134, 131, 127, 119, 114, 118, 118, 112, 112, 113, 116, 113, 107, 104, 103, 97, 84, 74, 0, 
    182, 105, 119, 117, 111, 117, 116, 112, 106, 103, 109, 120, 122, 117, 111, 107, 98, 92, 87, 83, 81, 81, 91, 97, 101, 105, 97, 88, 81, 69, 58, 0, 
    177, 97, 114, 117, 111, 117, 118, 112, 109, 112, 138, 146, 113, 104, 110, 109, 106, 85, 69, 77, 67, 59, 54, 65, 77, 88, 103, 95, 86, 76, 66, 0, 
    179, 100, 116, 120, 114, 120, 121, 113, 112, 124, 203, 215, 117, 98, 111, 101, 76, 62, 86, 101, 103, 92, 76, 60, 51, 67, 73, 91, 97, 85, 71, 0, 
    179, 100, 117, 128, 115, 116, 115, 109, 107, 120, 203, 217, 136, 83, 70, 60, 45, 45, 100, 150, 152, 138, 111, 92, 90, 54, 51, 80, 107, 97, 77, 0, 
    169, 60, 61, 125, 132, 114, 114, 109, 107, 109, 142, 137, 73, 58, 28, 23, 26, 56, 145, 195, 166, 133, 116, 119, 98, 54, 21, 45, 106, 116, 88, 0, 
    169, 17, 7, 93, 133, 118, 113, 116, 111, 100, 92, 98, 110, 95, 52, 62, 78, 76, 144, 214, 186, 117, 99, 113, 95, 46, 8, 30, 86, 120, 97, 0, 
    202, 20, 38, 147, 138, 112, 111, 120, 128, 99, 72, 125, 164, 139, 80, 75, 93, 79, 108, 185, 199, 126, 85, 88, 83, 47, 19, 1, 50, 116, 112, 0, 
    260, 75, 115, 206, 163, 109, 110, 160, 229, 185, 122, 156, 205, 158, 90, 70, 76, 56, 64, 156, 191, 139, 98, 73, 68, 65, 46, 12, 4, 73, 117, 0, 
    286, 125, 214, 246, 157, 108, 100, 199, 343, 321, 220, 230, 229, 153, 103, 78, 64, 42, 44, 173, 228, 173, 119, 74, 92, 93, 63, 32, 0, 32, 88, 0, 
    282, 145, 245, 271, 161, 107, 91, 155, 316, 354, 235, 223, 247, 168, 115, 92, 77, 17, 68, 251, 268, 192, 130, 71, 94, 111, 87, 47, 12, 17, 62, 0, 
    275, 133, 268, 261, 166, 126, 109, 87, 222, 273, 193, 212, 291, 208, 124, 108, 99, 35, 96, 304, 279, 176, 107, 60, 84, 108, 91, 76, 52, 43, 46, 0, 
    270, 132, 284, 231, 133, 136, 131, 59, 152, 237, 176, 218, 299, 256, 145, 128, 130, 62, 141, 315, 257, 135, 87, 58, 76, 90, 98, 98, 81, 71, 56, 0, 
    278, 154, 306, 204, 85, 115, 143, 63, 99, 193, 207, 259, 297, 246, 178, 167, 138, 63, 153, 310, 230, 137, 104, 70, 71, 87, 106, 123, 109, 81, 71, 0, 
    303, 184, 308, 202, 67, 110, 155, 77, 84, 166, 255, 341, 264, 178, 159, 156, 134, 84, 150, 274, 223, 141, 99, 80, 91, 115, 137, 147, 112, 82, 89, 0, 
    334, 205, 306, 238, 89, 105, 174, 117, 85, 155, 289, 329, 241, 167, 136, 135, 110, 86, 160, 240, 193, 150, 110, 55, 59, 107, 127, 125, 98, 92, 99, 0, 
    370, 223, 298, 275, 132, 96, 190, 181, 88, 129, 201, 218, 149, 89, 113, 103, 96, 121, 146, 128, 150, 174, 102, 49, 59, 89, 112, 109, 98, 108, 110, 0, 
    398, 245, 288, 287, 172, 87, 179, 209, 137, 110, 123, 126, 133, 98, 127, 109, 85, 153, 158, 95, 85, 99, 60, 20, 19, 63, 99, 122, 127, 130, 118, 0, 
    404, 256, 276, 284, 206, 97, 153, 212, 170, 150, 87, 90, 146, 146, 209, 164, 75, 142, 176, 128, 111, 75, 16, 0, 47, 89, 123, 146, 132, 121, 102, 0, 
    386, 270, 260, 272, 228, 119, 142, 229, 179, 119, 83, 110, 152, 192, 263, 208, 96, 103, 123, 104, 75, 31, 0, 14, 71, 119, 157, 162, 124, 103, 96, 0, 
    357, 289, 252, 267, 228, 119, 155, 319, 289, 159, 81, 119, 199, 246, 305, 257, 142, 103, 81, 19, 8, 3, 20, 48, 72, 108, 125, 133, 105, 86, 83, 0, 
    329, 313, 258, 265, 223, 121, 197, 391, 394, 283, 202, 177, 247, 287, 290, 243, 162, 115, 86, 50, 35, 53, 78, 102, 115, 114, 123, 126, 102, 87, 91, 0, 
    270, 304, 278, 280, 243, 175, 285, 440, 420, 276, 151, 154, 161, 162, 151, 133, 101, 78, 68, 65, 89, 103, 109, 111, 113, 114, 117, 122, 116, 106, 103, 0, 
    185, 206, 239, 293, 250, 231, 374, 450, 340, 172, 71, 52, 80, 83, 75, 78, 70, 69, 78, 82, 94, 98, 101, 107, 115, 122, 121, 120, 114, 107, 111, 0, 
    147, 116, 166, 240, 231, 265, 396, 397, 213, 83, 55, 78, 99, 98, 94, 93, 91, 82, 79, 84, 91, 96, 101, 114, 132, 135, 132, 129, 125, 132, 151, 2, 
    155, 93, 120, 176, 200, 310, 430, 323, 111, 42, 74, 107, 103, 96, 94, 90, 84, 80, 84, 91, 101, 113, 122, 130, 132, 131, 124, 130, 151, 169, 178, 16, 
    163, 88, 95, 121, 167, 317, 439, 252, 63, 52, 98, 109, 106, 86, 86, 94, 94, 95, 99, 107, 111, 115, 132, 138, 123, 103, 103, 139, 166, 163, 160, 8, 
    164, 92, 94, 105, 133, 256, 363, 210, 47, 85, 106, 118, 111, 96, 91, 88, 94, 102, 111, 114, 111, 110, 113, 112, 106, 103, 126, 152, 152, 118, 108, 0, 
    173, 91, 98, 109, 112, 159, 230, 135, 46, 68, 91, 116, 125, 116, 105, 100, 104, 108, 111, 113, 110, 101, 99, 103, 115, 137, 162, 161, 126, 57, 67, 0, 
    183, 99, 101, 111, 108, 107, 127, 88, 28, 50, 66, 83, 93, 101, 106, 111, 124, 132, 140, 133, 111, 96, 92, 105, 145, 192, 205, 164, 100, 63, 74, 0, 
    184, 100, 100, 109, 106, 99, 89, 85, 53, 47, 61, 69, 67, 65, 62, 81, 112, 132, 150, 150, 122, 103, 95, 118, 175, 222, 217, 153, 86, 70, 65, 0, 
    85, 52, 50, 53, 47, 43, 35, 31, 24, 13, 20, 22, 21, 19, 13, 16, 30, 49, 70, 73, 56, 46, 45, 62, 92, 118, 113, 69, 31, 27, 28, 0, 
    
    -- channel=14
    61, 63, 64, 58, 57, 61, 61, 60, 60, 64, 59, 58, 64, 66, 71, 72, 68, 65, 62, 56, 50, 49, 49, 52, 48, 45, 46, 49, 48, 43, 37, 0, 
    151, 175, 181, 176, 174, 176, 178, 175, 174, 171, 168, 172, 180, 185, 191, 191, 181, 172, 165, 161, 150, 148, 149, 151, 152, 147, 145, 147, 147, 139, 128, 21, 
    151, 171, 179, 177, 176, 180, 180, 178, 177, 172, 167, 156, 165, 180, 184, 180, 174, 156, 150, 130, 111, 100, 108, 124, 132, 151, 149, 146, 146, 141, 130, 20, 
    149, 166, 174, 179, 180, 186, 184, 182, 182, 183, 192, 151, 144, 162, 170, 162, 160, 149, 120, 92, 71, 54, 49, 59, 81, 103, 132, 144, 146, 142, 136, 23, 
    140, 162, 173, 183, 183, 187, 188, 183, 185, 190, 230, 225, 162, 145, 152, 148, 117, 100, 95, 87, 74, 59, 39, 39, 38, 52, 90, 128, 142, 137, 134, 24, 
    127, 133, 169, 189, 181, 183, 187, 182, 182, 190, 219, 226, 167, 115, 91, 84, 57, 58, 94, 99, 88, 82, 72, 60, 47, 40, 39, 90, 134, 137, 132, 25, 
    98, 76, 94, 156, 175, 181, 188, 186, 180, 178, 173, 168, 139, 89, 48, 42, 39, 45, 99, 126, 99, 83, 84, 82, 70, 38, 23, 43, 110, 140, 134, 25, 
    73, 32, 34, 91, 150, 177, 186, 183, 175, 147, 147, 136, 123, 95, 60, 58, 58, 48, 86, 153, 133, 80, 73, 89, 77, 42, 18, 16, 75, 136, 135, 22, 
    94, 19, 37, 89, 123, 162, 179, 183, 159, 107, 80, 118, 128, 109, 69, 60, 61, 54, 70, 128, 140, 98, 62, 61, 65, 48, 21, 1, 32, 116, 143, 21, 
    124, 65, 66, 121, 125, 154, 165, 204, 198, 151, 94, 126, 134, 105, 76, 47, 55, 38, 54, 101, 117, 108, 66, 52, 59, 52, 39, 11, 2, 62, 130, 29, 
    127, 100, 120, 141, 129, 148, 146, 195, 276, 227, 152, 147, 147, 95, 84, 63, 44, 22, 53, 113, 118, 117, 87, 64, 69, 69, 46, 25, 0, 16, 80, 24, 
    119, 100, 148, 151, 137, 152, 148, 146, 237, 229, 167, 175, 174, 109, 82, 78, 52, 6, 61, 146, 151, 124, 96, 61, 68, 82, 62, 39, 11, 8, 39, 0, 
    116, 89, 140, 140, 148, 165, 165, 116, 167, 195, 155, 162, 199, 145, 87, 83, 79, 24, 74, 168, 158, 114, 83, 58, 59, 77, 76, 53, 33, 29, 36, 0, 
    114, 89, 145, 115, 108, 160, 174, 120, 144, 172, 149, 151, 197, 187, 127, 96, 87, 53, 98, 169, 146, 106, 66, 45, 49, 54, 66, 67, 52, 54, 65, 0, 
    124, 98, 159, 104, 54, 124, 158, 120, 122, 141, 167, 170, 150, 167, 141, 123, 100, 60, 105, 174, 146, 98, 81, 60, 58, 60, 69, 86, 78, 81, 90, 0, 
    138, 107, 161, 116, 35, 83, 127, 116, 106, 149, 180, 225, 176, 125, 131, 121, 105, 76, 116, 162, 155, 109, 74, 52, 58, 77, 85, 101, 103, 99, 109, 10, 
    152, 112, 155, 140, 53, 58, 123, 111, 92, 129, 186, 219, 183, 122, 111, 92, 94, 90, 108, 158, 181, 134, 75, 57, 55, 77, 93, 93, 101, 113, 130, 20, 
    177, 119, 146, 155, 81, 41, 114, 124, 80, 87, 140, 151, 121, 101, 91, 66, 75, 102, 102, 103, 119, 137, 100, 53, 50, 60, 91, 97, 109, 138, 152, 28, 
    203, 140, 146, 156, 104, 37, 92, 132, 110, 80, 59, 105, 103, 103, 107, 62, 48, 114, 117, 80, 69, 84, 69, 31, 32, 46, 86, 119, 137, 154, 157, 30, 
    219, 160, 151, 158, 122, 53, 72, 111, 88, 101, 61, 76, 114, 111, 132, 96, 35, 77, 128, 121, 100, 52, 26, 24, 31, 72, 103, 145, 156, 160, 154, 33, 
    216, 170, 154, 160, 134, 75, 88, 125, 71, 35, 43, 45, 74, 101, 145, 122, 53, 40, 63, 82, 65, 26, 0, 0, 14, 55, 90, 128, 126, 120, 118, 18, 
    190, 172, 147, 156, 134, 76, 101, 166, 154, 60, 20, 64, 102, 140, 173, 152, 100, 63, 34, 10, 0, 0, 0, 0, 0, 18, 48, 68, 64, 56, 51, 0, 
    154, 178, 147, 149, 129, 75, 118, 204, 229, 163, 109, 99, 124, 142, 145, 133, 94, 55, 27, 3, 0, 0, 1, 8, 5, 3, 12, 19, 15, 6, 1, 0, 
    95, 135, 158, 155, 135, 130, 174, 231, 217, 173, 102, 52, 47, 46, 44, 41, 28, 10, 3, 4, 4, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    30, 33, 102, 154, 137, 158, 212, 231, 180, 114, 35, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 0, 20, 98, 126, 157, 221, 203, 127, 47, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 9, 7, 10, 3, 0, 4, 0, 
    32, 0, 0, 22, 82, 180, 227, 160, 70, 13, 6, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 3, 4, 14, 34, 0, 
    34, 0, 0, 0, 24, 151, 238, 128, 50, 17, 5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 12, 17, 27, 0, 
    27, 0, 0, 0, 0, 65, 177, 123, 33, 22, 14, 13, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    39, 0, 0, 0, 0, 0, 57, 66, 10, 0, 2, 10, 18, 18, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 0, 0, 0, 0, 0, 
    51, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 1, 8, 17, 24, 24, 22, 11, 0, 0, 0, 0, 20, 45, 43, 12, 0, 0, 0, 0, 
    91, 37, 29, 34, 33, 32, 28, 27, 22, 10, 12, 15, 14, 14, 15, 26, 45, 61, 76, 77, 59, 43, 38, 50, 82, 113, 117, 80, 33, 16, 9, 0, 
    
    -- channel=15
    45, 26, 30, 27, 23, 26, 27, 25, 25, 25, 27, 30, 28, 27, 31, 29, 26, 27, 27, 25, 23, 23, 22, 23, 22, 21, 23, 23, 22, 20, 16, 0, 
    129, 123, 134, 136, 129, 127, 128, 127, 124, 124, 127, 132, 133, 132, 135, 137, 134, 129, 125, 119, 113, 112, 112, 116, 117, 113, 110, 111, 112, 104, 95, 36, 
    125, 118, 129, 137, 135, 132, 130, 129, 129, 124, 123, 128, 130, 132, 138, 140, 134, 122, 105, 100, 92, 90, 97, 104, 114, 117, 113, 110, 110, 103, 93, 35, 
    127, 121, 129, 138, 136, 136, 133, 131, 130, 130, 138, 131, 109, 119, 134, 133, 127, 106, 97, 86, 68, 52, 49, 67, 75, 96, 109, 110, 108, 104, 97, 36, 
    130, 127, 126, 134, 134, 137, 136, 133, 133, 135, 166, 157, 105, 106, 119, 111, 95, 97, 91, 77, 58, 47, 37, 30, 44, 51, 70, 98, 108, 104, 99, 41, 
    122, 114, 117, 130, 131, 132, 136, 133, 132, 130, 134, 174, 137, 96, 80, 84, 72, 57, 69, 77, 64, 57, 47, 49, 41, 32, 39, 73, 105, 109, 99, 41, 
    109, 68, 74, 124, 131, 128, 135, 136, 132, 129, 118, 122, 117, 86, 47, 36, 36, 32, 66, 88, 68, 54, 62, 64, 51, 39, 22, 37, 88, 114, 104, 43, 
    92, 37, 22, 81, 114, 124, 133, 138, 137, 125, 106, 103, 102, 77, 44, 36, 41, 31, 55, 102, 96, 60, 56, 64, 63, 37, 25, 24, 61, 108, 108, 40, 
    96, 20, 33, 70, 87, 114, 131, 133, 138, 102, 81, 93, 95, 77, 50, 42, 51, 46, 41, 90, 123, 81, 47, 52, 59, 44, 21, 14, 36, 93, 112, 38, 
    128, 35, 41, 89, 89, 102, 123, 149, 160, 119, 58, 76, 101, 85, 63, 44, 39, 38, 45, 77, 103, 87, 59, 37, 44, 47, 34, 18, 10, 56, 110, 46, 
    123, 65, 76, 95, 94, 100, 108, 141, 186, 165, 114, 106, 118, 83, 71, 47, 38, 28, 37, 92, 99, 78, 65, 42, 53, 50, 36, 29, 17, 22, 73, 45, 
    121, 46, 101, 112, 98, 100, 109, 86, 170, 193, 136, 121, 138, 92, 57, 65, 41, 20, 40, 111, 108, 75, 71, 47, 52, 65, 46, 33, 23, 18, 37, 24, 
    121, 39, 103, 111, 104, 114, 124, 86, 109, 159, 118, 130, 152, 115, 56, 59, 62, 26, 38, 115, 118, 76, 65, 46, 45, 55, 56, 45, 35, 27, 34, 6, 
    124, 45, 102, 87, 86, 123, 132, 97, 88, 133, 121, 115, 136, 131, 78, 60, 64, 49, 51, 120, 108, 70, 53, 41, 39, 45, 57, 52, 41, 37, 46, 5, 
    130, 52, 111, 88, 48, 90, 126, 95, 73, 114, 125, 126, 103, 114, 109, 88, 62, 48, 65, 121, 103, 76, 59, 37, 39, 45, 47, 58, 52, 45, 67, 19, 
    143, 62, 112, 96, 35, 57, 111, 90, 64, 88, 133, 156, 92, 73, 87, 88, 82, 57, 58, 115, 114, 72, 54, 48, 48, 61, 61, 64, 65, 70, 83, 31, 
    151, 71, 111, 105, 43, 38, 96, 89, 46, 87, 124, 137, 140, 85, 79, 81, 68, 62, 78, 104, 111, 103, 60, 33, 35, 56, 66, 67, 81, 92, 98, 38, 
    159, 76, 103, 110, 63, 17, 87, 102, 63, 49, 92, 105, 106, 84, 74, 62, 53, 80, 69, 71, 103, 113, 65, 45, 43, 51, 69, 81, 89, 101, 108, 42, 
    169, 88, 93, 103, 78, 23, 57, 112, 87, 45, 52, 85, 93, 73, 78, 53, 29, 75, 95, 66, 39, 51, 64, 41, 36, 42, 58, 94, 98, 108, 112, 47, 
    170, 104, 93, 101, 89, 39, 40, 88, 92, 79, 38, 50, 91, 88, 106, 73, 16, 53, 101, 89, 62, 38, 33, 33, 39, 57, 70, 106, 115, 117, 114, 45, 
    166, 121, 93, 105, 97, 54, 45, 94, 57, 38, 59, 43, 79, 92, 100, 90, 43, 20, 57, 67, 66, 43, 14, 18, 25, 61, 86, 105, 104, 100, 96, 32, 
    150, 127, 93, 104, 94, 52, 61, 129, 118, 28, 16, 39, 61, 80, 104, 102, 70, 41, 22, 17, 16, 12, 9, 0, 2, 25, 45, 59, 58, 45, 46, 0, 
    119, 118, 94, 99, 91, 55, 71, 127, 147, 118, 38, 36, 74, 91, 103, 100, 75, 52, 41, 13, 0, 0, 0, 3, 1, 0, 5, 6, 3, 0, 0, 0, 
    68, 91, 102, 103, 96, 76, 96, 143, 137, 94, 63, 39, 38, 45, 45, 44, 36, 15, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 10, 72, 105, 88, 100, 140, 157, 107, 62, 29, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 0, 64, 91, 103, 147, 130, 68, 31, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 0, 0, 7, 69, 113, 148, 99, 37, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 0, 0, 0, 12, 97, 150, 89, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 0, 0, 0, 0, 28, 119, 84, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 0, 0, 0, 0, 0, 26, 58, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 6, 4, 0, 0, 0, 0, 0, 0, 11, 7, 0, 0, 0, 0, 0, 
    47, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 20, 25, 28, 24, 12, 5, 1, 9, 28, 41, 44, 20, 0, 0, 0, 0, 
    
    -- channel=16
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=17
    0, 56, 55, 55, 55, 55, 55, 55, 55, 55, 55, 56, 56, 56, 56, 56, 55, 55, 56, 55, 56, 58, 58, 55, 54, 55, 56, 55, 55, 55, 56, 59, 
    3, 50, 50, 50, 50, 50, 50, 50, 50, 49, 49, 50, 50, 50, 50, 50, 48, 46, 48, 49, 51, 53, 52, 50, 49, 49, 50, 50, 50, 50, 50, 55, 
    3, 51, 50, 50, 50, 50, 50, 50, 50, 49, 50, 49, 49, 49, 50, 49, 46, 44, 46, 45, 42, 45, 47, 49, 50, 49, 49, 49, 49, 50, 50, 55, 
    3, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 49, 50, 50, 49, 47, 47, 48, 41, 41, 46, 46, 50, 51, 50, 50, 50, 50, 50, 56, 
    3, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 46, 41, 42, 46, 52, 43, 39, 44, 50, 52, 51, 50, 50, 50, 51, 51, 56, 
    0, 47, 48, 48, 49, 50, 50, 50, 50, 50, 50, 49, 49, 50, 51, 48, 43, 41, 44, 46, 36, 32, 33, 45, 53, 51, 48, 49, 50, 51, 51, 57, 
    0, 49, 50, 50, 49, 50, 50, 49, 50, 51, 50, 48, 44, 46, 49, 52, 55, 56, 56, 57, 53, 46, 37, 37, 50, 53, 50, 51, 52, 52, 51, 57, 
    8, 56, 60, 60, 56, 53, 50, 48, 49, 50, 50, 52, 43, 38, 49, 54, 53, 61, 68, 70, 71, 71, 65, 57, 56, 57, 55, 55, 55, 54, 52, 57, 
    0, 26, 29, 35, 46, 53, 50, 46, 47, 49, 50, 54, 45, 39, 47, 52, 56, 58, 64, 68, 70, 69, 62, 55, 47, 38, 39, 47, 55, 55, 53, 58, 
    0, 20, 18, 17, 24, 41, 46, 43, 46, 49, 50, 54, 49, 49, 50, 52, 55, 57, 61, 58, 53, 51, 46, 40, 33, 25, 21, 28, 45, 55, 53, 58, 
    24, 62, 60, 56, 43, 43, 42, 33, 36, 44, 46, 45, 46, 50, 53, 55, 55, 58, 61, 63, 63, 60, 56, 52, 50, 45, 37, 34, 44, 55, 54, 59, 
    8, 65, 65, 67, 66, 61, 40, 22, 26, 33, 23, 8, 9, 14, 17, 21, 27, 39, 56, 69, 71, 67, 67, 65, 66, 70, 58, 49, 57, 57, 57, 62, 
    0, 30, 25, 26, 38, 50, 48, 44, 40, 43, 38, 13, 0, 0, 0, 2, 16, 32, 48, 61, 63, 64, 63, 56, 57, 60, 51, 47, 49, 48, 52, 62, 
    0, 16, 8, 9, 20, 22, 30, 40, 52, 63, 62, 42, 27, 32, 42, 48, 45, 41, 45, 46, 39, 34, 29, 23, 17, 15, 20, 28, 25, 27, 40, 56, 
    0, 14, 25, 22, 13, 12, 5, 11, 36, 55, 64, 60, 60, 59, 54, 48, 40, 33, 29, 22, 19, 14, 11, 10, 9, 9, 17, 26, 30, 33, 41, 53, 
    0, 0, 25, 39, 37, 18, 0, 8, 27, 44, 55, 58, 62, 61, 61, 52, 36, 29, 30, 35, 41, 40, 38, 37, 40, 41, 45, 50, 52, 47, 46, 52, 
    0, 0, 18, 60, 70, 42, 32, 37, 43, 51, 58, 57, 54, 60, 71, 71, 58, 54, 58, 62, 67, 71, 69, 65, 62, 57, 49, 45, 44, 43, 43, 42, 
    0, 2, 29, 60, 56, 53, 51, 51, 52, 58, 61, 58, 50, 45, 48, 46, 53, 55, 49, 46, 49, 53, 52, 47, 39, 35, 37, 34, 32, 33, 32, 33, 
    0, 26, 55, 53, 47, 50, 54, 55, 53, 54, 55, 55, 50, 53, 51, 42, 40, 44, 53, 45, 37, 40, 44, 41, 36, 33, 33, 30, 26, 27, 30, 34, 
    0, 24, 35, 34, 38, 44, 48, 50, 52, 54, 56, 57, 61, 70, 69, 60, 51, 51, 54, 48, 44, 46, 43, 37, 34, 34, 32, 27, 27, 28, 28, 29, 
    0, 0, 0, 0, 0, 2, 7, 10, 10, 11, 15, 19, 30, 41, 44, 44, 44, 42, 37, 32, 32, 32, 28, 23, 23, 30, 32, 27, 21, 19, 20, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 10, 13, 17, 16, 15, 15, 14, 14, 16, 23, 30, 32, 23, 14, 12, 14, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 8, 3, 0, 4, 7, 9, 13, 16, 20, 29, 33, 25, 16, 11, 8, 7, 9, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 52, 44, 34, 31, 29, 29, 29, 26, 24, 17, 4, 0, 0, 0, 0, 4, 12, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 34, 28, 24, 19, 12, 1, 0, 0, 0, 0, 0, 0, 0, 0, 9, 17, 32, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 14, 24, 37, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 20, 31, 40, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 20, 32, 42, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 13, 24, 32, 42, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 16, 27, 35, 44, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 8, 15, 24, 35, 43, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=18
    351, 49, 54, 53, 53, 53, 53, 53, 53, 54, 54, 53, 53, 53, 53, 52, 52, 54, 54, 53, 52, 50, 52, 55, 56, 54, 52, 53, 54, 54, 52, 0, 
    450, 143, 147, 147, 147, 147, 147, 147, 147, 148, 148, 148, 148, 148, 147, 146, 147, 150, 149, 144, 145, 143, 145, 148, 150, 148, 146, 147, 148, 148, 146, 0, 
    451, 143, 147, 147, 147, 147, 147, 147, 147, 148, 148, 148, 148, 149, 149, 147, 149, 152, 150, 132, 155, 166, 161, 163, 151, 148, 148, 148, 149, 149, 147, 0, 
    452, 144, 148, 147, 147, 147, 147, 146, 146, 148, 147, 146, 147, 148, 148, 146, 145, 140, 133, 100, 137, 185, 163, 171, 152, 144, 147, 147, 148, 148, 147, 0, 
    451, 144, 148, 147, 147, 147, 147, 146, 146, 148, 148, 145, 144, 148, 146, 141, 146, 144, 127, 91, 120, 186, 174, 166, 152, 145, 147, 148, 148, 147, 147, 0, 
    454, 150, 151, 151, 152, 149, 147, 146, 146, 148, 148, 140, 141, 153, 144, 114, 112, 131, 125, 100, 121, 176, 206, 201, 166, 147, 150, 150, 150, 149, 148, 0, 
    447, 155, 146, 145, 154, 154, 150, 149, 146, 146, 148, 127, 141, 172, 145, 98, 82, 94, 93, 77, 79, 113, 172, 220, 187, 146, 148, 149, 149, 149, 148, 0, 
    430, 147, 137, 134, 145, 152, 153, 152, 149, 146, 148, 107, 127, 191, 151, 97, 94, 103, 83, 64, 60, 66, 101, 157, 170, 145, 147, 147, 149, 150, 148, 0, 
    438, 195, 197, 203, 208, 178, 155, 153, 151, 149, 150, 108, 116, 182, 160, 120, 107, 125, 111, 92, 92, 89, 105, 133, 158, 170, 185, 192, 173, 154, 149, 0, 
    323, 150, 165, 203, 263, 223, 158, 159, 154, 149, 150, 126, 124, 158, 153, 140, 129, 134, 127, 111, 114, 117, 126, 136, 140, 151, 191, 245, 222, 161, 150, 0, 
    259, 44, 58, 89, 177, 192, 149, 169, 173, 160, 154, 149, 151, 156, 154, 149, 145, 140, 129, 96, 80, 91, 87, 88, 73, 59, 124, 218, 220, 163, 151, 0, 
    351, 77, 91, 92, 116, 124, 117, 160, 197, 167, 127, 165, 209, 211, 211, 209, 205, 206, 178, 109, 74, 87, 79, 77, 64, 21, 78, 166, 167, 160, 154, 0, 
    386, 153, 176, 183, 181, 154, 114, 117, 163, 115, 6, 58, 166, 177, 189, 207, 221, 235, 212, 141, 112, 116, 106, 110, 120, 89, 101, 139, 149, 179, 176, 0, 
    297, 129, 148, 192, 196, 185, 176, 162, 150, 71, 0, 0, 60, 81, 92, 98, 126, 170, 175, 145, 141, 151, 150, 153, 181, 188, 169, 147, 160, 211, 206, 0, 
    219, 104, 102, 131, 139, 149, 216, 236, 189, 109, 8, 0, 20, 53, 76, 86, 113, 145, 150, 143, 134, 138, 145, 141, 153, 170, 162, 131, 125, 174, 184, 0, 
    185, 170, 178, 92, 39, 88, 188, 211, 186, 150, 97, 69, 76, 100, 81, 63, 98, 122, 112, 96, 69, 58, 69, 75, 75, 89, 104, 94, 84, 114, 142, 0, 
    153, 233, 263, 92, 0, 53, 114, 134, 137, 142, 129, 117, 134, 145, 88, 34, 43, 74, 73, 61, 52, 36, 39, 48, 59, 77, 98, 115, 114, 115, 126, 0, 
    168, 239, 243, 114, 76, 98, 114, 128, 134, 140, 139, 127, 145, 161, 131, 114, 103, 102, 103, 110, 134, 119, 98, 93, 111, 129, 124, 127, 130, 118, 116, 0, 
    221, 188, 141, 113, 125, 133, 128, 128, 127, 128, 132, 122, 123, 116, 102, 121, 130, 120, 75, 79, 124, 120, 90, 77, 83, 101, 99, 102, 110, 111, 110, 0, 
    294, 157, 114, 113, 113, 108, 101, 99, 96, 90, 89, 86, 76, 50, 34, 49, 65, 69, 36, 32, 57, 59, 53, 51, 54, 67, 77, 91, 107, 111, 114, 0, 
    237, 148, 144, 130, 122, 113, 105, 107, 114, 117, 113, 110, 96, 71, 56, 61, 64, 59, 49, 46, 50, 51, 54, 57, 63, 70, 74, 85, 104, 117, 125, 0, 
    125, 75, 120, 103, 69, 65, 75, 88, 104, 119, 125, 129, 118, 92, 80, 87, 92, 75, 59, 56, 56, 61, 64, 66, 71, 76, 72, 73, 98, 124, 139, 0, 
    122, 44, 108, 133, 63, 10, 16, 39, 59, 78, 90, 105, 109, 45, 9, 32, 56, 53, 40, 43, 47, 53, 58, 61, 64, 66, 73, 84, 111, 138, 159, 0, 
    143, 84, 117, 180, 159, 72, 40, 39, 50, 70, 83, 102, 171, 109, 0, 0, 0, 0, 0, 1, 18, 37, 48, 61, 81, 99, 104, 108, 134, 158, 173, 0, 
    117, 84, 111, 157, 186, 142, 101, 82, 75, 83, 93, 102, 215, 291, 124, 3, 6, 17, 23, 32, 49, 77, 101, 109, 110, 126, 142, 141, 151, 171, 182, 0, 
    115, 40, 91, 119, 137, 136, 114, 98, 93, 96, 101, 101, 175, 315, 285, 160, 133, 132, 125, 120, 121, 125, 136, 145, 141, 145, 154, 155, 165, 175, 176, 0, 
    150, 9, 64, 103, 109, 113, 105, 97, 98, 100, 103, 103, 133, 241, 273, 184, 147, 142, 139, 140, 141, 141, 149, 161, 157, 148, 155, 169, 184, 179, 168, 0, 
    184, 6, 44, 100, 103, 106, 101, 97, 99, 101, 103, 103, 116, 195, 239, 163, 121, 130, 137, 141, 142, 147, 153, 158, 155, 149, 157, 173, 187, 186, 171, 0, 
    199, 24, 50, 96, 102, 103, 100, 99, 101, 102, 102, 103, 107, 157, 205, 155, 109, 127, 152, 167, 162, 154, 150, 151, 158, 159, 156, 166, 177, 179, 169, 0, 
    199, 47, 80, 96, 102, 102, 100, 99, 100, 100, 98, 98, 99, 119, 151, 139, 122, 140, 164, 180, 174, 158, 151, 157, 165, 171, 167, 168, 178, 177, 163, 0, 
    205, 74, 108, 110, 109, 108, 106, 102, 100, 99, 98, 99, 103, 115, 136, 146, 149, 156, 163, 178, 176, 157, 158, 165, 167, 169, 172, 174, 179, 182, 166, 0, 
    231, 148, 164, 161, 154, 152, 153, 152, 149, 150, 152, 156, 163, 177, 199, 211, 214, 221, 227, 235, 234, 221, 227, 235, 239, 245, 251, 259, 268, 278, 278, 88, 
    
    -- channel=19
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=20
    0, 200, 195, 196, 196, 196, 196, 196, 196, 195, 195, 197, 197, 197, 197, 198, 198, 196, 195, 194, 194, 196, 196, 196, 196, 197, 197, 196, 195, 195, 198, 433, 
    0, 34, 27, 28, 28, 28, 28, 28, 28, 26, 26, 27, 27, 27, 28, 31, 32, 30, 29, 27, 24, 22, 26, 26, 26, 28, 29, 28, 26, 26, 30, 507, 
    0, 33, 28, 28, 28, 28, 28, 28, 27, 25, 25, 26, 26, 25, 26, 31, 30, 25, 22, 20, 0, 0, 0, 0, 21, 28, 27, 26, 24, 25, 29, 508, 
    0, 32, 27, 28, 28, 28, 28, 29, 28, 27, 27, 28, 28, 25, 27, 33, 34, 33, 27, 46, 0, 0, 0, 0, 22, 31, 28, 28, 26, 27, 30, 509, 
    0, 33, 27, 28, 28, 28, 28, 30, 29, 27, 28, 31, 30, 25, 25, 26, 14, 4, 4, 60, 0, 0, 0, 0, 17, 31, 29, 28, 27, 27, 29, 511, 
    0, 21, 19, 22, 22, 26, 30, 31, 30, 27, 28, 33, 30, 13, 21, 38, 18, 0, 0, 24, 0, 0, 0, 0, 0, 29, 28, 26, 24, 26, 28, 512, 
    0, 10, 22, 24, 19, 23, 29, 31, 31, 29, 29, 40, 28, 0, 18, 74, 68, 27, 18, 33, 1, 0, 0, 0, 0, 25, 28, 26, 24, 25, 27, 513, 
    0, 7, 22, 25, 16, 18, 24, 27, 29, 30, 27, 73, 37, 0, 26, 89, 86, 43, 47, 73, 72, 58, 0, 0, 0, 18, 21, 20, 19, 21, 26, 514, 
    0, 0, 0, 0, 0, 0, 16, 24, 26, 27, 23, 102, 54, 0, 25, 79, 67, 28, 47, 58, 53, 42, 3, 0, 0, 0, 0, 0, 0, 10, 24, 513, 
    0, 0, 0, 0, 0, 0, 8, 17, 21, 25, 21, 84, 53, 0, 16, 50, 47, 15, 26, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 511, 
    0, 75, 57, 3, 0, 0, 7, 0, 0, 2, 5, 24, 7, 0, 0, 9, 15, 11, 18, 38, 36, 23, 27, 37, 43, 43, 0, 0, 0, 0, 16, 509, 
    0, 47, 42, 25, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 55, 94, 77, 81, 76, 94, 135, 37, 0, 0, 0, 6, 507, 
    0, 0, 0, 0, 0, 0, 35, 26, 0, 28, 99, 0, 0, 0, 0, 0, 0, 0, 0, 33, 57, 29, 33, 19, 27, 83, 12, 0, 0, 0, 0, 483, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 79, 248, 144, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 438, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 223, 197, 109, 73, 50, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 415, 
    0, 0, 0, 0, 49, 0, 0, 0, 0, 20, 118, 130, 88, 31, 17, 22, 0, 0, 0, 22, 55, 60, 47, 45, 39, 18, 16, 38, 35, 0, 0, 373, 
    0, 0, 0, 66, 193, 125, 31, 24, 25, 25, 39, 43, 13, 0, 73, 135, 110, 77, 68, 80, 96, 101, 82, 64, 50, 14, 0, 0, 0, 0, 0, 321, 
    0, 0, 0, 30, 109, 52, 11, 1, 0, 0, 0, 0, 0, 0, 0, 21, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 292, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 271, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 274, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 273, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 284, 
    0, 18, 0, 0, 7, 58, 38, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 309, 
    0, 6, 0, 0, 0, 37, 63, 49, 28, 3, 0, 0, 0, 0, 122, 126, 70, 56, 53, 42, 35, 28, 21, 5, 0, 0, 0, 1, 0, 0, 0, 338, 
    0, 21, 0, 0, 0, 0, 11, 26, 21, 2, 0, 0, 0, 0, 29, 148, 136, 118, 103, 90, 61, 24, 0, 0, 0, 0, 10, 13, 0, 0, 0, 359, 
    0, 76, 4, 0, 0, 0, 0, 15, 13, 0, 0, 0, 0, 0, 0, 46, 76, 62, 58, 50, 31, 8, 1, 22, 46, 30, 0, 0, 0, 0, 0, 371, 
    0, 133, 41, 0, 0, 0, 0, 9, 2, 0, 0, 0, 0, 0, 0, 89, 156, 136, 119, 98, 85, 81, 66, 41, 22, 1, 0, 0, 0, 0, 0, 379, 
    0, 165, 70, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 149, 225, 186, 147, 119, 104, 78, 38, 1, 0, 2, 0, 0, 0, 0, 0, 383, 
    0, 160, 79, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 108, 193, 157, 104, 63, 37, 18, 7, 0, 0, 2, 0, 0, 0, 0, 0, 389, 
    0, 138, 80, 35, 20, 12, 9, 7, 8, 9, 10, 6, 7, 0, 0, 77, 135, 89, 29, 0, 0, 10, 11, 0, 0, 0, 0, 0, 0, 0, 0, 394, 
    0, 113, 69, 53, 43, 37, 34, 35, 38, 41, 43, 40, 41, 26, 15, 43, 53, 27, 12, 2, 10, 26, 12, 0, 0, 0, 0, 0, 0, 0, 0, 393, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 143, 
    
    -- channel=21
    239, 190, 191, 191, 191, 191, 191, 191, 191, 192, 192, 192, 192, 192, 192, 191, 190, 192, 192, 192, 191, 191, 191, 191, 192, 191, 191, 191, 192, 192, 191, 10, 
    195, 33, 35, 34, 34, 34, 34, 34, 34, 35, 35, 34, 34, 35, 35, 33, 34, 36, 36, 33, 33, 34, 33, 35, 35, 34, 34, 34, 35, 35, 34, 0, 
    195, 30, 32, 32, 32, 32, 32, 32, 32, 32, 32, 31, 31, 32, 32, 30, 30, 31, 29, 10, 15, 28, 28, 38, 33, 31, 31, 32, 33, 33, 32, 0, 
    195, 32, 34, 33, 33, 33, 33, 33, 32, 33, 33, 32, 32, 33, 33, 33, 33, 27, 15, 0, 0, 23, 28, 34, 34, 33, 33, 33, 34, 34, 33, 0, 
    196, 31, 33, 33, 33, 33, 33, 32, 32, 34, 34, 33, 32, 33, 32, 22, 15, 13, 4, 0, 6, 36, 43, 48, 37, 33, 34, 34, 35, 35, 34, 0, 
    190, 31, 32, 32, 35, 35, 34, 33, 33, 35, 36, 30, 26, 34, 29, 5, 0, 0, 0, 0, 0, 21, 34, 52, 43, 31, 33, 34, 35, 34, 34, 0, 
    184, 30, 28, 27, 32, 34, 34, 35, 35, 35, 35, 16, 15, 39, 25, 1, 0, 3, 2, 0, 0, 1, 14, 41, 43, 31, 32, 33, 34, 34, 34, 0, 
    190, 32, 33, 32, 33, 32, 33, 34, 35, 34, 36, 5, 9, 40, 31, 12, 16, 43, 44, 36, 39, 47, 55, 58, 40, 30, 32, 33, 34, 34, 33, 0, 
    128, 3, 4, 19, 46, 47, 32, 32, 33, 33, 33, 9, 21, 48, 38, 28, 36, 49, 47, 49, 54, 51, 48, 41, 20, 5, 17, 39, 44, 35, 33, 0, 
    76, 0, 0, 0, 25, 41, 26, 32, 35, 32, 32, 22, 33, 51, 39, 31, 38, 46, 38, 22, 8, 0, 0, 0, 0, 0, 0, 28, 48, 36, 33, 0, 
    146, 24, 30, 36, 55, 34, 13, 23, 31, 32, 26, 21, 29, 39, 34, 32, 33, 36, 29, 3, 0, 0, 0, 0, 0, 0, 2, 56, 52, 35, 33, 0, 
    181, 80, 91, 96, 89, 43, 0, 0, 25, 14, 0, 0, 0, 0, 0, 0, 9, 31, 44, 23, 18, 34, 44, 56, 55, 38, 63, 84, 60, 37, 35, 0, 
    112, 0, 1, 10, 24, 26, 5, 15, 31, 0, 0, 0, 0, 0, 0, 0, 0, 26, 40, 31, 37, 50, 43, 38, 44, 43, 56, 49, 29, 32, 35, 0, 
    53, 0, 0, 0, 0, 0, 12, 57, 66, 11, 0, 0, 0, 0, 21, 34, 44, 59, 48, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 30, 0, 
    38, 0, 0, 17, 0, 0, 15, 38, 37, 8, 0, 21, 69, 91, 97, 86, 80, 58, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 24, 0, 
    13, 30, 102, 66, 0, 0, 17, 31, 23, 20, 29, 59, 93, 105, 68, 10, 0, 0, 0, 0, 0, 0, 0, 0, 10, 24, 34, 39, 40, 43, 27, 0, 
    15, 93, 141, 67, 24, 36, 71, 72, 61, 57, 54, 48, 56, 62, 25, 0, 0, 13, 31, 39, 49, 58, 63, 59, 56, 56, 49, 38, 27, 15, 4, 0, 
    83, 148, 122, 47, 33, 73, 84, 76, 63, 51, 33, 11, 12, 5, 0, 0, 29, 46, 26, 21, 36, 32, 17, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    150, 120, 57, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 
    109, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 14, 16, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 12, 20, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 9, 7, 14, 25, 31, 0, 
    5, 0, 0, 23, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 29, 28, 18, 15, 26, 31, 42, 0, 
    0, 0, 0, 14, 16, 5, 0, 0, 0, 0, 0, 0, 56, 93, 46, 11, 8, 5, 6, 15, 25, 39, 48, 41, 28, 25, 22, 13, 20, 41, 59, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 104, 100, 84, 83, 80, 77, 72, 63, 47, 34, 19, 2, 0, 2, 16, 41, 55, 59, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 44, 22, 12, 29, 34, 27, 13, 0, 0, 0, 0, 0, 14, 32, 40, 49, 52, 50, 0, 
    28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 13, 0, 0, 0, 0, 0, 0, 0, 0, 27, 39, 38, 33, 35, 48, 52, 45, 0, 
    35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 26, 0, 0, 0, 0, 0, 17, 36, 48, 46, 34, 21, 21, 32, 43, 44, 41, 0, 
    29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 16, 42, 60, 57, 39, 24, 19, 23, 29, 36, 44, 43, 37, 0, 
    24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 10, 36, 54, 62, 51, 27, 13, 12, 19, 27, 33, 39, 46, 48, 39, 0, 
    33, 0, 0, 2, 4, 4, 4, 5, 6, 8, 10, 13, 15, 24, 38, 44, 49, 55, 46, 36, 23, 9, 8, 16, 23, 27, 28, 32, 39, 41, 35, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=22
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=23
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 7, 9, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 11, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 13, 17, 14, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 13, 6, 5, 3, 3, 3, 2, 2, 1, 1, 3, 6, 0, 3, 15, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 11, 10, 8, 5, 4, 5, 5, 5, 4, 4, 3, 5, 8, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=24
    121, 263, 261, 261, 261, 261, 261, 261, 261, 261, 262, 262, 262, 262, 262, 261, 260, 260, 262, 263, 263, 262, 261, 261, 261, 262, 262, 261, 261, 262, 263, 331, 
    28, 266, 262, 262, 262, 262, 262, 262, 262, 262, 262, 263, 263, 263, 263, 262, 260, 260, 263, 267, 263, 264, 263, 262, 262, 262, 263, 262, 262, 262, 264, 367, 
    27, 265, 262, 262, 262, 262, 262, 263, 262, 262, 261, 262, 262, 261, 262, 261, 259, 259, 262, 271, 245, 246, 245, 250, 260, 262, 262, 262, 261, 262, 263, 368, 
    27, 265, 263, 263, 263, 263, 263, 263, 262, 261, 262, 263, 262, 261, 262, 262, 262, 266, 267, 269, 221, 216, 234, 246, 260, 263, 262, 262, 262, 263, 264, 369, 
    27, 265, 263, 263, 263, 263, 263, 264, 262, 261, 263, 265, 264, 261, 264, 269, 264, 258, 254, 251, 222, 202, 230, 238, 257, 264, 263, 263, 264, 264, 265, 370, 
    24, 259, 258, 258, 259, 262, 264, 264, 264, 262, 263, 269, 265, 257, 266, 275, 257, 237, 235, 238, 222, 185, 191, 213, 249, 264, 263, 263, 263, 265, 265, 371, 
    17, 253, 259, 258, 257, 261, 264, 264, 265, 263, 263, 276, 253, 243, 265, 276, 262, 244, 243, 242, 224, 196, 182, 195, 244, 266, 265, 265, 265, 266, 266, 372, 
    30, 263, 268, 268, 264, 262, 263, 263, 264, 264, 263, 280, 243, 230, 256, 279, 272, 259, 265, 265, 259, 246, 234, 226, 250, 271, 269, 269, 268, 267, 268, 373, 
    19, 211, 213, 213, 216, 245, 260, 261, 261, 263, 264, 277, 254, 228, 252, 277, 271, 264, 277, 283, 285, 287, 276, 254, 238, 242, 233, 233, 253, 268, 269, 374, 
    0, 159, 157, 153, 159, 224, 255, 252, 257, 262, 264, 272, 270, 244, 257, 270, 274, 268, 275, 290, 280, 264, 241, 222, 206, 194, 174, 173, 227, 265, 269, 375, 
    53, 207, 203, 196, 185, 222, 246, 237, 241, 252, 260, 263, 263, 250, 257, 262, 269, 272, 277, 289, 266, 244, 237, 225, 225, 214, 168, 163, 216, 262, 270, 375, 
    80, 253, 249, 251, 238, 231, 248, 216, 201, 238, 260, 214, 186, 187, 193, 201, 209, 213, 243, 281, 287, 275, 274, 262, 263, 261, 218, 211, 230, 258, 268, 375, 
    25, 205, 193, 200, 201, 215, 235, 214, 211, 256, 265, 169, 112, 112, 112, 113, 125, 157, 225, 279, 296, 282, 280, 269, 257, 270, 262, 239, 232, 232, 250, 365, 
    0, 139, 123, 109, 143, 185, 198, 223, 242, 272, 286, 205, 127, 114, 120, 145, 172, 202, 229, 258, 259, 240, 230, 214, 195, 203, 210, 198, 192, 181, 213, 339, 
    0, 99, 100, 119, 160, 141, 128, 173, 213, 252, 280, 256, 198, 196, 223, 238, 219, 201, 195, 202, 193, 173, 157, 151, 142, 138, 153, 173, 181, 172, 207, 322, 
    0, 33, 91, 192, 185, 136, 108, 132, 180, 229, 267, 279, 259, 258, 269, 247, 208, 186, 186, 187, 193, 187, 174, 177, 177, 173, 184, 208, 225, 218, 214, 296, 
    0, 0, 107, 235, 241, 204, 168, 183, 217, 244, 265, 277, 264, 265, 282, 280, 257, 228, 234, 242, 247, 249, 244, 239, 232, 229, 226, 223, 220, 210, 191, 263, 
    0, 45, 141, 236, 275, 247, 231, 232, 244, 246, 255, 262, 250, 257, 266, 270, 250, 238, 246, 231, 217, 235, 240, 229, 208, 193, 183, 173, 173, 179, 183, 239, 
    30, 132, 168, 223, 235, 228, 225, 222, 226, 226, 227, 231, 228, 221, 213, 200, 192, 203, 203, 186, 174, 186, 191, 181, 163, 151, 156, 159, 159, 162, 165, 222, 
    36, 117, 159, 175, 175, 180, 186, 186, 187, 191, 193, 202, 210, 210, 209, 192, 186, 187, 198, 190, 168, 163, 166, 161, 155, 147, 146, 141, 133, 140, 153, 225, 
    0, 60, 85, 93, 101, 107, 110, 111, 116, 124, 132, 144, 159, 172, 177, 168, 166, 165, 172, 163, 145, 139, 136, 131, 131, 127, 126, 125, 127, 137, 149, 220, 
    0, 31, 14, 37, 57, 56, 47, 41, 38, 37, 43, 52, 74, 92, 97, 96, 101, 112, 112, 105, 101, 101, 99, 98, 101, 112, 130, 141, 132, 127, 137, 222, 
    10, 36, 6, 17, 61, 72, 56, 34, 17, 2, 0, 0, 13, 66, 87, 75, 69, 73, 75, 73, 76, 80, 88, 99, 118, 139, 145, 133, 117, 122, 137, 239, 
    0, 24, 0, 0, 36, 72, 64, 43, 22, 0, 0, 0, 0, 66, 152, 148, 122, 113, 113, 110, 107, 111, 126, 141, 138, 117, 104, 111, 121, 128, 148, 258, 
    0, 11, 0, 0, 0, 14, 27, 23, 9, 0, 0, 0, 0, 4, 141, 179, 162, 149, 144, 139, 131, 120, 107, 91, 75, 74, 98, 121, 125, 138, 165, 274, 
    12, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 76, 76, 70, 69, 68, 60, 42, 28, 39, 70, 95, 105, 116, 134, 158, 179, 285, 
    22, 72, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 30, 60, 90, 104, 109, 123, 144, 168, 192, 294, 
    22, 98, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 46, 71, 84, 97, 114, 123, 131, 145, 171, 199, 300, 
    18, 93, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 59, 86, 100, 103, 109, 123, 134, 140, 154, 176, 203, 303, 
    10, 83, 37, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 25, 38, 47, 75, 101, 111, 114, 118, 126, 140, 151, 165, 186, 209, 305, 
    7, 83, 42, 25, 19, 17, 16, 15, 14, 14, 16, 18, 20, 14, 3, 21, 46, 54, 62, 67, 87, 105, 113, 118, 122, 129, 143, 157, 169, 187, 209, 305, 
    0, 34, 8, 2, 0, 0, 0, 0, 0, 0, 2, 4, 3, 1, 0, 0, 0, 4, 10, 14, 23, 36, 41, 41, 43, 48, 53, 60, 66, 73, 85, 133, 
    
    -- channel=25
    251, 316, 315, 315, 315, 315, 315, 315, 315, 315, 316, 316, 316, 316, 316, 314, 313, 313, 315, 316, 319, 320, 317, 314, 314, 315, 315, 315, 315, 316, 316, 284, 
    159, 96, 97, 96, 96, 96, 96, 96, 96, 96, 96, 95, 95, 95, 96, 93, 91, 92, 96, 100, 102, 102, 99, 95, 94, 95, 96, 96, 96, 97, 96, 53, 
    159, 94, 95, 95, 95, 95, 95, 95, 94, 94, 93, 93, 93, 93, 93, 89, 85, 87, 90, 83, 72, 72, 77, 83, 92, 93, 93, 94, 94, 94, 94, 51, 
    158, 94, 95, 96, 96, 96, 96, 96, 95, 95, 96, 96, 95, 95, 95, 94, 95, 98, 95, 84, 66, 77, 87, 94, 96, 96, 96, 97, 97, 97, 96, 53, 
    159, 94, 95, 94, 94, 95, 95, 95, 95, 96, 97, 98, 97, 97, 96, 88, 78, 77, 81, 87, 95, 110, 108, 109, 99, 96, 96, 96, 97, 98, 97, 54, 
    150, 85, 87, 88, 90, 94, 95, 95, 96, 96, 96, 96, 93, 94, 97, 93, 77, 71, 83, 94, 104, 95, 72, 82, 94, 95, 93, 94, 96, 96, 96, 53, 
    150, 91, 98, 96, 95, 95, 94, 95, 97, 96, 95, 88, 76, 82, 94, 99, 114, 138, 154, 159, 155, 137, 105, 95, 100, 100, 98, 100, 100, 99, 97, 53, 
    178, 127, 126, 120, 113, 101, 93, 92, 93, 94, 94, 89, 74, 84, 98, 107, 134, 173, 198, 206, 216, 226, 218, 183, 136, 109, 107, 108, 105, 103, 99, 53, 
    102, 20, 14, 26, 58, 84, 90, 87, 88, 90, 92, 92, 94, 109, 100, 112, 139, 157, 170, 181, 197, 196, 180, 144, 87, 47, 46, 68, 92, 103, 99, 53, 
    121, 36, 27, 22, 42, 75, 82, 79, 86, 91, 95, 97, 112, 127, 107, 105, 122, 139, 137, 132, 119, 93, 70, 53, 40, 24, 18, 40, 82, 102, 100, 53, 
    246, 247, 244, 229, 186, 127, 70, 57, 66, 78, 84, 83, 94, 104, 101, 102, 110, 121, 124, 126, 119, 116, 128, 144, 155, 148, 132, 131, 127, 108, 101, 54, 
    227, 227, 233, 234, 214, 143, 67, 40, 43, 57, 34, 0, 0, 0, 0, 0, 15, 45, 89, 130, 157, 187, 207, 216, 224, 225, 216, 209, 161, 110, 104, 58, 
    124, 49, 41, 39, 54, 65, 85, 105, 120, 119, 74, 12, 0, 0, 0, 0, 16, 60, 107, 129, 148, 164, 157, 143, 140, 151, 168, 154, 99, 77, 88, 50, 
    110, 32, 18, 19, 37, 45, 62, 116, 164, 154, 134, 151, 182, 187, 208, 228, 226, 199, 150, 91, 60, 42, 24, 11, 5, 9, 31, 36, 24, 43, 70, 37, 
    132, 108, 138, 155, 135, 70, 27, 51, 80, 95, 140, 232, 302, 309, 302, 267, 203, 131, 55, 7, 0, 0, 0, 9, 25, 31, 44, 71, 105, 125, 124, 58, 
    109, 111, 191, 246, 189, 97, 78, 82, 80, 105, 152, 215, 254, 257, 226, 149, 83, 62, 68, 94, 126, 150, 166, 181, 195, 199, 204, 211, 216, 197, 152, 60, 
    120, 153, 227, 249, 206, 204, 216, 199, 179, 173, 165, 158, 152, 154, 155, 153, 171, 193, 216, 236, 252, 268, 274, 263, 244, 226, 201, 164, 136, 120, 99, 40, 
    184, 254, 250, 160, 146, 197, 200, 175, 156, 140, 118, 101, 89, 85, 72, 88, 138, 162, 157, 135, 129, 139, 141, 121, 98, 87, 80, 70, 69, 84, 99, 62, 
    245, 296, 200, 97, 94, 110, 105, 95, 88, 83, 76, 75, 85, 90, 68, 64, 76, 101, 108, 93, 94, 94, 88, 86, 90, 97, 104, 114, 123, 128, 136, 89, 
    170, 147, 76, 66, 84, 93, 93, 97, 105, 115, 122, 129, 147, 162, 166, 176, 174, 168, 161, 171, 181, 163, 144, 148, 165, 173, 165, 151, 144, 140, 137, 94, 
    79, 0, 0, 19, 35, 47, 54, 55, 57, 64, 75, 91, 113, 131, 144, 157, 161, 154, 141, 144, 150, 147, 144, 148, 159, 165, 160, 150, 142, 136, 132, 88, 
    112, 66, 67, 90, 98, 85, 68, 54, 40, 28, 21, 32, 55, 72, 76, 79, 88, 97, 101, 107, 116, 128, 138, 147, 164, 180, 182, 171, 149, 127, 121, 84, 
    117, 112, 114, 138, 169, 175, 155, 127, 101, 81, 69, 79, 125, 170, 175, 155, 142, 138, 142, 152, 166, 178, 194, 212, 222, 210, 171, 133, 114, 111, 119, 92, 
    70, 58, 77, 77, 82, 102, 116, 113, 101, 91, 88, 95, 145, 251, 319, 316, 290, 272, 263, 260, 252, 244, 236, 209, 156, 106, 83, 81, 98, 118, 131, 97, 
    79, 56, 61, 54, 20, 0, 15, 39, 56, 67, 74, 82, 82, 108, 161, 205, 215, 216, 208, 192, 161, 122, 82, 51, 30, 28, 55, 91, 116, 125, 131, 88, 
    108, 92, 74, 67, 40, 9, 10, 27, 44, 60, 67, 74, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 77, 102, 108, 118, 128, 129, 77, 
    111, 96, 81, 70, 60, 47, 42, 48, 58, 65, 67, 68, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 65, 93, 98, 91, 93, 112, 126, 127, 77, 
    103, 78, 73, 71, 67, 65, 62, 63, 66, 68, 68, 69, 55, 0, 0, 0, 0, 0, 0, 0, 26, 76, 103, 103, 87, 78, 84, 97, 108, 114, 120, 77, 
    90, 52, 61, 76, 74, 76, 75, 73, 72, 71, 72, 75, 66, 11, 0, 0, 0, 0, 9, 65, 94, 102, 93, 76, 70, 82, 99, 110, 117, 122, 123, 76, 
    85, 41, 62, 85, 87, 90, 90, 87, 86, 87, 89, 95, 97, 74, 23, 0, 18, 69, 89, 82, 69, 62, 59, 64, 74, 84, 96, 107, 118, 126, 127, 75, 
    89, 54, 73, 88, 95, 101, 106, 110, 113, 116, 120, 125, 127, 121, 103, 88, 90, 92, 71, 46, 39, 45, 56, 73, 83, 87, 92, 100, 108, 111, 115, 69, 
    11, 0, 0, 2, 11, 18, 23, 27, 28, 27, 26, 25, 19, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=26
    73, 67, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 67, 66, 68, 69, 71, 71, 69, 66, 66, 68, 68, 68, 68, 68, 69, 107, 
    151, 115, 116, 116, 116, 116, 116, 116, 116, 116, 116, 116, 116, 116, 117, 115, 113, 113, 115, 119, 119, 123, 118, 116, 114, 115, 116, 116, 116, 117, 117, 148, 
    153, 116, 116, 116, 116, 116, 116, 116, 116, 116, 116, 116, 116, 116, 116, 114, 110, 111, 115, 121, 105, 125, 115, 120, 117, 115, 116, 116, 116, 117, 117, 148, 
    152, 116, 117, 116, 116, 116, 116, 117, 116, 116, 116, 116, 116, 116, 116, 114, 114, 117, 119, 124, 93, 117, 113, 115, 117, 116, 116, 116, 116, 117, 117, 149, 
    153, 115, 116, 116, 116, 116, 116, 117, 116, 116, 116, 117, 117, 116, 119, 116, 112, 119, 125, 124, 93, 108, 112, 121, 121, 116, 116, 116, 117, 118, 117, 150, 
    148, 114, 116, 114, 116, 116, 116, 116, 116, 115, 117, 119, 115, 117, 124, 123, 114, 114, 121, 117, 95, 103, 106, 123, 128, 117, 115, 116, 118, 119, 118, 151, 
    145, 119, 120, 116, 116, 117, 116, 116, 117, 117, 117, 122, 101, 116, 126, 121, 115, 115, 121, 118, 110, 104, 97, 107, 130, 121, 117, 119, 119, 120, 119, 151, 
    153, 128, 132, 127, 124, 120, 116, 115, 116, 118, 118, 126, 88, 106, 122, 120, 107, 117, 133, 127, 126, 119, 117, 119, 132, 127, 124, 124, 123, 123, 121, 152, 
    118, 121, 121, 119, 124, 132, 117, 114, 115, 118, 118, 123, 87, 104, 114, 117, 114, 121, 136, 135, 141, 137, 132, 131, 131, 120, 116, 123, 133, 126, 122, 153, 
    111, 91, 91, 83, 91, 127, 113, 110, 115, 116, 118, 121, 100, 112, 117, 119, 119, 128, 138, 139, 137, 137, 131, 121, 113, 100, 88, 97, 131, 128, 122, 153, 
    120, 90, 95, 88, 90, 117, 104, 99, 107, 115, 118, 116, 113, 121, 125, 126, 127, 133, 140, 145, 133, 128, 119, 105, 106, 91, 68, 92, 122, 128, 123, 154, 
    129, 116, 121, 121, 127, 130, 105, 81, 94, 117, 107, 82, 100, 107, 109, 111, 117, 121, 144, 147, 127, 120, 119, 113, 121, 115, 86, 110, 128, 128, 128, 157, 
    124, 117, 117, 121, 125, 129, 114, 93, 98, 122, 111, 54, 65, 72, 71, 74, 86, 100, 129, 133, 127, 129, 133, 123, 128, 127, 111, 125, 122, 124, 131, 159, 
    95, 94, 84, 83, 107, 97, 92, 101, 119, 141, 116, 51, 55, 59, 69, 77, 79, 91, 119, 125, 119, 116, 117, 104, 100, 101, 106, 115, 100, 102, 128, 154, 
    52, 66, 65, 70, 77, 65, 67, 90, 117, 135, 114, 77, 81, 83, 92, 93, 98, 112, 119, 108, 100, 87, 83, 74, 70, 72, 82, 87, 85, 90, 121, 141, 
    7, 24, 69, 99, 72, 46, 37, 71, 91, 110, 106, 101, 106, 117, 137, 122, 106, 102, 99, 94, 93, 79, 74, 72, 74, 76, 85, 94, 99, 101, 117, 131, 
    0, 4, 89, 126, 92, 53, 54, 77, 90, 109, 117, 123, 117, 140, 150, 129, 106, 95, 110, 109, 115, 115, 112, 112, 109, 109, 110, 112, 117, 115, 115, 116, 
    0, 36, 114, 141, 105, 103, 106, 115, 124, 136, 139, 138, 122, 136, 130, 120, 119, 125, 129, 123, 135, 145, 140, 134, 121, 120, 120, 113, 108, 101, 93, 95, 
    26, 94, 148, 144, 130, 141, 145, 148, 149, 150, 148, 144, 133, 144, 130, 125, 122, 132, 140, 121, 122, 133, 131, 122, 107, 102, 96, 86, 83, 82, 85, 95, 
    46, 125, 134, 125, 130, 141, 142, 143, 145, 147, 146, 146, 145, 151, 133, 126, 121, 129, 127, 110, 112, 117, 108, 99, 92, 91, 87, 79, 79, 82, 80, 89, 
    37, 63, 65, 78, 83, 94, 99, 102, 103, 105, 111, 120, 133, 140, 131, 125, 123, 126, 117, 106, 106, 104, 96, 89, 88, 91, 89, 78, 71, 68, 68, 84, 
    10, 0, 0, 29, 35, 33, 33, 34, 32, 34, 39, 53, 79, 96, 100, 99, 99, 101, 93, 88, 84, 80, 78, 75, 77, 79, 77, 64, 52, 54, 58, 83, 
    0, 0, 0, 0, 18, 6, 0, 0, 0, 0, 0, 0, 20, 67, 61, 59, 64, 68, 67, 63, 61, 61, 62, 65, 68, 65, 56, 47, 43, 43, 46, 85, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 62, 79, 53, 50, 53, 51, 49, 45, 44, 47, 47, 43, 42, 46, 39, 28, 35, 50, 96, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 66, 46, 30, 27, 25, 21, 18, 14, 14, 22, 24, 16, 12, 16, 27, 45, 60, 107, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 22, 37, 56, 73, 114, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 24, 41, 67, 83, 118, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 13, 26, 46, 70, 87, 121, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 12, 21, 32, 52, 72, 89, 122, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 15, 27, 40, 56, 76, 93, 122, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 9, 20, 30, 43, 59, 77, 94, 122, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 12, 23, 33, 54, 
    
    -- channel=27
    190, 423, 420, 420, 420, 420, 420, 420, 420, 420, 421, 422, 422, 422, 422, 421, 420, 418, 420, 421, 419, 419, 421, 423, 422, 422, 421, 420, 420, 421, 422, 423, 
    0, 181, 178, 178, 178, 178, 178, 178, 178, 177, 177, 177, 177, 177, 178, 178, 178, 177, 179, 180, 175, 173, 178, 179, 179, 178, 178, 178, 177, 178, 179, 331, 
    0, 179, 176, 176, 176, 176, 176, 176, 175, 174, 173, 173, 173, 173, 174, 177, 176, 173, 171, 169, 147, 129, 146, 151, 170, 175, 174, 174, 174, 174, 176, 330, 
    0, 179, 176, 177, 177, 177, 177, 177, 176, 175, 176, 177, 176, 175, 176, 178, 180, 179, 170, 156, 119, 100, 135, 154, 172, 177, 177, 177, 177, 177, 178, 332, 
    0, 179, 176, 176, 176, 177, 177, 177, 176, 176, 177, 179, 178, 175, 176, 180, 170, 151, 136, 144, 124, 122, 139, 154, 170, 178, 178, 178, 178, 178, 179, 333, 
    0, 168, 167, 169, 169, 175, 179, 179, 178, 176, 177, 180, 176, 167, 171, 173, 146, 116, 109, 134, 119, 93, 83, 102, 151, 180, 178, 177, 177, 178, 178, 333, 
    0, 156, 168, 171, 170, 175, 180, 180, 179, 177, 176, 180, 165, 142, 168, 182, 164, 153, 156, 159, 138, 109, 89, 98, 143, 182, 181, 179, 179, 179, 179, 334, 
    0, 175, 180, 182, 180, 180, 180, 178, 176, 175, 174, 184, 166, 136, 169, 199, 205, 197, 207, 218, 213, 212, 193, 174, 176, 185, 183, 183, 182, 182, 181, 335, 
    0, 56, 57, 67, 90, 138, 176, 174, 171, 171, 173, 198, 185, 159, 182, 202, 205, 200, 211, 221, 227, 235, 215, 167, 134, 116, 107, 116, 147, 179, 182, 337, 
    0, 5, 0, 10, 34, 107, 170, 163, 164, 172, 174, 201, 198, 182, 183, 194, 195, 187, 190, 189, 173, 136, 104, 76, 58, 47, 36, 46, 108, 174, 183, 337, 
    21, 204, 191, 177, 149, 156, 163, 144, 142, 152, 164, 177, 170, 162, 161, 168, 174, 176, 177, 174, 154, 131, 137, 146, 150, 148, 108, 84, 136, 176, 183, 338, 
    47, 243, 239, 230, 189, 174, 159, 123, 93, 118, 139, 81, 18, 19, 30, 42, 57, 74, 112, 180, 215, 231, 245, 246, 242, 244, 211, 167, 172, 170, 175, 338, 
    0, 54, 45, 43, 52, 90, 133, 137, 137, 162, 147, 38, 0, 0, 0, 0, 0, 22, 110, 198, 224, 221, 216, 199, 188, 209, 200, 166, 133, 116, 138, 318, 
    0, 0, 0, 0, 0, 58, 107, 141, 174, 204, 221, 157, 89, 77, 88, 125, 163, 166, 164, 159, 139, 110, 88, 68, 54, 66, 63, 57, 48, 43, 79, 282, 
    0, 0, 23, 60, 88, 62, 27, 52, 95, 151, 232, 251, 247, 254, 278, 275, 210, 125, 75, 47, 29, 11, 3, 6, 9, 12, 28, 62, 81, 84, 106, 284, 
    0, 0, 62, 175, 189, 102, 49, 50, 86, 148, 231, 273, 282, 264, 237, 182, 100, 60, 61, 78, 104, 122, 132, 145, 154, 154, 165, 190, 203, 175, 145, 261, 
    0, 0, 84, 230, 264, 232, 200, 190, 194, 208, 223, 228, 209, 184, 201, 209, 203, 194, 199, 223, 236, 248, 248, 240, 227, 209, 192, 167, 139, 103, 84, 214, 
    16, 50, 117, 195, 226, 230, 217, 196, 170, 153, 146, 149, 136, 128, 156, 164, 163, 159, 160, 130, 104, 117, 127, 110, 83, 55, 39, 30, 35, 57, 79, 207, 
    46, 99, 87, 79, 80, 75, 64, 53, 44, 41, 43, 61, 59, 52, 42, 26, 30, 32, 39, 19, 0, 8, 15, 12, 4, 8, 33, 57, 74, 87, 92, 205, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 28, 37, 55, 65, 69, 63, 63, 80, 77, 55, 45, 47, 57, 62, 69, 78, 74, 65, 71, 92, 210, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 23, 34, 31, 35, 44, 36, 23, 22, 28, 34, 34, 35, 44, 54, 66, 85, 100, 212, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 15, 40, 80, 109, 104, 94, 101, 220, 
    49, 78, 48, 43, 77, 101, 76, 47, 18, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 14, 35, 61, 96, 126, 131, 110, 89, 98, 120, 245, 
    32, 58, 34, 21, 50, 98, 106, 93, 74, 51, 35, 19, 3, 60, 178, 191, 145, 123, 116, 115, 120, 127, 141, 150, 132, 85, 56, 74, 101, 121, 139, 270, 
    36, 65, 29, 0, 0, 4, 31, 46, 49, 44, 40, 25, 0, 7, 126, 210, 208, 197, 186, 176, 160, 136, 94, 46, 17, 26, 70, 110, 122, 134, 146, 279, 
    76, 118, 62, 16, 0, 0, 2, 22, 35, 40, 40, 36, 0, 0, 0, 0, 14, 19, 21, 19, 0, 0, 0, 0, 60, 109, 123, 122, 128, 141, 149, 280, 
    86, 157, 89, 39, 26, 15, 19, 29, 37, 41, 40, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 95, 129, 131, 122, 122, 129, 141, 151, 285, 
    75, 172, 102, 49, 40, 33, 32, 37, 41, 43, 42, 43, 30, 0, 0, 0, 0, 0, 0, 0, 49, 111, 137, 134, 124, 124, 128, 126, 125, 135, 148, 287, 
    58, 161, 105, 69, 57, 53, 53, 51, 50, 48, 47, 48, 41, 0, 0, 0, 0, 0, 26, 88, 130, 148, 145, 130, 125, 134, 143, 140, 135, 143, 154, 290, 
    50, 158, 123, 103, 92, 87, 84, 78, 74, 72, 73, 73, 72, 39, 0, 0, 44, 102, 130, 130, 126, 130, 131, 129, 132, 138, 142, 145, 146, 151, 160, 293, 
    64, 173, 153, 142, 133, 128, 126, 125, 124, 123, 126, 130, 136, 128, 115, 124, 137, 141, 141, 130, 121, 125, 129, 135, 137, 137, 141, 142, 142, 144, 152, 288, 
    19, 55, 59, 59, 57, 58, 60, 59, 57, 55, 55, 56, 58, 54, 39, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 
    
    -- channel=28
    346, 471, 470, 471, 471, 471, 471, 471, 471, 471, 472, 473, 473, 473, 473, 472, 471, 470, 470, 471, 472, 472, 471, 471, 471, 472, 471, 471, 471, 472, 472, 349, 
    336, 397, 396, 396, 396, 396, 396, 396, 396, 396, 397, 397, 397, 397, 398, 397, 395, 394, 395, 395, 395, 397, 397, 398, 397, 397, 396, 396, 396, 398, 398, 304, 
    335, 395, 394, 394, 394, 394, 394, 394, 393, 393, 393, 393, 393, 393, 394, 394, 392, 391, 391, 380, 368, 375, 381, 389, 393, 393, 393, 393, 394, 395, 395, 303, 
    336, 396, 396, 396, 396, 396, 396, 395, 394, 394, 394, 394, 394, 394, 395, 395, 394, 389, 378, 349, 311, 329, 353, 378, 393, 395, 394, 394, 395, 396, 396, 304, 
    336, 395, 395, 396, 396, 396, 396, 395, 394, 395, 396, 396, 394, 394, 395, 391, 382, 372, 352, 321, 284, 321, 358, 388, 397, 396, 396, 397, 398, 399, 399, 306, 
    332, 393, 393, 393, 395, 396, 397, 396, 396, 397, 399, 397, 391, 391, 393, 374, 335, 307, 292, 282, 267, 294, 326, 369, 394, 397, 397, 397, 398, 400, 401, 308, 
    316, 381, 386, 386, 391, 397, 399, 399, 399, 400, 401, 391, 371, 376, 385, 362, 316, 290, 283, 274, 255, 248, 266, 325, 385, 399, 397, 397, 398, 400, 401, 309, 
    312, 386, 395, 393, 395, 398, 400, 400, 401, 401, 401, 383, 344, 359, 383, 365, 337, 338, 342, 332, 320, 315, 320, 351, 392, 401, 399, 400, 401, 403, 403, 310, 
    261, 328, 333, 344, 369, 393, 398, 397, 397, 397, 398, 388, 347, 367, 390, 385, 370, 373, 386, 384, 387, 390, 387, 379, 373, 359, 360, 376, 394, 403, 404, 310, 
    138, 154, 162, 191, 269, 359, 390, 391, 392, 393, 394, 394, 373, 389, 396, 397, 392, 395, 399, 386, 372, 348, 316, 283, 258, 238, 240, 291, 365, 401, 404, 311, 
    182, 223, 226, 237, 286, 359, 371, 368, 376, 382, 383, 384, 382, 390, 391, 392, 393, 396, 395, 370, 323, 282, 256, 244, 237, 217, 209, 267, 358, 398, 403, 311, 
    282, 365, 377, 385, 388, 386, 343, 319, 330, 344, 323, 287, 280, 289, 301, 315, 331, 351, 376, 377, 348, 340, 347, 349, 349, 324, 299, 338, 387, 396, 402, 311, 
    229, 279, 293, 311, 331, 342, 323, 297, 308, 322, 245, 119, 82, 93, 109, 134, 180, 250, 335, 387, 391, 396, 395, 379, 378, 372, 359, 372, 365, 366, 386, 306, 
    110, 123, 121, 142, 193, 245, 294, 329, 366, 362, 255, 114, 79, 90, 116, 156, 219, 294, 367, 380, 361, 343, 323, 295, 286, 296, 299, 289, 263, 284, 335, 278, 
    45, 75, 90, 127, 173, 195, 222, 281, 334, 337, 288, 225, 225, 249, 299, 342, 359, 352, 328, 282, 238, 200, 177, 159, 154, 165, 181, 192, 199, 236, 297, 250, 
    0, 58, 159, 230, 218, 161, 168, 228, 270, 306, 328, 341, 364, 385, 389, 337, 271, 233, 211, 197, 183, 166, 166, 175, 189, 204, 230, 261, 281, 292, 313, 238, 
    0, 49, 234, 339, 291, 239, 264, 302, 326, 364, 387, 396, 394, 402, 388, 326, 273, 262, 275, 290, 304, 307, 308, 308, 307, 306, 313, 317, 310, 286, 266, 189, 
    0, 139, 321, 385, 351, 364, 384, 393, 391, 395, 389, 375, 353, 356, 355, 340, 333, 327, 323, 312, 315, 322, 316, 293, 267, 252, 234, 212, 198, 195, 198, 155, 
    99, 246, 322, 300, 289, 307, 314, 309, 301, 298, 296, 294, 278, 269, 235, 214, 216, 224, 212, 169, 164, 181, 175, 150, 125, 121, 128, 139, 159, 182, 198, 154, 
    132, 232, 210, 188, 185, 187, 188, 191, 194, 196, 201, 208, 210, 208, 182, 173, 174, 185, 177, 153, 148, 145, 132, 124, 120, 130, 143, 151, 163, 178, 191, 152, 
    19, 33, 29, 46, 56, 65, 71, 78, 89, 104, 121, 138, 154, 168, 171, 174, 171, 168, 154, 137, 125, 111, 102, 102, 103, 109, 119, 124, 140, 167, 192, 156, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 22, 33, 42, 52, 58, 52, 41, 36, 38, 45, 56, 69, 91, 120, 140, 156, 177, 197, 159, 
    0, 0, 0, 0, 27, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 40, 72, 110, 146, 169, 171, 168, 180, 210, 179, 
    0, 0, 0, 0, 48, 60, 29, 0, 0, 0, 0, 0, 0, 80, 102, 66, 42, 36, 36, 47, 65, 91, 124, 154, 177, 181, 166, 153, 162, 198, 242, 209, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 131, 242, 241, 210, 196, 190, 186, 184, 184, 179, 160, 130, 110, 122, 155, 192, 230, 270, 230, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 158, 194, 191, 190, 181, 162, 134, 103, 73, 66, 84, 120, 160, 188, 213, 250, 285, 234, 
    36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 77, 97, 81, 69, 53, 34, 19, 21, 48, 97, 146, 170, 180, 194, 226, 268, 295, 236, 
    62, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 64, 87, 50, 21, 5, 12, 39, 83, 127, 159, 172, 170, 177, 198, 232, 268, 297, 240, 
    66, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 37, 0, 0, 5, 65, 122, 157, 169, 170, 170, 178, 194, 214, 240, 271, 299, 241, 
    57, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 11, 44, 90, 138, 164, 168, 163, 162, 172, 191, 210, 230, 256, 286, 309, 243, 
    59, 34, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 35, 70, 95, 126, 144, 156, 164, 160, 154, 164, 180, 196, 213, 233, 259, 286, 309, 242, 
    19, 12, 2, 0, 0, 0, 0, 0, 0, 0, 1, 4, 9, 19, 34, 54, 66, 74, 78, 77, 79, 73, 72, 83, 94, 103, 112, 123, 135, 150, 164, 138, 
    
    -- channel=29
    436, 401, 402, 402, 402, 402, 402, 402, 402, 403, 404, 404, 404, 404, 404, 404, 402, 402, 401, 401, 403, 404, 403, 401, 402, 402, 402, 402, 403, 404, 403, 114, 
    511, 372, 375, 374, 374, 374, 374, 374, 374, 375, 376, 376, 376, 376, 376, 375, 375, 374, 373, 370, 373, 377, 375, 375, 375, 375, 374, 374, 376, 377, 375, 42, 
    512, 372, 373, 373, 373, 373, 373, 373, 372, 373, 373, 372, 372, 374, 374, 371, 369, 369, 366, 343, 345, 365, 367, 380, 375, 372, 372, 373, 374, 375, 374, 40, 
    512, 373, 375, 375, 375, 375, 375, 374, 373, 373, 374, 373, 372, 374, 375, 373, 370, 361, 346, 296, 300, 340, 356, 373, 376, 373, 373, 374, 375, 376, 375, 41, 
    513, 372, 375, 375, 375, 375, 375, 373, 373, 375, 376, 374, 372, 374, 373, 358, 346, 337, 318, 272, 280, 336, 364, 388, 382, 375, 375, 376, 377, 378, 377, 42, 
    506, 372, 374, 374, 377, 377, 375, 374, 375, 378, 380, 371, 364, 374, 369, 328, 291, 279, 269, 246, 251, 303, 345, 389, 390, 375, 374, 376, 378, 379, 379, 43, 
    491, 368, 367, 368, 374, 378, 377, 377, 379, 380, 382, 353, 341, 374, 360, 309, 275, 270, 263, 246, 240, 252, 294, 362, 388, 375, 373, 375, 377, 379, 380, 43, 
    489, 370, 374, 372, 375, 377, 377, 379, 381, 381, 383, 333, 319, 366, 361, 318, 297, 319, 318, 300, 296, 302, 326, 369, 382, 373, 374, 376, 378, 380, 380, 43, 
    397, 315, 321, 340, 380, 392, 377, 377, 378, 378, 379, 333, 323, 370, 370, 345, 340, 358, 358, 354, 357, 353, 350, 354, 346, 331, 345, 374, 389, 382, 380, 43, 
    275, 166, 180, 223, 327, 380, 368, 373, 376, 374, 373, 350, 346, 378, 376, 366, 366, 378, 374, 351, 329, 305, 281, 258, 240, 226, 251, 334, 387, 382, 379, 43, 
    315, 217, 229, 256, 334, 361, 343, 353, 364, 366, 358, 349, 354, 372, 372, 372, 372, 376, 369, 325, 281, 255, 234, 227, 219, 190, 227, 333, 382, 380, 378, 42, 
    408, 335, 354, 370, 390, 366, 302, 296, 337, 331, 261, 238, 269, 284, 295, 309, 326, 357, 380, 340, 305, 308, 310, 320, 315, 277, 303, 369, 388, 380, 381, 43, 
    358, 272, 294, 315, 338, 339, 294, 290, 325, 284, 139, 72, 102, 116, 135, 173, 232, 318, 367, 360, 352, 364, 355, 347, 352, 334, 342, 356, 348, 365, 379, 46, 
    230, 141, 148, 197, 249, 258, 289, 338, 366, 298, 129, 58, 91, 121, 165, 210, 265, 335, 369, 348, 322, 310, 288, 270, 277, 284, 285, 272, 261, 312, 353, 38, 
    140, 107, 138, 187, 188, 198, 264, 319, 338, 295, 205, 178, 220, 262, 300, 318, 339, 344, 311, 258, 214, 186, 172, 163, 169, 185, 197, 199, 213, 277, 318, 22, 
    68, 134, 254, 247, 168, 160, 222, 278, 297, 302, 295, 304, 341, 373, 352, 284, 245, 227, 209, 194, 174, 158, 166, 177, 190, 213, 242, 260, 267, 291, 300, 24, 
    35, 202, 358, 308, 227, 223, 286, 320, 336, 357, 366, 358, 367, 386, 336, 267, 231, 243, 262, 269, 277, 279, 282, 280, 279, 286, 292, 291, 282, 266, 257, 7, 
    110, 300, 394, 345, 298, 335, 364, 374, 376, 380, 369, 337, 330, 328, 298, 281, 290, 306, 286, 280, 305, 305, 284, 258, 243, 240, 227, 211, 202, 196, 199, 0, 
    244, 331, 343, 286, 276, 297, 305, 305, 299, 295, 289, 273, 267, 248, 214, 206, 223, 229, 196, 169, 187, 190, 171, 143, 134, 140, 140, 148, 169, 190, 205, 8, 
    250, 268, 226, 202, 207, 209, 207, 213, 218, 220, 222, 221, 221, 206, 183, 183, 193, 194, 166, 152, 162, 153, 134, 125, 129, 143, 149, 160, 183, 200, 209, 6, 
    110, 69, 67, 84, 92, 101, 108, 117, 128, 141, 155, 169, 182, 185, 182, 187, 186, 177, 151, 140, 138, 125, 115, 117, 121, 133, 142, 150, 171, 191, 208, 8, 
    13, 0, 0, 11, 0, 0, 0, 0, 0, 6, 16, 35, 57, 68, 75, 84, 90, 85, 72, 67, 65, 66, 75, 89, 110, 136, 153, 156, 172, 198, 216, 9, 
    4, 0, 0, 45, 50, 8, 0, 0, 0, 0, 0, 0, 19, 28, 0, 0, 13, 18, 20, 29, 41, 60, 87, 124, 159, 176, 174, 171, 185, 202, 232, 17, 
    0, 0, 0, 37, 71, 48, 11, 0, 0, 0, 0, 0, 78, 163, 113, 63, 60, 61, 67, 82, 104, 134, 161, 177, 185, 189, 183, 170, 180, 218, 264, 27, 
    0, 0, 0, 0, 19, 10, 0, 0, 0, 0, 0, 0, 75, 242, 268, 226, 207, 202, 201, 198, 197, 194, 187, 172, 151, 142, 148, 167, 207, 250, 285, 33, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 188, 254, 232, 228, 229, 215, 186, 151, 126, 112, 108, 114, 137, 171, 197, 229, 263, 291, 29, 
    49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 112, 218, 195, 166, 143, 111, 83, 67, 67, 91, 131, 158, 171, 182, 203, 241, 275, 294, 26, 
    84, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 64, 190, 175, 118, 83, 70, 75, 91, 116, 146, 169, 172, 165, 174, 205, 244, 275, 295, 26, 
    91, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 114, 102, 55, 47, 70, 113, 149, 164, 163, 162, 164, 173, 189, 216, 249, 277, 295, 24, 
    83, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 61, 54, 82, 125, 164, 174, 158, 146, 149, 166, 186, 204, 228, 259, 288, 300, 24, 
    88, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 63, 95, 117, 142, 151, 160, 159, 143, 140, 153, 172, 191, 207, 230, 259, 285, 298, 23, 
    23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 33, 57, 70, 75, 71, 72, 71, 62, 65, 77, 89, 98, 110, 122, 137, 153, 162, 4, 
    
    -- channel=30
    82, 42, 43, 43, 43, 43, 43, 43, 43, 44, 44, 43, 43, 43, 43, 43, 43, 44, 43, 42, 41, 42, 43, 44, 44, 43, 43, 43, 44, 44, 43, 0, 
    253, 219, 219, 219, 219, 219, 219, 219, 219, 220, 221, 221, 221, 221, 220, 220, 221, 222, 220, 216, 218, 218, 220, 220, 221, 220, 219, 219, 220, 221, 220, 17, 
    255, 220, 221, 221, 221, 221, 221, 220, 221, 221, 222, 222, 222, 222, 222, 222, 223, 223, 222, 214, 230, 225, 228, 224, 222, 222, 221, 221, 222, 222, 221, 18, 
    255, 221, 221, 221, 221, 221, 221, 220, 220, 220, 220, 220, 220, 221, 221, 221, 218, 215, 213, 195, 211, 215, 214, 222, 220, 220, 220, 220, 220, 221, 221, 18, 
    255, 221, 221, 221, 221, 221, 221, 220, 220, 221, 220, 219, 219, 221, 220, 219, 222, 217, 204, 173, 173, 199, 207, 219, 221, 221, 221, 221, 221, 221, 221, 18, 
    258, 223, 223, 223, 223, 222, 222, 220, 220, 221, 222, 218, 220, 223, 217, 206, 203, 199, 182, 155, 158, 194, 222, 230, 224, 222, 222, 222, 223, 223, 223, 18, 
    255, 219, 217, 220, 223, 224, 223, 221, 221, 222, 224, 214, 224, 225, 214, 189, 164, 151, 140, 127, 126, 149, 189, 226, 226, 221, 221, 222, 223, 223, 223, 19, 
    238, 210, 210, 213, 219, 224, 224, 224, 224, 224, 225, 203, 211, 224, 212, 179, 158, 146, 131, 119, 107, 110, 137, 191, 219, 219, 220, 221, 223, 223, 223, 19, 
    258, 235, 239, 241, 239, 225, 224, 225, 226, 225, 226, 197, 191, 217, 216, 190, 176, 178, 168, 157, 150, 151, 167, 197, 223, 231, 237, 237, 226, 223, 224, 18, 
    189, 171, 181, 204, 236, 227, 224, 226, 225, 225, 225, 203, 191, 212, 219, 210, 199, 203, 201, 193, 200, 201, 200, 197, 192, 196, 215, 238, 231, 223, 224, 18, 
    88, 61, 68, 99, 171, 215, 220, 228, 230, 227, 224, 216, 211, 219, 221, 219, 215, 215, 210, 193, 182, 164, 141, 128, 109, 105, 141, 191, 224, 223, 224, 18, 
    144, 105, 111, 122, 164, 198, 198, 219, 232, 217, 210, 231, 237, 239, 240, 241, 240, 241, 221, 184, 150, 133, 119, 116, 104, 83, 110, 166, 212, 223, 223, 17, 
    219, 191, 205, 212, 220, 205, 176, 171, 190, 176, 133, 143, 161, 167, 179, 192, 202, 215, 215, 196, 176, 175, 171, 176, 176, 148, 152, 190, 216, 228, 228, 21, 
    169, 144, 159, 185, 189, 194, 186, 169, 180, 153, 60, 18, 32, 42, 48, 61, 99, 158, 206, 215, 216, 221, 215, 212, 220, 214, 206, 202, 205, 225, 227, 26, 
    87, 64, 63, 84, 119, 159, 191, 210, 215, 169, 73, 9, 8, 22, 46, 85, 136, 186, 212, 210, 198, 189, 176, 162, 163, 172, 166, 145, 139, 173, 194, 17, 
    50, 64, 60, 54, 82, 98, 145, 187, 198, 171, 126, 94, 96, 119, 139, 158, 170, 171, 155, 133, 103, 83, 75, 71, 72, 83, 93, 95, 100, 136, 172, 13, 
    18, 74, 116, 103, 62, 57, 99, 137, 159, 173, 178, 177, 192, 200, 177, 131, 106, 106, 93, 87, 76, 62, 63, 72, 82, 95, 118, 141, 147, 155, 163, 10, 
    0, 73, 172, 166, 124, 119, 143, 170, 187, 205, 213, 208, 214, 217, 200, 163, 140, 133, 139, 152, 158, 148, 144, 144, 150, 155, 157, 157, 149, 134, 127, 0, 
    23, 108, 178, 179, 176, 180, 187, 194, 196, 200, 201, 188, 182, 180, 172, 165, 159, 151, 136, 132, 144, 147, 135, 118, 110, 109, 101, 95, 96, 100, 105, 0, 
    114, 148, 150, 146, 146, 144, 142, 142, 140, 137, 136, 129, 120, 103, 85, 81, 90, 96, 72, 57, 68, 75, 65, 51, 43, 49, 57, 69, 82, 93, 102, 0, 
    119, 117, 109, 100, 98, 94, 94, 98, 102, 103, 105, 104, 98, 83, 71, 70, 74, 74, 63, 54, 54, 49, 42, 38, 40, 48, 52, 60, 74, 90, 104, 0, 
    15, 11, 27, 19, 14, 19, 27, 35, 45, 58, 67, 72, 70, 66, 66, 71, 69, 57, 48, 40, 35, 31, 27, 27, 31, 34, 35, 46, 72, 97, 113, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 3, 2, 0, 0, 0, 0, 0, 2, 12, 28, 52, 71, 87, 104, 122, 0, 
    3, 0, 0, 31, 23, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 56, 85, 93, 87, 96, 115, 134, 0, 
    0, 0, 0, 18, 48, 35, 11, 0, 0, 0, 0, 0, 44, 99, 40, 0, 0, 0, 0, 6, 23, 49, 79, 96, 100, 98, 95, 95, 110, 130, 152, 1, 
    0, 0, 0, 0, 5, 14, 4, 0, 0, 0, 0, 0, 29, 151, 170, 140, 130, 123, 121, 119, 118, 120, 118, 103, 82, 81, 97, 110, 123, 143, 164, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 85, 150, 158, 160, 156, 151, 137, 115, 89, 74, 76, 86, 98, 111, 122, 138, 153, 166, 4, 
    24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 103, 129, 135, 128, 109, 83, 65, 60, 70, 92, 106, 106, 111, 126, 148, 163, 169, 3, 
    45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 79, 106, 97, 80, 65, 61, 68, 81, 96, 105, 110, 108, 111, 127, 145, 162, 170, 4, 
    50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 52, 43, 41, 58, 83, 100, 108, 107, 106, 111, 118, 123, 133, 149, 163, 171, 4, 
    49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 30, 47, 63, 83, 106, 118, 116, 108, 106, 112, 122, 132, 141, 157, 172, 175, 4, 
    75, 37, 29, 24, 19, 15, 12, 11, 12, 14, 17, 21, 26, 38, 59, 84, 107, 124, 134, 142, 147, 141, 138, 143, 151, 162, 174, 188, 203, 221, 231, 91, 
    
    -- channel=31
    89, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    203, 136, 137, 137, 137, 137, 137, 137, 137, 138, 138, 138, 138, 138, 138, 138, 138, 139, 137, 135, 136, 137, 138, 137, 137, 137, 137, 137, 138, 138, 137, 47, 
    204, 138, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 140, 140, 140, 140, 141, 140, 135, 136, 140, 140, 142, 140, 139, 139, 139, 139, 140, 139, 49, 
    204, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 139, 139, 139, 138, 137, 134, 120, 126, 140, 140, 146, 141, 138, 138, 138, 138, 139, 139, 48, 
    204, 139, 139, 139, 139, 139, 139, 139, 138, 139, 139, 138, 138, 138, 139, 139, 136, 130, 123, 107, 104, 131, 129, 139, 141, 138, 138, 138, 139, 139, 139, 48, 
    204, 139, 140, 140, 140, 140, 138, 138, 139, 140, 140, 139, 136, 138, 137, 127, 122, 122, 114, 104, 92, 117, 134, 144, 143, 139, 139, 139, 140, 139, 140, 49, 
    201, 141, 140, 140, 142, 140, 139, 139, 139, 141, 142, 137, 133, 140, 135, 114, 98, 93, 89, 79, 76, 93, 125, 150, 146, 136, 137, 138, 139, 139, 140, 50, 
    193, 134, 133, 131, 135, 138, 139, 141, 142, 142, 143, 127, 126, 142, 132, 112, 95, 82, 74, 68, 64, 65, 82, 120, 138, 133, 134, 134, 135, 137, 139, 49, 
    183, 130, 135, 133, 134, 137, 138, 142, 144, 143, 143, 125, 114, 137, 137, 116, 104, 107, 99, 91, 89, 85, 85, 98, 124, 133, 135, 135, 136, 135, 137, 48, 
    144, 114, 123, 136, 155, 151, 138, 142, 144, 142, 139, 131, 115, 130, 137, 131, 120, 121, 123, 116, 113, 106, 105, 107, 114, 122, 133, 149, 147, 135, 137, 47, 
    91, 42, 51, 69, 117, 142, 135, 144, 146, 141, 136, 133, 125, 130, 133, 134, 131, 129, 127, 111, 99, 97, 91, 86, 81, 76, 90, 129, 146, 134, 135, 47, 
    122, 49, 56, 60, 82, 116, 124, 135, 147, 142, 129, 128, 136, 138, 140, 140, 139, 136, 130, 108, 87, 80, 68, 66, 61, 47, 65, 99, 126, 132, 134, 45, 
    165, 110, 121, 129, 128, 126, 108, 110, 134, 119, 78, 84, 111, 115, 121, 128, 135, 148, 147, 122, 99, 94, 94, 96, 101, 89, 86, 106, 122, 136, 138, 45, 
    134, 102, 112, 128, 146, 140, 123, 108, 105, 88, 33, 7, 30, 34, 45, 63, 88, 112, 129, 128, 124, 124, 124, 122, 132, 131, 115, 117, 125, 139, 144, 51, 
    79, 53, 52, 77, 85, 92, 126, 136, 123, 101, 49, 0, 4, 21, 38, 43, 59, 91, 121, 129, 124, 120, 119, 111, 112, 119, 117, 106, 99, 117, 129, 46, 
    50, 50, 56, 38, 30, 60, 103, 129, 131, 119, 88, 54, 49, 59, 66, 76, 98, 114, 115, 104, 88, 72, 70, 65, 59, 63, 72, 71, 64, 77, 95, 31, 
    27, 73, 106, 57, 31, 45, 75, 101, 111, 114, 107, 100, 100, 109, 97, 80, 76, 77, 72, 63, 52, 40, 38, 41, 44, 51, 63, 71, 71, 72, 88, 36, 
    28, 79, 114, 107, 76, 70, 84, 102, 110, 120, 124, 118, 123, 131, 119, 92, 68, 70, 72, 70, 80, 78, 72, 71, 76, 79, 79, 87, 92, 90, 88, 32, 
    58, 69, 107, 121, 116, 115, 116, 125, 128, 132, 131, 121, 111, 109, 104, 104, 106, 96, 83, 85, 102, 99, 87, 79, 77, 82, 77, 71, 72, 70, 66, 21, 
    80, 77, 97, 99, 97, 101, 103, 103, 101, 100, 102, 99, 87, 80, 65, 66, 71, 76, 62, 47, 51, 56, 50, 45, 39, 40, 41, 43, 53, 63, 70, 20, 
    82, 86, 85, 79, 75, 73, 72, 74, 75, 75, 74, 74, 71, 66, 56, 52, 47, 52, 51, 40, 38, 39, 37, 37, 37, 36, 38, 46, 60, 69, 70, 20, 
    29, 25, 40, 41, 38, 41, 45, 48, 52, 58, 62, 66, 70, 68, 67, 66, 63, 54, 48, 47, 43, 38, 36, 35, 36, 39, 40, 43, 53, 65, 72, 24, 
    4, 0, 3, 10, 0, 0, 0, 0, 3, 10, 17, 23, 29, 26, 21, 24, 32, 29, 25, 25, 21, 19, 21, 24, 30, 41, 46, 46, 59, 73, 81, 23, 
    22, 0, 0, 29, 29, 3, 0, 0, 0, 0, 0, 0, 21, 10, 0, 0, 0, 0, 0, 0, 2, 11, 22, 34, 44, 53, 65, 74, 78, 80, 86, 24, 
    16, 4, 0, 18, 52, 47, 30, 11, 0, 0, 0, 0, 46, 88, 41, 2, 0, 5, 12, 19, 30, 46, 57, 62, 74, 91, 97, 82, 75, 85, 91, 27, 
    4, 0, 0, 0, 26, 46, 39, 23, 6, 0, 0, 0, 20, 122, 172, 150, 134, 127, 123, 120, 115, 111, 113, 113, 102, 84, 74, 72, 78, 86, 94, 30, 
    20, 0, 0, 0, 6, 21, 23, 12, 2, 0, 0, 0, 5, 89, 199, 236, 237, 226, 207, 180, 154, 130, 111, 96, 76, 64, 68, 76, 81, 87, 93, 29, 
    42, 0, 0, 0, 0, 5, 8, 4, 0, 0, 0, 0, 7, 78, 192, 246, 242, 218, 184, 148, 113, 86, 70, 67, 68, 68, 69, 76, 84, 93, 95, 28, 
    52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 62, 162, 209, 191, 157, 122, 94, 73, 61, 58, 64, 71, 69, 66, 72, 82, 93, 97, 29, 
    51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 90, 127, 111, 76, 56, 62, 74, 71, 64, 63, 67, 71, 69, 74, 82, 90, 95, 28, 
    48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 31, 53, 53, 51, 60, 75, 84, 77, 66, 62, 63, 70, 75, 79, 86, 95, 97, 28, 
    55, 12, 11, 10, 7, 6, 5, 5, 6, 8, 9, 7, 9, 18, 33, 50, 68, 83, 89, 90, 89, 81, 74, 74, 79, 84, 89, 95, 103, 113, 119, 51, 
    
    -- channel=32
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=33
    8, 84, 73, 60, 67, 81, 83, 82, 82, 82, 79, 74, 70, 70, 68, 69, 64, 61, 66, 69, 70, 65, 63, 63, 64, 64, 62, 65, 65, 62, 63, 69, 
    27, 86, 76, 63, 70, 83, 83, 78, 77, 77, 73, 66, 62, 62, 62, 64, 59, 57, 59, 60, 57, 52, 51, 53, 59, 58, 58, 62, 60, 54, 57, 65, 
    23, 78, 67, 56, 61, 72, 75, 70, 66, 67, 64, 56, 54, 55, 56, 60, 57, 54, 56, 50, 39, 34, 41, 51, 56, 55, 54, 59, 57, 51, 53, 63, 
    20, 72, 60, 47, 53, 62, 64, 59, 55, 58, 55, 48, 46, 48, 48, 54, 54, 51, 53, 54, 43, 24, 33, 50, 56, 52, 50, 53, 53, 48, 51, 59, 
    16, 66, 54, 40, 45, 52, 55, 51, 46, 47, 46, 42, 40, 44, 37, 37, 41, 43, 48, 45, 27, 23, 40, 50, 54, 48, 43, 46, 44, 43, 50, 56, 
    9, 55, 44, 31, 36, 42, 45, 42, 38, 38, 36, 37, 39, 39, 29, 25, 26, 27, 38, 50, 24, 7, 24, 34, 44, 44, 36, 35, 33, 36, 46, 47, 
    5, 46, 37, 26, 30, 34, 33, 32, 30, 29, 27, 30, 32, 35, 34, 27, 16, 6, 2, 10, 2, 0, 0, 0, 0, 25, 31, 29, 24, 22, 28, 28, 
    0, 30, 26, 10, 9, 12, 11, 12, 13, 14, 12, 16, 20, 22, 20, 23, 24, 21, 22, 15, 12, 20, 13, 0, 0, 0, 3, 11, 6, 0, 0, 5, 
    0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 20, 27, 27, 29, 28, 28, 26, 24, 18, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 21, 23, 25, 26, 27, 22, 23, 26, 8, 0, 3, 6, 10, 0, 0, 0, 0, 
    0, 0, 7, 4, 9, 13, 4, 0, 0, 4, 5, 4, 12, 22, 34, 41, 36, 28, 27, 26, 24, 24, 31, 32, 29, 0, 0, 6, 3, 0, 0, 0, 
    0, 19, 20, 8, 13, 22, 18, 15, 17, 33, 38, 27, 30, 43, 51, 44, 35, 29, 25, 28, 31, 25, 24, 35, 43, 26, 0, 0, 3, 0, 0, 5, 
    0, 24, 29, 16, 7, 12, 13, 9, 18, 35, 44, 46, 46, 53, 57, 50, 43, 37, 34, 39, 40, 29, 25, 22, 22, 27, 1, 0, 0, 0, 0, 1, 
    0, 31, 31, 18, 16, 16, 15, 28, 40, 44, 50, 59, 64, 66, 67, 67, 66, 65, 61, 56, 45, 30, 25, 17, 10, 12, 2, 0, 0, 0, 0, 0, 
    2, 45, 43, 35, 38, 48, 53, 55, 62, 68, 69, 71, 74, 78, 77, 71, 69, 71, 65, 49, 27, 14, 10, 6, 6, 8, 10, 0, 0, 0, 0, 0, 
    6, 53, 54, 52, 47, 54, 66, 71, 76, 76, 77, 78, 78, 77, 74, 67, 57, 53, 50, 36, 14, 2, 0, 0, 6, 11, 20, 23, 18, 9, 7, 0, 
    7, 59, 54, 45, 40, 45, 61, 74, 77, 79, 78, 75, 71, 67, 60, 54, 47, 43, 44, 40, 23, 9, 7, 7, 12, 17, 23, 19, 6, 8, 21, 15, 
    6, 46, 43, 42, 43, 45, 51, 66, 71, 70, 68, 67, 66, 64, 58, 52, 45, 36, 37, 41, 31, 25, 25, 23, 23, 24, 21, 11, 1, 0, 0, 9, 
    0, 46, 48, 50, 54, 60, 63, 59, 61, 64, 65, 63, 62, 60, 56, 50, 46, 40, 36, 37, 34, 30, 30, 30, 28, 19, 10, 2, 0, 0, 0, 5, 
    16, 59, 47, 49, 60, 67, 68, 63, 61, 63, 62, 59, 56, 51, 45, 36, 28, 24, 30, 35, 35, 31, 28, 24, 15, 6, 3, 0, 0, 0, 0, 0, 
    10, 62, 65, 68, 67, 64, 62, 60, 52, 51, 56, 57, 54, 45, 28, 16, 9, 3, 15, 30, 29, 23, 16, 14, 10, 1, 0, 0, 0, 0, 0, 0, 
    1, 60, 67, 68, 64, 59, 51, 43, 36, 33, 36, 45, 50, 50, 38, 20, 13, 4, 4, 14, 16, 12, 11, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 42, 57, 59, 57, 52, 39, 27, 23, 25, 25, 32, 45, 51, 41, 24, 15, 7, 8, 11, 9, 6, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 37, 48, 51, 54, 57, 46, 31, 28, 33, 31, 27, 26, 23, 17, 15, 14, 11, 10, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 35, 43, 45, 45, 48, 41, 29, 24, 20, 12, 13, 12, 10, 9, 8, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 16, 20, 22, 19, 16, 11, 11, 13, 10, 4, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=34
    264, 0, 0, 45, 76, 33, 18, 24, 27, 24, 16, 34, 51, 43, 45, 24, 33, 63, 54, 47, 35, 41, 55, 52, 36, 38, 60, 45, 32, 53, 58, 0, 
    350, 38, 20, 99, 150, 107, 85, 98, 116, 106, 93, 116, 144, 136, 141, 117, 118, 151, 149, 144, 126, 146, 168, 158, 130, 130, 158, 136, 117, 152, 158, 0, 
    361, 54, 36, 111, 166, 129, 99, 105, 135, 124, 103, 126, 153, 143, 152, 132, 120, 153, 150, 125, 125, 190, 209, 169, 136, 133, 165, 142, 116, 156, 166, 0, 
    367, 60, 45, 124, 176, 145, 117, 116, 154, 141, 113, 131, 159, 144, 157, 154, 125, 154, 144, 82, 83, 204, 231, 176, 140, 133, 170, 150, 124, 158, 165, 0, 
    378, 70, 47, 132, 188, 158, 134, 123, 167, 157, 123, 135, 163, 137, 146, 178, 148, 174, 142, 46, 91, 228, 224, 175, 146, 133, 176, 159, 138, 168, 160, 0, 
    388, 85, 50, 139, 204, 171, 153, 137, 175, 164, 134, 145, 165, 129, 118, 175, 170, 191, 162, 20, 69, 241, 237, 207, 181, 140, 177, 174, 153, 180, 163, 0, 
    388, 90, 51, 138, 211, 169, 164, 155, 182, 166, 147, 158, 168, 134, 102, 126, 136, 162, 177, 103, 99, 207, 232, 268, 299, 221, 190, 179, 160, 199, 187, 0, 
    395, 113, 73, 145, 220, 175, 183, 191, 196, 180, 171, 178, 169, 153, 143, 114, 74, 84, 92, 83, 77, 98, 97, 153, 277, 296, 241, 198, 170, 227, 228, 0, 
    367, 147, 115, 151, 207, 185, 197, 223, 214, 205, 204, 206, 185, 176, 181, 121, 54, 57, 61, 54, 53, 65, 50, 80, 145, 202, 213, 170, 158, 228, 243, 0, 
    292, 145, 122, 137, 154, 140, 158, 183, 185, 180, 184, 190, 173, 165, 164, 112, 73, 78, 78, 63, 64, 88, 78, 108, 132, 147, 197, 94, 73, 157, 177, 0, 
    224, 117, 92, 112, 116, 76, 83, 129, 144, 117, 107, 133, 125, 106, 93, 68, 61, 77, 78, 63, 55, 102, 121, 91, 65, 89, 233, 143, 11, 88, 111, 0, 
    203, 94, 65, 108, 128, 59, 52, 101, 128, 81, 41, 77, 100, 74, 47, 48, 63, 78, 90, 78, 68, 131, 180, 132, 66, 17, 167, 221, 23, 53, 107, 0, 
    211, 93, 55, 86, 121, 80, 74, 116, 141, 112, 64, 52, 77, 65, 32, 33, 50, 65, 85, 82, 85, 150, 185, 167, 143, 52, 85, 214, 68, 22, 129, 0, 
    218, 79, 54, 68, 81, 65, 88, 103, 102, 97, 77, 47, 42, 39, 23, 26, 34, 34, 48, 59, 81, 142, 160, 156, 159, 114, 58, 134, 129, 45, 120, 26, 
    210, 50, 43, 45, 53, 30, 34, 57, 62, 57, 55, 50, 45, 39, 27, 41, 64, 55, 55, 60, 103, 161, 177, 170, 153, 133, 55, 32, 110, 92, 89, 9, 
    225, 46, 56, 43, 59, 63, 43, 49, 56, 60, 60, 62, 64, 64, 55, 53, 85, 99, 83, 58, 104, 173, 182, 181, 152, 134, 69, 11, 78, 75, 23, 0, 
    246, 54, 65, 65, 79, 113, 100, 67, 59, 60, 62, 66, 74, 82, 85, 78, 88, 113, 88, 38, 69, 144, 149, 150, 141, 129, 99, 76, 133, 128, 49, 0, 
    240, 57, 68, 74, 82, 104, 119, 88, 62, 59, 68, 75, 79, 82, 85, 85, 81, 110, 111, 62, 74, 124, 122, 116, 120, 115, 109, 111, 143, 157, 149, 0, 
    228, 37, 60, 67, 68, 66, 71, 83, 70, 65, 71, 74, 77, 78, 81, 88, 84, 101, 127, 103, 96, 120, 119, 105, 103, 108, 108, 111, 121, 151, 200, 0, 
    203, 4, 54, 79, 72, 66, 51, 55, 68, 71, 74, 77, 84, 87, 89, 96, 105, 141, 158, 123, 106, 111, 114, 101, 99, 114, 105, 100, 108, 125, 175, 41, 
    237, 33, 46, 58, 60, 65, 59, 43, 72, 98, 92, 93, 91, 72, 68, 92, 108, 174, 204, 135, 106, 109, 108, 103, 96, 102, 100, 94, 105, 105, 105, 43, 
    271, 84, 53, 48, 54, 57, 62, 65, 83, 108, 126, 129, 100, 42, 8, 49, 78, 136, 190, 145, 114, 112, 102, 93, 98, 100, 93, 99, 112, 98, 71, 42, 
    256, 127, 75, 61, 63, 41, 44, 75, 88, 88, 127, 155, 110, 41, 1, 34, 69, 106, 142, 123, 109, 102, 96, 92, 97, 97, 89, 96, 101, 86, 78, 50, 
    236, 127, 84, 71, 67, 17, 0, 50, 68, 63, 91, 128, 112, 83, 68, 78, 86, 96, 106, 99, 95, 99, 98, 90, 84, 80, 80, 85, 80, 80, 84, 51, 
    229, 116, 86, 72, 74, 37, 12, 48, 73, 82, 105, 114, 104, 91, 87, 92, 94, 95, 100, 96, 91, 89, 93, 105, 93, 64, 70, 85, 80, 78, 83, 46, 
    224, 123, 110, 94, 98, 88, 78, 85, 91, 92, 96, 99, 97, 93, 90, 93, 94, 97, 102, 93, 88, 91, 90, 102, 98, 69, 72, 85, 83, 79, 82, 42, 
    200, 113, 113, 104, 102, 96, 95, 97, 94, 93, 96, 97, 100, 103, 102, 98, 96, 96, 86, 77, 82, 88, 86, 92, 90, 77, 81, 86, 85, 84, 79, 42, 
    159, 86, 90, 98, 99, 95, 95, 104, 105, 102, 106, 106, 102, 97, 94, 89, 99, 122, 88, 48, 73, 89, 83, 83, 82, 82, 85, 86, 89, 84, 74, 51, 
    150, 82, 85, 95, 100, 100, 100, 105, 106, 99, 94, 95, 95, 93, 90, 85, 106, 144, 96, 39, 73, 91, 83, 80, 83, 86, 88, 88, 91, 77, 70, 74, 
    151, 91, 90, 96, 97, 94, 92, 94, 94, 94, 91, 91, 92, 91, 91, 87, 112, 155, 100, 42, 76, 88, 78, 81, 83, 86, 91, 94, 83, 67, 72, 92, 
    144, 92, 89, 93, 92, 91, 92, 94, 95, 97, 97, 96, 97, 95, 96, 96, 122, 168, 115, 51, 77, 84, 82, 82, 82, 85, 94, 94, 71, 62, 91, 98, 
    156, 125, 126, 127, 127, 126, 128, 130, 130, 131, 129, 125, 120, 114, 107, 102, 120, 165, 151, 101, 108, 115, 114, 113, 112, 112, 122, 122, 89, 82, 106, 106, 
    
    -- channel=35
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=36
    0, 153, 149, 77, 65, 122, 143, 145, 149, 161, 177, 166, 161, 180, 185, 208, 190, 166, 180, 189, 203, 199, 188, 191, 207, 199, 178, 196, 209, 186, 187, 450, 
    0, 20, 39, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 3, 45, 28, 0, 0, 5, 28, 12, 0, 10, 44, 33, 0, 29, 51, 8, 4, 531, 
    0, 17, 45, 0, 0, 0, 0, 0, 0, 0, 31, 0, 0, 0, 0, 35, 35, 0, 0, 6, 22, 0, 0, 1, 48, 34, 0, 30, 59, 0, 0, 535, 
    0, 28, 51, 0, 0, 0, 1, 2, 0, 0, 43, 12, 0, 5, 0, 13, 34, 0, 0, 66, 57, 0, 0, 0, 45, 38, 0, 26, 62, 0, 5, 534, 
    0, 39, 62, 0, 0, 0, 4, 17, 0, 4, 53, 24, 0, 21, 0, 0, 4, 0, 2, 123, 55, 0, 0, 0, 39, 42, 0, 20, 50, 0, 9, 527, 
    0, 40, 76, 0, 0, 0, 4, 29, 0, 13, 54, 27, 0, 46, 22, 0, 0, 0, 0, 156, 36, 0, 0, 0, 0, 32, 0, 14, 33, 0, 13, 517, 
    0, 53, 103, 0, 0, 0, 11, 26, 0, 31, 55, 26, 0, 67, 81, 14, 3, 0, 0, 54, 0, 0, 0, 0, 0, 0, 0, 11, 29, 0, 4, 503, 
    0, 29, 90, 0, 0, 0, 0, 0, 0, 25, 32, 10, 0, 52, 58, 44, 43, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 459, 
    0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 75, 53, 28, 18, 11, 0, 29, 0, 0, 0, 0, 0, 0, 0, 0, 356, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 102, 0, 0, 264, 
    0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 0, 0, 0, 0, 0, 0, 8, 71, 27, 0, 78, 170, 35, 0, 207, 
    0, 0, 0, 0, 0, 12, 19, 0, 0, 22, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 22, 129, 142, 0, 10, 176, 89, 0, 183, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 62, 188, 15, 0, 155, 112, 0, 151, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 2, 30, 31, 23, 28, 7, 13, 0, 0, 0, 0, 8, 129, 107, 0, 87, 84, 0, 124, 
    0, 0, 9, 13, 23, 37, 16, 0, 0, 0, 0, 14, 8, 10, 25, 10, 0, 5, 3, 2, 0, 0, 0, 0, 12, 58, 151, 78, 55, 74, 7, 140, 
    0, 0, 0, 12, 3, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 18, 31, 147, 190, 96, 119, 140, 229, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 90, 45, 0, 0, 0, 10, 13, 87, 124, 20, 56, 141, 297, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 86, 53, 0, 2, 6, 13, 10, 36, 22, 0, 0, 48, 309, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 13, 0, 2, 18, 19, 3, 1, 0, 0, 0, 0, 251, 
    0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 175, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 107, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 50, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 79, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 55, 104, 45, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 62, 
    0, 0, 0, 0, 0, 9, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51, 
    0, 0, 0, 0, 0, 18, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 55, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 54, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 13, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    
    -- channel=37
    196, 128, 112, 142, 172, 171, 169, 174, 180, 181, 174, 181, 192, 192, 195, 182, 184, 194, 199, 202, 194, 192, 199, 201, 190, 190, 201, 195, 187, 198, 204, 10, 
    165, 4, 0, 34, 62, 42, 26, 27, 37, 34, 22, 31, 41, 37, 40, 26, 27, 42, 40, 35, 18, 26, 43, 42, 30, 30, 47, 36, 22, 40, 48, 0, 
    163, 0, 0, 32, 60, 41, 25, 25, 37, 31, 17, 25, 38, 30, 35, 27, 23, 39, 35, 3, 0, 23, 52, 44, 28, 28, 47, 34, 18, 41, 45, 0, 
    165, 0, 0, 30, 59, 40, 24, 21, 43, 35, 15, 23, 37, 25, 32, 32, 23, 37, 30, 0, 0, 23, 54, 45, 29, 25, 44, 31, 19, 42, 41, 0, 
    168, 3, 0, 28, 58, 41, 26, 20, 41, 32, 14, 22, 37, 18, 14, 22, 16, 39, 24, 0, 0, 68, 73, 43, 26, 18, 38, 29, 21, 42, 38, 0, 
    164, 1, 0, 24, 58, 42, 31, 25, 46, 32, 15, 25, 39, 10, 0, 8, 6, 26, 13, 0, 0, 40, 44, 38, 33, 15, 30, 26, 22, 41, 32, 0, 
    163, 0, 0, 25, 61, 38, 28, 30, 44, 28, 17, 29, 35, 13, 6, 8, 0, 0, 0, 0, 0, 0, 0, 0, 21, 35, 37, 23, 10, 34, 32, 0, 
    143, 0, 0, 22, 51, 20, 17, 27, 30, 18, 18, 30, 25, 10, 18, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 10, 0, 18, 19, 0, 
    92, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 6, 0, 0, 5, 0, 0, 0, 0, 0, 3, 10, 0, 26, 43, 15, 0, 0, 0, 0, 0, 0, 
    53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 24, 31, 43, 52, 0, 0, 0, 0, 0, 
    48, 0, 0, 0, 9, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 50, 52, 14, 0, 42, 32, 0, 0, 0, 0, 
    67, 16, 0, 15, 30, 0, 0, 18, 36, 24, 6, 8, 20, 15, 0, 0, 0, 0, 6, 4, 6, 56, 88, 81, 54, 0, 31, 30, 0, 0, 0, 0, 
    81, 20, 0, 1, 0, 0, 0, 19, 38, 33, 18, 14, 12, 0, 0, 0, 0, 0, 6, 8, 17, 58, 66, 39, 26, 0, 9, 27, 0, 0, 0, 0, 
    80, 6, 0, 0, 0, 0, 0, 21, 20, 5, 2, 8, 16, 10, 4, 17, 29, 27, 29, 23, 29, 51, 43, 21, 8, 0, 0, 0, 0, 0, 0, 0, 
    88, 3, 0, 1, 19, 23, 30, 38, 40, 40, 34, 30, 36, 39, 29, 32, 44, 45, 34, 12, 12, 29, 26, 22, 13, 5, 0, 0, 0, 0, 0, 0, 
    100, 18, 28, 30, 40, 53, 63, 60, 51, 41, 36, 32, 27, 22, 14, 7, 7, 7, 0, 0, 0, 0, 9, 13, 13, 10, 0, 0, 37, 35, 5, 0, 
    102, 16, 12, 1, 8, 28, 35, 28, 19, 14, 9, 3, 0, 0, 0, 0, 0, 2, 0, 0, 0, 24, 25, 22, 13, 8, 0, 11, 61, 68, 45, 0, 
    93, 0, 0, 0, 0, 6, 12, 16, 8, 0, 0, 0, 0, 0, 0, 0, 0, 14, 21, 12, 28, 52, 38, 23, 12, 7, 1, 0, 6, 0, 0, 0, 
    72, 0, 0, 2, 17, 26, 18, 0, 0, 0, 0, 0, 1, 9, 15, 19, 14, 21, 24, 12, 18, 30, 23, 13, 6, 0, 0, 0, 0, 0, 5, 0, 
    86, 0, 10, 34, 41, 31, 12, 0, 0, 4, 10, 17, 21, 16, 4, 0, 0, 3, 28, 14, 9, 13, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    107, 25, 38, 25, 5, 0, 0, 0, 4, 18, 22, 18, 9, 0, 0, 0, 0, 0, 29, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    97, 23, 12, 5, 2, 0, 0, 0, 0, 0, 0, 11, 3, 0, 0, 0, 0, 3, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    84, 13, 3, 1, 0, 0, 0, 0, 0, 0, 0, 16, 10, 0, 0, 0, 5, 18, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    85, 21, 0, 0, 0, 0, 0, 0, 0, 0, 13, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    83, 25, 5, 0, 0, 0, 0, 1, 7, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    62, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=38
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=39
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    
    -- channel=40
    131, 257, 238, 202, 222, 258, 268, 267, 268, 272, 275, 261, 263, 271, 272, 281, 264, 262, 269, 276, 283, 275, 270, 275, 282, 270, 266, 279, 276, 262, 270, 350, 
    70, 283, 270, 217, 222, 269, 286, 277, 273, 284, 286, 268, 263, 273, 273, 287, 276, 260, 270, 280, 285, 261, 257, 272, 286, 277, 266, 283, 284, 262, 270, 389, 
    61, 276, 264, 213, 213, 258, 279, 270, 261, 275, 279, 263, 250, 266, 263, 280, 276, 259, 269, 283, 258, 211, 228, 260, 283, 276, 261, 281, 285, 256, 265, 387, 
    56, 271, 259, 205, 203, 244, 270, 265, 245, 264, 274, 254, 240, 260, 250, 264, 273, 255, 269, 285, 236, 181, 208, 253, 278, 273, 255, 275, 277, 255, 261, 384, 
    52, 268, 257, 194, 193, 233, 256, 254, 235, 256, 267, 248, 233, 255, 242, 235, 252, 234, 268, 295, 218, 151, 193, 247, 273, 271, 245, 262, 267, 253, 258, 375, 
    42, 258, 254, 181, 178, 219, 242, 246, 229, 247, 257, 242, 229, 254, 240, 200, 218, 213, 245, 280, 202, 141, 177, 214, 243, 259, 232, 244, 253, 240, 251, 364, 
    33, 248, 243, 168, 162, 211, 224, 229, 219, 234, 241, 231, 228, 243, 236, 215, 217, 202, 186, 205, 169, 99, 110, 118, 130, 193, 211, 227, 235, 210, 226, 345, 
    19, 220, 216, 159, 142, 188, 179, 187, 192, 206, 212, 208, 215, 221, 230, 236, 215, 177, 140, 146, 147, 103, 103, 78, 55, 114, 165, 191, 197, 156, 178, 295, 
    0, 163, 166, 135, 105, 131, 124, 132, 142, 152, 159, 161, 176, 177, 187, 209, 211, 182, 169, 162, 153, 144, 137, 94, 78, 83, 128, 160, 150, 107, 118, 218, 
    0, 112, 119, 100, 86, 108, 105, 94, 101, 112, 115, 117, 132, 142, 157, 181, 187, 167, 160, 159, 150, 128, 125, 127, 132, 101, 101, 170, 153, 107, 91, 170, 
    0, 94, 106, 99, 119, 139, 122, 90, 94, 124, 123, 115, 133, 159, 168, 172, 170, 155, 148, 155, 151, 114, 132, 163, 165, 159, 90, 178, 200, 133, 105, 155, 
    13, 109, 136, 117, 128, 155, 134, 102, 123, 162, 177, 161, 164, 183, 187, 180, 167, 148, 146, 158, 154, 124, 144, 192, 217, 214, 101, 133, 230, 145, 116, 149, 
    31, 131, 145, 122, 118, 139, 132, 125, 131, 160, 196, 187, 173, 187, 195, 184, 168, 162, 156, 165, 159, 140, 149, 185, 214, 231, 164, 94, 206, 154, 97, 135, 
    39, 133, 145, 135, 119, 127, 125, 120, 135, 166, 195, 209, 205, 210, 218, 207, 204, 206, 198, 196, 184, 163, 162, 176, 185, 204, 207, 111, 131, 134, 73, 114, 
    47, 152, 160, 156, 145, 164, 165, 175, 193, 205, 219, 235, 242, 240, 246, 238, 231, 235, 231, 217, 180, 147, 143, 161, 173, 179, 208, 151, 75, 113, 92, 111, 
    62, 177, 176, 187, 187, 202, 216, 218, 223, 234, 241, 246, 251, 254, 255, 244, 219, 216, 216, 203, 147, 114, 126, 149, 167, 176, 199, 182, 111, 147, 162, 154, 
    54, 187, 191, 200, 184, 170, 202, 229, 239, 244, 249, 251, 247, 239, 229, 222, 197, 185, 200, 205, 161, 130, 146, 153, 171, 177, 185, 192, 163, 165, 182, 206, 
    55, 192, 173, 158, 155, 163, 190, 225, 243, 242, 234, 227, 221, 216, 210, 209, 208, 190, 197, 214, 193, 160, 169, 177, 178, 179, 182, 180, 146, 131, 156, 228, 
    56, 162, 140, 160, 185, 201, 200, 213, 223, 216, 211, 213, 217, 220, 221, 217, 215, 191, 185, 206, 201, 179, 183, 195, 188, 186, 173, 152, 127, 105, 93, 195, 
    53, 183, 176, 189, 199, 205, 212, 205, 200, 212, 221, 223, 221, 219, 214, 201, 185, 158, 162, 191, 198, 189, 189, 196, 181, 156, 139, 127, 104, 87, 79, 134, 
    66, 208, 195, 190, 200, 206, 217, 215, 201, 206, 208, 209, 210, 216, 195, 155, 131, 103, 126, 182, 196, 187, 176, 162, 147, 131, 126, 108, 87, 92, 74, 69, 
    36, 187, 210, 212, 211, 213, 205, 197, 177, 164, 160, 175, 203, 218, 186, 137, 121, 101, 114, 161, 166, 154, 143, 138, 133, 118, 102, 88, 81, 75, 60, 52, 
    17, 164, 200, 206, 205, 210, 181, 149, 139, 133, 123, 148, 192, 214, 205, 162, 137, 119, 101, 122, 135, 134, 134, 124, 99, 89, 87, 79, 63, 51, 51, 46, 
    24, 135, 179, 192, 195, 207, 179, 140, 136, 143, 141, 146, 169, 178, 168, 139, 120, 114, 109, 123, 129, 119, 105, 92, 91, 89, 79, 65, 53, 48, 41, 39, 
    29, 129, 171, 184, 185, 197, 188, 154, 142, 142, 132, 115, 116, 121, 121, 118, 120, 120, 114, 109, 100, 91, 91, 85, 89, 83, 67, 54, 53, 46, 37, 42, 
    25, 116, 141, 148, 141, 142, 142, 121, 108, 104, 98, 97, 104, 110, 113, 109, 106, 97, 84, 86, 89, 90, 80, 65, 68, 73, 60, 48, 49, 47, 42, 47, 
    7, 79, 84, 89, 87, 88, 87, 84, 88, 93, 94, 92, 90, 87, 86, 85, 81, 76, 89, 97, 84, 70, 62, 59, 56, 59, 53, 46, 46, 47, 47, 44, 
    0, 56, 52, 55, 60, 65, 66, 66, 71, 74, 71, 69, 68, 72, 74, 76, 71, 74, 103, 99, 71, 58, 59, 55, 49, 50, 46, 45, 45, 49, 44, 31, 
    0, 47, 42, 39, 43, 49, 50, 49, 51, 58, 62, 65, 70, 75, 73, 70, 58, 57, 96, 101, 64, 53, 51, 46, 47, 45, 45, 45, 43, 48, 29, 12, 
    0, 38, 36, 35, 41, 46, 49, 51, 56, 62, 68, 69, 69, 70, 65, 57, 42, 38, 83, 95, 60, 45, 42, 44, 43, 43, 41, 41, 47, 36, 11, 0, 
    0, 39, 41, 44, 48, 52, 53, 55, 57, 59, 61, 60, 58, 57, 46, 33, 15, 14, 64, 84, 50, 37, 40, 40, 42, 41, 35, 42, 44, 18, 0, 0, 
    0, 11, 14, 14, 16, 17, 17, 18, 19, 19, 19, 18, 15, 14, 7, 0, 0, 0, 13, 33, 15, 10, 9, 10, 12, 12, 10, 10, 8, 1, 0, 0, 
    
    -- channel=41
    295, 365, 340, 328, 349, 369, 369, 365, 364, 364, 355, 344, 341, 342, 341, 340, 330, 330, 336, 341, 340, 330, 327, 332, 334, 330, 333, 337, 330, 326, 333, 301, 
    245, 213, 199, 202, 212, 206, 193, 179, 172, 167, 154, 138, 133, 125, 122, 121, 119, 124, 119, 113, 98, 84, 89, 103, 109, 111, 118, 118, 107, 106, 113, 63, 
    229, 185, 172, 178, 187, 175, 165, 156, 148, 142, 127, 117, 113, 106, 106, 109, 110, 115, 111, 87, 44, 34, 70, 95, 101, 101, 107, 106, 98, 97, 101, 50, 
    220, 174, 156, 157, 164, 150, 138, 128, 125, 119, 108, 102, 100, 96, 91, 96, 98, 106, 106, 91, 55, 55, 86, 94, 95, 92, 96, 92, 87, 94, 97, 45, 
    206, 157, 141, 138, 143, 129, 119, 108, 105, 100, 91, 90, 94, 90, 72, 65, 64, 82, 96, 72, 50, 90, 115, 96, 88, 80, 79, 74, 73, 88, 91, 39, 
    186, 129, 116, 113, 119, 104, 95, 89, 89, 81, 71, 82, 89, 82, 60, 46, 42, 55, 75, 76, 67, 85, 74, 51, 59, 64, 61, 55, 58, 73, 72, 27, 
    172, 110, 100, 101, 110, 86, 70, 60, 62, 54, 51, 67, 73, 71, 76, 87, 65, 27, 0, 0, 28, 43, 0, 0, 0, 2, 46, 48, 36, 36, 28, 2, 
    130, 65, 67, 74, 73, 34, 14, 10, 16, 10, 17, 40, 44, 40, 56, 94, 82, 64, 52, 54, 100, 127, 82, 19, 0, 0, 0, 0, 0, 0, 0, 0, 
    79, 2, 16, 30, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 56, 74, 111, 149, 179, 188, 184, 169, 162, 152, 89, 22, 0, 0, 0, 0, 0, 
    78, 18, 26, 42, 47, 27, 17, 5, 0, 0, 0, 0, 0, 19, 49, 62, 83, 129, 156, 160, 153, 151, 145, 140, 143, 103, 82, 66, 35, 21, 9, 0, 
    123, 104, 110, 123, 146, 142, 111, 86, 85, 97, 92, 92, 112, 140, 150, 139, 141, 156, 159, 159, 163, 169, 191, 211, 172, 90, 57, 75, 95, 101, 88, 52, 
    171, 182, 173, 158, 162, 153, 143, 151, 178, 200, 193, 185, 189, 201, 192, 169, 163, 163, 164, 172, 182, 186, 189, 182, 170, 140, 74, 41, 60, 93, 106, 86, 
    192, 199, 177, 149, 128, 112, 127, 156, 171, 168, 182, 200, 201, 200, 199, 196, 192, 187, 188, 189, 184, 179, 152, 92, 71, 86, 78, 41, 29, 63, 93, 77, 
    196, 189, 159, 151, 152, 138, 157, 190, 195, 184, 192, 219, 242, 246, 244, 253, 265, 267, 254, 232, 199, 168, 119, 65, 41, 38, 56, 23, 0, 28, 90, 68, 
    218, 215, 201, 203, 220, 248, 272, 274, 271, 263, 252, 250, 262, 267, 261, 251, 247, 242, 223, 181, 126, 85, 51, 39, 47, 50, 64, 55, 24, 53, 123, 95, 
    229, 231, 229, 233, 240, 256, 275, 279, 262, 245, 238, 235, 231, 224, 217, 200, 173, 151, 136, 102, 63, 48, 41, 47, 59, 70, 87, 116, 159, 193, 196, 135, 
    223, 223, 210, 187, 173, 173, 196, 223, 227, 221, 211, 201, 188, 171, 154, 145, 140, 138, 138, 131, 125, 126, 112, 95, 83, 85, 92, 110, 139, 147, 148, 127, 
    216, 190, 162, 141, 154, 178, 193, 205, 208, 196, 179, 169, 166, 163, 160, 163, 167, 161, 154, 155, 165, 164, 139, 118, 108, 101, 96, 88, 70, 26, 33, 69, 
    203, 176, 172, 202, 241, 259, 233, 192, 176, 172, 178, 185, 193, 198, 195, 185, 174, 157, 140, 134, 139, 135, 120, 117, 113, 95, 75, 51, 25, 6, 25, 39, 
    235, 234, 245, 256, 250, 231, 211, 191, 184, 198, 214, 213, 202, 182, 156, 123, 91, 88, 112, 125, 127, 125, 112, 96, 73, 55, 44, 36, 37, 47, 44, 15, 
    235, 257, 271, 250, 218, 200, 197, 196, 190, 194, 192, 181, 169, 141, 94, 57, 44, 59, 102, 123, 117, 102, 81, 60, 53, 56, 59, 67, 79, 90, 75, 11, 
    204, 213, 234, 228, 218, 204, 178, 155, 143, 129, 119, 137, 157, 154, 129, 116, 129, 140, 129, 96, 74, 67, 66, 65, 69, 79, 84, 85, 87, 82, 64, 42, 
    192, 191, 202, 201, 198, 179, 139, 111, 115, 125, 129, 150, 166, 164, 164, 177, 176, 162, 131, 84, 73, 83, 86, 86, 86, 87, 92, 94, 89, 69, 66, 72, 
    200, 199, 186, 188, 195, 191, 172, 170, 185, 200, 201, 176, 125, 92, 95, 122, 133, 133, 125, 110, 103, 99, 99, 104, 112, 114, 108, 108, 97, 87, 94, 86, 
    198, 200, 189, 187, 182, 177, 182, 196, 189, 166, 143, 113, 79, 75, 93, 114, 124, 126, 121, 108, 101, 102, 105, 111, 124, 122, 108, 106, 108, 110, 113, 96, 
    168, 149, 130, 116, 105, 94, 102, 121, 121, 112, 105, 98, 101, 117, 133, 133, 119, 106, 102, 101, 104, 111, 119, 114, 105, 98, 104, 114, 116, 119, 119, 99, 
    130, 95, 74, 66, 72, 79, 89, 105, 114, 117, 122, 124, 119, 116, 112, 104, 102, 119, 136, 134, 120, 113, 108, 107, 103, 99, 111, 121, 123, 124, 119, 89, 
    123, 101, 92, 92, 101, 109, 116, 118, 117, 110, 104, 102, 106, 115, 118, 112, 114, 140, 164, 143, 112, 106, 108, 112, 110, 112, 121, 124, 123, 118, 101, 69, 
    116, 110, 110, 113, 114, 113, 114, 113, 112, 113, 118, 122, 127, 135, 132, 118, 113, 129, 133, 111, 105, 109, 110, 109, 112, 118, 123, 124, 117, 100, 69, 51, 
    106, 102, 107, 115, 122, 125, 126, 130, 133, 135, 138, 139, 136, 131, 116, 95, 88, 109, 116, 104, 108, 113, 107, 110, 117, 119, 121, 120, 106, 77, 50, 53, 
    115, 116, 121, 128, 130, 131, 129, 129, 128, 125, 117, 109, 101, 93, 77, 58, 58, 87, 105, 102, 109, 108, 108, 115, 117, 118, 119, 114, 90, 55, 50, 67, 
    69, 49, 48, 49, 47, 44, 41, 39, 36, 34, 32, 33, 35, 39, 41, 38, 42, 47, 34, 27, 43, 48, 49, 51, 54, 56, 54, 51, 41, 39, 55, 65, 
    
    -- channel=42
    93, 108, 87, 70, 98, 109, 106, 104, 104, 104, 99, 85, 89, 86, 84, 89, 72, 80, 83, 87, 86, 76, 76, 80, 83, 74, 78, 85, 77, 72, 81, 119, 
    175, 177, 150, 128, 167, 179, 176, 165, 166, 168, 158, 141, 144, 141, 138, 145, 122, 134, 137, 140, 136, 117, 126, 127, 135, 122, 130, 141, 128, 118, 137, 164, 
    171, 166, 139, 116, 154, 164, 163, 149, 148, 155, 143, 127, 131, 136, 127, 142, 120, 128, 133, 137, 109, 94, 122, 123, 132, 118, 127, 139, 125, 114, 135, 161, 
    165, 154, 127, 100, 140, 145, 148, 129, 128, 141, 126, 114, 117, 127, 111, 136, 118, 121, 133, 136, 92, 74, 115, 120, 131, 114, 120, 134, 118, 112, 130, 155, 
    157, 142, 118, 84, 127, 126, 133, 114, 110, 125, 111, 104, 105, 123, 97, 116, 111, 109, 137, 123, 56, 78, 126, 120, 130, 108, 108, 124, 108, 109, 127, 149, 
    147, 127, 108, 65, 114, 107, 116, 97, 93, 110, 96, 95, 97, 116, 82, 90, 96, 91, 124, 122, 47, 66, 111, 109, 127, 107, 92, 107, 95, 101, 117, 138, 
    138, 111, 94, 48, 99, 89, 91, 79, 77, 89, 76, 83, 85, 100, 76, 84, 76, 74, 85, 83, 47, 59, 76, 57, 81, 104, 87, 92, 76, 74, 93, 117, 
    116, 94, 80, 37, 80, 75, 67, 68, 64, 68, 59, 69, 76, 78, 66, 87, 80, 76, 76, 65, 47, 58, 58, 17, 22, 51, 68, 76, 56, 38, 66, 86, 
    83, 69, 59, 33, 57, 56, 45, 46, 48, 46, 39, 50, 61, 59, 67, 93, 79, 72, 68, 70, 65, 63, 54, 21, 40, 34, 52, 51, 22, 8, 34, 53, 
    51, 48, 40, 28, 47, 41, 24, 33, 32, 33, 26, 37, 50, 54, 72, 86, 71, 74, 78, 83, 74, 68, 68, 30, 38, 26, 44, 64, 2, 3, 23, 34, 
    34, 42, 42, 29, 50, 46, 31, 24, 37, 48, 35, 42, 62, 75, 91, 92, 79, 73, 77, 77, 68, 52, 69, 63, 63, 17, 0, 70, 19, 9, 31, 32, 
    34, 58, 53, 31, 64, 68, 46, 41, 58, 78, 73, 64, 82, 107, 113, 100, 85, 78, 75, 76, 65, 48, 73, 78, 79, 46, 0, 48, 41, 0, 35, 39, 
    48, 72, 71, 50, 65, 61, 54, 51, 76, 99, 103, 100, 107, 125, 123, 108, 96, 85, 79, 85, 70, 59, 83, 76, 72, 61, 5, 19, 54, 0, 17, 38, 
    64, 86, 79, 55, 65, 59, 55, 77, 100, 106, 115, 119, 126, 132, 128, 117, 117, 109, 103, 101, 80, 71, 79, 66, 64, 54, 32, 1, 25, 0, 5, 23, 
    87, 95, 88, 72, 76, 87, 90, 102, 117, 128, 135, 137, 143, 149, 148, 133, 133, 135, 123, 107, 73, 68, 62, 54, 55, 50, 56, 8, 0, 0, 0, 10, 
    103, 106, 107, 104, 98, 114, 131, 142, 152, 154, 157, 158, 161, 160, 157, 146, 135, 132, 122, 99, 51, 47, 43, 41, 52, 51, 66, 23, 6, 22, 9, 9, 
    113, 127, 124, 114, 112, 126, 154, 165, 167, 168, 167, 163, 159, 153, 145, 134, 118, 113, 112, 87, 41, 39, 44, 47, 59, 58, 68, 36, 20, 43, 43, 43, 
    118, 122, 120, 117, 114, 122, 139, 160, 168, 164, 161, 155, 148, 138, 126, 114, 102, 90, 98, 90, 57, 61, 68, 65, 69, 68, 67, 48, 42, 45, 32, 59, 
    111, 117, 114, 116, 114, 128, 142, 147, 154, 150, 149, 140, 132, 124, 115, 106, 102, 92, 98, 95, 80, 80, 82, 79, 74, 68, 60, 47, 37, 19, 20, 70, 
    120, 115, 104, 118, 135, 147, 150, 142, 135, 137, 131, 129, 126, 122, 115, 104, 93, 77, 98, 99, 89, 88, 85, 82, 66, 58, 53, 35, 17, 11, 9, 38, 
    114, 128, 136, 147, 149, 146, 141, 133, 117, 124, 129, 130, 127, 124, 96, 78, 69, 48, 84, 100, 87, 85, 79, 71, 58, 45, 30, 18, 10, 10, 4, 6, 
    101, 148, 149, 147, 143, 139, 129, 119, 110, 114, 109, 123, 123, 119, 84, 54, 47, 34, 67, 82, 77, 73, 66, 55, 34, 26, 21, 10, 4, 4, 0, 0, 
    82, 132, 141, 138, 138, 136, 108, 97, 92, 94, 83, 104, 116, 112, 78, 51, 46, 40, 64, 69, 58, 53, 43, 33, 24, 23, 12, 3, 0, 0, 0, 0, 
    65, 117, 127, 125, 129, 131, 94, 76, 78, 80, 78, 94, 98, 90, 68, 59, 57, 49, 52, 46, 39, 32, 33, 30, 21, 10, 1, 0, 0, 0, 0, 0, 
    61, 104, 115, 112, 114, 114, 86, 72, 72, 71, 69, 81, 77, 68, 56, 48, 45, 40, 39, 36, 32, 27, 19, 8, 15, 12, 0, 0, 0, 0, 0, 0, 
    52, 81, 94, 90, 90, 85, 69, 66, 65, 59, 53, 47, 40, 37, 38, 37, 36, 32, 32, 31, 18, 9, 7, 6, 13, 5, 0, 0, 0, 0, 0, 0, 
    30, 52, 56, 53, 51, 46, 41, 40, 37, 29, 22, 21, 21, 26, 29, 28, 22, 22, 28, 15, 7, 6, 3, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    7, 13, 11, 8, 10, 11, 10, 11, 15, 15, 12, 12, 15, 18, 17, 12, 1, 8, 33, 21, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 5, 6, 4, 5, 7, 8, 3, 0, 6, 40, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 5, 8, 4, 0, 0, 0, 35, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=43
    146, 347, 333, 301, 310, 359, 378, 381, 384, 393, 400, 398, 399, 416, 422, 425, 418, 407, 417, 425, 435, 433, 426, 430, 434, 427, 418, 430, 432, 418, 422, 439, 
    0, 172, 170, 120, 106, 148, 165, 158, 151, 163, 174, 161, 158, 170, 173, 188, 183, 163, 169, 176, 181, 164, 157, 176, 190, 187, 171, 184, 192, 172, 171, 346, 
    0, 166, 168, 120, 106, 144, 163, 162, 152, 163, 176, 158, 147, 157, 161, 177, 183, 165, 166, 170, 149, 98, 114, 166, 188, 184, 165, 182, 191, 164, 161, 341, 
    0, 173, 174, 122, 104, 141, 166, 168, 150, 164, 183, 162, 146, 156, 153, 160, 178, 163, 163, 170, 141, 83, 107, 158, 183, 183, 161, 176, 185, 160, 165, 339, 
    0, 179, 178, 122, 103, 143, 164, 169, 153, 170, 186, 166, 149, 158, 146, 132, 143, 139, 155, 199, 143, 57, 104, 155, 178, 183, 156, 164, 177, 156, 166, 332, 
    0, 173, 174, 114, 92, 137, 160, 175, 160, 174, 183, 164, 154, 171, 149, 106, 108, 116, 135, 179, 134, 54, 77, 102, 133, 166, 152, 157, 166, 146, 158, 323, 
    0, 172, 173, 108, 89, 138, 155, 160, 154, 171, 174, 160, 157, 176, 167, 147, 142, 91, 64, 82, 51, 0, 0, 0, 0, 56, 123, 156, 161, 132, 139, 309, 
    0, 133, 147, 96, 77, 102, 102, 100, 119, 139, 142, 138, 140, 163, 172, 169, 142, 64, 23, 48, 51, 25, 17, 0, 0, 0, 53, 101, 110, 80, 91, 266, 
    0, 50, 76, 43, 14, 12, 12, 19, 37, 57, 64, 69, 76, 89, 89, 116, 121, 111, 117, 130, 130, 126, 135, 98, 53, 55, 44, 73, 62, 17, 27, 180, 
    0, 8, 35, 15, 1, 24, 19, 4, 5, 15, 22, 17, 25, 35, 46, 85, 99, 96, 100, 102, 93, 73, 95, 130, 129, 97, 69, 124, 135, 44, 32, 143, 
    0, 37, 63, 73, 90, 118, 93, 53, 41, 69, 80, 60, 68, 82, 86, 96, 101, 98, 96, 105, 105, 95, 124, 165, 187, 156, 106, 148, 208, 119, 77, 154, 
    0, 86, 125, 115, 102, 126, 109, 85, 101, 142, 156, 140, 118, 111, 110, 109, 104, 101, 108, 127, 141, 128, 151, 201, 236, 221, 126, 120, 189, 148, 78, 160, 
    10, 104, 118, 86, 69, 81, 85, 86, 83, 106, 131, 129, 103, 95, 107, 108, 109, 114, 118, 128, 145, 123, 124, 148, 178, 217, 152, 107, 145, 146, 67, 136, 
    0, 84, 100, 87, 72, 77, 71, 56, 64, 89, 119, 135, 137, 145, 157, 163, 172, 186, 181, 179, 172, 141, 129, 121, 125, 172, 157, 101, 89, 84, 55, 119, 
    0, 107, 122, 127, 127, 138, 150, 150, 154, 155, 164, 175, 178, 180, 186, 187, 181, 188, 188, 179, 138, 89, 90, 101, 117, 139, 161, 115, 78, 87, 102, 147, 
    5, 128, 135, 154, 164, 167, 170, 160, 151, 149, 151, 153, 156, 159, 161, 144, 121, 109, 117, 118, 79, 45, 73, 99, 119, 130, 170, 178, 165, 207, 227, 223, 
    0, 100, 118, 123, 88, 60, 70, 105, 116, 119, 124, 127, 124, 116, 113, 106, 93, 87, 115, 153, 139, 121, 128, 126, 124, 125, 155, 195, 198, 209, 209, 249, 
    0, 85, 57, 37, 31, 45, 71, 95, 111, 108, 95, 88, 88, 98, 113, 133, 144, 142, 149, 188, 185, 158, 149, 139, 129, 125, 140, 141, 101, 91, 116, 219, 
    0, 48, 29, 68, 120, 126, 112, 94, 84, 78, 81, 102, 126, 149, 164, 172, 166, 140, 129, 152, 152, 134, 134, 137, 139, 129, 117, 87, 62, 41, 35, 168, 
    0, 116, 125, 132, 127, 114, 101, 92, 88, 107, 142, 155, 155, 150, 137, 115, 96, 69, 73, 119, 131, 124, 123, 126, 113, 81, 64, 61, 52, 38, 27, 120, 
    10, 142, 124, 102, 88, 93, 107, 119, 120, 117, 124, 121, 119, 115, 91, 37, 16, 9, 33, 104, 128, 111, 90, 74, 62, 67, 76, 73, 71, 73, 37, 77, 
    0, 69, 106, 113, 112, 110, 107, 92, 64, 45, 39, 57, 103, 128, 113, 77, 73, 62, 61, 83, 77, 61, 53, 66, 81, 80, 76, 73, 70, 66, 46, 73, 
    0, 48, 92, 101, 99, 98, 72, 32, 17, 20, 25, 50, 105, 154, 170, 155, 141, 96, 52, 47, 54, 69, 85, 82, 64, 58, 70, 68, 53, 50, 57, 81, 
    0, 49, 78, 91, 96, 112, 105, 76, 79, 96, 89, 82, 83, 92, 95, 84, 81, 70, 69, 83, 92, 85, 67, 63, 73, 84, 78, 61, 60, 64, 65, 85, 
    0, 62, 88, 101, 101, 125, 136, 122, 111, 103, 67, 28, 13, 21, 41, 64, 84, 90, 87, 79, 66, 61, 73, 84, 85, 86, 69, 59, 66, 69, 66, 88, 
    0, 41, 45, 45, 34, 47, 53, 44, 37, 34, 31, 37, 53, 71, 83, 87, 81, 60, 42, 50, 74, 85, 81, 63, 59, 66, 59, 59, 65, 66, 66, 91, 
    0, 0, 0, 0, 0, 4, 13, 22, 43, 68, 81, 84, 77, 64, 55, 54, 54, 52, 75, 101, 89, 69, 63, 53, 55, 61, 62, 62, 66, 68, 68, 87, 
    0, 20, 17, 22, 33, 47, 54, 56, 60, 62, 59, 53, 49, 51, 59, 71, 78, 83, 104, 111, 74, 57, 63, 60, 58, 62, 63, 65, 68, 70, 68, 73, 
    23, 62, 59, 54, 56, 61, 59, 52, 50, 52, 59, 68, 77, 83, 84, 85, 73, 54, 81, 99, 68, 60, 60, 56, 59, 63, 64, 65, 67, 70, 62, 53, 
    24, 61, 64, 62, 65, 71, 73, 74, 78, 85, 90, 89, 84, 79, 72, 68, 49, 27, 66, 97, 69, 55, 53, 55, 59, 61, 59, 60, 65, 67, 49, 48, 
    29, 71, 75, 78, 80, 81, 81, 80, 80, 77, 73, 67, 61, 55, 47, 39, 19, 2, 50, 87, 60, 52, 53, 56, 58, 58, 55, 59, 64, 59, 47, 53, 
    17, 23, 21, 19, 16, 14, 11, 8, 7, 7, 8, 7, 8, 9, 11, 15, 6, 0, 0, 14, 12, 11, 11, 13, 15, 17, 15, 12, 23, 37, 41, 45, 
    
    -- channel=44
    265, 366, 331, 324, 373, 416, 429, 437, 447, 455, 454, 451, 463, 474, 479, 475, 460, 468, 483, 492, 492, 485, 485, 490, 486, 476, 480, 489, 482, 477, 488, 367, 
    257, 317, 279, 266, 319, 356, 363, 363, 373, 385, 382, 374, 389, 399, 404, 404, 384, 392, 402, 412, 406, 391, 399, 410, 411, 398, 407, 416, 403, 399, 418, 325, 
    258, 314, 279, 267, 320, 358, 366, 359, 369, 384, 377, 366, 379, 388, 393, 401, 384, 390, 397, 390, 356, 343, 380, 407, 411, 397, 407, 418, 402, 396, 415, 321, 
    263, 316, 279, 267, 319, 354, 366, 358, 369, 385, 374, 361, 369, 378, 378, 395, 383, 386, 390, 359, 290, 284, 363, 404, 412, 395, 402, 414, 398, 392, 412, 316, 
    271, 323, 282, 262, 316, 350, 364, 354, 361, 381, 371, 356, 362, 369, 350, 366, 363, 371, 378, 331, 253, 280, 367, 398, 407, 388, 390, 401, 388, 390, 409, 310, 
    272, 320, 277, 249, 308, 342, 361, 354, 362, 379, 364, 352, 357, 360, 317, 313, 314, 331, 354, 295, 200, 240, 333, 367, 389, 375, 370, 381, 372, 380, 396, 298, 
    272, 312, 267, 236, 301, 334, 353, 352, 360, 370, 351, 347, 352, 354, 310, 290, 277, 264, 263, 223, 157, 171, 200, 217, 283, 331, 350, 365, 351, 356, 374, 283, 
    259, 296, 257, 228, 293, 315, 322, 327, 341, 346, 332, 335, 338, 335, 319, 311, 260, 186, 132, 98, 74, 81, 69, 47, 107, 215, 293, 326, 304, 299, 327, 249, 
    190, 216, 197, 178, 215, 218, 218, 239, 264, 270, 267, 280, 283, 277, 273, 270, 210, 162, 144, 147, 142, 143, 140, 117, 130, 172, 214, 231, 203, 197, 236, 177, 
    100, 119, 117, 107, 121, 119, 119, 141, 156, 164, 167, 178, 186, 188, 199, 202, 165, 151, 153, 149, 130, 127, 137, 147, 187, 200, 223, 218, 153, 124, 147, 97, 
    52, 83, 89, 96, 125, 133, 114, 110, 125, 140, 135, 137, 154, 166, 175, 166, 141, 135, 138, 129, 111, 121, 173, 208, 215, 171, 212, 266, 199, 136, 127, 80, 
    52, 107, 118, 127, 165, 163, 125, 118, 153, 190, 178, 168, 185, 198, 188, 167, 152, 150, 153, 154, 151, 174, 259, 317, 315, 240, 199, 259, 210, 133, 111, 79, 
    71, 138, 142, 119, 133, 126, 114, 133, 183, 218, 215, 197, 188, 187, 173, 154, 146, 145, 156, 169, 179, 210, 280, 313, 322, 290, 212, 236, 202, 108, 86, 69, 
    85, 140, 133, 110, 111, 97, 98, 128, 158, 179, 200, 204, 204, 208, 205, 202, 207, 210, 210, 217, 223, 249, 286, 285, 284, 278, 218, 181, 159, 77, 57, 40, 
    99, 145, 145, 138, 146, 147, 158, 184, 218, 241, 255, 261, 270, 276, 272, 267, 280, 287, 278, 262, 240, 246, 262, 265, 267, 262, 224, 130, 91, 56, 58, 37, 
    131, 184, 197, 202, 216, 243, 263, 274, 285, 290, 294, 294, 295, 294, 291, 272, 263, 262, 254, 217, 170, 175, 206, 235, 254, 252, 238, 165, 143, 159, 140, 76, 
    139, 194, 210, 214, 210, 224, 249, 267, 275, 280, 282, 279, 274, 266, 257, 237, 219, 221, 226, 201, 163, 186, 221, 241, 249, 245, 243, 222, 244, 287, 248, 139, 
    131, 177, 176, 162, 149, 167, 215, 255, 268, 265, 257, 246, 234, 224, 218, 218, 217, 231, 255, 254, 235, 252, 263, 252, 245, 238, 235, 222, 221, 221, 210, 157, 
    114, 136, 122, 135, 171, 208, 231, 237, 234, 221, 213, 214, 222, 237, 247, 257, 257, 248, 257, 261, 255, 261, 265, 255, 244, 231, 216, 188, 159, 135, 154, 142, 
    111, 134, 150, 201, 239, 250, 236, 216, 204, 206, 226, 246, 259, 265, 259, 240, 219, 207, 232, 251, 250, 251, 252, 241, 214, 187, 156, 118, 91, 77, 92, 97, 
    147, 203, 212, 218, 212, 213, 215, 212, 211, 229, 250, 254, 249, 230, 188, 141, 111, 117, 188, 237, 240, 231, 215, 189, 148, 118, 96, 78, 69, 66, 52, 23, 
    124, 196, 211, 213, 212, 212, 209, 197, 183, 182, 188, 210, 224, 206, 140, 83, 70, 91, 163, 203, 194, 171, 144, 119, 98, 89, 75, 58, 56, 55, 19, 0, 
    82, 167, 202, 206, 206, 190, 151, 120, 106, 105, 119, 175, 220, 217, 167, 131, 129, 129, 147, 141, 120, 109, 99, 87, 72, 57, 42, 31, 28, 15, 0, 0, 
    69, 154, 178, 182, 187, 169, 114, 85, 93, 109, 130, 174, 195, 184, 155, 135, 124, 109, 108, 103, 97, 88, 75, 59, 45, 38, 29, 19, 9, 0, 0, 0, 
    73, 150, 173, 179, 184, 178, 141, 128, 133, 137, 137, 138, 116, 90, 74, 77, 88, 95, 99, 94, 75, 52, 38, 44, 58, 47, 19, 7, 2, 0, 0, 0, 
    64, 123, 143, 139, 131, 122, 105, 98, 90, 73, 60, 55, 57, 68, 78, 85, 83, 71, 61, 50, 41, 37, 37, 35, 40, 23, 2, 0, 0, 0, 0, 0, 
    20, 44, 44, 35, 30, 25, 22, 27, 38, 47, 54, 61, 63, 63, 61, 53, 40, 33, 40, 44, 41, 34, 24, 14, 13, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 11, 21, 36, 42, 41, 37, 32, 27, 26, 26, 27, 50, 79, 62, 28, 16, 12, 7, 2, 0, 0, 0, 2, 2, 0, 0, 
    0, 0, 0, 0, 0, 1, 3, 6, 10, 11, 11, 13, 20, 29, 35, 34, 29, 51, 78, 44, 10, 8, 7, 1, 0, 0, 0, 2, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 6, 11, 19, 27, 33, 34, 31, 26, 19, 8, 28, 56, 26, 2, 3, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 
    0, 0, 0, 3, 8, 13, 18, 22, 25, 26, 25, 21, 14, 5, 0, 0, 0, 0, 37, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=45
    343, 299, 264, 301, 359, 372, 374, 382, 394, 398, 388, 393, 409, 410, 414, 395, 392, 410, 421, 428, 417, 411, 417, 420, 406, 403, 420, 416, 402, 415, 427, 124, 
    416, 282, 239, 288, 359, 361, 350, 354, 374, 376, 357, 365, 384, 384, 390, 369, 359, 385, 393, 394, 369, 369, 391, 393, 378, 373, 400, 391, 368, 390, 408, 50, 
    420, 279, 237, 287, 360, 363, 349, 348, 372, 371, 348, 352, 377, 374, 383, 372, 356, 379, 384, 349, 302, 348, 397, 398, 378, 372, 402, 393, 364, 390, 407, 46, 
    423, 279, 233, 283, 356, 360, 346, 339, 371, 371, 340, 343, 368, 360, 371, 376, 356, 375, 370, 293, 241, 320, 394, 401, 381, 368, 398, 388, 362, 389, 401, 42, 
    429, 282, 229, 278, 351, 356, 345, 332, 364, 363, 332, 334, 360, 342, 335, 353, 342, 370, 353, 229, 204, 345, 407, 397, 378, 356, 384, 377, 358, 387, 394, 39, 
    428, 279, 216, 265, 346, 349, 345, 332, 362, 354, 325, 331, 355, 321, 283, 307, 305, 337, 325, 195, 170, 299, 360, 375, 376, 345, 362, 361, 347, 379, 381, 33, 
    427, 272, 204, 259, 345, 340, 338, 336, 358, 342, 318, 330, 344, 310, 274, 274, 243, 239, 222, 146, 136, 205, 215, 242, 322, 347, 354, 346, 323, 356, 366, 26, 
    400, 260, 204, 251, 330, 313, 316, 331, 340, 322, 311, 325, 323, 297, 286, 262, 199, 151, 124, 84, 72, 108, 81, 82, 184, 264, 315, 310, 274, 311, 326, 11, 
    313, 202, 170, 194, 241, 222, 235, 259, 269, 262, 263, 278, 268, 258, 264, 223, 152, 129, 131, 131, 129, 137, 114, 136, 195, 223, 245, 211, 170, 219, 238, 0, 
    206, 129, 111, 122, 149, 129, 136, 164, 172, 173, 174, 189, 187, 194, 204, 168, 129, 141, 148, 136, 121, 135, 142, 165, 187, 221, 265, 193, 103, 135, 151, 0, 
    142, 102, 95, 116, 142, 118, 103, 121, 154, 147, 133, 150, 167, 174, 173, 149, 130, 135, 139, 120, 102, 150, 212, 228, 193, 150, 249, 237, 121, 110, 126, 0, 
    141, 129, 109, 137, 174, 135, 105, 143, 187, 185, 158, 161, 189, 196, 174, 150, 140, 146, 149, 141, 137, 214, 300, 311, 269, 171, 226, 253, 121, 84, 114, 0, 
    167, 151, 124, 129, 139, 106, 111, 155, 208, 221, 195, 184, 193, 189, 163, 144, 141, 142, 156, 164, 179, 254, 314, 309, 287, 207, 194, 244, 123, 49, 90, 0, 
    181, 149, 119, 109, 112, 94, 112, 165, 195, 201, 200, 198, 208, 206, 191, 193, 203, 199, 206, 207, 222, 273, 295, 282, 271, 225, 158, 167, 100, 38, 69, 0, 
    201, 152, 140, 134, 152, 158, 175, 206, 233, 251, 254, 253, 260, 265, 252, 252, 268, 269, 255, 226, 221, 256, 268, 267, 256, 238, 152, 82, 74, 45, 60, 0, 
    232, 186, 200, 200, 218, 244, 265, 279, 289, 290, 289, 287, 284, 280, 267, 252, 254, 255, 233, 174, 159, 201, 227, 242, 245, 238, 177, 111, 160, 152, 97, 0, 
    251, 208, 214, 200, 211, 251, 277, 280, 281, 282, 277, 268, 258, 249, 237, 217, 217, 232, 217, 157, 153, 207, 229, 241, 239, 234, 208, 186, 242, 253, 195, 0, 
    246, 175, 174, 168, 176, 213, 249, 270, 268, 257, 248, 238, 228, 218, 211, 207, 206, 230, 242, 213, 213, 255, 255, 243, 234, 230, 216, 201, 213, 207, 191, 3, 
    212, 135, 150, 169, 197, 227, 246, 242, 229, 220, 219, 218, 223, 228, 232, 237, 229, 238, 254, 238, 237, 257, 257, 240, 227, 210, 187, 163, 138, 131, 185, 12, 
    216, 136, 170, 217, 247, 253, 236, 216, 208, 216, 225, 238, 247, 247, 233, 213, 189, 210, 253, 245, 238, 246, 243, 215, 183, 161, 134, 96, 76, 86, 124, 0, 
    250, 199, 224, 232, 223, 221, 212, 201, 211, 232, 245, 246, 239, 201, 146, 119, 104, 157, 238, 240, 221, 214, 195, 162, 127, 102, 73, 59, 68, 65, 51, 0, 
    244, 222, 217, 213, 213, 208, 195, 179, 183, 189, 203, 230, 222, 163, 93, 72, 76, 135, 204, 196, 175, 156, 132, 101, 76, 68, 55, 48, 56, 39, 4, 0, 
    212, 205, 206, 204, 204, 167, 125, 117, 118, 121, 160, 217, 223, 172, 114, 107, 114, 140, 167, 142, 114, 99, 80, 61, 58, 50, 31, 27, 24, 6, 0, 0, 
    191, 196, 189, 186, 188, 138, 85, 91, 109, 122, 162, 199, 186, 149, 120, 122, 120, 115, 117, 98, 79, 66, 59, 52, 44, 27, 18, 16, 6, 0, 0, 0, 
    183, 187, 183, 178, 180, 144, 110, 121, 132, 132, 142, 149, 123, 94, 79, 83, 86, 89, 91, 80, 61, 45, 31, 42, 53, 31, 11, 9, 1, 0, 0, 0, 
    156, 150, 150, 139, 132, 109, 91, 100, 97, 82, 72, 65, 64, 70, 78, 82, 71, 63, 64, 52, 34, 28, 29, 43, 39, 10, 1, 5, 1, 0, 5, 0, 
    95, 70, 62, 53, 48, 38, 36, 46, 52, 50, 53, 57, 59, 63, 63, 51, 37, 45, 50, 31, 30, 30, 24, 21, 14, 0, 0, 6, 5, 6, 3, 0, 
    46, 7, 3, 4, 11, 14, 20, 34, 42, 42, 40, 38, 37, 35, 32, 23, 28, 70, 75, 34, 18, 20, 14, 9, 5, 0, 4, 7, 11, 8, 0, 0, 
    29, 0, 0, 2, 5, 6, 9, 16, 20, 18, 18, 19, 24, 30, 34, 27, 36, 84, 70, 8, 6, 15, 9, 6, 0, 2, 7, 11, 16, 0, 0, 0, 
    20, 0, 0, 1, 4, 5, 7, 12, 17, 22, 27, 32, 33, 29, 24, 10, 19, 70, 51, 0, 1, 10, 6, 0, 0, 1, 6, 15, 5, 0, 0, 0, 
    19, 0, 3, 9, 13, 16, 21, 26, 29, 29, 26, 20, 13, 1, 0, 0, 0, 49, 41, 0, 0, 6, 2, 2, 0, 0, 6, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=46
    36, 0, 0, 8, 17, 12, 14, 18, 21, 22, 21, 31, 35, 36, 38, 29, 35, 42, 43, 41, 39, 43, 46, 43, 37, 40, 45, 39, 38, 44, 44, 0, 
    176, 111, 94, 128, 160, 163, 163, 175, 184, 185, 184, 195, 208, 211, 218, 202, 204, 216, 221, 224, 221, 229, 229, 227, 214, 214, 225, 218, 211, 224, 227, 17, 
    187, 127, 107, 138, 173, 180, 174, 181, 197, 197, 191, 200, 216, 215, 226, 210, 207, 218, 223, 219, 225, 239, 236, 234, 220, 219, 232, 224, 212, 230, 235, 21, 
    191, 131, 113, 148, 180, 191, 184, 188, 209, 205, 195, 201, 215, 212, 229, 218, 208, 220, 218, 192, 183, 216, 235, 238, 223, 221, 236, 229, 217, 228, 235, 22, 
    197, 138, 116, 154, 185, 198, 192, 193, 215, 212, 200, 199, 215, 205, 220, 229, 216, 228, 209, 161, 159, 199, 227, 238, 225, 221, 239, 231, 220, 230, 233, 24, 
    206, 149, 117, 159, 190, 204, 200, 197, 218, 217, 203, 201, 214, 196, 199, 219, 212, 227, 210, 131, 128, 197, 234, 248, 234, 218, 236, 231, 222, 235, 233, 25, 
    207, 152, 116, 155, 188, 201, 207, 206, 223, 218, 207, 205, 215, 194, 171, 171, 181, 203, 214, 145, 113, 179, 221, 256, 269, 230, 227, 225, 221, 243, 237, 28, 
    215, 163, 124, 153, 197, 206, 221, 220, 231, 225, 214, 213, 214, 201, 178, 156, 144, 136, 125, 89, 66, 82, 91, 136, 208, 233, 231, 227, 220, 248, 241, 43, 
    207, 166, 133, 149, 194, 200, 209, 222, 230, 225, 220, 221, 213, 206, 197, 160, 110, 74, 48, 34, 30, 30, 21, 38, 86, 164, 194, 194, 190, 217, 227, 57, 
    151, 125, 109, 114, 128, 127, 141, 163, 174, 172, 179, 184, 175, 168, 164, 133, 91, 67, 60, 51, 48, 57, 42, 53, 79, 124, 155, 113, 111, 136, 157, 29, 
    81, 67, 57, 62, 59, 55, 66, 92, 97, 90, 100, 109, 100, 97, 100, 84, 64, 62, 61, 47, 37, 56, 53, 64, 77, 99, 174, 110, 60, 80, 83, 0, 
    47, 31, 28, 55, 66, 46, 40, 52, 62, 58, 46, 61, 72, 70, 66, 58, 55, 58, 59, 47, 38, 70, 106, 117, 92, 68, 159, 164, 66, 70, 60, 0, 
    47, 39, 36, 56, 77, 60, 41, 58, 89, 90, 63, 59, 74, 70, 53, 44, 45, 47, 58, 56, 59, 101, 154, 179, 163, 98, 116, 180, 83, 56, 67, 0, 
    60, 50, 40, 41, 49, 39, 42, 59, 77, 88, 78, 60, 56, 55, 42, 37, 33, 35, 47, 57, 75, 121, 161, 181, 183, 143, 99, 149, 113, 46, 57, 0, 
    58, 37, 29, 25, 23, 7, 16, 35, 53, 66, 74, 73, 70, 69, 62, 68, 78, 76, 80, 88, 116, 151, 172, 172, 168, 155, 94, 82, 88, 34, 28, 0, 
    66, 41, 43, 34, 45, 49, 49, 66, 84, 94, 100, 106, 108, 108, 103, 104, 123, 127, 120, 106, 122, 144, 156, 164, 157, 149, 97, 41, 38, 17, 8, 0, 
    90, 57, 69, 75, 92, 114, 108, 103, 107, 113, 118, 122, 126, 130, 127, 116, 118, 126, 109, 75, 76, 105, 125, 146, 147, 144, 113, 74, 90, 97, 58, 0, 
    91, 69, 86, 87, 82, 96, 115, 113, 110, 116, 121, 122, 118, 114, 108, 99, 92, 112, 111, 80, 77, 107, 122, 130, 136, 132, 122, 118, 146, 156, 129, 0, 
    88, 59, 58, 44, 47, 65, 95, 114, 113, 111, 105, 99, 94, 92, 92, 98, 100, 117, 130, 116, 112, 129, 132, 127, 127, 125, 125, 124, 124, 132, 146, 8, 
    65, 15, 29, 50, 72, 87, 87, 94, 96, 85, 85, 90, 100, 107, 114, 123, 126, 136, 138, 129, 124, 129, 134, 131, 128, 126, 111, 95, 83, 80, 112, 30, 
    76, 30, 48, 74, 87, 90, 84, 74, 86, 96, 104, 111, 116, 110, 113, 115, 105, 128, 139, 127, 126, 128, 132, 127, 108, 91, 75, 59, 48, 40, 62, 14, 
    115, 70, 67, 71, 74, 79, 87, 85, 95, 112, 125, 120, 109, 80, 55, 49, 40, 75, 123, 131, 126, 119, 107, 87, 71, 59, 47, 38, 36, 34, 20, 0, 
    105, 84, 79, 77, 79, 72, 78, 79, 75, 76, 96, 110, 103, 67, 25, 18, 27, 58, 101, 107, 94, 80, 67, 56, 50, 39, 26, 22, 26, 16, 0, 0, 
    80, 81, 79, 77, 74, 47, 29, 30, 29, 29, 54, 95, 110, 92, 65, 54, 52, 57, 65, 63, 57, 57, 49, 33, 18, 14, 10, 7, 2, 0, 0, 0, 
    71, 70, 69, 71, 73, 46, 15, 19, 34, 46, 69, 92, 93, 76, 59, 52, 46, 45, 50, 51, 45, 35, 24, 20, 12, 4, 2, 0, 0, 0, 0, 0, 
    72, 74, 81, 82, 85, 71, 51, 49, 55, 54, 55, 53, 45, 37, 35, 38, 40, 43, 45, 35, 23, 14, 11, 18, 19, 4, 0, 0, 0, 0, 0, 0, 
    63, 60, 67, 62, 56, 48, 40, 35, 31, 26, 24, 26, 30, 34, 39, 37, 30, 21, 11, 10, 11, 11, 8, 9, 9, 0, 0, 0, 0, 0, 0, 0, 
    27, 13, 15, 15, 13, 9, 9, 14, 19, 22, 26, 27, 24, 20, 19, 14, 12, 16, 7, 3, 7, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 1, 8, 13, 11, 8, 7, 5, 4, 5, 4, 13, 37, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 6, 8, 4, 17, 43, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 6, 7, 9, 7, 6, 1, 13, 40, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 6, 7, 10, 13, 14, 16, 19, 22, 22, 20, 16, 12, 4, 0, 0, 0, 29, 32, 4, 0, 1, 1, 1, 0, 0, 3, 6, 0, 0, 0, 0, 
    
    -- channel=47
    63, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 3, 0, 
    139, 62, 48, 66, 96, 95, 93, 100, 110, 113, 111, 118, 129, 129, 131, 126, 119, 132, 137, 139, 134, 133, 140, 139, 133, 129, 138, 136, 130, 138, 144, 47, 
    146, 73, 58, 72, 104, 106, 100, 105, 119, 120, 117, 121, 134, 136, 138, 133, 123, 134, 137, 137, 131, 143, 153, 147, 138, 132, 143, 142, 131, 142, 151, 52, 
    149, 76, 64, 78, 109, 114, 112, 109, 123, 127, 118, 122, 136, 137, 138, 140, 125, 135, 135, 114, 110, 144, 163, 150, 141, 134, 147, 146, 134, 143, 153, 53, 
    155, 79, 65, 83, 115, 118, 117, 113, 130, 132, 121, 124, 135, 133, 134, 146, 131, 137, 133, 102, 85, 123, 152, 150, 144, 134, 146, 147, 139, 145, 151, 52, 
    160, 88, 70, 86, 121, 122, 125, 118, 130, 133, 124, 125, 133, 127, 118, 140, 136, 142, 129, 79, 77, 129, 147, 147, 147, 132, 143, 147, 139, 148, 149, 54, 
    165, 95, 73, 88, 129, 128, 134, 129, 137, 137, 128, 130, 132, 122, 101, 118, 121, 124, 131, 89, 57, 100, 134, 154, 165, 143, 140, 146, 137, 149, 153, 56, 
    170, 102, 81, 94, 138, 135, 144, 148, 151, 145, 135, 137, 135, 131, 113, 95, 82, 77, 88, 87, 55, 58, 75, 101, 161, 169, 151, 146, 133, 151, 165, 65, 
    163, 115, 97, 98, 137, 139, 151, 161, 158, 156, 147, 147, 141, 135, 124, 101, 68, 56, 42, 29, 21, 22, 13, 14, 63, 120, 141, 140, 129, 149, 164, 73, 
    126, 101, 88, 79, 100, 108, 110, 125, 132, 135, 132, 133, 129, 122, 115, 93, 59, 45, 37, 28, 26, 31, 37, 50, 50, 69, 101, 95, 89, 106, 123, 61, 
    79, 60, 52, 51, 57, 47, 50, 66, 81, 82, 79, 83, 86, 80, 73, 58, 45, 39, 37, 30, 22, 38, 51, 46, 61, 73, 117, 88, 42, 52, 65, 25, 
    51, 33, 27, 31, 40, 27, 21, 41, 59, 48, 35, 45, 50, 43, 39, 36, 29, 30, 34, 27, 17, 41, 76, 69, 56, 34, 99, 129, 46, 37, 43, 9, 
    53, 28, 17, 26, 53, 41, 35, 44, 53, 55, 33, 26, 39, 40, 32, 28, 31, 33, 36, 34, 33, 57, 98, 116, 108, 62, 63, 130, 67, 31, 46, 6, 
    56, 31, 30, 24, 35, 39, 36, 38, 55, 66, 58, 37, 35, 39, 30, 23, 22, 18, 23, 32, 43, 70, 100, 115, 128, 111, 65, 103, 89, 24, 39, 13, 
    61, 29, 29, 21, 26, 19, 24, 36, 40, 43, 49, 46, 37, 36, 35, 37, 38, 35, 34, 42, 57, 85, 108, 115, 117, 115, 76, 51, 82, 41, 24, 7, 
    70, 27, 30, 27, 37, 35, 27, 35, 48, 54, 55, 56, 56, 57, 52, 52, 66, 72, 66, 58, 71, 99, 117, 120, 114, 106, 80, 28, 43, 37, 12, 0, 
    82, 38, 51, 45, 48, 68, 68, 64, 67, 72, 71, 68, 66, 64, 63, 58, 64, 78, 75, 55, 56, 84, 94, 103, 106, 97, 86, 60, 61, 54, 22, 0, 
    90, 45, 47, 49, 53, 73, 83, 74, 68, 68, 67, 63, 60, 59, 58, 58, 57, 70, 73, 56, 47, 69, 80, 87, 92, 89, 89, 79, 86, 107, 94, 12, 
    76, 30, 43, 50, 47, 42, 58, 69, 64, 58, 60, 59, 56, 54, 52, 54, 51, 60, 80, 75, 68, 82, 90, 84, 83, 83, 81, 77, 85, 92, 104, 41, 
    69, 23, 37, 38, 37, 41, 44, 53, 57, 54, 50, 49, 52, 57, 60, 64, 67, 71, 83, 83, 79, 86, 94, 87, 78, 75, 72, 69, 63, 64, 86, 46, 
    78, 14, 19, 37, 49, 59, 55, 47, 53, 53, 49, 54, 59, 63, 63, 64, 65, 80, 94, 84, 79, 82, 84, 78, 66, 66, 57, 42, 40, 38, 36, 39, 
    87, 41, 36, 39, 43, 46, 50, 47, 49, 63, 68, 70, 63, 44, 31, 38, 38, 53, 87, 80, 71, 71, 67, 65, 53, 38, 29, 27, 29, 24, 17, 13, 
    81, 55, 42, 39, 42, 39, 39, 47, 47, 51, 66, 76, 63, 42, 16, 14, 17, 22, 52, 65, 61, 56, 48, 34, 27, 25, 19, 17, 17, 21, 15, 0, 
    59, 48, 45, 43, 42, 26, 15, 26, 30, 26, 37, 62, 66, 57, 35, 24, 25, 29, 43, 45, 39, 29, 19, 16, 20, 18, 10, 6, 10, 10, 5, 0, 
    55, 42, 43, 40, 42, 27, 5, 10, 17, 20, 25, 42, 54, 55, 50, 42, 36, 31, 31, 26, 18, 16, 17, 17, 9, 5, 5, 8, 4, 1, 2, 0, 
    59, 44, 45, 41, 43, 43, 27, 22, 24, 24, 33, 42, 43, 36, 28, 21, 19, 21, 24, 23, 19, 12, 3, 10, 17, 9, 4, 7, 4, 0, 3, 0, 
    48, 35, 43, 41, 40, 37, 33, 30, 29, 23, 18, 16, 17, 18, 19, 17, 13, 14, 20, 13, 6, 6, 8, 12, 14, 8, 3, 1, 0, 0, 1, 0, 
    30, 15, 21, 21, 17, 11, 9, 12, 14, 13, 12, 12, 13, 14, 15, 13, 11, 15, 5, 0, 3, 10, 10, 7, 6, 2, 1, 1, 1, 1, 0, 0, 
    19, 1, 1, 3, 3, 1, 0, 4, 9, 9, 9, 10, 9, 4, 3, 2, 7, 21, 17, 0, 3, 10, 7, 6, 4, 1, 1, 0, 4, 2, 0, 0, 
    20, 4, 2, 2, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 3, 6, 12, 27, 21, 0, 2, 7, 8, 7, 2, 0, 1, 3, 5, 0, 0, 0, 
    18, 3, 1, 1, 0, 0, 0, 0, 0, 0, 2, 4, 5, 3, 4, 7, 14, 29, 22, 0, 0, 8, 7, 5, 1, 0, 1, 6, 1, 0, 0, 0, 
    17, 8, 7, 7, 8, 9, 11, 13, 13, 12, 12, 10, 8, 4, 4, 6, 11, 28, 28, 5, 8, 11, 12, 9, 6, 4, 7, 7, 3, 0, 0, 0, 
    
    -- channel=48
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=49
    0, 31, 53, 59, 63, 52, 40, 36, 33, 34, 40, 41, 37, 36, 34, 35, 35, 34, 33, 34, 36, 37, 36, 36, 36, 39, 44, 47, 49, 52, 58, 40, 
    0, 37, 62, 69, 74, 68, 53, 39, 32, 37, 50, 53, 49, 47, 45, 43, 46, 47, 47, 47, 46, 47, 46, 46, 47, 47, 48, 54, 56, 53, 55, 40, 
    0, 48, 68, 71, 74, 71, 53, 12, 0, 15, 26, 35, 33, 30, 29, 30, 34, 34, 33, 35, 36, 36, 37, 30, 40, 54, 57, 57, 56, 55, 59, 43, 
    0, 54, 66, 68, 75, 71, 53, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 54, 60, 53, 52, 55, 61, 43, 
    0, 53, 64, 67, 74, 70, 48, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 50, 62, 58, 55, 57, 60, 42, 
    0, 50, 61, 67, 77, 68, 31, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 7, 13, 11, 10, 10, 9, 13, 20, 32, 50, 58, 57, 56, 61, 45, 
    0, 51, 61, 68, 78, 58, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 34, 58, 57, 55, 61, 45, 
    0, 55, 63, 68, 73, 51, 12, 0, 0, 0, 4, 5, 1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 10, 9, 7, 33, 56, 58, 59, 63, 46, 
    0, 58, 63, 65, 71, 59, 35, 24, 25, 24, 23, 20, 23, 26, 23, 21, 24, 28, 25, 20, 13, 14, 20, 30, 32, 42, 57, 61, 61, 63, 66, 48, 
    0, 62, 65, 65, 72, 66, 60, 58, 47, 42, 41, 39, 44, 44, 43, 41, 41, 44, 46, 43, 36, 37, 38, 42, 50, 61, 66, 64, 62, 64, 68, 48, 
    0, 62, 67, 68, 72, 65, 67, 70, 64, 59, 59, 59, 57, 59, 60, 59, 61, 62, 60, 58, 56, 54, 54, 55, 60, 62, 61, 59, 59, 62, 67, 48, 
    0, 57, 61, 58, 55, 44, 49, 63, 68, 69, 67, 65, 65, 65, 65, 66, 65, 65, 65, 65, 63, 61, 61, 64, 65, 63, 63, 63, 62, 63, 67, 47, 
    0, 53, 58, 57, 47, 18, 0, 7, 35, 57, 66, 66, 64, 64, 66, 67, 68, 67, 66, 66, 64, 63, 65, 65, 64, 63, 63, 62, 61, 61, 63, 46, 
    0, 53, 69, 77, 71, 45, 12, 0, 0, 0, 32, 55, 62, 63, 64, 66, 66, 64, 63, 61, 60, 59, 59, 60, 61, 61, 60, 60, 58, 59, 63, 46, 
    0, 53, 64, 68, 71, 68, 61, 31, 0, 0, 0, 16, 44, 58, 62, 63, 61, 59, 59, 58, 57, 56, 57, 60, 61, 61, 61, 60, 59, 61, 65, 48, 
    0, 55, 66, 68, 68, 61, 60, 58, 33, 0, 0, 0, 0, 18, 43, 55, 58, 59, 58, 57, 56, 56, 57, 59, 60, 61, 63, 63, 62, 63, 68, 52, 
    0, 57, 64, 63, 66, 62, 55, 55, 52, 20, 0, 0, 0, 0, 0, 10, 33, 48, 56, 57, 56, 58, 61, 61, 61, 62, 63, 63, 63, 64, 68, 53, 
    0, 54, 59, 57, 61, 58, 56, 55, 52, 27, 0, 0, 0, 0, 0, 0, 0, 0, 7, 26, 39, 51, 61, 64, 63, 63, 61, 61, 60, 60, 66, 52, 
    0, 51, 55, 52, 56, 55, 56, 54, 47, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 35, 43, 51, 57, 60, 60, 61, 66, 51, 
    0, 47, 55, 51, 54, 56, 58, 49, 38, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 34, 48, 57, 63, 52, 
    0, 41, 58, 55, 53, 57, 58, 53, 42, 19, 3, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 9, 15, 26, 43, 52, 48, 
    0, 40, 60, 58, 55, 56, 57, 63, 56, 40, 45, 49, 29, 13, 6, 4, 23, 45, 48, 28, 15, 29, 36, 24, 10, 14, 36, 45, 45, 47, 48, 45, 
    0, 36, 55, 51, 47, 46, 44, 42, 37, 39, 46, 51, 45, 39, 34, 32, 36, 43, 52, 48, 42, 43, 48, 50, 43, 42, 43, 44, 50, 53, 52, 49, 
    0, 0, 15, 11, 7, 6, 4, 1, 0, 0, 0, 0, 0, 3, 8, 17, 26, 28, 28, 28, 35, 35, 33, 35, 42, 47, 46, 44, 43, 43, 44, 43, 
    0, 0, 11, 12, 12, 14, 12, 11, 11, 9, 9, 10, 9, 9, 8, 10, 19, 24, 23, 24, 23, 22, 22, 23, 26, 28, 30, 30, 25, 21, 22, 14, 
    0, 0, 7, 6, 8, 8, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=50
    283, 80, 51, 31, 0, 12, 48, 54, 61, 63, 56, 48, 52, 49, 52, 58, 51, 55, 61, 60, 61, 56, 55, 57, 58, 63, 63, 55, 44, 42, 26, 0, 
    352, 147, 109, 96, 49, 39, 83, 99, 107, 111, 105, 96, 94, 91, 87, 105, 99, 91, 97, 97, 103, 99, 92, 99, 105, 119, 128, 120, 113, 118, 96, 0, 
    344, 136, 98, 95, 68, 52, 62, 93, 144, 147, 123, 118, 110, 110, 110, 123, 119, 111, 112, 111, 112, 109, 104, 119, 112, 104, 107, 107, 108, 115, 95, 0, 
    340, 134, 100, 101, 87, 78, 50, 55, 140, 164, 146, 157, 148, 141, 155, 163, 156, 149, 157, 154, 148, 150, 139, 169, 176, 119, 102, 112, 113, 117, 97, 0, 
    337, 130, 100, 99, 87, 83, 45, 43, 107, 95, 97, 120, 105, 108, 120, 126, 112, 99, 112, 108, 95, 109, 103, 129, 172, 124, 97, 108, 107, 109, 91, 0, 
    332, 132, 106, 98, 86, 84, 60, 95, 141, 88, 94, 112, 92, 107, 124, 127, 117, 102, 105, 101, 93, 104, 108, 118, 153, 146, 118, 112, 111, 117, 92, 0, 
    328, 123, 104, 98, 86, 72, 54, 114, 173, 122, 117, 132, 107, 110, 135, 145, 139, 135, 148, 124, 142, 148, 140, 128, 135, 186, 159, 112, 108, 117, 92, 0, 
    327, 111, 96, 98, 80, 50, 33, 81, 121, 108, 91, 99, 98, 83, 100, 104, 95, 95, 106, 84, 105, 123, 119, 104, 76, 146, 158, 116, 106, 109, 87, 0, 
    331, 96, 87, 97, 76, 56, 48, 56, 77, 95, 90, 91, 99, 98, 104, 100, 92, 85, 85, 78, 93, 112, 121, 121, 84, 95, 113, 104, 98, 101, 82, 0, 
    348, 88, 75, 93, 77, 82, 76, 47, 62, 92, 89, 96, 92, 96, 99, 93, 96, 95, 89, 84, 99, 105, 116, 139, 116, 90, 98, 102, 96, 100, 81, 0, 
    365, 99, 72, 92, 71, 85, 85, 50, 48, 70, 64, 66, 72, 73, 73, 67, 61, 61, 65, 67, 73, 82, 87, 106, 109, 95, 99, 102, 101, 105, 83, 0, 
    381, 116, 77, 94, 79, 109, 144, 106, 67, 68, 72, 77, 79, 81, 82, 76, 72, 71, 76, 80, 85, 90, 91, 92, 95, 96, 96, 97, 98, 103, 83, 0, 
    389, 127, 65, 60, 63, 99, 186, 215, 167, 124, 93, 85, 88, 92, 91, 87, 82, 81, 83, 84, 90, 95, 91, 89, 95, 99, 100, 104, 104, 107, 86, 0, 
    395, 135, 61, 24, 9, 10, 54, 156, 223, 225, 182, 127, 101, 96, 94, 91, 89, 92, 91, 87, 93, 101, 101, 97, 99, 101, 102, 103, 103, 108, 85, 0, 
    400, 144, 86, 71, 52, 24, 0, 0, 83, 181, 227, 211, 163, 121, 99, 94, 96, 101, 101, 94, 97, 104, 101, 96, 96, 96, 95, 96, 96, 102, 79, 0, 
    401, 150, 99, 96, 90, 91, 59, 0, 0, 50, 169, 222, 238, 214, 160, 117, 98, 95, 97, 97, 99, 104, 102, 98, 98, 96, 91, 92, 92, 95, 74, 0, 
    402, 152, 107, 108, 98, 106, 107, 67, 0, 0, 94, 163, 196, 242, 250, 215, 166, 129, 105, 95, 96, 103, 100, 95, 97, 97, 94, 96, 95, 96, 74, 0, 
    406, 155, 116, 124, 110, 113, 113, 104, 0, 0, 46, 133, 136, 167, 201, 232, 241, 226, 197, 155, 131, 128, 108, 89, 90, 92, 94, 99, 99, 99, 77, 0, 
    411, 157, 117, 131, 118, 118, 115, 109, 16, 0, 50, 145, 140, 145, 142, 147, 169, 197, 217, 214, 213, 231, 208, 161, 136, 117, 102, 96, 94, 96, 73, 0, 
    414, 162, 115, 128, 121, 119, 116, 90, 14, 0, 33, 132, 151, 149, 143, 133, 121, 122, 123, 122, 148, 210, 245, 238, 238, 224, 191, 160, 130, 108, 75, 0, 
    415, 165, 112, 120, 120, 120, 111, 57, 0, 1, 0, 13, 103, 134, 154, 167, 110, 59, 39, 69, 89, 88, 118, 154, 215, 226, 176, 163, 158, 136, 93, 0, 
    410, 164, 108, 113, 115, 117, 107, 52, 7, 36, 0, 0, 0, 40, 76, 151, 130, 42, 0, 5, 85, 46, 0, 20, 109, 165, 121, 96, 108, 115, 93, 0, 
    407, 170, 112, 117, 122, 125, 124, 111, 101, 108, 85, 20, 11, 46, 69, 120, 135, 100, 48, 38, 86, 87, 55, 38, 73, 112, 114, 109, 107, 108, 93, 0, 
    391, 210, 164, 160, 167, 170, 174, 175, 174, 179, 172, 152, 148, 150, 155, 154, 133, 120, 118, 113, 110, 114, 116, 110, 98, 90, 90, 94, 100, 109, 103, 0, 
    295, 143, 119, 104, 105, 103, 104, 102, 101, 107, 105, 99, 100, 101, 108, 119, 101, 79, 85, 91, 89, 88, 95, 99, 94, 85, 79, 72, 77, 93, 105, 0, 
    271, 118, 99, 89, 83, 81, 90, 96, 102, 107, 107, 106, 103, 104, 105, 111, 114, 100, 104, 116, 116, 113, 116, 124, 125, 125, 123, 114, 107, 119, 138, 8, 
    267, 146, 146, 136, 130, 121, 119, 131, 138, 137, 137, 140, 136, 135, 135, 134, 136, 128, 123, 130, 135, 134, 132, 130, 130, 133, 133, 128, 126, 142, 154, 19, 
    221, 119, 133, 127, 128, 122, 120, 132, 136, 131, 130, 128, 126, 128, 130, 133, 135, 131, 124, 124, 129, 133, 133, 129, 126, 126, 125, 130, 139, 151, 152, 15, 
    212, 113, 125, 122, 129, 122, 123, 134, 133, 128, 129, 129, 125, 124, 131, 139, 139, 132, 128, 130, 130, 131, 132, 131, 127, 126, 132, 142, 151, 154, 146, 34, 
    206, 110, 122, 115, 121, 118, 119, 126, 124, 124, 128, 120, 110, 107, 115, 128, 123, 114, 112, 115, 115, 120, 130, 131, 138, 146, 151, 148, 140, 130, 139, 60, 
    206, 112, 131, 128, 128, 121, 119, 123, 126, 130, 147, 148, 127, 123, 131, 146, 145, 135, 132, 128, 116, 116, 134, 139, 152, 167, 166, 145, 118, 127, 151, 64, 
    216, 150, 163, 164, 166, 161, 156, 156, 161, 163, 173, 181, 172, 170, 171, 177, 182, 179, 177, 174, 164, 156, 167, 181, 215, 232, 196, 160, 158, 165, 175, 116, 
    
    -- channel=51
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=52
    0, 103, 120, 146, 176, 150, 120, 117, 114, 115, 127, 137, 139, 136, 135, 129, 134, 131, 123, 126, 127, 131, 135, 134, 133, 135, 139, 156, 170, 170, 196, 372, 
    0, 0, 0, 0, 62, 56, 24, 17, 5, 0, 5, 28, 34, 45, 41, 27, 37, 39, 33, 32, 27, 35, 38, 32, 27, 10, 2, 13, 21, 14, 68, 441, 
    0, 0, 0, 0, 32, 58, 44, 45, 0, 0, 0, 2, 9, 25, 18, 0, 10, 26, 22, 21, 15, 23, 28, 20, 9, 2, 0, 8, 15, 5, 61, 442, 
    0, 0, 0, 0, 0, 17, 89, 119, 39, 10, 7, 0, 1, 18, 10, 0, 2, 6, 0, 0, 0, 2, 17, 0, 0, 0, 4, 10, 12, 6, 61, 445, 
    0, 0, 0, 0, 0, 0, 128, 170, 111, 121, 123, 103, 121, 134, 106, 94, 117, 129, 114, 117, 124, 106, 137, 52, 0, 19, 15, 13, 17, 11, 66, 452, 
    0, 0, 0, 0, 0, 0, 95, 87, 57, 121, 115, 102, 117, 113, 96, 83, 99, 109, 91, 111, 111, 85, 110, 37, 0, 0, 0, 2, 8, 2, 60, 450, 
    0, 0, 0, 0, 0, 17, 119, 63, 46, 69, 49, 42, 80, 86, 71, 35, 34, 20, 13, 38, 27, 19, 20, 21, 3, 0, 0, 0, 0, 0, 51, 444, 
    0, 0, 0, 0, 0, 75, 182, 150, 120, 99, 100, 86, 123, 125, 114, 100, 114, 97, 96, 134, 105, 103, 76, 122, 111, 4, 0, 0, 0, 0, 47, 435, 
    0, 0, 0, 0, 0, 67, 118, 125, 98, 57, 68, 42, 52, 50, 44, 55, 73, 76, 74, 103, 77, 63, 30, 64, 93, 37, 2, 1, 4, 0, 45, 427, 
    0, 0, 0, 0, 0, 0, 12, 52, 38, 4, 2, 0, 0, 0, 0, 0, 1, 1, 4, 19, 11, 3, 0, 0, 0, 21, 1, 0, 0, 0, 44, 424, 
    0, 8, 0, 0, 0, 0, 0, 57, 51, 33, 39, 35, 38, 30, 31, 40, 42, 45, 45, 47, 36, 35, 15, 0, 0, 4, 1, 0, 0, 0, 46, 426, 
    0, 0, 0, 0, 0, 0, 0, 0, 36, 30, 33, 25, 19, 17, 21, 32, 41, 39, 27, 23, 18, 15, 12, 0, 0, 0, 6, 9, 10, 0, 52, 435, 
    0, 0, 17, 7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 16, 18, 17, 14, 8, 3, 7, 12, 4, 0, 0, 0, 0, 0, 47, 432, 
    0, 0, 62, 103, 131, 114, 0, 0, 0, 0, 0, 0, 0, 0, 5, 11, 16, 15, 18, 18, 7, 0, 0, 2, 0, 0, 0, 0, 0, 0, 46, 428, 
    0, 0, 41, 75, 106, 171, 201, 116, 0, 0, 0, 0, 0, 0, 6, 13, 11, 7, 10, 18, 13, 2, 3, 7, 5, 3, 5, 4, 1, 0, 47, 421, 
    0, 0, 3, 11, 30, 82, 176, 237, 189, 20, 0, 0, 0, 0, 0, 0, 16, 16, 16, 20, 15, 7, 9, 10, 5, 5, 9, 9, 5, 0, 47, 418, 
    0, 0, 2, 10, 16, 17, 47, 162, 270, 182, 0, 0, 0, 0, 0, 0, 0, 0, 7, 19, 14, 2, 3, 8, 2, 2, 5, 3, 2, 0, 45, 419, 
    0, 0, 0, 1, 15, 15, 15, 64, 239, 269, 68, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 13, 10, 6, 0, 0, 0, 41, 418, 
    0, 0, 3, 2, 16, 16, 25, 30, 186, 270, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 12, 12, 1, 49, 423, 
    0, 0, 9, 6, 14, 12, 18, 27, 175, 240, 75, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 426, 
    0, 0, 8, 8, 9, 8, 10, 80, 205, 243, 187, 100, 1, 0, 0, 0, 61, 122, 123, 86, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 418, 
    0, 0, 10, 11, 12, 10, 25, 145, 223, 209, 260, 277, 169, 112, 67, 15, 72, 166, 231, 172, 109, 140, 165, 141, 18, 0, 10, 12, 0, 0, 37, 413, 
    0, 0, 0, 0, 0, 0, 0, 55, 72, 32, 94, 207, 163, 116, 56, 0, 0, 47, 148, 99, 22, 60, 121, 117, 12, 0, 0, 0, 0, 0, 8, 382, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 319, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 246, 
    0, 0, 0, 1, 9, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 173, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 175, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 1, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 170, 
    0, 34, 0, 0, 0, 0, 1, 0, 0, 6, 4, 0, 0, 0, 0, 0, 0, 0, 4, 3, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 132, 
    0, 40, 0, 4, 0, 5, 2, 0, 3, 9, 9, 10, 24, 27, 21, 11, 19, 32, 31, 25, 20, 12, 1, 1, 0, 0, 0, 0, 0, 0, 0, 131, 
    0, 40, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 3, 13, 6, 0, 0, 10, 12, 12, 22, 17, 2, 3, 0, 0, 0, 0, 0, 0, 0, 121, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 
    
    -- channel=53
    171, 151, 152, 151, 128, 118, 128, 133, 136, 142, 145, 142, 141, 138, 136, 141, 138, 137, 140, 141, 145, 144, 141, 142, 145, 153, 164, 164, 161, 165, 145, 0, 
    145, 46, 34, 31, 11, 2, 7, 10, 20, 28, 24, 17, 18, 13, 11, 18, 20, 19, 18, 18, 19, 16, 14, 14, 19, 31, 38, 36, 34, 38, 13, 0, 
    145, 41, 26, 26, 16, 16, 6, 0, 35, 53, 43, 38, 34, 31, 35, 48, 44, 39, 47, 45, 43, 40, 32, 46, 61, 49, 39, 31, 25, 29, 5, 0, 
    145, 41, 27, 27, 19, 10, 0, 0, 10, 3, 0, 5, 0, 0, 0, 9, 8, 3, 9, 9, 4, 8, 0, 23, 59, 43, 25, 25, 24, 29, 7, 0, 
    143, 39, 24, 24, 16, 9, 0, 0, 42, 13, 0, 7, 0, 0, 8, 17, 9, 0, 4, 0, 0, 3, 0, 19, 46, 29, 22, 26, 26, 31, 6, 0, 
    140, 36, 25, 25, 17, 0, 0, 13, 61, 30, 38, 52, 34, 33, 47, 61, 57, 57, 65, 48, 54, 60, 50, 61, 66, 55, 41, 26, 25, 31, 7, 0, 
    142, 35, 24, 25, 15, 0, 0, 0, 27, 10, 15, 23, 7, 1, 15, 23, 15, 15, 16, 3, 11, 19, 22, 8, 0, 34, 42, 25, 22, 26, 2, 0, 
    146, 33, 23, 26, 12, 0, 0, 12, 25, 13, 9, 13, 6, 13, 23, 20, 11, 8, 2, 0, 0, 5, 16, 10, 7, 37, 36, 18, 16, 23, 0, 0, 
    153, 30, 20, 26, 12, 5, 19, 31, 35, 32, 26, 32, 26, 26, 31, 35, 42, 41, 32, 24, 37, 40, 49, 52, 47, 64, 50, 25, 21, 26, 2, 0, 
    161, 32, 19, 25, 16, 17, 18, 3, 1, 11, 6, 6, 10, 9, 13, 13, 12, 9, 7, 4, 8, 15, 19, 33, 36, 38, 33, 24, 23, 27, 2, 0, 
    168, 33, 23, 31, 15, 14, 18, 8, 12, 22, 20, 24, 25, 32, 33, 30, 27, 20, 18, 20, 26, 29, 34, 37, 27, 19, 18, 18, 20, 26, 4, 0, 
    170, 36, 15, 10, 0, 0, 33, 41, 37, 39, 37, 42, 46, 45, 44, 41, 38, 38, 40, 39, 40, 41, 39, 39, 32, 23, 23, 24, 25, 29, 7, 0, 
    170, 35, 0, 0, 0, 0, 0, 13, 37, 43, 33, 24, 24, 27, 28, 25, 23, 24, 24, 21, 22, 26, 27, 24, 23, 23, 24, 26, 26, 31, 6, 0, 
    173, 40, 13, 7, 0, 0, 0, 0, 0, 5, 32, 37, 31, 28, 27, 25, 25, 26, 25, 22, 23, 26, 25, 23, 23, 22, 21, 19, 18, 22, 0, 0, 
    174, 44, 24, 33, 46, 46, 26, 0, 0, 0, 0, 21, 42, 41, 31, 25, 23, 22, 21, 18, 18, 21, 21, 17, 17, 18, 17, 15, 17, 22, 0, 0, 
    176, 45, 25, 28, 24, 27, 37, 32, 0, 0, 0, 0, 9, 35, 42, 33, 23, 18, 15, 16, 20, 24, 23, 23, 25, 25, 23, 22, 22, 25, 2, 0, 
    179, 47, 27, 33, 28, 27, 25, 16, 0, 0, 0, 0, 0, 0, 0, 21, 34, 34, 29, 21, 19, 24, 25, 21, 22, 21, 20, 21, 22, 26, 4, 0, 
    180, 46, 25, 33, 27, 27, 24, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 21, 23, 35, 32, 24, 22, 20, 19, 20, 20, 24, 3, 0, 
    180, 46, 23, 29, 25, 25, 25, 20, 0, 0, 0, 0, 0, 4, 1, 0, 0, 0, 0, 0, 0, 3, 27, 31, 33, 33, 28, 23, 21, 24, 3, 0, 
    179, 46, 21, 28, 27, 26, 25, 0, 0, 0, 0, 0, 0, 0, 0, 5, 2, 0, 0, 0, 0, 0, 0, 0, 0, 9, 22, 33, 36, 33, 9, 0, 
    175, 46, 19, 25, 25, 25, 19, 0, 0, 0, 0, 0, 0, 0, 6, 44, 47, 16, 0, 0, 20, 2, 0, 0, 0, 2, 0, 0, 10, 23, 8, 0, 
    172, 45, 19, 26, 26, 25, 20, 0, 1, 38, 51, 29, 24, 22, 37, 76, 89, 70, 26, 25, 56, 65, 44, 25, 53, 74, 63, 48, 31, 22, 2, 0, 
    164, 43, 18, 19, 19, 17, 14, 13, 30, 61, 57, 43, 69, 89, 95, 102, 72, 40, 34, 60, 78, 65, 64, 78, 88, 75, 42, 31, 34, 31, 6, 0, 
    103, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 15, 19, 0, 0, 0, 0, 4, 0, 0, 0, 9, 2, 0, 0, 0, 0, 0, 0, 
    77, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    83, 9, 8, 5, 6, 4, 4, 6, 9, 9, 8, 7, 8, 10, 10, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 41, 20, 0, 
    34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 36, 38, 17, 0, 0, 
    33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 6, 5, 0, 0, 0, 0, 0, 0, 0, 0, 22, 42, 31, 1, 0, 0, 0, 
    34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 14, 10, 5, 4, 8, 9, 8, 9, 9, 0, 0, 0, 2, 25, 39, 24, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=54
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=55
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=56
    73, 195, 211, 229, 239, 211, 192, 192, 192, 195, 199, 205, 203, 205, 199, 195, 200, 197, 197, 199, 199, 205, 205, 203, 201, 199, 207, 221, 229, 233, 237, 267, 
    15, 197, 223, 238, 260, 240, 206, 199, 194, 198, 207, 217, 217, 220, 216, 207, 214, 215, 212, 212, 214, 219, 218, 214, 213, 213, 225, 235, 240, 244, 250, 314, 
    21, 203, 234, 247, 266, 259, 221, 181, 149, 171, 203, 208, 213, 208, 204, 197, 206, 212, 211, 214, 214, 216, 214, 209, 225, 235, 237, 241, 247, 249, 253, 319, 
    25, 204, 234, 247, 259, 254, 219, 151, 109, 123, 133, 128, 136, 134, 129, 130, 138, 141, 142, 150, 149, 149, 155, 146, 185, 233, 244, 241, 244, 245, 249, 318, 
    26, 204, 233, 247, 255, 245, 218, 168, 132, 120, 114, 109, 119, 119, 108, 109, 120, 131, 127, 139, 139, 135, 144, 139, 170, 233, 251, 246, 248, 251, 253, 320, 
    25, 200, 230, 246, 254, 240, 200, 153, 142, 157, 151, 146, 147, 128, 119, 131, 158, 166, 170, 178, 172, 174, 175, 178, 172, 207, 244, 249, 246, 250, 252, 319, 
    29, 202, 227, 244, 250, 227, 154, 100, 105, 142, 144, 133, 139, 124, 109, 118, 134, 142, 147, 147, 138, 145, 145, 164, 146, 154, 214, 247, 251, 249, 249, 316, 
    33, 209, 228, 241, 248, 219, 158, 127, 110, 138, 147, 141, 154, 150, 134, 133, 137, 144, 137, 142, 126, 129, 145, 158, 159, 155, 200, 240, 247, 247, 249, 314, 
    38, 222, 231, 239, 247, 234, 218, 202, 176, 177, 180, 183, 181, 185, 178, 175, 181, 192, 189, 182, 169, 167, 179, 180, 211, 209, 220, 245, 252, 252, 253, 313, 
    37, 235, 241, 241, 249, 249, 247, 237, 215, 202, 202, 198, 196, 202, 200, 202, 206, 211, 207, 203, 196, 193, 201, 202, 230, 243, 247, 250, 253, 254, 253, 313, 
    33, 244, 251, 248, 261, 250, 244, 253, 243, 227, 228, 223, 226, 226, 227, 230, 229, 231, 233, 234, 226, 223, 226, 224, 233, 249, 250, 246, 248, 251, 253, 315, 
    29, 241, 264, 250, 245, 216, 204, 241, 262, 253, 251, 248, 243, 244, 246, 250, 253, 252, 250, 248, 245, 241, 244, 241, 242, 252, 251, 250, 252, 254, 255, 319, 
    24, 237, 267, 240, 214, 182, 147, 158, 196, 227, 249, 253, 250, 249, 251, 256, 257, 256, 257, 255, 252, 249, 250, 253, 253, 252, 253, 253, 252, 252, 252, 314, 
    21, 237, 265, 257, 239, 216, 156, 104, 113, 145, 186, 222, 240, 249, 254, 257, 258, 258, 259, 257, 250, 246, 250, 252, 250, 248, 248, 246, 246, 247, 248, 309, 
    19, 237, 271, 277, 270, 257, 231, 174, 114, 86, 107, 155, 202, 237, 254, 257, 255, 252, 250, 251, 245, 241, 244, 249, 248, 249, 249, 247, 246, 248, 250, 308, 
    19, 235, 263, 263, 265, 268, 273, 266, 212, 117, 65, 84, 125, 168, 212, 242, 253, 252, 249, 248, 245, 243, 246, 248, 249, 251, 252, 250, 251, 252, 253, 310, 
    20, 234, 262, 263, 267, 260, 259, 273, 282, 189, 77, 53, 63, 88, 127, 168, 203, 227, 241, 249, 248, 243, 246, 249, 249, 250, 252, 251, 253, 254, 255, 314, 
    18, 233, 257, 257, 263, 259, 255, 253, 293, 244, 101, 59, 59, 49, 60, 85, 114, 143, 172, 200, 211, 219, 240, 251, 251, 251, 252, 248, 249, 253, 252, 311, 
    14, 229, 253, 249, 256, 257, 256, 255, 285, 246, 104, 43, 50, 50, 52, 51, 57, 69, 87, 108, 117, 126, 159, 199, 221, 236, 248, 250, 250, 252, 251, 311, 
    11, 229, 253, 245, 252, 256, 254, 266, 255, 204, 103, 28, 28, 40, 48, 59, 64, 61, 60, 60, 55, 44, 68, 107, 125, 151, 181, 203, 224, 242, 249, 312, 
    8, 224, 252, 243, 249, 252, 255, 263, 225, 186, 150, 93, 44, 32, 24, 38, 94, 133, 135, 85, 65, 68, 60, 49, 36, 80, 146, 176, 198, 221, 239, 308, 
    7, 222, 251, 245, 249, 251, 254, 256, 252, 225, 227, 206, 127, 99, 93, 103, 165, 208, 208, 156, 140, 158, 154, 133, 108, 131, 179, 195, 203, 219, 235, 303, 
    7, 214, 242, 240, 241, 240, 239, 246, 253, 229, 234, 255, 224, 188, 182, 166, 188, 224, 240, 224, 188, 202, 221, 215, 194, 178, 200, 214, 210, 213, 225, 285, 
    0, 156, 180, 176, 173, 169, 163, 162, 159, 153, 161, 175, 172, 151, 146, 146, 161, 179, 189, 194, 176, 175, 186, 196, 191, 182, 185, 187, 187, 189, 193, 245, 
    0, 119, 134, 134, 135, 131, 129, 128, 124, 123, 123, 123, 121, 120, 123, 129, 146, 155, 148, 146, 151, 153, 146, 148, 157, 164, 165, 164, 153, 150, 144, 191, 
    9, 123, 123, 132, 134, 133, 126, 120, 117, 115, 113, 114, 112, 108, 106, 102, 110, 119, 112, 106, 105, 104, 101, 100, 101, 104, 106, 106, 97, 93, 83, 136, 
    0, 86, 81, 87, 90, 92, 85, 77, 77, 74, 71, 67, 64, 64, 64, 66, 65, 70, 67, 57, 54, 54, 56, 55, 55, 54, 53, 54, 52, 49, 70, 141, 
    0, 63, 49, 52, 54, 58, 55, 49, 50, 49, 48, 44, 45, 45, 44, 44, 46, 53, 52, 44, 40, 39, 40, 42, 41, 40, 42, 40, 46, 83, 117, 147, 
    0, 59, 41, 44, 43, 44, 43, 40, 41, 42, 40, 38, 39, 40, 39, 37, 43, 46, 46, 43, 41, 40, 40, 39, 42, 44, 47, 63, 103, 129, 101, 118, 
    0, 57, 42, 46, 45, 46, 45, 42, 43, 43, 40, 48, 57, 57, 51, 48, 56, 59, 58, 56, 57, 50, 44, 44, 41, 44, 75, 122, 128, 94, 66, 99, 
    0, 56, 39, 44, 42, 45, 46, 42, 41, 42, 40, 49, 55, 57, 54, 49, 53, 59, 59, 58, 59, 48, 41, 43, 50, 84, 121, 116, 88, 72, 52, 75, 
    0, 9, 0, 2, 1, 3, 4, 2, 1, 0, 0, 0, 9, 10, 8, 3, 4, 8, 9, 10, 13, 11, 4, 10, 23, 37, 43, 40, 36, 19, 0, 15, 
    
    -- channel=57
    209, 291, 317, 330, 322, 293, 273, 268, 267, 271, 276, 275, 272, 268, 264, 264, 267, 266, 264, 264, 267, 270, 269, 267, 269, 278, 294, 306, 312, 317, 300, 247, 
    160, 159, 173, 177, 179, 168, 147, 125, 120, 132, 142, 146, 141, 140, 137, 137, 142, 146, 145, 142, 141, 140, 137, 134, 135, 139, 143, 140, 133, 135, 112, 55, 
    176, 180, 191, 187, 182, 176, 123, 55, 28, 62, 89, 82, 82, 76, 76, 90, 89, 93, 99, 100, 105, 102, 87, 108, 136, 159, 162, 139, 131, 135, 113, 55, 
    181, 179, 185, 183, 179, 161, 92, 27, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 70, 127, 139, 125, 126, 131, 111, 53, 
    185, 176, 182, 188, 184, 156, 84, 43, 67, 56, 29, 32, 29, 21, 16, 34, 45, 51, 57, 64, 60, 60, 61, 75, 123, 144, 141, 139, 135, 139, 115, 54, 
    183, 170, 178, 189, 188, 137, 36, 0, 22, 41, 45, 69, 40, 18, 16, 37, 54, 70, 74, 76, 71, 69, 74, 72, 91, 97, 116, 139, 136, 140, 114, 52, 
    189, 176, 179, 188, 177, 106, 0, 0, 0, 0, 12, 29, 4, 0, 0, 3, 4, 0, 0, 0, 0, 0, 7, 12, 7, 30, 91, 128, 127, 133, 111, 50, 
    195, 182, 184, 188, 175, 123, 49, 52, 81, 76, 83, 81, 79, 78, 80, 78, 79, 79, 73, 52, 47, 58, 71, 85, 78, 104, 135, 138, 142, 146, 121, 55, 
    201, 187, 185, 187, 179, 152, 129, 128, 121, 117, 114, 112, 110, 105, 109, 108, 115, 124, 116, 97, 92, 100, 111, 119, 135, 175, 175, 153, 152, 158, 131, 61, 
    201, 189, 189, 190, 182, 172, 167, 151, 133, 136, 131, 129, 131, 135, 139, 134, 130, 129, 127, 121, 121, 125, 130, 136, 145, 159, 162, 153, 151, 158, 134, 65, 
    195, 181, 189, 196, 188, 177, 174, 178, 188, 195, 195, 195, 196, 201, 199, 196, 193, 190, 187, 189, 188, 183, 186, 185, 165, 149, 151, 147, 147, 156, 134, 67, 
    185, 164, 166, 158, 127, 107, 119, 157, 190, 199, 193, 194, 194, 190, 187, 183, 182, 184, 186, 184, 180, 176, 177, 179, 167, 154, 155, 154, 156, 162, 135, 67, 
    178, 153, 156, 135, 92, 54, 28, 34, 78, 132, 162, 168, 165, 163, 163, 163, 164, 164, 167, 165, 162, 162, 162, 161, 160, 157, 153, 151, 150, 153, 124, 58, 
    173, 153, 175, 191, 190, 172, 116, 29, 0, 14, 73, 124, 150, 159, 160, 159, 157, 156, 156, 153, 149, 147, 146, 147, 147, 147, 145, 140, 137, 142, 118, 53, 
    172, 151, 164, 182, 198, 211, 223, 188, 106, 38, 21, 53, 105, 142, 153, 150, 143, 139, 136, 136, 136, 139, 142, 146, 148, 150, 150, 147, 147, 154, 130, 63, 
    175, 152, 160, 163, 153, 146, 165, 202, 191, 124, 61, 20, 11, 42, 90, 124, 138, 139, 135, 135, 140, 143, 146, 149, 152, 155, 157, 157, 159, 166, 142, 72, 
    177, 151, 151, 155, 152, 143, 127, 132, 153, 136, 92, 54, 10, 0, 0, 15, 65, 105, 130, 138, 140, 143, 147, 149, 150, 151, 152, 153, 156, 164, 143, 76, 
    174, 141, 134, 135, 134, 131, 126, 117, 113, 108, 90, 71, 58, 37, 0, 0, 0, 0, 13, 55, 89, 119, 144, 154, 154, 151, 149, 147, 147, 156, 138, 72, 
    168, 133, 124, 123, 122, 123, 126, 120, 92, 49, 38, 40, 40, 54, 60, 45, 9, 0, 0, 0, 0, 0, 26, 65, 98, 125, 144, 151, 153, 159, 139, 71, 
    161, 127, 121, 120, 121, 126, 126, 102, 52, 16, 32, 38, 34, 46, 50, 58, 68, 65, 53, 26, 0, 0, 0, 0, 0, 0, 30, 73, 112, 142, 135, 73, 
    153, 123, 122, 121, 121, 127, 122, 98, 57, 80, 155, 146, 88, 57, 52, 88, 143, 165, 141, 119, 135, 139, 86, 18, 2, 39, 71, 77, 89, 114, 114, 65, 
    152, 129, 131, 127, 128, 129, 127, 129, 147, 200, 256, 275, 250, 221, 203, 204, 222, 238, 233, 211, 223, 252, 250, 227, 211, 210, 201, 184, 163, 146, 124, 67, 
    143, 122, 121, 111, 105, 102, 95, 91, 114, 145, 152, 175, 225, 251, 246, 224, 171, 135, 155, 201, 221, 196, 203, 232, 244, 209, 151, 133, 137, 134, 119, 66, 
    72, 13, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 39, 50, 65, 63, 51, 53, 79, 99, 89, 84, 98, 120, 121, 109, 101, 93, 92, 82, 39, 
    104, 57, 55, 53, 56, 61, 64, 66, 67, 68, 69, 70, 75, 80, 81, 83, 92, 100, 100, 95, 92, 93, 92, 89, 90, 97, 109, 110, 96, 82, 57, 16, 
    113, 103, 113, 112, 118, 116, 109, 101, 96, 94, 90, 91, 97, 100, 102, 93, 79, 69, 63, 58, 54, 53, 51, 48, 44, 41, 41, 37, 29, 34, 33, 16, 
    64, 23, 27, 26, 29, 34, 31, 24, 21, 17, 12, 16, 20, 24, 27, 28, 27, 24, 26, 24, 20, 23, 30, 34, 32, 29, 26, 22, 27, 66, 98, 79, 
    69, 36, 40, 33, 33, 35, 35, 35, 35, 31, 36, 45, 49, 51, 49, 49, 49, 48, 51, 54, 55, 56, 57, 58, 59, 60, 63, 76, 110, 154, 155, 94, 
    65, 51, 63, 56, 59, 60, 56, 56, 53, 48, 52, 62, 69, 66, 60, 57, 59, 58, 55, 59, 65, 67, 65, 60, 60, 70, 99, 137, 162, 150, 85, 20, 
    67, 52, 68, 66, 69, 68, 67, 67, 61, 60, 73, 89, 94, 88, 81, 80, 83, 84, 85, 86, 81, 71, 64, 59, 70, 105, 152, 167, 129, 65, 9, 7, 
    64, 46, 58, 57, 64, 66, 64, 61, 56, 53, 56, 67, 70, 64, 59, 56, 55, 58, 65, 68, 67, 58, 54, 68, 101, 135, 142, 106, 44, 13, 21, 36, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=58
    28, 58, 71, 84, 80, 56, 50, 49, 47, 52, 55, 55, 50, 53, 47, 49, 51, 45, 48, 49, 51, 54, 50, 50, 49, 50, 57, 61, 64, 67, 64, 67, 
    88, 113, 136, 150, 148, 122, 99, 88, 85, 101, 110, 113, 104, 104, 98, 95, 102, 99, 99, 100, 100, 103, 101, 99, 98, 99, 107, 114, 117, 119, 113, 103, 
    100, 130, 155, 165, 161, 136, 100, 53, 38, 73, 86, 89, 88, 80, 78, 80, 88, 83, 87, 88, 91, 93, 86, 90, 112, 124, 134, 134, 131, 128, 121, 108, 
    103, 128, 151, 159, 162, 145, 105, 40, 9, 31, 34, 37, 41, 33, 28, 32, 37, 35, 36, 43, 45, 46, 44, 42, 93, 129, 135, 128, 129, 126, 121, 109, 
    108, 131, 152, 158, 164, 149, 108, 33, 18, 33, 19, 25, 31, 13, 14, 24, 42, 40, 37, 51, 46, 43, 49, 40, 87, 130, 134, 130, 130, 132, 125, 110, 
    107, 124, 147, 156, 161, 143, 85, 14, 33, 46, 23, 30, 26, 6, 5, 16, 37, 40, 46, 49, 42, 45, 47, 45, 71, 112, 133, 136, 135, 135, 127, 111, 
    109, 124, 146, 154, 153, 126, 47, 0, 8, 35, 30, 35, 39, 13, 13, 22, 38, 36, 41, 44, 22, 40, 44, 57, 46, 69, 118, 133, 133, 134, 130, 113, 
    114, 126, 145, 153, 153, 130, 57, 15, 26, 48, 59, 55, 59, 42, 44, 49, 58, 56, 61, 53, 30, 50, 47, 69, 55, 60, 111, 135, 140, 138, 133, 114, 
    122, 131, 144, 153, 156, 137, 94, 75, 66, 79, 81, 80, 83, 75, 78, 76, 80, 83, 82, 71, 56, 68, 69, 93, 91, 97, 128, 138, 141, 141, 135, 115, 
    127, 140, 143, 152, 154, 145, 138, 131, 104, 107, 105, 101, 107, 103, 106, 106, 107, 111, 111, 106, 92, 99, 99, 111, 127, 130, 139, 139, 141, 143, 137, 115, 
    128, 141, 142, 151, 154, 147, 152, 149, 127, 125, 124, 122, 120, 122, 126, 126, 129, 129, 124, 121, 116, 115, 118, 128, 143, 142, 142, 140, 141, 143, 135, 115, 
    125, 138, 142, 139, 137, 121, 129, 148, 137, 137, 133, 132, 135, 135, 138, 139, 137, 135, 134, 133, 128, 129, 131, 137, 145, 142, 140, 137, 138, 139, 132, 115, 
    122, 134, 145, 130, 114, 85, 72, 103, 131, 146, 150, 146, 145, 147, 149, 150, 149, 146, 145, 143, 139, 140, 142, 141, 140, 140, 139, 137, 138, 139, 132, 114, 
    119, 133, 148, 136, 112, 79, 47, 38, 56, 92, 127, 145, 145, 145, 146, 147, 145, 143, 142, 139, 137, 138, 140, 140, 140, 141, 140, 140, 139, 140, 132, 112, 
    118, 135, 146, 136, 125, 106, 77, 45, 19, 34, 70, 105, 133, 144, 145, 143, 140, 138, 137, 136, 131, 132, 137, 138, 138, 140, 139, 138, 139, 141, 134, 113, 
    119, 136, 147, 148, 141, 124, 98, 82, 46, 5, 25, 54, 77, 110, 135, 141, 140, 136, 134, 132, 130, 131, 134, 136, 138, 140, 141, 140, 142, 144, 138, 117, 
    120, 137, 143, 144, 143, 136, 123, 109, 87, 18, 0, 19, 28, 45, 72, 102, 122, 130, 133, 132, 129, 131, 137, 137, 138, 141, 141, 140, 143, 145, 140, 120, 
    120, 133, 135, 135, 137, 133, 129, 122, 114, 34, 0, 0, 0, 4, 20, 33, 54, 77, 99, 118, 122, 132, 142, 139, 138, 139, 138, 137, 140, 143, 138, 121, 
    116, 129, 128, 128, 130, 130, 128, 124, 122, 35, 0, 0, 0, 0, 0, 1, 8, 15, 30, 49, 63, 85, 115, 125, 128, 133, 137, 135, 137, 140, 136, 118, 
    112, 126, 126, 124, 128, 131, 129, 128, 100, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 5, 16, 41, 52, 63, 88, 106, 120, 133, 139, 136, 121, 
    108, 125, 129, 124, 127, 132, 132, 129, 79, 23, 3, 0, 0, 0, 0, 0, 12, 5, 0, 0, 0, 2, 0, 0, 4, 51, 76, 82, 106, 125, 131, 120, 
    105, 126, 133, 129, 129, 131, 132, 128, 85, 52, 57, 41, 8, 8, 0, 10, 48, 64, 58, 12, 16, 34, 35, 13, 6, 46, 81, 98, 108, 116, 123, 116, 
    99, 121, 133, 127, 123, 123, 122, 114, 96, 96, 106, 88, 62, 61, 57, 75, 101, 105, 98, 75, 81, 86, 83, 77, 76, 99, 111, 114, 122, 125, 127, 114, 
    67, 85, 107, 99, 94, 90, 88, 87, 86, 85, 90, 79, 70, 78, 82, 100, 117, 113, 108, 102, 112, 114, 112, 112, 120, 129, 129, 129, 126, 122, 119, 103, 
    60, 56, 74, 72, 68, 64, 63, 61, 58, 56, 57, 56, 57, 60, 65, 72, 89, 92, 93, 97, 96, 95, 96, 102, 105, 106, 108, 110, 102, 99, 88, 74, 
    35, 27, 53, 50, 50, 47, 41, 36, 31, 28, 28, 28, 31, 34, 42, 48, 55, 53, 47, 47, 48, 49, 48, 49, 52, 54, 56, 55, 48, 44, 37, 42, 
    15, 0, 23, 24, 26, 28, 23, 13, 10, 4, 0, 0, 2, 3, 4, 5, 6, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 20, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 12, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=59
    136, 296, 323, 336, 345, 329, 304, 303, 304, 303, 311, 321, 323, 320, 317, 310, 314, 316, 313, 314, 314, 320, 324, 321, 321, 323, 334, 355, 367, 368, 379, 376, 
    0, 102, 117, 131, 155, 157, 141, 128, 113, 105, 119, 135, 143, 144, 143, 137, 141, 146, 142, 140, 141, 143, 142, 139, 138, 141, 148, 155, 156, 155, 181, 303, 
    0, 97, 111, 124, 156, 171, 163, 127, 65, 61, 95, 107, 115, 120, 109, 107, 118, 130, 129, 131, 129, 131, 131, 125, 126, 146, 146, 138, 142, 145, 175, 302, 
    0, 101, 117, 120, 136, 152, 146, 108, 41, 42, 37, 10, 20, 29, 25, 21, 23, 30, 29, 30, 31, 33, 41, 46, 46, 105, 140, 135, 140, 141, 171, 301, 
    0, 98, 117, 123, 130, 133, 147, 131, 80, 88, 71, 50, 72, 73, 57, 56, 64, 82, 79, 83, 89, 85, 97, 91, 80, 119, 144, 142, 145, 141, 172, 302, 
    0, 100, 116, 125, 131, 127, 129, 75, 44, 98, 100, 94, 101, 89, 64, 72, 88, 107, 108, 122, 117, 108, 125, 101, 82, 85, 117, 147, 148, 141, 167, 298, 
    0, 104, 116, 124, 132, 122, 95, 22, 11, 51, 52, 53, 63, 70, 42, 33, 34, 43, 37, 46, 40, 32, 52, 47, 51, 29, 66, 125, 134, 131, 157, 290, 
    0, 112, 117, 122, 132, 137, 133, 94, 87, 87, 84, 93, 105, 113, 93, 83, 84, 81, 83, 90, 77, 78, 90, 95, 103, 83, 100, 133, 136, 131, 156, 288, 
    0, 124, 123, 119, 130, 147, 152, 139, 119, 103, 108, 102, 109, 112, 109, 105, 106, 113, 121, 120, 104, 106, 102, 121, 145, 135, 129, 138, 141, 136, 162, 290, 
    0, 136, 138, 126, 136, 144, 140, 137, 119, 102, 107, 99, 97, 105, 106, 105, 104, 104, 104, 110, 107, 106, 105, 107, 124, 136, 138, 142, 141, 136, 164, 292, 
    0, 147, 154, 144, 151, 141, 132, 151, 159, 158, 156, 156, 159, 159, 159, 156, 149, 148, 157, 163, 164, 162, 153, 135, 130, 135, 140, 139, 136, 134, 165, 295, 
    0, 145, 155, 143, 123, 91, 75, 124, 170, 177, 177, 171, 166, 162, 160, 163, 166, 168, 167, 169, 168, 165, 160, 143, 135, 138, 142, 144, 148, 146, 173, 299, 
    0, 142, 150, 126, 96, 64, 22, 7, 40, 88, 128, 143, 138, 131, 132, 136, 140, 143, 146, 149, 147, 142, 142, 146, 147, 148, 149, 150, 149, 143, 166, 292, 
    0, 141, 163, 172, 192, 182, 109, 17, 0, 0, 25, 80, 118, 132, 138, 142, 146, 149, 152, 150, 142, 136, 137, 139, 137, 135, 133, 130, 128, 125, 153, 283, 
    0, 138, 177, 202, 233, 261, 254, 194, 91, 0, 0, 2, 61, 115, 141, 144, 142, 140, 139, 139, 136, 131, 132, 134, 135, 136, 137, 135, 132, 128, 157, 284, 
    0, 135, 154, 154, 170, 211, 263, 285, 247, 119, 0, 0, 0, 15, 68, 115, 135, 138, 138, 139, 139, 140, 142, 143, 142, 143, 145, 143, 142, 137, 160, 286, 
    0, 136, 159, 158, 162, 167, 187, 233, 265, 209, 74, 0, 0, 0, 0, 12, 59, 99, 124, 139, 139, 132, 133, 138, 136, 137, 140, 141, 141, 137, 160, 287, 
    0, 136, 157, 153, 158, 160, 155, 177, 242, 238, 128, 61, 40, 0, 0, 0, 0, 0, 19, 52, 74, 89, 118, 140, 141, 140, 140, 138, 137, 134, 155, 282, 
    0, 135, 156, 149, 152, 155, 158, 163, 215, 216, 104, 48, 58, 52, 36, 8, 0, 0, 0, 0, 0, 0, 0, 53, 93, 118, 137, 146, 145, 137, 154, 282, 
    0, 134, 155, 148, 147, 150, 156, 158, 178, 153, 85, 38, 27, 47, 64, 70, 71, 51, 23, 0, 0, 0, 0, 0, 0, 0, 33, 65, 95, 118, 150, 281, 
    0, 122, 145, 143, 142, 144, 147, 151, 170, 175, 179, 159, 85, 38, 34, 50, 125, 192, 195, 141, 85, 76, 44, 0, 0, 0, 41, 72, 78, 95, 131, 269, 
    0, 118, 141, 142, 143, 147, 147, 180, 227, 265, 299, 287, 220, 169, 160, 170, 218, 262, 266, 240, 220, 233, 235, 211, 170, 157, 165, 151, 133, 127, 140, 269, 
    0, 107, 127, 128, 128, 127, 129, 163, 187, 183, 210, 256, 261, 255, 224, 173, 154, 170, 211, 213, 199, 208, 229, 240, 201, 153, 131, 114, 102, 101, 118, 249, 
    0, 14, 13, 14, 9, 7, 1, 0, 0, 0, 0, 34, 42, 38, 22, 1, 1, 13, 41, 49, 40, 36, 49, 60, 50, 34, 23, 17, 19, 27, 51, 189, 
    0, 9, 3, 2, 5, 10, 12, 14, 15, 14, 18, 18, 14, 10, 7, 7, 16, 23, 13, 8, 13, 12, 3, 0, 7, 16, 21, 18, 8, 0, 13, 140, 
    5, 89, 80, 85, 90, 95, 94, 93, 95, 94, 92, 89, 85, 75, 56, 39, 36, 40, 33, 24, 19, 15, 10, 5, 1, 0, 0, 0, 0, 0, 4, 118, 
    0, 41, 19, 20, 18, 18, 20, 21, 25, 31, 27, 19, 15, 14, 16, 13, 16, 25, 29, 22, 15, 17, 18, 19, 18, 15, 13, 19, 25, 32, 75, 185, 
    0, 48, 24, 25, 26, 35, 41, 44, 54, 63, 56, 53, 53, 56, 59, 61, 67, 78, 84, 80, 78, 78, 79, 79, 77, 75, 78, 85, 105, 147, 187, 220, 
    36, 93, 72, 75, 70, 76, 82, 80, 86, 90, 86, 81, 80, 88, 89, 89, 92, 94, 94, 94, 94, 95, 94, 92, 89, 90, 97, 127, 179, 187, 146, 157, 
    33, 93, 75, 78, 75, 79, 82, 81, 85, 87, 85, 91, 105, 107, 106, 105, 109, 115, 115, 116, 115, 107, 99, 103, 102, 104, 139, 182, 167, 109, 90, 136, 
    38, 98, 82, 85, 79, 80, 83, 84, 86, 90, 91, 93, 101, 104, 105, 102, 104, 108, 110, 109, 108, 101, 94, 100, 116, 152, 175, 140, 97, 92, 98, 136, 
    0, 6, 5, 7, 5, 2, 1, 3, 5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 7, 10, 19, 25, 15, 0, 2, 15, 17, 13, 45, 
    
    -- channel=60
    214, 332, 365, 381, 367, 339, 327, 328, 334, 346, 356, 359, 358, 355, 350, 349, 347, 345, 349, 353, 357, 360, 359, 359, 358, 363, 376, 391, 400, 405, 397, 274, 
    201, 278, 309, 328, 317, 285, 269, 264, 263, 272, 287, 295, 292, 288, 279, 280, 287, 285, 283, 283, 287, 292, 290, 287, 290, 304, 328, 346, 350, 350, 346, 241, 
    197, 271, 302, 321, 328, 319, 302, 274, 251, 270, 295, 307, 310, 307, 300, 303, 312, 316, 317, 317, 322, 320, 310, 315, 322, 335, 349, 349, 347, 345, 342, 239, 
    200, 272, 301, 317, 326, 328, 307, 252, 202, 225, 238, 238, 242, 232, 231, 241, 250, 253, 252, 256, 262, 258, 249, 262, 293, 331, 344, 342, 348, 347, 344, 241, 
    197, 270, 295, 310, 317, 327, 320, 276, 245, 248, 221, 207, 220, 212, 214, 226, 230, 234, 232, 235, 236, 237, 235, 245, 280, 323, 342, 340, 349, 347, 346, 243, 
    194, 266, 294, 307, 310, 315, 303, 265, 262, 281, 268, 273, 279, 264, 255, 274, 289, 304, 307, 310, 305, 305, 307, 304, 314, 326, 340, 347, 355, 353, 351, 245, 
    196, 265, 290, 306, 308, 303, 268, 202, 207, 239, 243, 246, 241, 233, 227, 238, 244, 251, 258, 263, 246, 251, 260, 256, 252, 262, 305, 338, 341, 343, 342, 241, 
    205, 270, 289, 305, 308, 302, 279, 237, 230, 239, 244, 246, 247, 254, 248, 248, 246, 239, 246, 243, 228, 233, 248, 266, 254, 253, 295, 330, 334, 335, 334, 236, 
    218, 279, 289, 304, 308, 315, 318, 308, 283, 273, 277, 281, 280, 277, 281, 290, 296, 294, 297, 294, 281, 285, 288, 313, 325, 323, 325, 334, 336, 333, 333, 234, 
    233, 294, 294, 303, 307, 314, 317, 301, 265, 255, 253, 251, 251, 248, 258, 267, 270, 269, 269, 262, 255, 263, 263, 292, 334, 339, 332, 335, 339, 334, 332, 232, 
    243, 311, 309, 316, 313, 310, 314, 304, 282, 281, 278, 278, 280, 288, 298, 300, 296, 287, 284, 285, 288, 293, 294, 305, 329, 332, 329, 330, 332, 331, 332, 234, 
    249, 322, 318, 315, 296, 279, 294, 324, 330, 332, 330, 331, 336, 339, 344, 345, 343, 339, 336, 335, 334, 336, 335, 333, 333, 331, 333, 332, 334, 336, 337, 239, 
    251, 324, 313, 278, 225, 184, 193, 252, 298, 322, 330, 330, 331, 334, 338, 340, 339, 336, 333, 330, 329, 331, 335, 333, 332, 335, 340, 342, 345, 346, 343, 240, 
    255, 330, 328, 294, 248, 194, 135, 116, 151, 221, 284, 318, 329, 334, 340, 343, 345, 344, 345, 340, 335, 334, 338, 337, 336, 335, 334, 333, 334, 333, 330, 230, 
    256, 336, 351, 355, 356, 336, 265, 170, 104, 105, 165, 246, 307, 340, 350, 349, 346, 344, 342, 335, 327, 326, 327, 326, 325, 326, 326, 325, 325, 326, 325, 227, 
    256, 338, 350, 354, 353, 361, 359, 313, 209, 112, 98, 145, 216, 286, 329, 343, 343, 338, 334, 331, 329, 331, 332, 333, 333, 336, 334, 332, 330, 330, 327, 228, 
    258, 343, 356, 362, 359, 360, 364, 358, 284, 152, 79, 79, 98, 143, 213, 277, 315, 331, 334, 332, 329, 331, 333, 332, 331, 333, 332, 332, 333, 332, 329, 232, 
    260, 346, 357, 365, 363, 363, 358, 357, 315, 186, 93, 78, 72, 70, 86, 124, 177, 232, 275, 298, 306, 318, 334, 338, 335, 332, 329, 328, 330, 329, 327, 232, 
    261, 347, 355, 359, 358, 359, 358, 354, 318, 181, 75, 68, 69, 73, 76, 71, 67, 79, 107, 138, 168, 217, 275, 309, 322, 330, 332, 331, 331, 330, 326, 230, 
    262, 348, 355, 358, 357, 358, 361, 344, 281, 138, 30, 17, 32, 55, 75, 86, 86, 71, 50, 25, 7, 33, 94, 152, 201, 247, 285, 311, 327, 332, 331, 233, 
    257, 345, 351, 354, 351, 355, 355, 321, 237, 143, 89, 44, 22, 38, 56, 98, 135, 138, 113, 79, 62, 52, 45, 37, 56, 122, 183, 229, 275, 306, 321, 231, 
    250, 335, 348, 351, 348, 351, 350, 333, 280, 266, 268, 201, 122, 96, 107, 178, 266, 289, 237, 168, 176, 203, 182, 139, 145, 221, 279, 288, 291, 300, 305, 222, 
    242, 325, 340, 342, 338, 337, 338, 343, 343, 356, 361, 326, 285, 283, 283, 307, 337, 338, 324, 290, 301, 314, 313, 303, 296, 313, 316, 313, 317, 312, 302, 216, 
    185, 246, 259, 256, 246, 239, 232, 227, 221, 217, 220, 216, 215, 228, 232, 239, 239, 225, 229, 235, 245, 242, 246, 254, 257, 249, 232, 225, 231, 237, 239, 176, 
    108, 121, 127, 125, 115, 110, 106, 102, 97, 93, 93, 87, 83, 86, 96, 119, 139, 141, 138, 140, 141, 141, 144, 149, 156, 161, 165, 164, 161, 156, 153, 115, 
    121, 146, 160, 160, 159, 157, 154, 152, 148, 146, 144, 138, 136, 135, 133, 132, 131, 124, 113, 110, 109, 105, 99, 98, 100, 102, 104, 100, 90, 79, 81, 68, 
    88, 92, 102, 105, 102, 96, 86, 77, 74, 70, 62, 57, 54, 51, 51, 50, 53, 48, 37, 30, 25, 24, 24, 24, 22, 22, 22, 20, 17, 26, 56, 60, 
    49, 26, 31, 31, 28, 30, 28, 29, 34, 32, 24, 21, 21, 25, 28, 30, 36, 39, 35, 29, 25, 26, 31, 34, 33, 31, 30, 33, 50, 84, 124, 102, 
    55, 42, 47, 46, 43, 44, 41, 43, 48, 43, 37, 38, 40, 41, 40, 43, 46, 46, 40, 37, 37, 37, 36, 36, 36, 36, 44, 71, 112, 139, 133, 68, 
    49, 34, 38, 37, 36, 38, 37, 38, 39, 35, 37, 45, 52, 52, 50, 54, 59, 56, 51, 50, 49, 45, 42, 40, 41, 54, 86, 126, 142, 108, 61, 18, 
    52, 38, 40, 40, 44, 46, 44, 44, 43, 42, 52, 71, 81, 76, 71, 74, 81, 82, 82, 80, 71, 53, 46, 44, 57, 92, 132, 134, 92, 46, 36, 25, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 8, 8, 6, 5, 7, 7, 10, 11, 9, 0, 0, 5, 24, 56, 60, 25, 0, 0, 3, 0, 
    
    -- channel=61
    289, 302, 329, 331, 297, 277, 281, 283, 291, 306, 314, 310, 306, 302, 297, 303, 298, 296, 301, 304, 311, 310, 306, 305, 307, 318, 336, 344, 347, 353, 327, 73, 
    345, 300, 323, 332, 294, 266, 264, 260, 269, 288, 299, 294, 289, 279, 272, 281, 285, 282, 283, 284, 289, 288, 283, 283, 290, 312, 333, 343, 342, 342, 307, 10, 
    347, 299, 317, 328, 311, 296, 285, 254, 279, 310, 309, 318, 311, 301, 301, 316, 321, 315, 319, 320, 323, 318, 310, 317, 337, 346, 349, 347, 339, 339, 304, 6, 
    349, 300, 311, 321, 319, 314, 276, 232, 251, 263, 258, 275, 271, 258, 262, 279, 282, 281, 282, 283, 286, 284, 269, 292, 337, 348, 340, 339, 341, 344, 312, 9, 
    348, 295, 304, 312, 316, 318, 282, 261, 285, 274, 249, 258, 248, 233, 255, 271, 273, 260, 266, 265, 260, 266, 251, 284, 332, 335, 335, 340, 342, 346, 314, 10, 
    343, 290, 302, 309, 309, 309, 269, 268, 310, 288, 285, 297, 287, 280, 292, 310, 316, 320, 331, 319, 317, 321, 313, 332, 352, 352, 347, 343, 344, 347, 318, 13, 
    344, 286, 300, 307, 306, 287, 247, 245, 260, 262, 270, 279, 265, 256, 268, 281, 281, 284, 292, 282, 275, 282, 292, 282, 273, 311, 336, 335, 334, 342, 313, 12, 
    352, 286, 298, 309, 304, 282, 262, 259, 267, 265, 268, 274, 260, 260, 275, 283, 277, 270, 276, 256, 257, 266, 279, 277, 269, 303, 326, 326, 325, 333, 306, 9, 
    369, 287, 295, 309, 303, 297, 298, 296, 292, 287, 283, 287, 280, 274, 288, 301, 307, 303, 300, 286, 292, 298, 304, 331, 329, 340, 342, 331, 329, 332, 302, 9, 
    390, 296, 293, 307, 303, 306, 306, 278, 258, 261, 256, 255, 258, 257, 269, 277, 277, 273, 268, 261, 262, 269, 274, 317, 341, 339, 333, 330, 330, 332, 301, 7, 
    406, 306, 302, 315, 301, 301, 308, 284, 270, 276, 271, 275, 278, 290, 299, 299, 296, 285, 279, 276, 283, 288, 297, 322, 334, 328, 324, 324, 324, 329, 302, 9, 
    415, 317, 300, 296, 268, 270, 315, 330, 316, 318, 315, 320, 330, 335, 339, 338, 332, 327, 323, 320, 320, 326, 329, 333, 333, 326, 326, 326, 327, 335, 308, 10, 
    418, 321, 282, 246, 197, 175, 219, 285, 324, 337, 332, 326, 329, 336, 340, 339, 335, 331, 327, 322, 322, 328, 331, 327, 325, 327, 330, 333, 336, 341, 310, 12, 
    422, 331, 300, 266, 218, 156, 124, 141, 195, 268, 321, 339, 337, 338, 341, 341, 339, 338, 335, 328, 327, 331, 331, 328, 328, 329, 328, 328, 327, 332, 301, 7, 
    425, 341, 328, 323, 312, 274, 204, 136, 107, 152, 229, 299, 344, 354, 349, 343, 339, 337, 334, 324, 321, 325, 324, 320, 321, 322, 320, 319, 320, 326, 296, 7, 
    428, 347, 341, 344, 334, 322, 295, 229, 129, 95, 152, 213, 271, 330, 354, 349, 337, 330, 325, 321, 322, 326, 326, 325, 327, 328, 325, 324, 323, 327, 298, 9, 
    433, 354, 347, 352, 346, 343, 336, 292, 170, 72, 90, 131, 154, 199, 259, 310, 335, 340, 336, 325, 320, 327, 330, 326, 327, 327, 324, 325, 325, 329, 301, 12, 
    437, 355, 347, 355, 349, 347, 342, 328, 208, 64, 69, 96, 94, 115, 139, 171, 217, 264, 298, 309, 315, 337, 343, 334, 331, 326, 322, 322, 323, 326, 302, 14, 
    439, 355, 343, 351, 346, 345, 343, 335, 213, 40, 37, 78, 77, 92, 103, 108, 109, 119, 139, 159, 199, 268, 319, 331, 334, 334, 328, 325, 323, 327, 302, 13, 
    438, 353, 340, 347, 346, 347, 347, 307, 170, 28, 0, 28, 58, 77, 90, 99, 94, 86, 71, 47, 47, 101, 157, 186, 229, 275, 303, 326, 337, 338, 309, 17, 
    430, 351, 340, 345, 344, 347, 342, 264, 151, 84, 50, 16, 25, 58, 90, 150, 161, 121, 66, 55, 85, 83, 66, 64, 126, 204, 229, 255, 296, 322, 303, 17, 
    422, 347, 340, 346, 343, 344, 337, 285, 230, 233, 210, 132, 105, 106, 141, 229, 277, 252, 169, 141, 178, 187, 154, 125, 184, 265, 291, 300, 306, 309, 288, 11, 
    407, 340, 336, 335, 329, 326, 322, 310, 306, 334, 318, 252, 240, 257, 277, 327, 336, 304, 263, 260, 292, 288, 271, 268, 293, 319, 309, 307, 318, 315, 285, 16, 
    314, 259, 262, 254, 244, 236, 232, 228, 223, 225, 216, 194, 199, 225, 244, 267, 258, 233, 227, 233, 253, 252, 248, 253, 263, 262, 248, 245, 249, 253, 240, 7, 
    230, 151, 151, 146, 137, 131, 129, 122, 117, 117, 113, 107, 109, 117, 134, 158, 170, 165, 167, 172, 169, 168, 176, 184, 186, 188, 193, 192, 189, 187, 176, 0, 
    207, 152, 171, 167, 164, 158, 154, 152, 150, 146, 141, 136, 137, 142, 148, 156, 151, 133, 126, 127, 127, 123, 122, 124, 126, 128, 128, 121, 112, 105, 112, 0, 
    157, 98, 121, 121, 117, 109, 98, 92, 88, 77, 69, 68, 71, 72, 72, 73, 73, 60, 47, 43, 42, 42, 42, 43, 40, 39, 39, 33, 30, 55, 83, 0, 
    107, 32, 52, 48, 47, 42, 36, 42, 39, 29, 25, 28, 30, 33, 36, 37, 41, 35, 27, 25, 24, 27, 32, 32, 33, 33, 32, 38, 65, 99, 100, 0, 
    93, 31, 52, 45, 48, 45, 40, 45, 43, 34, 32, 38, 44, 41, 38, 43, 43, 36, 30, 29, 32, 34, 35, 34, 34, 35, 52, 87, 108, 99, 83, 0, 
    91, 27, 43, 39, 41, 39, 38, 41, 37, 33, 44, 56, 54, 49, 49, 57, 57, 49, 45, 45, 39, 35, 37, 32, 37, 65, 100, 109, 91, 64, 34, 0, 
    90, 25, 42, 39, 47, 48, 46, 45, 42, 41, 58, 77, 77, 68, 64, 71, 74, 73, 74, 72, 56, 42, 40, 40, 65, 99, 107, 87, 51, 17, 23, 0, 
    25, 0, 0, 0, 0, 4, 4, 2, 0, 0, 9, 16, 11, 9, 7, 10, 11, 11, 13, 12, 3, 0, 0, 3, 25, 50, 40, 0, 0, 0, 0, 0, 
    
    -- channel=62
    44, 17, 15, 8, 0, 6, 15, 16, 19, 21, 22, 21, 24, 21, 23, 23, 19, 23, 24, 26, 26, 24, 25, 25, 24, 26, 24, 23, 22, 25, 21, 0, 
    162, 148, 149, 151, 127, 114, 125, 131, 139, 143, 148, 145, 145, 141, 138, 144, 140, 138, 141, 143, 146, 145, 144, 145, 148, 155, 165, 173, 176, 181, 169, 0, 
    158, 147, 146, 152, 136, 120, 123, 141, 161, 158, 160, 159, 156, 157, 151, 157, 157, 154, 154, 154, 156, 158, 156, 158, 152, 158, 170, 178, 177, 181, 170, 0, 
    157, 148, 144, 153, 151, 144, 130, 129, 163, 178, 178, 186, 184, 181, 179, 183, 188, 187, 190, 190, 186, 191, 184, 189, 189, 179, 176, 181, 179, 184, 173, 0, 
    158, 148, 139, 149, 150, 148, 124, 111, 145, 150, 147, 155, 147, 148, 150, 161, 155, 149, 159, 152, 148, 160, 146, 158, 193, 182, 170, 174, 177, 182, 171, 0, 
    156, 147, 140, 146, 149, 146, 131, 149, 169, 138, 132, 148, 144, 144, 148, 158, 156, 152, 155, 150, 149, 156, 151, 162, 203, 198, 180, 178, 179, 183, 172, 0, 
    151, 143, 138, 145, 146, 137, 135, 156, 184, 152, 154, 169, 148, 147, 162, 172, 173, 175, 181, 171, 182, 178, 175, 172, 189, 203, 191, 180, 179, 185, 173, 0, 
    149, 137, 135, 144, 144, 121, 107, 128, 156, 143, 139, 145, 132, 131, 143, 147, 146, 149, 153, 141, 156, 152, 157, 151, 136, 175, 192, 175, 168, 175, 167, 0, 
    152, 134, 133, 144, 139, 116, 111, 129, 145, 142, 137, 141, 145, 140, 138, 141, 143, 142, 141, 137, 146, 151, 164, 156, 130, 159, 177, 169, 165, 170, 161, 0, 
    165, 134, 130, 141, 140, 136, 136, 128, 130, 133, 130, 135, 133, 131, 131, 135, 144, 144, 139, 133, 138, 143, 150, 159, 159, 166, 167, 163, 164, 169, 158, 0, 
    179, 144, 132, 141, 138, 144, 142, 120, 110, 114, 109, 110, 111, 113, 116, 118, 121, 120, 118, 115, 119, 123, 127, 148, 166, 167, 166, 166, 165, 169, 158, 0, 
    191, 159, 138, 154, 150, 160, 166, 140, 125, 127, 127, 128, 131, 137, 141, 140, 138, 136, 136, 136, 137, 140, 144, 154, 162, 163, 163, 164, 163, 168, 158, 0, 
    198, 167, 138, 144, 136, 138, 181, 199, 182, 163, 151, 151, 155, 159, 162, 161, 159, 157, 156, 154, 155, 157, 159, 160, 161, 162, 164, 167, 167, 172, 165, 0, 
    202, 172, 133, 107, 79, 61, 95, 158, 194, 202, 187, 168, 162, 163, 165, 165, 165, 164, 162, 160, 162, 166, 166, 165, 166, 167, 169, 171, 171, 175, 165, 0, 
    206, 178, 148, 132, 110, 71, 33, 38, 95, 154, 189, 194, 182, 172, 169, 171, 172, 174, 173, 167, 166, 169, 167, 165, 164, 163, 163, 164, 163, 167, 157, 0, 
    206, 183, 167, 170, 164, 146, 105, 41, 16, 67, 130, 178, 209, 211, 194, 179, 172, 171, 171, 168, 166, 166, 166, 164, 162, 161, 160, 159, 158, 162, 151, 0, 
    207, 188, 174, 177, 175, 176, 171, 128, 38, 19, 71, 111, 158, 202, 221, 214, 195, 180, 169, 164, 165, 167, 165, 164, 165, 165, 163, 163, 161, 162, 151, 0, 
    210, 193, 182, 189, 186, 184, 185, 173, 87, 18, 43, 63, 82, 117, 158, 194, 213, 215, 205, 187, 178, 173, 165, 161, 163, 164, 164, 165, 163, 163, 153, 0, 
    213, 195, 184, 194, 191, 187, 185, 180, 116, 40, 46, 61, 61, 66, 77, 100, 133, 164, 187, 195, 200, 212, 208, 193, 182, 172, 164, 162, 160, 162, 152, 0, 
    216, 196, 182, 193, 191, 187, 187, 175, 128, 41, 21, 49, 54, 57, 62, 60, 62, 71, 81, 92, 113, 160, 195, 208, 217, 212, 201, 188, 173, 167, 154, 0, 
    216, 196, 181, 189, 189, 188, 186, 158, 103, 26, 0, 0, 30, 46, 65, 67, 40, 23, 14, 25, 16, 32, 76, 113, 152, 161, 161, 174, 179, 179, 160, 0, 
    211, 191, 179, 183, 185, 187, 181, 138, 76, 46, 4, 0, 0, 0, 18, 64, 74, 50, 9, 8, 20, 8, 0, 2, 48, 97, 115, 127, 149, 167, 156, 0, 
    208, 191, 180, 185, 189, 190, 186, 166, 141, 143, 125, 63, 27, 31, 52, 109, 149, 138, 86, 60, 86, 91, 66, 46, 73, 125, 146, 148, 155, 164, 152, 0, 
    211, 210, 197, 201, 203, 203, 202, 201, 202, 204, 195, 169, 149, 147, 154, 165, 169, 165, 150, 138, 142, 148, 145, 136, 135, 139, 143, 144, 150, 157, 149, 9, 
    142, 138, 130, 125, 122, 118, 114, 112, 109, 109, 107, 102, 98, 98, 105, 116, 111, 104, 108, 110, 109, 109, 115, 119, 116, 109, 104, 102, 110, 121, 127, 8, 
    96, 83, 75, 71, 68, 65, 68, 69, 68, 70, 68, 63, 61, 63, 69, 83, 90, 84, 84, 88, 89, 88, 90, 95, 98, 100, 100, 96, 92, 97, 106, 0, 
    106, 100, 96, 97, 95, 88, 87, 89, 89, 88, 84, 82, 80, 79, 79, 80, 84, 75, 69, 71, 72, 69, 66, 65, 67, 69, 70, 66, 61, 64, 66, 0, 
    71, 64, 65, 66, 65, 61, 56, 58, 57, 54, 48, 46, 44, 45, 46, 48, 49, 45, 39, 36, 35, 36, 35, 34, 33, 33, 33, 33, 32, 37, 57, 0, 
    48, 37, 35, 36, 39, 37, 35, 38, 39, 35, 30, 30, 29, 30, 35, 38, 38, 38, 33, 30, 28, 30, 32, 32, 28, 29, 31, 32, 40, 66, 85, 0, 
    47, 36, 33, 29, 32, 30, 30, 34, 35, 32, 29, 23, 24, 24, 28, 33, 32, 28, 23, 23, 23, 30, 32, 32, 35, 36, 35, 48, 74, 78, 65, 0, 
    44, 37, 36, 32, 31, 30, 29, 33, 33, 33, 40, 44, 42, 41, 42, 50, 50, 45, 43, 41, 34, 35, 37, 37, 41, 49, 67, 82, 67, 47, 45, 0, 
    64, 51, 50, 48, 50, 50, 49, 50, 50, 51, 60, 71, 70, 68, 67, 71, 75, 74, 74, 72, 62, 53, 54, 60, 79, 101, 101, 78, 53, 47, 56, 9, 
    
    -- channel=63
    64, 8, 2, 0, 0, 0, 0, 0, 0, 4, 4, 1, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 0, 0, 0, 0, 3, 3, 1, 1, 0, 0, 
    135, 105, 102, 104, 86, 78, 91, 97, 102, 109, 111, 107, 106, 104, 103, 108, 104, 102, 104, 106, 110, 108, 106, 109, 109, 115, 119, 118, 116, 117, 113, 23, 
    131, 99, 94, 103, 96, 80, 86, 104, 122, 124, 118, 116, 112, 110, 105, 112, 112, 108, 109, 107, 110, 112, 105, 108, 109, 107, 113, 119, 122, 119, 114, 24, 
    131, 94, 89, 99, 96, 95, 95, 119, 158, 155, 149, 156, 150, 148, 150, 159, 156, 154, 157, 151, 151, 155, 140, 151, 155, 125, 118, 123, 126, 122, 115, 26, 
    129, 93, 86, 94, 95, 103, 125, 135, 155, 152, 156, 173, 170, 166, 167, 169, 173, 169, 167, 165, 162, 165, 160, 155, 168, 139, 115, 121, 122, 123, 119, 29, 
    129, 96, 86, 91, 89, 97, 138, 148, 161, 151, 151, 161, 145, 156, 168, 171, 168, 155, 153, 152, 149, 146, 154, 133, 140, 140, 120, 117, 118, 122, 120, 29, 
    127, 93, 87, 89, 87, 96, 128, 164, 183, 160, 146, 149, 143, 149, 166, 164, 162, 154, 151, 152, 155, 147, 152, 144, 146, 163, 145, 123, 119, 121, 121, 31, 
    129, 90, 84, 91, 87, 104, 143, 157, 170, 152, 142, 151, 156, 141, 153, 155, 160, 152, 161, 159, 160, 169, 158, 153, 142, 156, 144, 116, 115, 116, 117, 30, 
    133, 89, 83, 92, 96, 117, 139, 138, 135, 133, 134, 130, 135, 122, 129, 138, 145, 138, 140, 141, 141, 148, 131, 141, 128, 121, 124, 113, 113, 111, 109, 25, 
    139, 89, 80, 92, 93, 97, 97, 98, 98, 101, 101, 99, 100, 98, 101, 108, 112, 108, 102, 104, 107, 107, 109, 127, 123, 112, 108, 106, 106, 107, 105, 23, 
    148, 94, 78, 89, 85, 88, 93, 86, 78, 82, 77, 81, 83, 82, 87, 88, 90, 92, 91, 84, 85, 87, 88, 104, 114, 110, 108, 108, 109, 110, 106, 22, 
    153, 102, 86, 94, 87, 92, 107, 101, 84, 83, 84, 84, 89, 93, 97, 99, 97, 93, 90, 88, 86, 92, 93, 96, 107, 108, 109, 109, 108, 108, 107, 22, 
    156, 109, 86, 88, 81, 88, 120, 129, 114, 104, 99, 100, 104, 108, 111, 111, 110, 107, 104, 102, 103, 106, 106, 105, 105, 106, 107, 107, 107, 108, 110, 25, 
    160, 111, 85, 74, 61, 44, 68, 121, 145, 141, 125, 112, 111, 113, 114, 114, 112, 110, 108, 106, 107, 111, 111, 109, 107, 109, 110, 113, 115, 116, 115, 30, 
    162, 116, 100, 91, 68, 39, 11, 27, 74, 121, 146, 140, 126, 118, 115, 116, 116, 116, 114, 112, 112, 113, 114, 112, 111, 110, 110, 111, 112, 113, 110, 25, 
    162, 119, 103, 112, 111, 103, 71, 19, 5, 41, 95, 135, 147, 140, 128, 122, 119, 119, 118, 115, 112, 113, 111, 109, 108, 107, 106, 106, 106, 106, 105, 23, 
    162, 121, 106, 114, 111, 112, 119, 92, 25, 6, 46, 81, 118, 150, 155, 142, 129, 121, 117, 115, 114, 113, 112, 111, 111, 111, 108, 107, 104, 104, 104, 22, 
    164, 125, 112, 121, 118, 117, 119, 122, 73, 9, 28, 54, 59, 85, 121, 145, 150, 144, 135, 124, 118, 120, 117, 112, 111, 110, 108, 107, 107, 106, 106, 25, 
    166, 128, 115, 126, 124, 122, 121, 121, 92, 27, 29, 54, 50, 51, 57, 77, 104, 126, 141, 141, 139, 143, 138, 124, 118, 114, 109, 108, 108, 108, 108, 28, 
    168, 131, 117, 126, 125, 123, 123, 118, 85, 33, 29, 53, 56, 59, 59, 56, 52, 55, 64, 80, 98, 128, 149, 146, 142, 137, 127, 119, 116, 112, 109, 29, 
    167, 135, 120, 125, 127, 124, 123, 103, 79, 43, 9, 21, 40, 52, 60, 67, 57, 41, 26, 17, 19, 37, 66, 88, 114, 132, 133, 135, 134, 125, 116, 34, 
    164, 133, 122, 124, 123, 123, 119, 102, 76, 63, 23, 0, 0, 28, 50, 83, 73, 37, 9, 22, 38, 14, 7, 19, 55, 86, 81, 89, 112, 119, 114, 35, 
    161, 129, 122, 125, 123, 123, 124, 123, 99, 90, 84, 41, 15, 26, 35, 70, 101, 94, 62, 36, 59, 67, 46, 30, 41, 79, 100, 100, 103, 106, 104, 30, 
    154, 132, 128, 130, 130, 127, 128, 129, 129, 131, 131, 117, 93, 91, 94, 104, 118, 123, 119, 98, 94, 105, 109, 99, 90, 97, 108, 116, 121, 118, 109, 37, 
    115, 108, 111, 110, 109, 103, 102, 100, 98, 99, 95, 90, 90, 94, 103, 109, 101, 91, 91, 95, 95, 93, 96, 101, 101, 95, 90, 89, 94, 99, 98, 41, 
    90, 59, 65, 65, 62, 58, 55, 53, 51, 48, 47, 46, 45, 46, 49, 61, 68, 61, 62, 66, 65, 65, 66, 69, 72, 74, 75, 71, 73, 76, 76, 33, 
    88, 67, 73, 74, 73, 68, 66, 67, 66, 63, 64, 65, 63, 64, 65, 64, 66, 62, 57, 59, 60, 59, 57, 58, 59, 60, 61, 63, 58, 54, 59, 12, 
    69, 53, 62, 63, 65, 61, 55, 54, 53, 48, 44, 45, 46, 43, 43, 43, 45, 42, 34, 31, 33, 34, 35, 33, 32, 32, 32, 31, 29, 26, 19, 0, 
    58, 30, 37, 37, 38, 34, 34, 36, 35, 31, 30, 29, 30, 30, 30, 32, 32, 30, 27, 25, 24, 25, 25, 26, 29, 29, 24, 22, 21, 4, 0, 0, 
    58, 33, 36, 33, 37, 36, 32, 34, 34, 31, 29, 32, 32, 29, 29, 31, 29, 27, 25, 25, 25, 24, 24, 25, 24, 23, 26, 20, 1, 2, 26, 8, 
    59, 31, 33, 28, 31, 33, 31, 31, 31, 31, 35, 35, 33, 32, 33, 36, 37, 34, 32, 30, 27, 27, 32, 28, 25, 25, 14, 0, 8, 25, 30, 5, 
    59, 36, 39, 37, 39, 41, 41, 41, 41, 39, 45, 54, 54, 51, 49, 51, 55, 54, 54, 53, 47, 40, 41, 39, 34, 23, 13, 25, 33, 32, 40, 17, 
    
    -- channel=64
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=65
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 11, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 8, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=66
    196, 96, 56, 82, 128, 133, 118, 113, 96, 53, 79, 166, 158, 113, 103, 133, 165, 158, 137, 142, 129, 84, 91, 183, 177, 32, 70, 175, 124, 112, 128, 35, 
    245, 141, 76, 113, 178, 163, 143, 156, 124, 71, 115, 212, 210, 154, 135, 192, 228, 200, 201, 224, 211, 137, 139, 263, 257, 64, 87, 216, 179, 160, 148, 49, 
    249, 150, 94, 130, 193, 161, 147, 158, 109, 68, 134, 212, 208, 165, 135, 208, 238, 164, 155, 207, 212, 132, 135, 276, 266, 61, 63, 194, 175, 140, 109, 42, 
    258, 148, 112, 135, 192, 155, 156, 157, 93, 67, 143, 198, 193, 172, 144, 194, 233, 176, 148, 186, 205, 139, 147, 277, 270, 83, 68, 189, 184, 135, 98, 15, 
    272, 170, 159, 144, 183, 158, 154, 156, 94, 68, 139, 179, 178, 167, 162, 175, 194, 182, 163, 172, 220, 177, 156, 279, 281, 119, 89, 179, 198, 158, 121, 15, 
    265, 158, 187, 200, 182, 160, 130, 138, 106, 81, 156, 186, 186, 178, 167, 158, 188, 211, 146, 115, 224, 226, 161, 274, 296, 136, 98, 172, 200, 166, 129, 46, 
    248, 127, 168, 221, 182, 164, 116, 107, 101, 117, 206, 217, 211, 202, 165, 143, 188, 254, 163, 63, 202, 245, 175, 270, 315, 156, 112, 176, 193, 130, 68, 64, 
    226, 119, 177, 222, 141, 125, 134, 109, 74, 143, 250, 237, 221, 195, 138, 138, 197, 220, 173, 116, 182, 222, 195, 268, 300, 195, 138, 182, 180, 81, 19, 67, 
    219, 118, 220, 253, 149, 68, 104, 156, 109, 161, 243, 219, 199, 153, 119, 181, 231, 186, 149, 186, 211, 211, 214, 279, 290, 204, 163, 179, 159, 48, 17, 78, 
    228, 114, 236, 279, 189, 89, 41, 128, 196, 228, 236, 214, 165, 88, 111, 208, 241, 201, 186, 216, 235, 212, 200, 299, 319, 202, 174, 173, 134, 21, 24, 93, 
    228, 102, 237, 287, 214, 145, 41, 50, 193, 260, 228, 220, 168, 107, 132, 173, 184, 196, 224, 230, 239, 209, 167, 275, 310, 197, 186, 175, 121, 12, 20, 101, 
    229, 92, 236, 287, 236, 200, 105, 49, 151, 219, 199, 203, 163, 156, 223, 212, 178, 187, 208, 216, 207, 196, 189, 267, 277, 181, 193, 203, 132, 16, 23, 82, 
    218, 81, 206, 256, 230, 240, 179, 129, 155, 188, 190, 192, 163, 151, 206, 228, 209, 205, 202, 191, 168, 167, 191, 244, 270, 189, 174, 212, 150, 30, 53, 55, 
    231, 97, 181, 219, 196, 243, 235, 177, 162, 178, 205, 197, 186, 177, 173, 171, 175, 184, 197, 196, 177, 178, 176, 184, 215, 202, 191, 207, 155, 58, 109, 61, 
    255, 123, 198, 213, 176, 215, 252, 187, 162, 124, 130, 212, 237, 211, 204, 180, 157, 144, 155, 182, 175, 202, 217, 175, 143, 153, 208, 201, 136, 82, 168, 88, 
    260, 133, 196, 219, 183, 184, 223, 193, 210, 175, 32, 124, 255, 216, 197, 203, 195, 175, 155, 155, 141, 146, 212, 228, 165, 105, 158, 202, 100, 57, 197, 97, 
    265, 151, 175, 210, 196, 190, 202, 196, 210, 255, 108, 40, 186, 215, 189, 174, 174, 199, 210, 196, 186, 164, 158, 208, 216, 152, 126, 179, 103, 39, 208, 112, 
    272, 178, 180, 181, 172, 184, 212, 202, 199, 225, 244, 111, 97, 192, 205, 184, 176, 162, 178, 190, 176, 196, 186, 177, 179, 157, 162, 177, 172, 90, 168, 76, 
    283, 184, 181, 176, 158, 161, 218, 210, 210, 163, 247, 256, 105, 140, 193, 171, 189, 180, 169, 162, 150, 182, 203, 177, 158, 113, 121, 169, 195, 194, 193, 20, 
    298, 167, 165, 169, 172, 147, 210, 216, 216, 195, 153, 268, 246, 158, 179, 167, 149, 183, 202, 151, 128, 173, 194, 166, 159, 110, 89, 137, 148, 215, 244, 13, 
    303, 130, 161, 189, 165, 134, 195, 203, 160, 233, 165, 139, 280, 255, 180, 169, 154, 150, 184, 179, 144, 167, 193, 168, 154, 136, 118, 142, 160, 187, 202, 22, 
    298, 103, 170, 236, 163, 132, 188, 210, 147, 168, 219, 137, 195, 273, 219, 163, 168, 154, 132, 162, 176, 170, 178, 175, 153, 146, 133, 168, 209, 187, 175, 32, 
    286, 131, 180, 194, 148, 128, 163, 229, 208, 140, 173, 227, 207, 223, 230, 191, 167, 168, 138, 135, 170, 180, 175, 176, 165, 161, 164, 186, 206, 190, 194, 38, 
    291, 179, 223, 184, 130, 133, 145, 202, 221, 175, 150, 203, 253, 215, 211, 206, 169, 172, 148, 135, 185, 170, 149, 174, 172, 177, 199, 224, 202, 203, 215, 28, 
    332, 244, 288, 260, 199, 163, 166, 193, 184, 171, 207, 196, 195, 212, 199, 193, 185, 207, 175, 136, 187, 188, 127, 150, 176, 165, 162, 239, 247, 218, 216, 45, 
    325, 226, 298, 350, 304, 236, 196, 200, 194, 165, 209, 252, 213, 203, 196, 165, 200, 261, 234, 168, 166, 188, 150, 133, 162, 146, 107, 227, 284, 214, 206, 60, 
    292, 160, 215, 359, 384, 318, 268, 218, 199, 195, 191, 220, 238, 222, 186, 129, 150, 259, 269, 196, 168, 159, 162, 157, 145, 106, 122, 229, 262, 196, 193, 73, 
    276, 124, 116, 258, 390, 386, 328, 285, 218, 191, 204, 211, 226, 229, 206, 158, 119, 188, 253, 198, 184, 189, 143, 144, 139, 97, 159, 234, 243, 220, 164, 17, 
    279, 113, 87, 140, 276, 404, 379, 334, 276, 210, 189, 213, 232, 227, 236, 230, 192, 198, 222, 198, 189, 194, 152, 132, 113, 110, 186, 208, 243, 323, 196, 0, 
    287, 123, 140, 137, 149, 302, 404, 382, 333, 284, 225, 202, 214, 213, 230, 225, 184, 205, 237, 211, 204, 211, 188, 173, 127, 104, 152, 157, 223, 320, 214, 0, 
    272, 136, 201, 207, 115, 177, 316, 410, 375, 332, 308, 265, 220, 198, 226, 232, 149, 107, 179, 200, 181, 203, 200, 211, 167, 118, 139, 173, 209, 245, 200, 0, 
    238, 145, 215, 252, 172, 150, 212, 325, 374, 351, 357, 362, 334, 306, 321, 343, 294, 213, 201, 207, 200, 243, 266, 291, 277, 240, 251, 274, 288, 295, 280, 112, 
    
    -- channel=67
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=68
    0, 66, 88, 53, 3, 4, 28, 17, 27, 67, 22, 0, 0, 43, 47, 17, 0, 29, 50, 42, 55, 84, 62, 0, 20, 170, 84, 0, 36, 35, 15, 110, 
    0, 24, 83, 39, 0, 0, 0, 0, 0, 62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 6, 0, 0, 180, 74, 0, 0, 0, 0, 122, 
    0, 10, 76, 22, 0, 0, 0, 0, 10, 71, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 4, 0, 0, 219, 135, 0, 0, 2, 25, 122, 
    0, 1, 69, 16, 0, 0, 0, 0, 36, 69, 0, 0, 0, 0, 0, 0, 0, 2, 10, 0, 0, 39, 0, 0, 0, 220, 152, 0, 0, 19, 81, 155, 
    0, 0, 25, 0, 0, 0, 0, 0, 44, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 164, 126, 0, 0, 29, 74, 197, 
    0, 0, 0, 0, 0, 0, 0, 0, 38, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 122, 121, 0, 0, 3, 23, 161, 
    0, 0, 0, 0, 0, 0, 14, 0, 43, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 85, 0, 0, 1, 0, 0, 87, 110, 0, 0, 15, 63, 118, 
    0, 46, 0, 0, 8, 21, 36, 30, 86, 0, 0, 0, 0, 0, 31, 19, 0, 0, 11, 83, 0, 0, 3, 0, 0, 42, 68, 0, 0, 88, 143, 82, 
    0, 35, 0, 0, 33, 87, 47, 20, 81, 0, 0, 0, 0, 24, 69, 0, 0, 0, 17, 18, 0, 0, 0, 0, 0, 11, 38, 0, 0, 144, 148, 48, 
    0, 18, 0, 0, 0, 129, 100, 10, 0, 0, 0, 0, 17, 119, 92, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 14, 16, 0, 12, 178, 129, 27, 
    0, 36, 0, 0, 0, 75, 165, 93, 0, 0, 0, 0, 48, 149, 69, 0, 0, 0, 0, 0, 0, 0, 35, 0, 0, 30, 0, 0, 41, 205, 125, 13, 
    0, 47, 0, 0, 0, 0, 137, 163, 0, 0, 0, 0, 57, 68, 0, 0, 3, 0, 0, 0, 0, 25, 40, 0, 0, 32, 0, 0, 33, 217, 144, 28, 
    0, 83, 0, 0, 0, 0, 26, 97, 15, 0, 18, 22, 82, 55, 0, 0, 0, 0, 4, 20, 56, 61, 21, 0, 0, 36, 0, 0, 32, 219, 141, 87, 
    0, 85, 0, 0, 0, 0, 0, 1, 27, 29, 26, 31, 80, 95, 45, 35, 42, 33, 26, 16, 53, 49, 48, 13, 0, 39, 0, 0, 27, 172, 62, 106, 
    0, 34, 0, 0, 0, 0, 0, 0, 66, 100, 98, 24, 0, 33, 61, 82, 99, 104, 71, 42, 43, 13, 17, 57, 83, 62, 0, 0, 30, 102, 0, 84, 
    0, 15, 0, 0, 0, 0, 0, 0, 3, 98, 195, 70, 0, 9, 46, 53, 73, 99, 114, 111, 122, 65, 0, 5, 86, 123, 36, 0, 62, 114, 0, 103, 
    0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 221, 166, 3, 15, 45, 58, 65, 59, 66, 57, 87, 88, 30, 0, 8, 113, 52, 8, 108, 143, 0, 87, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 63, 150, 85, 9, 15, 67, 71, 70, 59, 59, 70, 81, 80, 18, 5, 52, 55, 0, 40, 104, 0, 122, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 120, 66, 39, 54, 61, 85, 78, 88, 97, 43, 44, 59, 74, 75, 67, 0, 0, 19, 0, 198, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 18, 53, 54, 60, 65, 59, 50, 90, 121, 60, 40, 74, 78, 142, 106, 28, 0, 0, 0, 224, 
    0, 0, 0, 0, 11, 27, 0, 0, 0, 0, 9, 0, 0, 0, 26, 69, 94, 59, 37, 76, 102, 52, 35, 69, 74, 119, 84, 30, 0, 0, 0, 223, 
    0, 55, 0, 0, 17, 40, 0, 0, 19, 0, 6, 28, 0, 0, 14, 63, 76, 88, 70, 67, 72, 53, 50, 86, 94, 92, 79, 5, 0, 0, 0, 209, 
    0, 83, 0, 0, 97, 88, 0, 0, 0, 0, 0, 0, 0, 0, 0, 55, 58, 71, 96, 88, 56, 67, 67, 74, 95, 95, 86, 0, 0, 0, 0, 206, 
    0, 37, 0, 60, 133, 146, 67, 0, 0, 9, 0, 0, 0, 0, 0, 44, 77, 56, 85, 100, 47, 60, 91, 74, 82, 80, 36, 0, 0, 0, 0, 209, 
    0, 0, 0, 0, 92, 142, 116, 9, 0, 2, 0, 0, 0, 7, 17, 43, 51, 11, 50, 94, 29, 64, 108, 89, 78, 81, 36, 0, 0, 0, 0, 195, 
    0, 0, 0, 0, 0, 69, 96, 62, 59, 37, 0, 0, 0, 0, 9, 38, 0, 0, 0, 78, 32, 48, 108, 119, 81, 104, 94, 0, 0, 0, 0, 158, 
    0, 0, 0, 0, 0, 0, 30, 63, 80, 80, 0, 0, 0, 0, 31, 96, 28, 0, 0, 38, 70, 54, 101, 105, 72, 115, 113, 0, 0, 0, 0, 161, 
    0, 46, 0, 0, 0, 0, 0, 9, 65, 86, 69, 11, 0, 0, 40, 106, 90, 0, 0, 15, 55, 57, 89, 87, 91, 127, 35, 0, 0, 0, 26, 237, 
    0, 79, 102, 0, 0, 0, 0, 0, 18, 91, 94, 60, 14, 1, 0, 1, 29, 0, 0, 19, 24, 30, 99, 97, 114, 131, 0, 0, 0, 0, 52, 289, 
    0, 62, 64, 37, 0, 0, 0, 0, 0, 11, 71, 67, 47, 40, 2, 0, 29, 0, 0, 0, 0, 0, 23, 69, 135, 130, 9, 32, 0, 0, 38, 317, 
    0, 35, 0, 0, 52, 0, 0, 0, 0, 0, 0, 10, 42, 69, 36, 50, 132, 129, 21, 0, 0, 0, 15, 27, 92, 115, 60, 39, 0, 0, 51, 320, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 113, 
    
    -- channel=69
    66, 40, 9, 7, 34, 40, 34, 39, 28, 0, 0, 39, 48, 36, 28, 46, 69, 69, 67, 73, 71, 44, 37, 89, 100, 24, 18, 49, 39, 47, 50, 0, 
    66, 5, 0, 0, 32, 23, 4, 2, 0, 0, 0, 35, 29, 0, 0, 14, 30, 0, 0, 1, 5, 0, 0, 54, 50, 0, 0, 8, 0, 2, 0, 0, 
    68, 0, 0, 2, 35, 6, 0, 2, 0, 0, 0, 25, 9, 0, 0, 14, 31, 0, 0, 0, 6, 0, 0, 60, 51, 0, 0, 35, 29, 11, 0, 0, 
    69, 10, 0, 1, 21, 0, 0, 2, 0, 0, 0, 6, 0, 0, 0, 19, 25, 0, 1, 15, 12, 0, 0, 70, 59, 0, 0, 49, 43, 6, 0, 0, 
    61, 1, 0, 6, 4, 0, 0, 0, 0, 0, 0, 7, 5, 7, 11, 23, 17, 0, 0, 0, 1, 0, 0, 68, 74, 0, 0, 33, 26, 6, 0, 0, 
    49, 0, 0, 0, 4, 0, 0, 0, 0, 0, 10, 41, 39, 34, 19, 0, 0, 13, 0, 0, 2, 16, 1, 71, 81, 0, 0, 17, 28, 1, 0, 0, 
    42, 0, 0, 5, 0, 2, 0, 0, 0, 0, 50, 61, 42, 23, 0, 0, 0, 19, 0, 0, 22, 36, 9, 65, 75, 2, 0, 19, 32, 0, 0, 0, 
    40, 0, 20, 59, 16, 0, 0, 0, 0, 1, 69, 50, 22, 0, 0, 0, 10, 27, 0, 0, 58, 46, 18, 50, 58, 0, 0, 16, 19, 0, 0, 0, 
    45, 0, 46, 82, 34, 0, 0, 0, 1, 48, 74, 31, 0, 0, 0, 5, 67, 43, 10, 15, 51, 47, 13, 39, 52, 0, 0, 11, 0, 0, 0, 0, 
    48, 0, 47, 70, 28, 0, 0, 0, 1, 62, 56, 20, 0, 0, 0, 47, 63, 29, 23, 40, 45, 14, 0, 21, 49, 8, 2, 10, 0, 0, 0, 0, 
    44, 0, 42, 65, 26, 2, 0, 0, 14, 37, 13, 3, 0, 1, 54, 73, 41, 10, 14, 27, 23, 0, 0, 32, 42, 0, 8, 10, 0, 0, 0, 0, 
    32, 0, 34, 53, 24, 21, 0, 0, 42, 37, 8, 7, 0, 4, 57, 73, 41, 22, 16, 8, 0, 0, 7, 66, 64, 0, 0, 14, 0, 0, 0, 0, 
    38, 0, 25, 37, 12, 21, 15, 13, 41, 39, 16, 14, 14, 10, 15, 0, 0, 7, 11, 16, 12, 14, 18, 41, 38, 0, 0, 16, 0, 0, 0, 0, 
    56, 0, 39, 39, 6, 23, 27, 4, 0, 0, 5, 21, 21, 28, 37, 13, 0, 0, 0, 18, 22, 33, 39, 32, 10, 0, 18, 25, 0, 0, 0, 0, 
    55, 0, 26, 36, 7, 23, 28, 4, 4, 0, 0, 0, 30, 28, 33, 45, 38, 18, 11, 9, 0, 14, 49, 48, 20, 0, 12, 24, 0, 0, 0, 0, 
    53, 0, 13, 28, 18, 23, 28, 0, 19, 45, 0, 0, 26, 29, 23, 19, 25, 41, 43, 39, 26, 14, 17, 40, 47, 7, 10, 14, 0, 0, 8, 0, 
    63, 4, 25, 31, 20, 17, 25, 0, 2, 24, 9, 10, 30, 38, 39, 26, 12, 9, 24, 41, 40, 43, 35, 22, 11, 7, 16, 1, 0, 0, 23, 0, 
    74, 24, 36, 28, 0, 0, 0, 0, 0, 6, 25, 37, 27, 28, 28, 26, 37, 27, 17, 10, 0, 4, 21, 30, 7, 0, 0, 0, 0, 0, 39, 0, 
    88, 29, 12, 0, 0, 0, 0, 10, 11, 0, 8, 28, 20, 19, 29, 21, 19, 35, 45, 26, 8, 21, 20, 11, 7, 0, 0, 0, 0, 5, 66, 0, 
    96, 8, 0, 0, 0, 0, 11, 7, 2, 5, 0, 0, 16, 46, 49, 41, 25, 18, 33, 23, 0, 13, 23, 6, 1, 0, 0, 0, 0, 30, 43, 0, 
    89, 0, 0, 6, 0, 0, 18, 11, 0, 0, 0, 0, 6, 43, 51, 26, 27, 23, 11, 7, 6, 16, 23, 9, 0, 0, 0, 20, 47, 52, 26, 0, 
    71, 0, 0, 29, 11, 0, 12, 32, 8, 10, 4, 18, 46, 48, 40, 30, 21, 19, 10, 0, 0, 16, 15, 6, 5, 0, 0, 23, 47, 31, 11, 0, 
    64, 0, 53, 52, 0, 0, 0, 27, 31, 12, 2, 8, 61, 58, 33, 23, 20, 16, 3, 4, 16, 16, 21, 23, 9, 5, 13, 39, 31, 3, 0, 0, 
    96, 46, 95, 85, 36, 9, 12, 25, 10, 0, 6, 18, 27, 42, 33, 18, 11, 18, 3, 0, 35, 38, 10, 6, 1, 0, 3, 33, 25, 0, 5, 0, 
    102, 49, 80, 69, 42, 24, 17, 34, 9, 0, 14, 54, 36, 13, 20, 2, 0, 24, 24, 11, 36, 32, 6, 0, 6, 0, 0, 10, 20, 6, 0, 0, 
    72, 0, 0, 25, 34, 29, 26, 18, 12, 2, 11, 25, 29, 17, 0, 0, 0, 17, 33, 26, 27, 17, 4, 2, 2, 0, 0, 12, 29, 0, 0, 0, 
    64, 0, 0, 0, 27, 29, 30, 33, 14, 6, 17, 6, 0, 0, 0, 0, 0, 9, 41, 23, 21, 20, 0, 4, 3, 0, 0, 40, 23, 0, 0, 0, 
    70, 0, 0, 0, 7, 32, 35, 39, 36, 16, 6, 18, 15, 1, 7, 11, 14, 38, 41, 20, 18, 25, 10, 0, 0, 0, 0, 24, 20, 41, 8, 0, 
    75, 0, 0, 0, 0, 26, 48, 45, 39, 34, 18, 15, 26, 16, 12, 14, 16, 40, 42, 16, 20, 14, 0, 0, 0, 0, 5, 7, 29, 74, 40, 0, 
    67, 0, 0, 4, 0, 10, 25, 47, 41, 38, 42, 37, 26, 14, 19, 13, 0, 0, 5, 4, 0, 0, 0, 0, 1, 1, 25, 25, 40, 69, 3, 0, 
    34, 0, 0, 11, 0, 0, 2, 24, 33, 18, 25, 43, 41, 24, 35, 52, 23, 0, 0, 0, 0, 0, 0, 33, 38, 34, 51, 59, 73, 66, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=70
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=71
    0, 3, 5, 7, 12, 9, 10, 9, 6, 0, 10, 10, 9, 12, 9, 11, 13, 13, 14, 16, 13, 10, 11, 16, 5, 5, 21, 6, 5, 14, 8, 0, 
    0, 0, 0, 6, 3, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 1, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 23, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 25, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 2, 4, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 12, 0, 0, 0, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 4, 4, 4, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 10, 7, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 11, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 3, 6, 0, 0, 9, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 1, 0, 0, 0, 0, 0, 0, 4, 11, 0, 0, 0, 0, 1, 18, 4, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 17, 9, 0, 0, 11, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 3, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 
    0, 0, 0, 0, 0, 0, 0, 13, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 
    0, 6, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 25, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 14, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 2, 1, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 0, 0, 0, 5, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 4, 5, 4, 8, 13, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 
    0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 5, 0, 0, 0, 0, 0, 
    0, 0, 16, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 12, 0, 0, 6, 0, 0, 7, 
    0, 0, 11, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=72
    9, 74, 74, 36, 15, 45, 67, 72, 79, 73, 17, 0, 37, 67, 63, 45, 58, 88, 99, 93, 102, 108, 78, 42, 94, 149, 69, 37, 59, 51, 60, 89, 
    0, 85, 97, 47, 33, 67, 76, 78, 90, 77, 23, 0, 33, 74, 66, 34, 49, 76, 74, 61, 81, 114, 79, 23, 75, 167, 83, 0, 40, 69, 77, 92, 
    8, 89, 105, 59, 52, 82, 88, 85, 99, 72, 17, 0, 26, 60, 53, 18, 39, 87, 78, 61, 80, 112, 77, 18, 72, 174, 99, 21, 67, 100, 94, 84, 
    14, 90, 118, 84, 71, 91, 90, 88, 104, 69, 11, 0, 14, 33, 44, 34, 48, 94, 95, 73, 74, 105, 76, 21, 74, 181, 141, 62, 89, 120, 104, 114, 
    3, 97, 99, 92, 77, 91, 89, 79, 99, 64, 4, 0, 17, 41, 66, 67, 63, 88, 101, 79, 44, 80, 84, 30, 79, 193, 169, 90, 98, 129, 134, 153, 
    0, 91, 52, 66, 66, 91, 94, 72, 83, 53, 0, 10, 52, 78, 94, 96, 66, 55, 99, 78, 9, 61, 98, 35, 86, 199, 180, 122, 113, 148, 143, 116, 
    0, 83, 29, 41, 78, 86, 93, 79, 67, 28, 0, 50, 86, 103, 115, 79, 22, 17, 91, 89, 18, 51, 97, 62, 90, 197, 189, 139, 131, 161, 122, 71, 
    6, 80, 44, 54, 113, 107, 83, 81, 68, 23, 19, 76, 102, 121, 98, 33, 5, 37, 76, 89, 52, 63, 112, 96, 97, 183, 184, 142, 141, 169, 118, 45, 
    21, 86, 49, 73, 145, 155, 99, 65, 65, 43, 49, 98, 127, 117, 61, 15, 33, 79, 78, 84, 88, 97, 134, 95, 102, 160, 175, 146, 153, 171, 104, 28, 
    27, 96, 37, 72, 151, 188, 146, 64, 36, 49, 72, 107, 125, 110, 66, 39, 61, 94, 113, 101, 102, 133, 129, 54, 90, 159, 167, 154, 160, 168, 89, 14, 
    31, 100, 29, 64, 144, 178, 195, 106, 25, 59, 88, 91, 108, 110, 94, 94, 103, 121, 127, 116, 109, 124, 111, 60, 96, 163, 158, 156, 163, 174, 86, 0, 
    22, 88, 21, 53, 121, 159, 195, 160, 94, 90, 99, 81, 92, 97, 87, 103, 131, 132, 112, 100, 101, 97, 116, 88, 99, 170, 154, 137, 164, 173, 78, 11, 
    10, 98, 34, 51, 105, 131, 172, 186, 143, 101, 100, 78, 74, 79, 64, 85, 105, 99, 94, 89, 97, 90, 102, 82, 98, 166, 149, 128, 167, 164, 85, 63, 
    23, 112, 58, 66, 108, 99, 145, 167, 138, 97, 76, 60, 71, 87, 83, 77, 79, 84, 80, 78, 87, 88, 92, 95, 106, 134, 147, 138, 159, 162, 95, 86, 
    20, 108, 68, 77, 110, 96, 120, 149, 123, 123, 100, 48, 46, 73, 84, 89, 101, 99, 81, 71, 83, 73, 82, 121, 127, 129, 133, 142, 165, 144, 46, 79, 
    6, 105, 69, 80, 115, 126, 118, 150, 119, 131, 155, 60, 25, 66, 82, 100, 103, 96, 104, 99, 108, 101, 88, 102, 135, 165, 126, 140, 169, 111, 16, 99, 
    2, 104, 94, 94, 129, 132, 125, 132, 109, 88, 165, 134, 56, 71, 96, 100, 95, 103, 108, 109, 112, 113, 96, 90, 130, 144, 141, 125, 154, 131, 33, 90, 
    5, 103, 117, 120, 133, 111, 114, 110, 113, 76, 100, 179, 118, 71, 93, 100, 109, 112, 98, 104, 112, 109, 117, 108, 100, 118, 134, 92, 109, 133, 50, 105, 
    10, 113, 132, 129, 116, 105, 79, 97, 106, 118, 61, 105, 147, 100, 92, 114, 120, 120, 126, 132, 125, 95, 102, 119, 108, 126, 87, 85, 77, 86, 91, 165, 
    19, 137, 121, 100, 109, 111, 57, 97, 93, 105, 94, 39, 95, 124, 112, 135, 129, 119, 127, 144, 134, 108, 103, 119, 112, 124, 111, 97, 73, 72, 117, 191, 
    26, 146, 85, 91, 114, 110, 70, 84, 101, 72, 125, 72, 36, 101, 132, 146, 148, 142, 121, 129, 136, 113, 97, 112, 108, 116, 135, 94, 96, 122, 125, 195, 
    20, 130, 73, 79, 110, 120, 85, 75, 125, 104, 105, 130, 58, 74, 135, 150, 152, 157, 138, 121, 113, 102, 96, 107, 110, 113, 122, 99, 122, 148, 145, 193, 
    6, 112, 87, 105, 146, 146, 105, 83, 123, 151, 100, 99, 95, 89, 113, 149, 150, 144, 156, 125, 101, 110, 104, 103, 112, 106, 108, 115, 128, 141, 158, 193, 
    3, 122, 135, 166, 188, 176, 144, 109, 120, 140, 119, 83, 92, 107, 104, 128, 144, 136, 148, 137, 102, 115, 120, 107, 104, 98, 98, 100, 122, 144, 154, 196, 
    11, 119, 110, 150, 199, 204, 185, 145, 134, 127, 115, 116, 105, 111, 116, 116, 120, 108, 127, 137, 107, 125, 137, 104, 89, 103, 95, 61, 107, 140, 149, 181, 
    0, 92, 65, 87, 153, 192, 195, 177, 154, 145, 114, 116, 121, 101, 111, 100, 73, 51, 89, 130, 129, 108, 130, 116, 103, 106, 94, 38, 83, 140, 119, 148, 
    0, 100, 56, 18, 60, 133, 173, 183, 180, 172, 137, 102, 108, 105, 102, 106, 76, 26, 59, 121, 127, 117, 130, 118, 110, 105, 73, 40, 85, 119, 98, 141, 
    0, 110, 70, 0, 0, 51, 124, 171, 193, 186, 168, 138, 116, 115, 113, 136, 131, 71, 62, 104, 111, 125, 126, 116, 108, 88, 47, 73, 58, 87, 146, 167, 
    5, 112, 87, 28, 0, 0, 62, 123, 175, 202, 193, 172, 153, 140, 130, 136, 134, 98, 65, 91, 105, 112, 131, 111, 91, 79, 62, 59, 29, 84, 168, 201, 
    8, 120, 72, 60, 24, 0, 1, 66, 128, 180, 203, 196, 182, 171, 146, 134, 135, 101, 58, 77, 89, 74, 77, 85, 113, 117, 87, 74, 88, 81, 155, 220, 
    4, 85, 28, 54, 77, 13, 0, 0, 75, 130, 163, 190, 197, 194, 171, 159, 176, 142, 85, 78, 56, 45, 70, 101, 153, 166, 137, 134, 139, 113, 162, 220, 
    0, 22, 3, 2, 36, 8, 0, 0, 4, 31, 42, 64, 83, 84, 70, 60, 79, 78, 34, 18, 23, 15, 26, 34, 54, 73, 66, 57, 54, 58, 70, 101, 
    
    -- channel=73
    120, 149, 141, 118, 122, 142, 156, 160, 156, 134, 106, 108, 133, 142, 139, 137, 140, 147, 144, 142, 152, 154, 143, 141, 167, 159, 109, 97, 110, 124, 139, 136, 
    99, 94, 85, 81, 98, 118, 110, 107, 100, 72, 65, 85, 84, 74, 67, 58, 59, 39, 12, 15, 41, 52, 55, 65, 68, 32, 17, 41, 49, 78, 94, 61, 
    110, 89, 75, 85, 100, 100, 95, 108, 95, 65, 63, 75, 53, 41, 40, 45, 62, 61, 51, 52, 62, 57, 58, 69, 59, 33, 52, 104, 115, 116, 90, 45, 
    113, 90, 85, 86, 92, 83, 88, 106, 86, 56, 53, 55, 38, 42, 60, 80, 76, 65, 76, 80, 65, 47, 59, 80, 68, 53, 89, 132, 119, 102, 92, 78, 
    90, 53, 62, 58, 70, 70, 86, 88, 67, 51, 59, 67, 78, 92, 103, 110, 90, 57, 52, 41, 23, 35, 67, 85, 71, 60, 89, 111, 91, 88, 94, 97, 
    80, 27, 3, 8, 57, 80, 91, 70, 50, 48, 78, 109, 126, 128, 111, 74, 43, 49, 63, 39, 21, 47, 78, 85, 76, 65, 73, 97, 96, 81, 53, 23, 
    84, 42, 28, 43, 72, 86, 85, 69, 48, 47, 97, 124, 114, 84, 50, 11, 0, 29, 75, 71, 75, 78, 71, 75, 71, 55, 63, 95, 99, 74, 14, 0, 
    98, 68, 85, 132, 129, 93, 66, 73, 76, 73, 108, 104, 67, 32, 2, 0, 56, 94, 72, 66, 115, 104, 67, 77, 56, 28, 46, 82, 85, 59, 10, 17, 
    113, 84, 99, 134, 136, 117, 69, 47, 74, 108, 125, 83, 40, 11, 0, 42, 120, 139, 91, 71, 105, 93, 47, 38, 38, 30, 45, 76, 76, 45, 12, 46, 
    110, 80, 87, 105, 97, 109, 99, 50, 28, 75, 93, 56, 45, 37, 53, 108, 121, 84, 75, 90, 78, 46, 4, 0, 17, 40, 58, 84, 82, 45, 23, 57, 
    105, 61, 74, 90, 83, 93, 110, 103, 67, 68, 48, 15, 18, 54, 131, 175, 129, 65, 51, 51, 24, 10, 16, 31, 52, 39, 61, 92, 80, 48, 37, 59, 
    85, 39, 61, 73, 63, 75, 104, 134, 144, 111, 45, 9, 2, 7, 50, 78, 69, 49, 27, 13, 2, 0, 22, 64, 60, 29, 51, 75, 66, 48, 51, 79, 
    92, 63, 89, 84, 54, 63, 79, 98, 110, 69, 16, 1, 0, 13, 13, 0, 0, 0, 0, 9, 22, 21, 31, 30, 7, 18, 64, 77, 63, 55, 79, 122, 
    105, 87, 110, 105, 69, 58, 63, 58, 27, 0, 0, 0, 0, 7, 35, 22, 0, 0, 0, 0, 0, 9, 34, 34, 9, 4, 53, 87, 68, 48, 72, 99, 
    94, 58, 77, 88, 78, 66, 71, 51, 37, 28, 0, 0, 0, 0, 0, 14, 31, 30, 8, 0, 0, 0, 7, 38, 49, 24, 45, 71, 51, 10, 21, 44, 
    89, 56, 76, 85, 93, 99, 93, 50, 17, 42, 48, 0, 0, 0, 0, 0, 0, 0, 25, 42, 48, 32, 2, 0, 30, 53, 53, 54, 48, 19, 34, 72, 
    95, 81, 104, 101, 85, 84, 70, 52, 5, 0, 28, 78, 58, 12, 7, 8, 0, 0, 0, 0, 0, 17, 29, 3, 0, 0, 27, 51, 53, 50, 70, 75, 
    104, 90, 111, 108, 73, 41, 35, 36, 30, 0, 0, 57, 77, 7, 0, 0, 8, 18, 0, 0, 0, 0, 0, 19, 5, 0, 0, 0, 24, 67, 112, 80, 
    117, 101, 85, 62, 43, 33, 42, 40, 59, 41, 0, 0, 21, 27, 21, 12, 3, 4, 20, 20, 0, 0, 0, 0, 4, 0, 0, 0, 16, 47, 119, 126, 
    123, 88, 54, 21, 29, 48, 57, 51, 36, 43, 26, 0, 0, 24, 50, 45, 28, 0, 1, 14, 0, 0, 2, 0, 0, 17, 49, 84, 87, 84, 111, 89, 
    116, 59, 25, 35, 72, 68, 73, 81, 46, 28, 66, 50, 0, 0, 40, 30, 24, 22, 0, 0, 0, 0, 0, 0, 0, 7, 51, 97, 118, 151, 124, 40, 
    99, 40, 26, 57, 73, 66, 80, 87, 99, 91, 68, 82, 76, 24, 16, 20, 11, 23, 16, 0, 0, 0, 0, 0, 0, 12, 39, 74, 110, 125, 89, 42, 
    90, 57, 111, 131, 87, 76, 82, 77, 88, 112, 67, 32, 65, 55, 0, 0, 2, 2, 8, 10, 0, 0, 0, 0, 0, 0, 24, 80, 107, 77, 60, 53, 
    121, 108, 147, 148, 104, 86, 96, 102, 72, 54, 74, 61, 35, 29, 0, 0, 0, 4, 13, 5, 13, 26, 3, 0, 0, 0, 0, 45, 72, 65, 77, 64, 
    97, 58, 46, 23, 34, 58, 77, 96, 84, 40, 59, 114, 80, 16, 0, 0, 0, 0, 7, 13, 13, 16, 0, 0, 0, 0, 0, 1, 38, 68, 67, 35, 
    76, 0, 0, 0, 0, 3, 39, 54, 60, 67, 59, 52, 35, 0, 0, 0, 0, 0, 0, 6, 16, 0, 0, 0, 0, 0, 0, 10, 51, 57, 39, 7, 
    83, 21, 0, 0, 0, 0, 0, 36, 49, 56, 70, 46, 2, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 47, 86, 50, 24, 25, 
    95, 49, 9, 0, 0, 0, 0, 0, 39, 44, 42, 57, 48, 25, 21, 64, 108, 85, 31, 0, 0, 0, 1, 0, 0, 0, 4, 67, 76, 68, 99, 79, 
    104, 58, 45, 46, 0, 0, 0, 0, 0, 39, 57, 54, 56, 48, 33, 34, 43, 43, 15, 0, 0, 0, 0, 0, 0, 0, 49, 76, 30, 53, 97, 63, 
    87, 30, 27, 69, 68, 0, 0, 0, 0, 0, 37, 64, 66, 55, 50, 49, 17, 0, 0, 0, 0, 0, 0, 0, 48, 97, 132, 122, 96, 87, 21, 0, 
    52, 0, 0, 52, 73, 46, 0, 0, 0, 0, 0, 10, 54, 59, 56, 75, 86, 58, 11, 0, 0, 0, 10, 64, 111, 137, 143, 140, 140, 93, 35, 21, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=74
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 7, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 23, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 38, 0, 0, 0, 20, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 1, 5, 32, 0, 0, 
    0, 0, 0, 0, 7, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 8, 14, 24, 0, 0, 
    7, 0, 0, 12, 19, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 19, 15, 0, 0, 
    17, 0, 0, 11, 22, 26, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 19, 3, 0, 0, 
    15, 0, 0, 3, 12, 27, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 23, 0, 0, 0, 
    16, 0, 0, 0, 0, 11, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 19, 0, 0, 0, 
    16, 0, 0, 0, 0, 0, 25, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 
    15, 0, 0, 0, 0, 0, 14, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 14, 0, 0, 0, 
    11, 0, 0, 0, 2, 0, 8, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 16, 0, 0, 4, 
    4, 0, 0, 0, 3, 0, 12, 8, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 11, 
    5, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 
    14, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 
    27, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 
    38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 39, 
    38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 13, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 10, 30, 
    28, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 0, 6, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 14, 0, 21, 
    24, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 22, 
    14, 0, 2, 18, 0, 0, 0, 0, 0, 0, 0, 5, 1, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=75
    105, 188, 193, 152, 132, 160, 190, 190, 189, 173, 127, 105, 159, 197, 189, 179, 199, 240, 253, 248, 243, 241, 213, 190, 240, 291, 224, 153, 174, 172, 174, 182, 
    54, 156, 178, 152, 134, 158, 166, 152, 155, 157, 111, 88, 133, 155, 145, 118, 121, 154, 144, 126, 146, 180, 158, 102, 153, 248, 167, 67, 115, 147, 145, 160, 
    57, 166, 177, 168, 146, 172, 164, 155, 166, 159, 101, 79, 102, 115, 118, 93, 113, 165, 164, 142, 156, 186, 156, 93, 149, 256, 198, 121, 169, 187, 167, 148, 
    55, 165, 190, 193, 156, 171, 154, 152, 168, 156, 88, 65, 71, 93, 118, 125, 144, 180, 182, 159, 154, 181, 157, 94, 154, 275, 253, 176, 180, 191, 188, 186, 
    51, 153, 169, 163, 154, 150, 141, 138, 153, 145, 81, 75, 99, 140, 170, 161, 145, 153, 159, 140, 114, 144, 167, 110, 150, 274, 260, 180, 172, 199, 235, 237, 
    38, 116, 115, 97, 134, 144, 143, 126, 132, 132, 96, 129, 187, 212, 205, 181, 131, 104, 139, 143, 80, 129, 187, 120, 139, 259, 256, 196, 192, 216, 209, 174, 
    40, 121, 104, 100, 156, 151, 146, 131, 129, 113, 110, 184, 236, 231, 206, 143, 69, 67, 134, 169, 109, 138, 200, 146, 147, 237, 253, 210, 197, 193, 154, 104, 
    56, 163, 140, 152, 206, 192, 157, 134, 154, 132, 135, 205, 233, 220, 181, 111, 86, 116, 168, 166, 143, 183, 233, 193, 164, 212, 222, 198, 178, 189, 158, 87, 
    75, 187, 141, 163, 232, 230, 190, 136, 156, 158, 168, 221, 233, 207, 157, 122, 159, 195, 200, 197, 193, 224, 245, 203, 159, 204, 203, 186, 174, 196, 149, 74, 
    80, 179, 109, 121, 214, 251, 220, 154, 126, 132, 178, 203, 200, 204, 182, 164, 185, 221, 232, 226, 217, 226, 217, 149, 143, 215, 202, 183, 182, 205, 145, 70, 
    76, 174, 83, 99, 180, 240, 258, 205, 131, 135, 174, 158, 168, 203, 211, 221, 233, 244, 238, 213, 198, 197, 198, 159, 186, 229, 190, 176, 201, 227, 154, 65, 
    63, 150, 67, 81, 147, 196, 261, 272, 225, 207, 193, 153, 149, 160, 151, 170, 213, 221, 203, 181, 162, 180, 207, 184, 197, 228, 190, 164, 199, 240, 157, 84, 
    59, 165, 98, 91, 133, 155, 223, 277, 250, 219, 196, 165, 140, 117, 101, 109, 129, 139, 148, 156, 155, 169, 179, 159, 171, 209, 193, 177, 207, 242, 183, 151, 
    83, 200, 135, 129, 142, 138, 166, 215, 200, 169, 134, 118, 139, 158, 151, 139, 127, 124, 124, 112, 122, 129, 146, 154, 167, 188, 189, 196, 211, 237, 181, 163, 
    66, 180, 132, 132, 152, 141, 148, 179, 182, 172, 165, 99, 82, 132, 150, 155, 172, 171, 140, 112, 109, 98, 106, 149, 179, 189, 183, 179, 212, 196, 99, 123, 
    53, 164, 139, 136, 172, 172, 172, 181, 183, 175, 196, 133, 59, 99, 135, 151, 154, 153, 166, 177, 171, 152, 122, 105, 153, 203, 195, 164, 196, 169, 83, 154, 
    58, 174, 172, 172, 182, 176, 158, 162, 124, 127, 181, 200, 143, 122, 131, 132, 130, 141, 151, 154, 170, 157, 128, 108, 120, 153, 159, 169, 192, 212, 128, 154, 
    57, 179, 187, 196, 178, 148, 119, 150, 123, 100, 132, 184, 193, 119, 99, 128, 134, 143, 133, 122, 136, 150, 149, 126, 95, 117, 120, 106, 158, 197, 137, 177, 
    57, 177, 190, 183, 155, 136, 116, 133, 159, 130, 94, 87, 147, 142, 108, 133, 150, 150, 155, 172, 157, 126, 132, 139, 133, 116, 105, 80, 130, 159, 164, 254, 
    58, 179, 155, 131, 148, 155, 126, 128, 158, 132, 91, 66, 69, 128, 155, 146, 149, 142, 135, 149, 156, 134, 133, 146, 142, 147, 155, 147, 145, 159, 186, 264, 
    51, 169, 132, 125, 183, 181, 135, 134, 143, 148, 132, 114, 69, 83, 141, 163, 153, 144, 136, 127, 138, 133, 123, 129, 131, 159, 168, 165, 174, 195, 204, 250, 
    38, 166, 141, 140, 196, 204, 150, 149, 181, 189, 194, 167, 125, 104, 131, 153, 157, 147, 137, 130, 119, 109, 122, 136, 146, 161, 159, 158, 176, 213, 212, 251, 
    37, 180, 169, 219, 275, 252, 194, 153, 190, 203, 187, 158, 130, 129, 132, 141, 141, 138, 144, 138, 124, 133, 139, 142, 164, 171, 173, 167, 172, 203, 214, 263, 
    59, 223, 249, 295, 330, 324, 272, 203, 180, 190, 154, 149, 138, 127, 126, 129, 135, 123, 142, 156, 128, 135, 158, 140, 146, 155, 163, 142, 162, 211, 223, 276, 
    63, 180, 159, 203, 279, 342, 340, 276, 222, 202, 172, 156, 167, 153, 124, 125, 109, 90, 118, 146, 132, 140, 152, 131, 126, 146, 146, 106, 140, 213, 224, 254, 
    12, 98, 67, 83, 182, 279, 321, 319, 289, 247, 202, 164, 140, 135, 109, 90, 46, 21, 73, 135, 132, 127, 125, 143, 149, 153, 138, 97, 134, 211, 191, 205, 
    21, 123, 87, 28, 64, 171, 254, 294, 328, 314, 241, 184, 155, 136, 126, 120, 97, 54, 64, 125, 125, 125, 152, 146, 128, 139, 123, 98, 160, 196, 183, 218, 
    46, 173, 131, 32, 4, 65, 179, 251, 303, 333, 316, 268, 235, 214, 205, 215, 212, 155, 106, 104, 122, 127, 148, 141, 120, 108, 108, 125, 159, 174, 254, 298, 
    56, 199, 185, 109, 52, 37, 102, 188, 254, 306, 340, 331, 298, 282, 261, 244, 225, 152, 102, 97, 100, 123, 148, 130, 124, 142, 128, 125, 146, 191, 285, 311, 
    61, 195, 185, 162, 131, 58, 57, 108, 183, 246, 300, 329, 330, 316, 278, 248, 235, 170, 89, 76, 81, 55, 67, 104, 175, 226, 190, 202, 210, 207, 254, 283, 
    50, 146, 117, 160, 197, 109, 45, 50, 111, 181, 220, 256, 299, 323, 308, 302, 311, 270, 173, 97, 64, 48, 100, 167, 246, 280, 264, 272, 248, 230, 248, 293, 
    0, 47, 35, 53, 78, 54, 7, 0, 0, 0, 0, 0, 1, 24, 25, 27, 54, 61, 26, 10, 13, 11, 11, 0, 5, 18, 20, 11, 5, 0, 27, 82, 
    
    -- channel=76
    41, 81, 53, 13, 10, 35, 56, 68, 66, 35, 0, 0, 44, 66, 59, 63, 95, 132, 146, 146, 148, 126, 90, 104, 172, 154, 67, 64, 81, 66, 71, 52, 
    55, 93, 59, 19, 36, 67, 64, 61, 52, 14, 0, 0, 63, 73, 50, 48, 86, 103, 90, 89, 105, 96, 58, 86, 175, 140, 17, 19, 46, 53, 68, 37, 
    68, 106, 80, 46, 71, 86, 69, 71, 57, 10, 0, 7, 49, 51, 27, 28, 82, 93, 68, 69, 100, 98, 55, 90, 188, 150, 28, 43, 89, 102, 80, 18, 
    85, 116, 101, 74, 93, 89, 73, 81, 60, 3, 0, 0, 12, 22, 21, 37, 94, 116, 100, 96, 109, 96, 58, 104, 202, 182, 85, 107, 143, 132, 90, 24, 
    87, 117, 125, 95, 93, 78, 74, 78, 54, 0, 0, 0, 1, 31, 57, 77, 97, 98, 88, 77, 79, 86, 70, 120, 223, 222, 139, 136, 147, 146, 129, 81, 
    66, 78, 75, 63, 79, 73, 74, 57, 35, 0, 0, 15, 61, 91, 105, 91, 73, 80, 81, 40, 29, 82, 93, 134, 237, 245, 166, 149, 160, 171, 143, 80, 
    46, 49, 20, 46, 79, 89, 84, 45, 16, 0, 15, 82, 124, 131, 107, 46, 6, 40, 90, 46, 28, 102, 115, 143, 246, 264, 186, 177, 186, 176, 90, 0, 
    38, 46, 36, 102, 127, 101, 83, 57, 20, 0, 59, 130, 142, 121, 61, 0, 0, 43, 93, 73, 83, 133, 138, 160, 235, 251, 194, 194, 191, 159, 40, 0, 
    51, 62, 73, 163, 196, 146, 83, 66, 60, 51, 116, 152, 138, 94, 18, 0, 61, 118, 109, 100, 142, 178, 169, 178, 217, 229, 189, 196, 182, 131, 7, 0, 
    69, 69, 80, 166, 215, 190, 107, 53, 58, 99, 160, 170, 147, 80, 14, 45, 125, 155, 137, 154, 183, 184, 148, 138, 199, 222, 196, 197, 177, 107, 0, 0, 
    78, 64, 68, 158, 207, 215, 155, 71, 45, 97, 146, 156, 152, 117, 111, 146, 167, 157, 161, 177, 176, 165, 119, 111, 204, 218, 195, 197, 178, 103, 0, 0, 
    79, 49, 50, 138, 189, 215, 203, 143, 111, 140, 145, 147, 147, 129, 165, 217, 214, 188, 177, 167, 152, 143, 130, 159, 240, 211, 174, 191, 184, 109, 0, 0, 
    75, 40, 45, 114, 155, 190, 220, 213, 204, 193, 167, 167, 160, 119, 124, 152, 169, 169, 167, 172, 169, 158, 155, 169, 216, 198, 161, 177, 184, 119, 19, 2, 
    94, 83, 83, 125, 142, 166, 207, 225, 212, 177, 161, 167, 166, 158, 162, 153, 143, 138, 150, 170, 181, 182, 196, 185, 191, 182, 170, 188, 192, 128, 62, 59, 
    98, 96, 95, 133, 143, 148, 191, 214, 215, 182, 137, 125, 157, 178, 192, 200, 195, 177, 158, 150, 150, 160, 207, 229, 220, 177, 167, 186, 176, 101, 48, 49, 
    86, 85, 87, 126, 155, 160, 192, 204, 232, 257, 187, 96, 125, 171, 187, 201, 219, 220, 206, 197, 185, 165, 183, 228, 258, 219, 180, 172, 149, 57, 15, 50, 
    85, 107, 113, 141, 172, 180, 189, 185, 189, 239, 232, 152, 151, 192, 212, 212, 200, 200, 222, 239, 242, 222, 199, 193, 231, 243, 194, 159, 138, 62, 43, 90, 
    93, 136, 158, 165, 161, 143, 143, 155, 156, 183, 233, 235, 212, 194, 207, 219, 223, 218, 207, 204, 203, 201, 210, 204, 197, 182, 153, 129, 125, 92, 76, 82, 
    110, 157, 179, 167, 146, 103, 110, 131, 157, 156, 177, 233, 233, 193, 199, 213, 231, 246, 244, 244, 224, 203, 206, 204, 194, 148, 99, 58, 79, 99, 132, 133, 
    129, 167, 158, 125, 107, 85, 96, 121, 148, 154, 129, 155, 205, 226, 241, 250, 247, 235, 250, 255, 220, 197, 208, 205, 188, 158, 99, 81, 85, 102, 164, 168, 
    136, 145, 112, 101, 112, 94, 90, 123, 108, 120, 132, 116, 145, 217, 260, 268, 261, 246, 241, 239, 220, 207, 210, 202, 179, 162, 121, 126, 136, 158, 185, 138, 
    127, 117, 82, 118, 144, 107, 96, 137, 132, 125, 155, 153, 161, 215, 263, 274, 262, 259, 235, 209, 198, 198, 195, 193, 178, 160, 127, 124, 162, 203, 187, 120, 
    110, 120, 125, 173, 170, 131, 104, 127, 175, 168, 150, 158, 197, 234, 257, 268, 258, 254, 236, 212, 197, 203, 209, 211, 192, 173, 148, 142, 174, 186, 162, 115, 
    122, 179, 246, 300, 264, 200, 146, 134, 161, 169, 137, 144, 193, 241, 246, 256, 243, 235, 232, 213, 213, 232, 218, 206, 189, 162, 146, 149, 170, 166, 166, 124, 
    144, 221, 285, 326, 312, 270, 215, 186, 168, 145, 146, 181, 215, 234, 235, 237, 215, 217, 238, 222, 220, 253, 231, 197, 176, 149, 115, 102, 135, 161, 167, 115, 
    108, 144, 163, 221, 287, 301, 270, 228, 200, 161, 151, 188, 217, 228, 207, 175, 132, 154, 216, 235, 228, 242, 222, 193, 174, 156, 97, 55, 116, 152, 138, 75, 
    83, 98, 65, 100, 197, 265, 284, 271, 237, 203, 170, 155, 152, 170, 167, 116, 68, 103, 194, 234, 231, 224, 213, 202, 181, 132, 59, 47, 120, 130, 105, 56, 
    82, 103, 31, 5, 73, 173, 249, 290, 288, 249, 204, 181, 166, 163, 170, 159, 136, 145, 201, 225, 222, 228, 225, 180, 142, 78, 32, 62, 122, 138, 140, 91, 
    90, 113, 37, 0, 0, 87, 191, 269, 308, 295, 255, 224, 208, 195, 183, 190, 187, 181, 201, 204, 201, 220, 211, 163, 107, 45, 36, 76, 93, 171, 244, 144, 
    92, 106, 54, 38, 11, 29, 106, 207, 278, 311, 311, 283, 255, 231, 202, 191, 159, 134, 150, 169, 167, 172, 158, 137, 127, 98, 91, 107, 111, 206, 245, 127, 
    68, 56, 22, 58, 47, 12, 30, 107, 196, 253, 288, 308, 303, 275, 252, 263, 237, 163, 113, 104, 90, 85, 106, 153, 205, 202, 194, 202, 224, 254, 231, 124, 
    0, 0, 0, 21, 20, 0, 0, 5, 63, 103, 123, 153, 177, 173, 161, 183, 192, 143, 79, 43, 17, 36, 80, 121, 151, 138, 126, 129, 142, 139, 138, 79, 
    
    -- channel=77
    81, 50, 0, 0, 18, 32, 26, 37, 26, 0, 0, 19, 44, 32, 25, 52, 89, 93, 91, 98, 96, 58, 40, 118, 157, 41, 4, 53, 42, 43, 56, 0, 
    116, 58, 0, 0, 44, 43, 26, 30, 2, 0, 0, 33, 55, 29, 6, 45, 80, 56, 38, 63, 74, 21, 9, 128, 171, 0, 0, 33, 34, 36, 35, 0, 
    128, 66, 16, 21, 65, 40, 27, 38, 0, 0, 0, 26, 39, 13, 0, 39, 86, 45, 22, 53, 74, 19, 12, 141, 184, 5, 0, 65, 81, 64, 20, 0, 
    140, 88, 44, 36, 64, 35, 38, 48, 0, 0, 0, 2, 10, 6, 4, 46, 86, 63, 48, 68, 79, 23, 21, 158, 203, 55, 8, 106, 121, 75, 29, 0, 
    139, 88, 67, 53, 49, 36, 43, 46, 0, 0, 0, 0, 11, 25, 35, 59, 74, 55, 36, 30, 58, 44, 35, 164, 236, 110, 49, 111, 118, 91, 65, 0, 
    120, 38, 32, 42, 51, 44, 34, 25, 0, 0, 0, 40, 54, 62, 57, 26, 29, 68, 36, 0, 43, 73, 47, 176, 261, 142, 68, 104, 129, 108, 51, 0, 
    93, 0, 7, 51, 51, 60, 39, 7, 0, 0, 54, 86, 79, 68, 12, 0, 0, 71, 49, 0, 54, 104, 70, 171, 260, 169, 94, 126, 152, 92, 0, 0, 
    77, 0, 38, 115, 86, 49, 36, 23, 0, 0, 97, 98, 73, 23, 0, 0, 12, 70, 44, 31, 107, 123, 91, 149, 228, 164, 118, 147, 154, 50, 0, 0, 
    83, 1, 85, 178, 137, 62, 20, 33, 23, 63, 124, 98, 48, 0, 0, 0, 90, 89, 66, 81, 130, 134, 90, 136, 203, 157, 125, 151, 133, 4, 0, 0, 
    95, 8, 107, 193, 166, 88, 19, 6, 45, 115, 138, 112, 65, 0, 0, 63, 119, 99, 86, 117, 140, 109, 42, 119, 197, 151, 135, 151, 113, 0, 0, 0, 
    104, 0, 104, 191, 175, 135, 43, 0, 54, 106, 107, 117, 96, 60, 99, 138, 124, 95, 93, 111, 123, 84, 38, 125, 190, 134, 139, 156, 108, 0, 0, 0, 
    99, 0, 88, 170, 168, 169, 103, 56, 91, 106, 97, 127, 112, 98, 161, 197, 158, 122, 116, 116, 108, 84, 74, 160, 210, 124, 119, 159, 114, 0, 0, 0, 
    105, 0, 71, 138, 143, 166, 158, 129, 141, 140, 127, 142, 134, 114, 135, 141, 132, 131, 138, 150, 137, 130, 122, 157, 183, 117, 110, 150, 105, 0, 0, 0, 
    128, 21, 89, 131, 119, 155, 180, 161, 143, 130, 135, 156, 151, 144, 154, 142, 128, 124, 138, 163, 166, 178, 186, 176, 156, 116, 126, 150, 107, 9, 22, 0, 
    132, 36, 88, 129, 110, 144, 176, 170, 175, 146, 86, 111, 168, 170, 175, 189, 181, 154, 145, 149, 143, 167, 221, 224, 182, 133, 126, 148, 79, 0, 34, 0, 
    128, 36, 79, 122, 125, 141, 171, 159, 204, 222, 108, 74, 162, 184, 185, 188, 194, 202, 193, 187, 168, 160, 188, 234, 244, 167, 134, 132, 47, 0, 43, 0, 
    137, 69, 95, 124, 136, 138, 162, 141, 177, 231, 166, 117, 165, 202, 213, 202, 190, 187, 201, 218, 212, 201, 197, 209, 220, 192, 156, 118, 46, 0, 58, 8, 
    154, 110, 129, 134, 105, 101, 116, 122, 134, 189, 223, 201, 180, 198, 212, 211, 220, 207, 202, 199, 185, 179, 188, 201, 191, 150, 95, 104, 70, 16, 86, 0, 
    179, 137, 134, 111, 86, 63, 90, 117, 131, 131, 194, 237, 201, 187, 211, 217, 219, 229, 237, 220, 187, 193, 196, 183, 173, 105, 53, 45, 47, 61, 142, 0, 
    201, 126, 100, 84, 60, 32, 89, 104, 113, 117, 126, 171, 210, 228, 243, 245, 232, 227, 246, 227, 184, 189, 202, 177, 161, 102, 60, 52, 59, 107, 154, 0, 
    203, 73, 68, 90, 59, 31, 86, 100, 71, 100, 98, 112, 181, 245, 267, 247, 239, 235, 229, 216, 192, 194, 202, 179, 153, 117, 77, 95, 128, 150, 146, 0, 
    184, 38, 62, 113, 90, 40, 73, 124, 90, 99, 107, 116, 189, 252, 266, 257, 244, 234, 216, 189, 181, 193, 192, 174, 156, 126, 81, 109, 160, 152, 121, 0, 
    166, 71, 139, 163, 95, 48, 54, 114, 138, 106, 107, 129, 211, 253, 259, 251, 239, 234, 203, 186, 195, 195, 198, 197, 163, 130, 105, 132, 150, 121, 90, 0, 
    199, 165, 246, 247, 167, 90, 67, 101, 123, 97, 100, 145, 198, 240, 250, 244, 221, 227, 207, 182, 218, 231, 196, 184, 152, 115, 106, 133, 132, 100, 98, 0, 
    220, 207, 282, 285, 223, 152, 102, 115, 104, 78, 114, 181, 214, 216, 229, 212, 192, 224, 230, 199, 232, 242, 198, 168, 149, 109, 63, 92, 112, 100, 88, 0, 
    185, 123, 162, 226, 244, 206, 161, 124, 103, 84, 113, 160, 195, 210, 180, 131, 121, 196, 239, 224, 227, 231, 198, 166, 149, 102, 26, 60, 112, 78, 56, 0, 
    153, 47, 35, 126, 209, 223, 200, 174, 129, 95, 103, 118, 118, 141, 126, 67, 55, 152, 238, 230, 218, 222, 181, 170, 151, 61, 0, 76, 97, 48, 46, 0, 
    150, 26, 0, 14, 119, 192, 213, 218, 190, 133, 96, 101, 108, 106, 113, 100, 92, 160, 227, 222, 216, 220, 194, 146, 87, 8, 21, 66, 86, 118, 80, 0, 
    155, 31, 0, 0, 24, 131, 205, 239, 233, 191, 139, 111, 113, 106, 107, 117, 115, 160, 213, 204, 209, 213, 164, 117, 51, 0, 31, 47, 100, 187, 148, 0, 
    143, 9, 0, 0, 0, 58, 138, 213, 240, 236, 211, 177, 148, 119, 118, 118, 81, 80, 145, 167, 153, 161, 136, 119, 83, 49, 69, 77, 117, 204, 140, 0, 
    95, 0, 7, 28, 0, 0, 54, 138, 196, 207, 219, 229, 211, 164, 162, 187, 142, 77, 74, 79, 78, 98, 116, 156, 158, 132, 142, 156, 183, 211, 135, 0, 
    3, 0, 0, 0, 0, 0, 0, 25, 46, 65, 89, 108, 109, 94, 100, 126, 103, 49, 33, 10, 0, 31, 73, 117, 117, 89, 82, 98, 101, 96, 71, 0, 
    
    -- channel=78
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 15, 19, 17, 20, 9, 0, 0, 29, 22, 0, 0, 15, 0, 0, 0, 0, 
    63, 42, 5, 9, 28, 32, 37, 35, 17, 0, 0, 38, 50, 34, 36, 64, 83, 88, 95, 102, 88, 50, 47, 109, 119, 34, 33, 63, 47, 38, 39, 0, 
    70, 59, 17, 28, 50, 49, 41, 39, 13, 0, 1, 46, 61, 47, 37, 68, 83, 62, 62, 83, 86, 46, 43, 118, 133, 33, 10, 39, 43, 44, 35, 0, 
    79, 64, 29, 47, 63, 55, 45, 45, 9, 0, 7, 43, 49, 44, 24, 53, 86, 66, 52, 74, 88, 47, 48, 120, 141, 45, 16, 58, 75, 60, 29, 0, 
    94, 77, 68, 61, 69, 53, 47, 54, 9, 0, 3, 26, 27, 29, 29, 51, 80, 79, 64, 73, 99, 57, 49, 126, 152, 79, 55, 84, 100, 71, 37, 0, 
    93, 77, 97, 78, 63, 49, 40, 51, 13, 0, 4, 22, 32, 44, 49, 58, 78, 79, 43, 44, 89, 70, 57, 134, 166, 109, 82, 87, 102, 80, 73, 2, 
    79, 47, 66, 68, 59, 57, 33, 30, 9, 0, 30, 54, 74, 78, 63, 55, 64, 84, 41, 3, 65, 87, 76, 135, 185, 130, 96, 93, 107, 81, 62, 2, 
    60, 24, 40, 60, 48, 53, 48, 21, 0, 14, 69, 95, 101, 83, 51, 28, 31, 61, 62, 21, 55, 100, 93, 137, 187, 150, 112, 110, 116, 62, 15, 0, 
    49, 22, 67, 92, 69, 33, 46, 48, 6, 32, 91, 103, 94, 64, 25, 19, 43, 59, 62, 62, 84, 114, 115, 153, 170, 150, 123, 117, 112, 42, 0, 0, 
    55, 29, 94, 130, 110, 49, 17, 49, 64, 82, 109, 107, 78, 26, 5, 40, 91, 91, 76, 95, 126, 127, 122, 164, 166, 143, 124, 114, 101, 16, 0, 0, 
    56, 33, 99, 141, 134, 90, 15, 14, 75, 110, 119, 116, 81, 36, 21, 58, 97, 103, 109, 119, 139, 125, 93, 135, 164, 140, 127, 117, 90, 0, 0, 0, 
    63, 33, 95, 141, 147, 126, 60, 10, 52, 97, 100, 103, 92, 90, 114, 118, 110, 112, 119, 119, 120, 112, 86, 135, 166, 131, 133, 132, 86, 0, 0, 0, 
    60, 19, 75, 122, 138, 149, 108, 68, 82, 105, 94, 105, 108, 104, 134, 149, 143, 133, 117, 112, 108, 105, 104, 150, 173, 129, 120, 131, 90, 10, 0, 0, 
    62, 27, 62, 99, 112, 151, 141, 121, 115, 122, 125, 128, 123, 111, 109, 116, 122, 123, 125, 130, 125, 124, 119, 134, 153, 140, 117, 126, 94, 25, 21, 0, 
    83, 52, 79, 98, 96, 129, 151, 131, 115, 93, 111, 147, 144, 137, 135, 121, 108, 107, 117, 130, 127, 146, 148, 134, 128, 124, 137, 126, 88, 48, 70, 0, 
    89, 56, 83, 101, 91, 106, 142, 129, 142, 117, 60, 109, 145, 141, 144, 148, 150, 135, 114, 115, 106, 118, 159, 174, 139, 106, 133, 130, 68, 33, 67, 0, 
    85, 59, 72, 101, 102, 117, 132, 133, 149, 179, 85, 48, 115, 142, 143, 148, 152, 159, 159, 153, 145, 131, 135, 168, 174, 147, 116, 131, 59, 0, 68, 0, 
    87, 82, 82, 97, 105, 121, 126, 126, 121, 165, 166, 81, 100, 151, 156, 155, 143, 145, 158, 162, 158, 162, 143, 146, 162, 150, 137, 133, 85, 14, 63, 0, 
    95, 98, 101, 113, 96, 93, 116, 111, 111, 110, 184, 175, 108, 130, 150, 148, 161, 156, 146, 146, 145, 158, 157, 145, 136, 109, 112, 100, 96, 72, 64, 0, 
    108, 104, 110, 111, 85, 69, 101, 101, 124, 106, 111, 196, 164, 126, 149, 148, 153, 170, 172, 152, 140, 148, 152, 141, 135, 92, 60, 57, 66, 86, 111, 0, 
    117, 95, 101, 85, 72, 55, 83, 94, 94, 123, 73, 106, 180, 168, 159, 164, 155, 153, 180, 168, 140, 147, 159, 141, 131, 101, 71, 68, 59, 84, 129, 3, 
    121, 71, 80, 100, 79, 52, 80, 95, 62, 89, 105, 62, 124, 183, 181, 168, 169, 156, 153, 162, 154, 144, 151, 141, 125, 112, 90, 87, 99, 119, 120, 0, 
    113, 63, 68, 94, 87, 61, 75, 107, 94, 74, 107, 113, 114, 164, 196, 177, 174, 169, 144, 139, 144, 143, 148, 143, 137, 128, 98, 98, 131, 133, 112, 0, 
    102, 80, 108, 124, 106, 85, 69, 99, 119, 100, 82, 112, 150, 159, 186, 185, 173, 168, 148, 132, 148, 139, 144, 151, 152, 134, 120, 138, 133, 121, 109, 0, 
    128, 149, 201, 206, 165, 122, 98, 105, 105, 99, 99, 99, 137, 163, 172, 182, 177, 176, 154, 133, 157, 157, 139, 148, 146, 113, 114, 157, 133, 115, 113, 0, 
    141, 161, 219, 248, 223, 182, 141, 131, 114, 87, 115, 144, 144, 159, 166, 165, 172, 186, 169, 146, 155, 177, 147, 128, 128, 109, 84, 132, 128, 112, 117, 0, 
    114, 95, 141, 219, 248, 226, 193, 153, 131, 113, 111, 139, 151, 149, 141, 107, 103, 154, 169, 164, 162, 155, 149, 137, 123, 101, 79, 99, 113, 106, 91, 0, 
    94, 55, 54, 130, 218, 231, 220, 195, 159, 136, 123, 120, 129, 132, 120, 79, 55, 104, 161, 168, 168, 158, 140, 138, 124, 80, 68, 87, 119, 88, 52, 0, 
    95, 46, 15, 29, 125, 209, 223, 227, 202, 158, 136, 131, 130, 127, 130, 123, 102, 108, 149, 159, 162, 166, 144, 126, 94, 52, 61, 86, 112, 130, 97, 0, 
    102, 52, 42, 2, 36, 142, 216, 234, 234, 211, 172, 144, 140, 135, 135, 130, 113, 123, 149, 149, 165, 173, 153, 122, 66, 34, 54, 55, 89, 175, 145, 0, 
    97, 58, 68, 37, 8, 60, 156, 222, 234, 241, 226, 191, 165, 147, 142, 130, 90, 79, 118, 129, 133, 128, 117, 115, 83, 63, 68, 75, 113, 166, 136, 0, 
    81, 35, 61, 79, 40, 28, 72, 155, 206, 224, 244, 253, 243, 217, 211, 222, 193, 132, 112, 107, 91, 110, 137, 172, 178, 159, 154, 168, 188, 194, 176, 45, 
    
    -- channel=79
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    47, 16, 0, 0, 4, 0, 0, 0, 0, 0, 0, 6, 8, 0, 0, 10, 21, 20, 21, 25, 23, 4, 0, 35, 53, 1, 0, 26, 23, 12, 9, 0, 
    46, 18, 0, 0, 8, 0, 0, 0, 0, 0, 0, 10, 16, 8, 0, 15, 28, 10, 12, 25, 24, 0, 0, 44, 65, 4, 0, 22, 21, 3, 0, 0, 
    46, 18, 10, 0, 9, 0, 0, 0, 0, 0, 0, 10, 14, 11, 2, 14, 32, 12, 0, 10, 18, 3, 0, 47, 73, 16, 0, 16, 19, 2, 0, 0, 
    58, 26, 19, 0, 9, 1, 1, 3, 0, 0, 0, 6, 5, 10, 5, 0, 20, 21, 8, 9, 24, 11, 0, 49, 82, 34, 0, 14, 25, 14, 5, 0, 
    62, 24, 38, 19, 13, 6, 2, 7, 0, 0, 0, 1, 0, 0, 0, 0, 6, 13, 4, 0, 31, 31, 0, 48, 91, 49, 0, 14, 24, 26, 10, 0, 
    49, 3, 16, 34, 18, 9, 2, 2, 0, 0, 8, 3, 0, 0, 0, 0, 6, 35, 11, 0, 22, 38, 0, 43, 93, 58, 11, 19, 28, 22, 6, 14, 
    33, 0, 0, 19, 5, 11, 14, 0, 0, 0, 20, 5, 0, 0, 0, 0, 5, 27, 30, 0, 9, 36, 9, 27, 83, 69, 27, 33, 37, 22, 0, 2, 
    24, 0, 4, 31, 3, 0, 13, 17, 0, 0, 20, 12, 0, 0, 0, 0, 12, 0, 6, 22, 20, 35, 13, 21, 58, 65, 41, 43, 41, 15, 0, 0, 
    30, 0, 20, 51, 35, 0, 0, 24, 31, 19, 26, 21, 2, 0, 0, 10, 17, 9, 0, 19, 31, 30, 13, 38, 63, 50, 42, 45, 28, 0, 0, 0, 
    42, 0, 26, 61, 45, 27, 0, 0, 32, 39, 32, 43, 43, 11, 0, 6, 15, 18, 13, 20, 33, 19, 5, 40, 71, 47, 43, 41, 23, 0, 0, 0, 
    50, 0, 29, 63, 50, 44, 3, 0, 0, 19, 21, 51, 74, 66, 51, 34, 28, 18, 20, 34, 43, 42, 23, 30, 56, 39, 37, 41, 26, 0, 0, 0, 
    55, 0, 22, 53, 53, 52, 38, 5, 0, 19, 35, 63, 75, 68, 86, 93, 75, 60, 54, 64, 65, 62, 48, 57, 72, 33, 22, 46, 32, 0, 0, 0, 
    55, 0, 7, 38, 36, 53, 55, 36, 42, 66, 78, 89, 96, 75, 66, 80, 87, 92, 95, 94, 95, 88, 77, 76, 86, 55, 26, 31, 27, 3, 0, 0, 
    57, 4, 15, 34, 26, 43, 62, 50, 63, 80, 96, 104, 106, 101, 92, 84, 82, 80, 90, 103, 106, 113, 115, 94, 78, 70, 49, 32, 25, 4, 11, 6, 
    59, 7, 22, 34, 35, 29, 54, 60, 83, 81, 51, 79, 117, 108, 112, 117, 106, 94, 87, 91, 85, 96, 127, 124, 100, 63, 60, 46, 9, 0, 30, 13, 
    60, 10, 14, 29, 37, 29, 40, 48, 78, 128, 71, 38, 96, 113, 107, 107, 120, 129, 117, 107, 99, 76, 87, 132, 139, 88, 60, 56, 11, 0, 23, 9, 
    61, 26, 14, 22, 26, 40, 44, 46, 54, 110, 135, 63, 66, 112, 124, 116, 109, 106, 120, 125, 127, 123, 97, 95, 116, 129, 80, 54, 36, 0, 3, 22, 
    63, 34, 37, 24, 21, 25, 44, 40, 49, 53, 128, 129, 79, 100, 124, 125, 125, 115, 110, 113, 103, 111, 116, 98, 101, 85, 73, 57, 47, 17, 8, 0, 
    71, 31, 34, 34, 36, 6, 37, 39, 47, 36, 57, 145, 127, 96, 116, 109, 115, 131, 127, 115, 107, 108, 113, 103, 99, 68, 41, 28, 15, 42, 33, 0, 
    76, 19, 32, 33, 25, 0, 24, 32, 27, 60, 22, 60, 143, 124, 115, 124, 114, 116, 132, 127, 107, 107, 113, 103, 95, 84, 34, 20, 17, 18, 26, 0, 
    74, 10, 34, 38, 13, 3, 12, 34, 5, 28, 47, 8, 74, 137, 123, 120, 129, 114, 112, 124, 116, 111, 117, 110, 95, 77, 42, 43, 42, 15, 10, 0, 
    74, 18, 21, 45, 23, 0, 7, 40, 31, 0, 35, 48, 54, 106, 134, 126, 121, 129, 108, 100, 114, 118, 108, 111, 98, 69, 53, 46, 36, 24, 9, 0, 
    70, 41, 48, 40, 19, 0, 0, 18, 43, 22, 10, 62, 86, 99, 127, 138, 123, 125, 114, 103, 106, 114, 113, 117, 102, 81, 70, 48, 29, 18, 2, 0, 
    85, 57, 83, 91, 55, 20, 0, 0, 12, 33, 38, 36, 75, 110, 126, 136, 126, 123, 115, 103, 121, 126, 108, 110, 103, 86, 62, 60, 36, 8, 7, 0, 
    84, 66, 104, 128, 106, 58, 22, 7, 3, 3, 40, 63, 60, 94, 119, 120, 116, 130, 134, 116, 116, 132, 114, 104, 104, 81, 41, 45, 40, 3, 0, 0, 
    70, 35, 55, 107, 119, 99, 62, 31, 21, 0, 0, 44, 74, 79, 90, 80, 77, 111, 139, 132, 111, 122, 124, 106, 93, 78, 39, 27, 30, 0, 2, 0, 
    62, 12, 0, 51, 105, 106, 95, 72, 34, 15, 4, 1, 30, 47, 53, 43, 19, 60, 119, 125, 129, 115, 104, 108, 92, 54, 42, 22, 7, 7, 1, 0, 
    55, 10, 0, 0, 57, 98, 90, 94, 79, 42, 16, 5, 6, 14, 23, 29, 22, 38, 97, 121, 123, 129, 106, 83, 68, 42, 27, 4, 25, 48, 8, 0, 
    58, 11, 0, 0, 0, 65, 91, 95, 104, 86, 41, 18, 16, 7, 6, 19, 35, 59, 95, 116, 115, 116, 109, 86, 49, 13, 0, 11, 25, 55, 54, 0, 
    53, 3, 10, 2, 0, 3, 66, 93, 91, 97, 92, 60, 36, 22, 19, 28, 12, 21, 69, 84, 80, 99, 96, 82, 50, 7, 4, 18, 14, 43, 44, 0, 
    44, 10, 21, 32, 0, 0, 19, 74, 88, 87, 110, 118, 97, 73, 70, 86, 72, 30, 27, 50, 53, 70, 71, 77, 75, 59, 54, 56, 66, 71, 65, 0, 
    
    -- channel=80
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=81
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=82
    252, 69, 100, 163, 170, 140, 136, 142, 148, 135, 138, 155, 143, 124, 126, 149, 132, 90, 91, 122, 129, 115, 108, 112, 124, 124, 130, 140, 106, 72, 96, 34, 
    309, 153, 189, 196, 198, 202, 213, 210, 208, 203, 199, 207, 205, 201, 186, 199, 183, 135, 131, 157, 169, 154, 143, 132, 133, 146, 159, 167, 146, 120, 133, 47, 
    330, 191, 221, 192, 186, 206, 225, 212, 217, 215, 201, 208, 197, 198, 200, 196, 187, 141, 122, 159, 182, 170, 163, 151, 144, 146, 143, 144, 143, 145, 143, 40, 
    349, 215, 229, 210, 190, 213, 230, 209, 221, 224, 208, 215, 205, 197, 215, 212, 186, 151, 101, 127, 175, 175, 164, 170, 182, 170, 153, 140, 132, 156, 163, 38, 
    351, 197, 224, 229, 196, 222, 239, 222, 225, 225, 223, 223, 215, 204, 211, 238, 219, 175, 115, 91, 148, 165, 134, 140, 171, 175, 166, 155, 141, 150, 163, 38, 
    343, 170, 216, 241, 200, 215, 233, 235, 232, 228, 223, 227, 227, 204, 190, 232, 252, 220, 173, 115, 135, 173, 136, 129, 158, 158, 167, 174, 166, 157, 160, 38, 
    332, 167, 230, 240, 211, 220, 226, 233, 235, 232, 224, 226, 237, 216, 190, 209, 240, 238, 220, 181, 155, 183, 169, 142, 161, 153, 159, 185, 180, 168, 167, 39, 
    326, 169, 236, 225, 223, 226, 229, 242, 236, 230, 235, 235, 231, 218, 210, 210, 226, 237, 235, 219, 176, 177, 177, 135, 152, 156, 150, 168, 170, 165, 167, 40, 
    318, 188, 219, 221, 221, 222, 225, 242, 251, 234, 226, 227, 217, 200, 205, 199, 191, 207, 238, 238, 200, 197, 185, 116, 137, 168, 166, 160, 161, 161, 164, 42, 
    311, 211, 232, 224, 218, 222, 221, 225, 244, 241, 233, 219, 206, 189, 196, 181, 141, 153, 212, 240, 214, 212, 199, 120, 139, 184, 175, 171, 174, 169, 162, 42, 
    292, 254, 265, 210, 235, 248, 229, 231, 230, 239, 250, 233, 189, 152, 189, 203, 136, 122, 180, 214, 198, 196, 175, 131, 156, 189, 163, 166, 178, 177, 171, 41, 
    244, 308, 268, 172, 213, 230, 219, 224, 210, 222, 268, 267, 198, 122, 142, 201, 203, 166, 182, 205, 170, 156, 127, 109, 159, 185, 171, 166, 176, 176, 170, 46, 
    205, 313, 277, 208, 227, 206, 197, 200, 187, 219, 272, 267, 205, 143, 130, 105, 165, 192, 164, 193, 156, 118, 107, 101, 138, 168, 178, 172, 175, 173, 165, 51, 
    201, 236, 267, 270, 251, 199, 206, 191, 167, 218, 253, 219, 191, 193, 190, 111, 109, 160, 138, 149, 129, 96, 92, 95, 121, 152, 173, 165, 165, 160, 159, 58, 
    231, 161, 229, 295, 250, 186, 194, 210, 195, 222, 230, 183, 156, 196, 232, 180, 147, 162, 157, 147, 106, 83, 75, 88, 117, 150, 186, 159, 126, 140, 153, 58, 
    254, 121, 201, 289, 251, 188, 173, 216, 248, 236, 212, 197, 174, 187, 241, 215, 179, 183, 195, 173, 124, 77, 63, 95, 125, 173, 219, 185, 95, 94, 154, 63, 
    276, 135, 172, 247, 238, 187, 146, 191, 281, 240, 198, 232, 220, 181, 223, 239, 215, 200, 203, 206, 172, 101, 76, 111, 133, 202, 248, 215, 110, 50, 131, 78, 
    287, 155, 191, 241, 220, 185, 132, 151, 301, 242, 148, 234, 226, 150, 195, 228, 244, 227, 191, 205, 183, 133, 113, 118, 134, 197, 253, 226, 130, 32, 89, 81, 
    291, 148, 203, 274, 233, 175, 115, 82, 272, 295, 149, 222, 207, 114, 171, 182, 142, 176, 146, 153, 147, 127, 131, 112, 125, 188, 248, 247, 138, 11, 44, 80, 
    290, 133, 177, 267, 246, 183, 118, 22, 159, 349, 260, 221, 193, 136, 223, 233, 94, 78, 96, 125, 126, 112, 133, 105, 116, 195, 259, 274, 172, 0, 0, 64, 
    296, 141, 172, 247, 246, 186, 128, 22, 56, 248, 295, 259, 219, 170, 237, 280, 176, 94, 77, 122, 152, 136, 150, 119, 105, 174, 262, 298, 213, 25, 0, 41, 
    309, 143, 161, 235, 246, 180, 115, 53, 58, 115, 148, 190, 206, 182, 195, 216, 177, 152, 121, 116, 146, 143, 168, 170, 134, 156, 227, 302, 256, 77, 0, 26, 
    311, 149, 155, 203, 228, 182, 113, 86, 101, 99, 82, 105, 128, 147, 153, 138, 114, 145, 157, 136, 135, 121, 139, 185, 185, 181, 197, 264, 289, 139, 10, 6, 
    302, 171, 186, 167, 186, 208, 158, 119, 103, 118, 135, 134, 126, 133, 135, 90, 69, 98, 119, 125, 123, 109, 110, 141, 178, 199, 178, 206, 291, 225, 58, 0, 
    285, 174, 205, 171, 152, 211, 244, 189, 99, 117, 155, 130, 152, 151, 127, 96, 73, 74, 84, 93, 100, 98, 112, 120, 151, 192, 154, 159, 250, 272, 169, 0, 
    293, 182, 189, 179, 153, 158, 215, 257, 181, 143, 184, 144, 157, 170, 131, 108, 97, 86, 85, 84, 82, 77, 102, 116, 125, 157, 136, 139, 190, 184, 203, 59, 
    298, 174, 181, 208, 187, 142, 135, 215, 246, 142, 155, 181, 187, 196, 150, 118, 121, 123, 111, 103, 98, 91, 112, 123, 107, 115, 127, 150, 180, 126, 125, 74, 
    292, 148, 154, 218, 207, 155, 143, 171, 209, 170, 148, 165, 175, 195, 169, 133, 128, 150, 139, 127, 127, 131, 150, 149, 125, 124, 137, 151, 175, 155, 133, 34, 
    302, 152, 142, 190, 183, 148, 152, 169, 154, 143, 179, 170, 157, 182, 177, 153, 144, 160, 151, 148, 159, 162, 176, 173, 151, 151, 154, 145, 145, 164, 186, 24, 
    288, 176, 165, 167, 154, 157, 159, 173, 162, 147, 174, 164, 158, 176, 178, 182, 173, 165, 151, 156, 180, 178, 184, 188, 166, 158, 162, 145, 141, 175, 195, 26, 
    296, 192, 182, 158, 150, 186, 193, 184, 174, 186, 199, 180, 170, 163, 157, 185, 197, 179, 162, 158, 177, 182, 183, 192, 175, 157, 167, 156, 149, 167, 178, 23, 
    300, 255, 245, 216, 192, 210, 237, 238, 222, 222, 242, 233, 229, 216, 192, 203, 225, 227, 221, 212, 223, 231, 231, 241, 232, 215, 219, 225, 218, 218, 220, 118, 
    
    -- channel=83
    0, 8, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=84
    0, 228, 147, 85, 112, 155, 162, 154, 157, 168, 154, 139, 152, 154, 138, 102, 107, 131, 105, 71, 69, 87, 94, 76, 67, 65, 59, 59, 109, 125, 91, 130, 
    0, 222, 143, 89, 94, 127, 120, 123, 129, 150, 146, 129, 134, 144, 131, 85, 96, 135, 107, 42, 33, 65, 88, 89, 84, 72, 58, 36, 87, 111, 78, 171, 
    0, 152, 111, 132, 151, 131, 95, 122, 126, 146, 158, 153, 157, 160, 156, 125, 136, 156, 128, 41, 8, 37, 63, 88, 95, 86, 81, 71, 89, 90, 74, 197, 
    0, 100, 92, 137, 170, 128, 105, 137, 123, 144, 158, 156, 175, 171, 147, 144, 159, 205, 189, 85, 9, 19, 44, 52, 45, 64, 91, 106, 107, 81, 69, 212, 
    0, 109, 90, 110, 164, 121, 109, 137, 127, 139, 149, 146, 165, 173, 143, 135, 159, 213, 237, 160, 62, 52, 99, 88, 51, 68, 86, 111, 120, 84, 70, 226, 
    0, 150, 79, 85, 154, 121, 113, 128, 128, 138, 142, 154, 160, 185, 176, 121, 123, 164, 211, 209, 121, 87, 139, 127, 77, 75, 80, 81, 92, 88, 77, 237, 
    0, 155, 42, 72, 130, 123, 123, 121, 127, 134, 149, 154, 152, 177, 192, 138, 109, 127, 155, 187, 145, 102, 134, 136, 92, 87, 79, 53, 63, 81, 76, 240, 
    0, 121, 42, 71, 108, 119, 119, 112, 119, 127, 144, 145, 148, 158, 170, 143, 106, 98, 108, 142, 182, 153, 159, 175, 110, 101, 96, 70, 75, 79, 78, 241, 
    0, 96, 53, 76, 111, 124, 119, 103, 109, 133, 153, 157, 165, 157, 158, 150, 134, 102, 90, 106, 176, 153, 153, 196, 131, 83, 85, 79, 80, 81, 81, 238, 
    0, 58, 38, 82, 112, 120, 138, 124, 118, 138, 155, 149, 151, 148, 143, 157, 188, 148, 88, 73, 129, 105, 121, 188, 116, 36, 52, 65, 62, 76, 80, 240, 
    0, 0, 0, 82, 77, 89, 134, 137, 123, 120, 124, 133, 144, 146, 94, 98, 179, 187, 106, 72, 112, 93, 101, 158, 66, 18, 59, 66, 54, 63, 73, 237, 
    0, 0, 0, 148, 106, 116, 142, 128, 139, 125, 91, 75, 111, 144, 61, 21, 70, 111, 87, 65, 105, 116, 139, 144, 41, 4, 50, 60, 50, 52, 67, 233, 
    0, 0, 0, 129, 90, 117, 136, 131, 159, 115, 41, 16, 78, 140, 126, 104, 74, 87, 95, 66, 108, 142, 159, 122, 28, 0, 29, 52, 48, 52, 64, 219, 
    0, 0, 0, 11, 47, 116, 123, 134, 168, 95, 34, 47, 101, 112, 132, 213, 133, 105, 135, 88, 142, 164, 152, 118, 48, 17, 26, 54, 61, 58, 65, 204, 
    0, 3, 0, 0, 44, 129, 107, 118, 132, 69, 59, 130, 170, 130, 84, 156, 119, 93, 113, 116, 172, 187, 179, 119, 55, 19, 14, 73, 106, 87, 62, 190, 
    0, 122, 12, 0, 25, 126, 116, 75, 53, 45, 81, 145, 177, 135, 57, 75, 86, 75, 68, 109, 171, 202, 186, 94, 38, 0, 0, 71, 154, 130, 56, 168, 
    0, 166, 58, 0, 36, 128, 161, 80, 0, 16, 83, 56, 101, 136, 62, 45, 57, 55, 48, 58, 93, 159, 142, 67, 18, 0, 0, 21, 174, 179, 60, 144, 
    0, 152, 77, 0, 48, 123, 185, 99, 0, 2, 132, 39, 82, 157, 78, 17, 22, 22, 35, 8, 25, 107, 98, 61, 27, 0, 0, 0, 163, 226, 94, 120, 
    0, 144, 52, 0, 35, 107, 202, 163, 0, 0, 148, 51, 79, 194, 127, 115, 121, 92, 85, 48, 55, 93, 78, 76, 40, 0, 0, 0, 140, 264, 145, 104, 
    0, 186, 80, 0, 13, 89, 186, 248, 0, 0, 0, 0, 78, 187, 56, 95, 199, 189, 162, 85, 72, 79, 53, 81, 42, 0, 0, 0, 114, 296, 210, 115, 
    0, 190, 99, 0, 0, 62, 140, 288, 80, 0, 0, 0, 3, 79, 0, 0, 144, 210, 180, 76, 22, 18, 9, 79, 77, 0, 0, 0, 51, 291, 258, 139, 
    0, 169, 110, 0, 0, 66, 142, 275, 188, 0, 0, 0, 0, 31, 0, 0, 87, 135, 130, 56, 0, 0, 0, 29, 66, 17, 0, 0, 0, 237, 272, 170, 
    0, 172, 128, 36, 16, 82, 180, 239, 180, 135, 108, 64, 46, 71, 57, 73, 92, 41, 35, 22, 0, 3, 0, 0, 0, 0, 0, 0, 0, 164, 277, 211, 
    0, 143, 112, 92, 59, 72, 157, 201, 184, 161, 127, 119, 106, 89, 86, 137, 147, 67, 16, 9, 0, 12, 0, 0, 0, 0, 3, 0, 0, 64, 256, 267, 
    0, 126, 92, 128, 102, 39, 41, 115, 226, 208, 144, 143, 127, 108, 140, 190, 180, 114, 62, 37, 18, 19, 3, 0, 0, 0, 23, 0, 0, 0, 144, 278, 
    0, 117, 92, 135, 158, 82, 3, 29, 157, 156, 104, 122, 115, 121, 175, 190, 175, 137, 112, 94, 81, 75, 38, 30, 1, 0, 54, 48, 0, 0, 42, 221, 
    0, 111, 110, 91, 125, 151, 102, 1, 52, 115, 99, 104, 82, 78, 151, 179, 169, 137, 130, 123, 119, 118, 82, 75, 82, 70, 96, 66, 24, 74, 46, 182, 
    0, 133, 114, 38, 75, 149, 165, 53, 19, 132, 109, 100, 85, 69, 135, 186, 170, 126, 121, 121, 116, 122, 94, 97, 133, 130, 112, 70, 22, 107, 97, 209, 
    0, 137, 132, 52, 103, 154, 159, 119, 97, 139, 108, 115, 114, 94, 124, 172, 162, 113, 111, 116, 112, 116, 97, 109, 140, 138, 120, 116, 98, 97, 83, 255, 
    0, 145, 137, 106, 142, 161, 147, 118, 149, 145, 94, 133, 147, 118, 110, 121, 124, 118, 133, 123, 105, 109, 104, 112, 139, 141, 128, 152, 148, 87, 40, 273, 
    0, 116, 117, 138, 138, 102, 94, 96, 118, 109, 78, 124, 140, 137, 124, 89, 91, 118, 140, 126, 100, 110, 115, 106, 136, 142, 132, 150, 148, 97, 73, 291, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 141, 
    
    -- channel=85
    95, 53, 68, 77, 78, 79, 85, 87, 83, 78, 78, 78, 77, 71, 63, 71, 67, 47, 36, 39, 44, 43, 38, 35, 33, 41, 52, 62, 49, 38, 37, 0, 
    79, 9, 42, 51, 31, 16, 30, 29, 27, 20, 16, 17, 12, 11, 15, 23, 12, 0, 0, 0, 9, 6, 6, 2, 1, 4, 10, 17, 4, 0, 5, 0, 
    91, 29, 48, 31, 5, 14, 29, 19, 23, 23, 19, 24, 17, 14, 19, 23, 14, 0, 0, 0, 5, 7, 12, 17, 26, 30, 25, 10, 0, 0, 10, 0, 
    97, 24, 31, 13, 3, 24, 36, 25, 26, 27, 26, 26, 21, 21, 27, 29, 23, 1, 0, 0, 1, 6, 0, 2, 18, 23, 17, 6, 0, 5, 15, 0, 
    102, 5, 9, 13, 3, 23, 37, 29, 31, 30, 24, 26, 22, 13, 14, 27, 32, 28, 9, 3, 19, 26, 6, 0, 6, 5, 6, 5, 6, 14, 17, 0, 
    101, 0, 18, 25, 12, 27, 28, 25, 32, 30, 22, 21, 27, 18, 11, 21, 28, 34, 33, 25, 36, 40, 20, 12, 18, 8, 1, 9, 13, 17, 20, 0, 
    81, 0, 31, 26, 18, 24, 29, 32, 30, 30, 24, 25, 29, 25, 20, 26, 29, 26, 27, 25, 25, 26, 10, 0, 5, 0, 0, 8, 10, 10, 14, 0, 
    73, 1, 21, 23, 15, 20, 26, 33, 34, 22, 18, 27, 26, 14, 12, 20, 23, 23, 26, 25, 12, 20, 8, 0, 0, 0, 7, 12, 10, 10, 10, 0, 
    78, 2, 31, 25, 19, 22, 20, 24, 27, 25, 22, 20, 16, 9, 13, 15, 4, 2, 13, 27, 19, 34, 32, 0, 0, 11, 18, 22, 18, 11, 11, 0, 
    63, 8, 39, 25, 27, 28, 25, 29, 26, 23, 26, 28, 23, 17, 36, 35, 6, 0, 8, 22, 18, 24, 14, 0, 0, 13, 8, 7, 10, 11, 12, 0, 
    24, 24, 38, 11, 23, 35, 31, 33, 28, 20, 31, 46, 36, 7, 26, 43, 13, 0, 14, 24, 11, 6, 0, 0, 0, 7, 0, 0, 3, 8, 12, 0, 
    10, 51, 55, 17, 31, 27, 19, 25, 9, 8, 38, 67, 49, 10, 0, 0, 0, 0, 16, 33, 15, 0, 0, 0, 0, 4, 1, 4, 11, 11, 8, 0, 
    34, 75, 60, 44, 67, 50, 32, 16, 0, 22, 60, 58, 21, 0, 0, 0, 0, 0, 8, 26, 9, 0, 0, 0, 0, 0, 0, 2, 9, 7, 5, 0, 
    65, 53, 31, 46, 48, 20, 18, 18, 10, 41, 60, 28, 0, 0, 32, 31, 50, 50, 39, 38, 0, 0, 0, 0, 0, 0, 9, 8, 4, 1, 0, 0, 
    69, 23, 29, 52, 44, 11, 8, 17, 34, 59, 59, 24, 0, 13, 50, 50, 56, 63, 50, 34, 8, 0, 0, 0, 0, 8, 33, 26, 0, 0, 0, 0, 
    65, 2, 25, 67, 49, 13, 1, 17, 45, 61, 43, 22, 20, 34, 59, 49, 27, 26, 27, 28, 11, 0, 0, 0, 0, 15, 47, 43, 3, 0, 0, 0, 
    70, 16, 47, 66, 41, 16, 0, 6, 57, 40, 0, 16, 25, 12, 21, 20, 19, 13, 8, 6, 0, 0, 0, 0, 0, 15, 53, 49, 2, 0, 0, 0, 
    77, 14, 43, 80, 55, 23, 0, 0, 59, 29, 0, 18, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 55, 52, 3, 0, 0, 0, 
    76, 0, 27, 70, 59, 29, 0, 0, 19, 40, 5, 39, 29, 0, 13, 17, 0, 0, 0, 0, 0, 0, 0, 0, 3, 34, 63, 70, 27, 0, 0, 0, 
    78, 4, 27, 62, 55, 26, 0, 0, 0, 17, 21, 37, 0, 0, 39, 74, 28, 0, 0, 0, 0, 0, 11, 0, 0, 27, 67, 84, 42, 0, 0, 0, 
    87, 13, 31, 71, 58, 12, 0, 0, 0, 0, 0, 0, 0, 0, 5, 25, 0, 0, 0, 0, 0, 1, 14, 0, 0, 16, 53, 83, 51, 0, 0, 0, 
    92, 7, 12, 45, 42, 2, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 22, 40, 64, 50, 0, 0, 0, 
    83, 2, 16, 32, 33, 3, 0, 0, 6, 22, 24, 18, 4, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 24, 35, 41, 0, 0, 0, 
    64, 5, 34, 32, 17, 19, 24, 19, 4, 9, 24, 38, 45, 39, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 1, 3, 33, 16, 0, 0, 
    67, 13, 31, 25, 12, 16, 37, 46, 11, 10, 24, 11, 11, 22, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 16, 0, 0, 11, 10, 0, 0, 
    77, 28, 34, 24, 16, 11, 0, 13, 12, 7, 25, 18, 22, 29, 17, 8, 7, 8, 7, 7, 2, 0, 0, 7, 8, 7, 0, 0, 28, 1, 0, 0, 
    79, 15, 8, 31, 35, 18, 0, 3, 7, 0, 0, 0, 21, 41, 26, 8, 4, 17, 22, 20, 18, 20, 35, 38, 23, 15, 6, 23, 54, 17, 0, 0, 
    82, 1, 0, 26, 22, 0, 0, 21, 13, 0, 13, 20, 21, 30, 16, 2, 9, 21, 21, 18, 22, 26, 43, 45, 32, 29, 32, 31, 23, 3, 19, 0, 
    74, 12, 14, 32, 14, 0, 2, 22, 21, 0, 14, 32, 30, 27, 15, 9, 14, 19, 8, 10, 20, 26, 36, 35, 24, 23, 27, 14, 3, 9, 25, 0, 
    73, 18, 34, 38, 20, 13, 24, 34, 30, 32, 40, 22, 11, 13, 5, 7, 12, 11, 3, 6, 21, 27, 29, 30, 22, 18, 17, 6, 8, 29, 42, 0, 
    89, 44, 37, 17, 0, 6, 25, 28, 13, 12, 27, 18, 14, 6, 0, 0, 6, 13, 13, 18, 28, 24, 24, 29, 19, 13, 16, 16, 18, 29, 25, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=86
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=87
    0, 7, 15, 10, 2, 3, 4, 3, 3, 3, 7, 4, 3, 5, 6, 5, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 11, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 5, 10, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 5, 9, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 2, 7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 3, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 3, 
    0, 0, 0, 0, 0, 0, 0, 8, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 6, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 5, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=88
    12, 66, 29, 21, 38, 42, 31, 32, 38, 41, 31, 29, 31, 35, 32, 27, 46, 53, 34, 12, 11, 17, 20, 18, 15, 8, 7, 15, 41, 38, 23, 53, 
    0, 54, 50, 30, 15, 10, 6, 13, 6, 13, 11, 0, 0, 4, 5, 0, 16, 41, 28, 0, 0, 0, 6, 11, 0, 1, 4, 3, 18, 33, 16, 61, 
    0, 63, 46, 45, 34, 8, 6, 12, 9, 17, 15, 2, 4, 0, 0, 2, 7, 32, 23, 0, 0, 0, 1, 9, 12, 15, 12, 13, 14, 15, 11, 71, 
    0, 63, 40, 52, 38, 10, 9, 17, 16, 14, 18, 13, 13, 4, 0, 0, 0, 28, 40, 3, 0, 0, 0, 0, 0, 4, 15, 20, 15, 5, 11, 77, 
    0, 67, 35, 40, 42, 18, 9, 21, 18, 15, 22, 15, 12, 13, 0, 0, 0, 25, 58, 38, 0, 0, 11, 0, 0, 0, 7, 14, 19, 11, 6, 82, 
    0, 75, 32, 37, 47, 25, 15, 16, 21, 25, 22, 14, 15, 20, 11, 0, 0, 16, 46, 61, 25, 11, 29, 17, 0, 0, 0, 0, 11, 14, 8, 86, 
    0, 62, 38, 36, 43, 32, 19, 19, 29, 29, 27, 18, 16, 18, 24, 2, 0, 6, 27, 47, 40, 4, 18, 20, 0, 0, 0, 0, 0, 7, 11, 84, 
    0, 63, 43, 29, 38, 29, 24, 24, 30, 30, 18, 14, 13, 14, 18, 11, 0, 0, 1, 13, 33, 10, 26, 38, 4, 0, 0, 0, 0, 6, 9, 83, 
    0, 72, 25, 32, 38, 31, 31, 20, 22, 23, 16, 22, 25, 19, 11, 20, 20, 1, 0, 0, 25, 26, 40, 61, 17, 0, 4, 5, 3, 11, 7, 82, 
    0, 27, 19, 43, 38, 36, 31, 27, 22, 27, 30, 36, 39, 40, 31, 53, 60, 30, 0, 0, 11, 24, 43, 74, 17, 0, 0, 1, 2, 6, 8, 83, 
    0, 0, 19, 40, 20, 23, 36, 42, 36, 23, 21, 47, 83, 94, 66, 68, 88, 63, 8, 0, 15, 28, 41, 48, 4, 0, 0, 0, 0, 0, 8, 81, 
    0, 0, 6, 45, 35, 47, 56, 47, 47, 25, 21, 66, 125, 127, 93, 65, 52, 49, 22, 12, 35, 40, 43, 34, 5, 0, 0, 0, 0, 0, 3, 76, 
    0, 0, 0, 57, 66, 70, 69, 68, 58, 32, 36, 80, 117, 119, 102, 76, 29, 45, 52, 36, 64, 62, 53, 38, 0, 0, 0, 0, 0, 0, 0, 67, 
    0, 0, 0, 27, 62, 86, 82, 81, 70, 52, 64, 93, 92, 83, 87, 116, 85, 80, 94, 83, 93, 80, 60, 36, 6, 0, 0, 0, 0, 0, 0, 59, 
    0, 1, 0, 3, 57, 96, 84, 73, 80, 76, 82, 102, 97, 71, 72, 118, 135, 110, 120, 125, 110, 105, 79, 45, 20, 0, 0, 13, 27, 8, 0, 55, 
    0, 26, 0, 0, 52, 95, 88, 55, 66, 86, 106, 112, 108, 76, 60, 99, 126, 116, 118, 118, 133, 135, 89, 48, 9, 0, 0, 24, 67, 35, 0, 51, 
    0, 36, 11, 1, 53, 90, 103, 61, 39, 102, 113, 71, 78, 86, 63, 72, 88, 98, 92, 95, 114, 110, 70, 23, 0, 0, 0, 19, 88, 74, 3, 42, 
    0, 35, 19, 15, 65, 101, 116, 78, 12, 88, 91, 48, 81, 107, 45, 33, 38, 56, 62, 45, 45, 43, 25, 1, 0, 0, 0, 22, 91, 113, 25, 28, 
    0, 31, 0, 8, 77, 113, 126, 118, 0, 30, 102, 70, 80, 92, 27, 51, 57, 41, 42, 15, 9, 0, 0, 7, 0, 0, 0, 22, 104, 147, 55, 22, 
    0, 32, 12, 10, 76, 126, 138, 149, 11, 0, 53, 53, 63, 74, 26, 45, 94, 59, 41, 9, 7, 7, 0, 11, 0, 0, 0, 16, 117, 176, 93, 29, 
    0, 49, 32, 10, 66, 119, 128, 138, 36, 0, 0, 5, 14, 25, 0, 0, 60, 62, 38, 6, 0, 0, 0, 2, 1, 0, 0, 6, 103, 189, 129, 43, 
    0, 51, 27, 11, 54, 101, 110, 96, 48, 0, 0, 0, 0, 0, 0, 0, 12, 22, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 68, 165, 142, 59, 
    0, 42, 27, 20, 38, 84, 96, 74, 64, 39, 14, 0, 0, 0, 0, 7, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 119, 144, 76, 
    0, 17, 21, 39, 42, 53, 81, 96, 78, 24, 22, 19, 16, 9, 13, 19, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 125, 109, 
    0, 14, 15, 41, 48, 34, 53, 78, 84, 42, 32, 30, 10, 4, 12, 38, 49, 25, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 65, 136, 
    0, 18, 7, 24, 54, 48, 30, 25, 84, 83, 29, 25, 0, 9, 36, 46, 45, 35, 24, 16, 14, 11, 0, 0, 0, 0, 0, 0, 0, 0, 17, 104, 
    0, 22, 15, 8, 43, 64, 42, 4, 35, 77, 24, 18, 7, 11, 35, 46, 35, 28, 31, 37, 33, 24, 8, 13, 19, 3, 3, 4, 0, 40, 6, 60, 
    0, 38, 15, 0, 26, 52, 45, 17, 12, 51, 22, 15, 13, 5, 24, 42, 30, 25, 36, 33, 21, 18, 15, 21, 32, 28, 19, 13, 8, 19, 20, 77, 
    0, 27, 20, 8, 20, 36, 30, 28, 29, 27, 30, 27, 20, 9, 17, 30, 33, 24, 23, 9, 5, 10, 8, 14, 30, 29, 22, 22, 7, 0, 21, 107, 
    0, 18, 34, 33, 27, 34, 30, 25, 39, 42, 25, 26, 29, 19, 14, 9, 18, 13, 11, 5, 0, 3, 5, 10, 29, 27, 25, 26, 20, 10, 5, 105, 
    0, 16, 35, 42, 36, 10, 6, 16, 32, 32, 17, 18, 21, 22, 17, 0, 0, 4, 14, 11, 0, 7, 11, 12, 28, 31, 21, 25, 30, 17, 12, 105, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    
    -- channel=89
    65, 72, 75, 74, 59, 44, 42, 44, 43, 37, 29, 26, 30, 36, 40, 46, 64, 73, 67, 60, 60, 62, 62, 57, 53, 54, 62, 72, 85, 84, 83, 95, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 15, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    76, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 70, 66, 51, 34, 0, 0, 0, 1, 18, 7, 0, 0, 0, 0, 0, 0, 
    54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 40, 48, 24, 26, 8, 0, 9, 19, 28, 14, 0, 2, 0, 0, 0, 0, 
    19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 8, 12, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 13, 0, 0, 0, 7, 2, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 37, 25, 0, 0, 20, 27, 11, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 36, 33, 14, 0, 0, 0, 27, 43, 27, 35, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 10, 7, 2, 7, 0, 0, 0, 5, 21, 23, 44, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 61, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 32, 
    0, 0, 0, 0, 0, 0, 0, 0, 21, 61, 56, 51, 28, 0, 0, 0, 0, 0, 0, 0, 18, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 
    0, 0, 0, 0, 0, 0, 0, 2, 5, 0, 0, 14, 22, 2, 0, 0, 0, 14, 25, 26, 35, 43, 44, 25, 0, 0, 0, 0, 0, 0, 0, 37, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 61, 70, 64, 59, 54, 55, 56, 32, 10, 0, 0, 0, 0, 0, 27, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 37, 58, 71, 81, 80, 76, 74, 58, 26, 0, 0, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 48, 58, 60, 67, 73, 64, 39, 13, 16, 31, 24, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 17, 11, 8, 9, 0, 0, 0, 0, 29, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=90
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=91
    146, 238, 189, 196, 217, 217, 205, 209, 219, 217, 209, 201, 199, 194, 191, 178, 178, 180, 159, 137, 129, 137, 138, 136, 129, 120, 121, 137, 156, 157, 139, 139, 
    31, 170, 170, 164, 130, 100, 86, 96, 102, 107, 108, 95, 93, 94, 92, 79, 85, 107, 91, 54, 40, 54, 69, 73, 72, 71, 73, 60, 71, 81, 76, 112, 
    31, 160, 160, 158, 136, 99, 77, 94, 98, 108, 116, 107, 105, 103, 96, 95, 103, 105, 92, 46, 27, 44, 60, 76, 89, 93, 86, 70, 67, 59, 63, 123, 
    19, 131, 132, 136, 136, 108, 96, 112, 109, 111, 116, 122, 124, 113, 101, 89, 103, 122, 121, 80, 36, 34, 44, 46, 40, 53, 69, 72, 71, 65, 67, 127, 
    11, 128, 113, 110, 138, 117, 108, 118, 111, 113, 119, 116, 116, 113, 96, 84, 100, 142, 159, 136, 85, 69, 80, 61, 36, 41, 49, 67, 78, 73, 66, 126, 
    20, 144, 104, 116, 145, 119, 110, 109, 110, 115, 120, 118, 112, 122, 114, 91, 91, 116, 150, 165, 141, 114, 113, 92, 52, 44, 42, 46, 63, 70, 68, 130, 
    16, 136, 92, 124, 134, 118, 109, 110, 117, 120, 122, 123, 112, 118, 123, 103, 88, 95, 122, 147, 132, 100, 87, 83, 54, 42, 36, 26, 41, 56, 58, 126, 
    3, 123, 107, 114, 113, 113, 112, 111, 114, 117, 114, 102, 96, 99, 103, 96, 85, 76, 76, 95, 107, 104, 111, 117, 74, 51, 51, 53, 56, 56, 57, 123, 
    19, 124, 103, 103, 119, 122, 116, 106, 100, 106, 111, 109, 102, 94, 91, 94, 94, 73, 55, 65, 105, 118, 133, 146, 98, 64, 71, 71, 66, 62, 59, 120, 
    4, 79, 74, 114, 124, 122, 125, 113, 116, 127, 127, 113, 105, 106, 112, 130, 149, 112, 64, 46, 73, 85, 111, 130, 88, 47, 55, 51, 48, 53, 57, 124, 
    0, 11, 57, 110, 86, 92, 130, 135, 131, 122, 107, 113, 139, 161, 130, 117, 155, 146, 85, 54, 70, 71, 82, 85, 47, 39, 50, 50, 45, 51, 54, 122, 
    0, 0, 66, 125, 111, 139, 151, 131, 123, 113, 108, 138, 176, 176, 111, 72, 65, 79, 82, 67, 83, 85, 75, 79, 49, 41, 49, 54, 48, 46, 50, 114, 
    3, 4, 80, 139, 142, 158, 146, 135, 134, 112, 113, 135, 148, 149, 111, 86, 71, 79, 111, 99, 103, 108, 96, 81, 46, 32, 43, 52, 50, 48, 43, 104, 
    33, 41, 45, 56, 98, 136, 133, 132, 145, 132, 132, 135, 128, 117, 134, 175, 175, 175, 175, 152, 150, 125, 102, 83, 60, 55, 57, 67, 62, 49, 42, 96, 
    38, 60, 20, 25, 94, 136, 129, 126, 142, 147, 147, 155, 161, 144, 129, 176, 186, 179, 181, 173, 171, 156, 138, 104, 78, 64, 62, 90, 102, 71, 43, 97, 
    12, 83, 46, 29, 85, 130, 120, 105, 105, 131, 157, 175, 176, 152, 109, 122, 136, 137, 133, 145, 173, 181, 150, 88, 57, 37, 52, 102, 131, 109, 50, 92, 
    10, 93, 65, 51, 87, 125, 140, 114, 79, 121, 142, 89, 96, 122, 98, 82, 85, 95, 98, 103, 114, 117, 88, 42, 28, 18, 26, 81, 136, 133, 66, 82, 
    0, 90, 71, 53, 102, 143, 160, 122, 51, 77, 120, 65, 101, 133, 67, 28, 39, 37, 48, 22, 7, 23, 23, 35, 42, 24, 26, 64, 139, 158, 91, 76, 
    0, 67, 35, 27, 89, 135, 169, 143, 28, 25, 137, 128, 115, 113, 68, 79, 116, 69, 30, 3, 0, 23, 43, 75, 73, 37, 35, 64, 143, 194, 123, 74, 
    0, 72, 56, 45, 84, 130, 173, 166, 26, 0, 26, 64, 77, 100, 71, 101, 147, 126, 76, 38, 48, 76, 75, 83, 63, 22, 12, 58, 145, 219, 165, 95, 
    0, 103, 82, 46, 65, 112, 139, 153, 34, 0, 0, 0, 0, 18, 0, 0, 52, 85, 83, 60, 49, 48, 36, 53, 56, 31, 14, 32, 116, 220, 195, 118, 
    0, 88, 62, 29, 49, 92, 114, 137, 93, 35, 7, 0, 0, 0, 0, 0, 7, 28, 43, 39, 23, 18, 9, 26, 55, 51, 16, 0, 57, 181, 191, 132, 
    0, 73, 56, 43, 53, 89, 128, 155, 160, 147, 103, 71, 62, 63, 53, 47, 23, 0, 13, 25, 29, 31, 13, 3, 12, 17, 5, 0, 10, 125, 186, 151, 
    0, 50, 45, 67, 74, 79, 135, 194, 184, 129, 94, 112, 108, 99, 71, 66, 67, 51, 42, 41, 39, 43, 31, 12, 0, 3, 28, 3, 0, 60, 161, 183, 
    0, 56, 56, 67, 68, 72, 94, 135, 171, 153, 119, 117, 82, 55, 70, 104, 121, 114, 95, 77, 56, 54, 51, 45, 36, 25, 39, 6, 0, 2, 90, 172, 
    0, 66, 50, 60, 83, 85, 62, 57, 119, 158, 108, 67, 49, 56, 102, 123, 125, 119, 112, 104, 100, 99, 86, 85, 78, 48, 42, 31, 10, 27, 60, 109, 
    0, 55, 51, 42, 78, 105, 75, 41, 54, 85, 80, 53, 50, 58, 89, 105, 105, 97, 113, 129, 134, 130, 118, 123, 119, 97, 97, 91, 85, 84, 58, 92, 
    0, 60, 43, 13, 42, 83, 85, 47, 55, 80, 68, 77, 72, 50, 65, 84, 90, 90, 105, 105, 100, 109, 111, 118, 130, 128, 121, 100, 70, 69, 61, 136, 
    0, 45, 51, 39, 55, 62, 77, 75, 69, 91, 84, 91, 79, 57, 57, 75, 85, 81, 71, 58, 62, 83, 85, 89, 105, 107, 102, 92, 61, 59, 79, 162, 
    0, 64, 85, 79, 78, 75, 80, 82, 98, 103, 85, 87, 79, 63, 51, 48, 54, 59, 57, 55, 56, 65, 68, 72, 84, 89, 84, 92, 92, 76, 61, 144, 
    0, 80, 87, 83, 65, 37, 31, 44, 73, 74, 56, 62, 61, 63, 55, 34, 31, 52, 70, 69, 59, 63, 67, 66, 77, 80, 71, 83, 94, 79, 61, 139, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    
    -- channel=92
    145, 140, 89, 100, 146, 164, 157, 154, 160, 158, 146, 145, 144, 130, 112, 113, 122, 105, 72, 61, 69, 72, 66, 57, 56, 57, 64, 86, 100, 77, 57, 22, 
    167, 136, 130, 156, 160, 142, 140, 149, 150, 142, 127, 123, 115, 108, 97, 90, 93, 70, 41, 35, 48, 55, 54, 46, 38, 37, 53, 73, 84, 61, 55, 26, 
    177, 170, 189, 187, 155, 131, 134, 147, 148, 151, 143, 137, 127, 114, 107, 106, 106, 75, 30, 12, 32, 53, 64, 74, 79, 87, 89, 81, 71, 57, 60, 30, 
    176, 185, 199, 185, 160, 139, 148, 156, 155, 163, 157, 154, 152, 136, 127, 128, 120, 87, 37, 3, 17, 41, 52, 61, 78, 98, 97, 87, 67, 58, 73, 49, 
    175, 182, 170, 172, 161, 150, 165, 169, 169, 171, 167, 168, 160, 141, 126, 131, 140, 129, 89, 45, 39, 60, 64, 54, 60, 78, 85, 86, 78, 73, 83, 51, 
    185, 180, 155, 175, 175, 166, 169, 169, 175, 177, 176, 170, 164, 155, 131, 123, 147, 151, 140, 110, 96, 110, 109, 84, 77, 78, 74, 79, 86, 90, 94, 59, 
    184, 164, 150, 186, 184, 174, 174, 174, 180, 186, 187, 178, 173, 173, 154, 134, 145, 148, 156, 153, 136, 125, 110, 80, 71, 66, 55, 60, 77, 87, 93, 61, 
    166, 142, 153, 183, 174, 171, 174, 181, 189, 186, 187, 179, 172, 166, 155, 140, 143, 149, 156, 158, 142, 118, 111, 83, 63, 59, 52, 61, 77, 84, 90, 57, 
    153, 147, 169, 172, 174, 175, 173, 174, 181, 184, 182, 174, 168, 159, 149, 137, 131, 125, 134, 151, 158, 146, 155, 114, 69, 67, 76, 88, 91, 90, 91, 56, 
    133, 141, 157, 176, 188, 186, 183, 173, 176, 188, 192, 185, 173, 170, 175, 178, 162, 126, 118, 136, 152, 145, 156, 112, 62, 65, 76, 79, 81, 89, 89, 56, 
    73, 91, 147, 176, 173, 185, 194, 191, 194, 188, 183, 185, 190, 194, 197, 216, 202, 150, 119, 129, 138, 131, 120, 71, 32, 54, 61, 57, 63, 81, 89, 59, 
    1, 56, 168, 172, 161, 191, 203, 200, 189, 168, 172, 211, 245, 231, 181, 163, 160, 142, 122, 140, 146, 126, 86, 29, 9, 48, 57, 57, 62, 76, 83, 52, 
    0, 74, 195, 206, 228, 247, 228, 203, 182, 163, 189, 230, 248, 216, 164, 114, 83, 106, 121, 144, 154, 125, 77, 27, 13, 27, 39, 49, 56, 72, 76, 43, 
    22, 91, 158, 183, 228, 234, 218, 209, 186, 177, 217, 233, 212, 183, 190, 186, 166, 190, 189, 186, 171, 121, 68, 24, 11, 21, 42, 54, 55, 63, 61, 32, 
    77, 98, 108, 155, 223, 224, 206, 207, 207, 221, 253, 244, 207, 182, 207, 241, 243, 262, 248, 235, 204, 138, 83, 40, 25, 34, 63, 85, 72, 57, 52, 26, 
    104, 91, 83, 158, 226, 226, 198, 186, 209, 248, 270, 265, 252, 225, 226, 248, 246, 247, 241, 246, 220, 170, 100, 41, 20, 28, 79, 129, 111, 61, 43, 25, 
    122, 112, 109, 161, 213, 220, 192, 161, 199, 250, 248, 234, 242, 219, 206, 215, 220, 217, 212, 215, 202, 154, 62, 2, 0, 8, 84, 148, 143, 73, 32, 16, 
    131, 129, 133, 184, 230, 235, 212, 153, 176, 236, 198, 173, 217, 204, 163, 148, 148, 165, 151, 128, 99, 49, 0, 0, 0, 7, 85, 149, 160, 91, 27, 2, 
    140, 125, 114, 171, 236, 248, 222, 132, 111, 205, 200, 201, 237, 189, 132, 135, 120, 104, 69, 31, 4, 0, 0, 0, 0, 28, 96, 166, 189, 121, 25, 0, 
    143, 123, 104, 159, 228, 252, 238, 135, 30, 114, 179, 207, 204, 157, 149, 225, 204, 126, 42, 3, 4, 8, 25, 29, 6, 30, 94, 179, 220, 166, 36, 0, 
    154, 147, 139, 174, 217, 234, 214, 118, 0, 0, 46, 95, 116, 97, 93, 161, 167, 116, 39, 0, 11, 25, 39, 35, 3, 18, 82, 176, 235, 199, 67, 0, 
    165, 157, 134, 148, 189, 204, 166, 83, 0, 0, 0, 0, 3, 26, 38, 66, 64, 39, 14, 0, 0, 0, 0, 21, 26, 39, 75, 146, 213, 201, 83, 0, 
    164, 152, 130, 136, 166, 178, 150, 95, 60, 69, 44, 15, 13, 33, 53, 57, 12, 0, 0, 0, 0, 0, 0, 0, 9, 35, 56, 95, 165, 186, 97, 2, 
    144, 133, 141, 154, 150, 162, 178, 164, 135, 98, 75, 85, 96, 97, 89, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 40, 52, 108, 160, 127, 27, 
    129, 118, 147, 165, 140, 138, 185, 221, 186, 116, 112, 116, 108, 103, 91, 58, 20, 0, 0, 0, 0, 0, 0, 0, 0, 11, 36, 15, 41, 102, 134, 70, 
    139, 142, 156, 157, 144, 129, 135, 171, 192, 159, 160, 136, 109, 117, 120, 98, 69, 42, 24, 4, 0, 0, 0, 0, 0, 13, 17, 0, 28, 59, 80, 62, 
    137, 142, 141, 152, 174, 163, 126, 109, 146, 135, 103, 88, 101, 144, 156, 124, 90, 75, 70, 60, 54, 42, 34, 47, 46, 38, 31, 40, 88, 98, 61, 26, 
    137, 134, 114, 125, 161, 155, 127, 103, 124, 120, 106, 108, 112, 142, 152, 131, 100, 96, 105, 100, 90, 82, 88, 107, 105, 91, 87, 87, 94, 97, 71, 49, 
    132, 131, 109, 125, 152, 133, 118, 117, 124, 111, 112, 149, 141, 141, 145, 140, 117, 116, 113, 98, 96, 104, 116, 131, 128, 119, 117, 105, 79, 70, 92, 93, 
    114, 124, 138, 162, 162, 145, 143, 148, 156, 146, 153, 162, 140, 131, 127, 128, 119, 112, 101, 90, 104, 120, 128, 139, 141, 133, 127, 115, 95, 94, 127, 102, 
    133, 159, 172, 174, 143, 133, 143, 148, 149, 142, 158, 161, 141, 122, 99, 92, 100, 106, 108, 107, 118, 127, 131, 142, 149, 139, 131, 127, 114, 115, 128, 89, 
    67, 88, 91, 76, 43, 29, 41, 59, 61, 47, 50, 58, 58, 54, 36, 24, 33, 43, 53, 53, 56, 64, 65, 70, 75, 65, 59, 63, 65, 64, 65, 36, 
    
    -- channel=93
    183, 77, 81, 118, 141, 144, 147, 149, 145, 134, 131, 133, 126, 110, 94, 106, 105, 72, 52, 61, 75, 71, 59, 52, 49, 59, 79, 104, 88, 60, 55, 0, 
    229, 107, 130, 155, 152, 139, 156, 160, 156, 141, 128, 128, 119, 106, 99, 110, 99, 48, 23, 50, 77, 76, 69, 57, 55, 62, 79, 103, 91, 61, 65, 0, 
    251, 161, 183, 165, 130, 132, 158, 155, 158, 152, 139, 142, 130, 118, 116, 121, 104, 51, 6, 26, 67, 79, 86, 89, 99, 107, 108, 98, 76, 70, 82, 0, 
    266, 177, 188, 159, 131, 146, 167, 160, 163, 165, 158, 157, 144, 132, 137, 141, 124, 63, 5, 4, 51, 76, 76, 85, 112, 125, 115, 94, 74, 79, 96, 0, 
    274, 159, 161, 162, 137, 154, 176, 169, 172, 175, 166, 165, 153, 132, 128, 150, 149, 113, 53, 29, 67, 98, 80, 77, 101, 110, 108, 98, 87, 95, 107, 0, 
    276, 136, 159, 178, 153, 165, 173, 172, 179, 179, 174, 164, 163, 145, 123, 142, 159, 150, 122, 90, 106, 130, 105, 88, 106, 105, 96, 103, 105, 108, 118, 0, 
    255, 124, 171, 184, 167, 169, 177, 183, 182, 186, 181, 173, 173, 166, 141, 140, 159, 161, 157, 138, 126, 131, 107, 77, 89, 82, 77, 97, 107, 109, 117, 0, 
    234, 132, 163, 180, 166, 169, 177, 187, 191, 183, 179, 179, 176, 164, 145, 138, 150, 162, 172, 166, 132, 127, 108, 62, 69, 75, 81, 96, 104, 109, 113, 0, 
    233, 135, 175, 178, 171, 174, 170, 176, 186, 187, 183, 173, 165, 157, 151, 143, 130, 135, 158, 177, 152, 151, 143, 71, 59, 88, 100, 109, 113, 110, 113, 0, 
    206, 142, 186, 181, 185, 185, 175, 175, 184, 187, 182, 174, 168, 168, 187, 183, 140, 115, 139, 168, 161, 158, 140, 55, 50, 93, 96, 97, 105, 110, 114, 0, 
    134, 146, 188, 165, 180, 197, 188, 184, 187, 178, 179, 187, 189, 172, 196, 221, 170, 114, 130, 161, 153, 140, 97, 21, 45, 86, 80, 76, 90, 106, 114, 0, 
    71, 164, 214, 165, 185, 196, 186, 190, 167, 153, 181, 225, 228, 186, 164, 150, 140, 125, 131, 168, 156, 119, 57, 3, 26, 76, 75, 75, 90, 105, 108, 0, 
    63, 189, 232, 205, 238, 231, 209, 186, 148, 159, 215, 245, 221, 174, 141, 98, 95, 119, 128, 164, 150, 97, 43, 9, 31, 59, 64, 68, 83, 96, 100, 0, 
    107, 162, 193, 224, 244, 214, 202, 190, 160, 189, 236, 224, 181, 165, 183, 157, 175, 193, 179, 189, 138, 83, 38, 11, 27, 48, 71, 73, 74, 83, 84, 0, 
    149, 116, 160, 228, 246, 203, 191, 192, 199, 233, 257, 224, 177, 174, 222, 227, 232, 248, 232, 209, 161, 94, 41, 25, 30, 57, 104, 103, 70, 61, 75, 0, 
    177, 91, 133, 237, 252, 205, 174, 186, 227, 263, 259, 236, 214, 209, 249, 255, 234, 233, 232, 226, 183, 105, 40, 19, 21, 68, 137, 148, 87, 40, 62, 0, 
    202, 116, 158, 234, 240, 210, 158, 158, 242, 256, 205, 228, 237, 205, 215, 221, 220, 213, 207, 203, 166, 82, 9, 0, 0, 65, 154, 181, 107, 29, 41, 0, 
    223, 138, 171, 250, 255, 223, 159, 126, 235, 240, 160, 208, 227, 161, 156, 163, 158, 170, 141, 120, 78, 6, 0, 0, 0, 72, 162, 195, 130, 21, 14, 0, 
    231, 128, 160, 245, 262, 240, 167, 65, 162, 241, 183, 221, 230, 140, 154, 161, 116, 92, 52, 28, 2, 0, 0, 0, 15, 86, 175, 219, 171, 27, 0, 0, 
    236, 129, 153, 231, 260, 244, 182, 25, 44, 184, 202, 226, 188, 117, 188, 248, 175, 88, 10, 8, 20, 25, 51, 30, 21, 86, 182, 246, 210, 59, 0, 0, 
    252, 149, 163, 236, 259, 226, 157, 0, 0, 66, 93, 122, 126, 97, 155, 219, 151, 77, 11, 1, 28, 42, 69, 46, 20, 72, 166, 255, 245, 89, 0, 0, 
    266, 157, 153, 206, 231, 195, 111, 0, 0, 23, 12, 9, 39, 58, 107, 129, 61, 21, 0, 0, 1, 0, 25, 47, 48, 76, 143, 229, 250, 113, 0, 0, 
    261, 153, 156, 184, 203, 174, 104, 57, 50, 53, 46, 45, 50, 68, 91, 59, 0, 0, 0, 0, 0, 0, 0, 18, 40, 75, 109, 173, 225, 142, 0, 0, 
    231, 152, 184, 184, 170, 174, 170, 142, 96, 79, 89, 104, 115, 118, 100, 39, 0, 0, 0, 0, 0, 0, 0, 0, 13, 65, 72, 102, 184, 169, 58, 0, 
    221, 157, 190, 180, 150, 161, 204, 214, 140, 107, 130, 120, 121, 130, 104, 45, 0, 0, 0, 0, 0, 0, 0, 0, 12, 62, 46, 44, 115, 148, 116, 0, 
    231, 174, 194, 182, 155, 146, 154, 187, 164, 128, 151, 136, 141, 158, 130, 88, 55, 35, 19, 7, 0, 0, 0, 0, 16, 42, 27, 36, 95, 104, 89, 0, 
    235, 165, 162, 193, 196, 158, 125, 143, 158, 114, 96, 98, 142, 187, 166, 116, 84, 81, 74, 60, 49, 39, 53, 65, 54, 51, 44, 71, 131, 99, 78, 0, 
    239, 142, 133, 187, 194, 148, 115, 134, 150, 99, 121, 136, 148, 183, 171, 129, 107, 115, 113, 103, 99, 94, 112, 124, 104, 93, 96, 106, 116, 92, 98, 0, 
    227, 147, 143, 184, 177, 144, 130, 144, 145, 119, 141, 169, 166, 175, 170, 148, 129, 133, 122, 118, 126, 128, 145, 152, 134, 125, 127, 109, 89, 99, 130, 2, 
    222, 158, 174, 193, 178, 162, 165, 177, 166, 162, 187, 178, 153, 150, 145, 147, 139, 130, 117, 118, 139, 149, 157, 167, 155, 144, 139, 114, 99, 126, 170, 3, 
    239, 198, 200, 177, 145, 157, 179, 184, 162, 156, 184, 175, 155, 132, 106, 116, 130, 132, 127, 131, 153, 156, 158, 173, 165, 150, 147, 138, 127, 145, 162, 0, 
    121, 107, 103, 76, 48, 56, 71, 79, 69, 63, 67, 68, 66, 55, 36, 40, 52, 59, 63, 64, 73, 77, 78, 86, 83, 70, 71, 70, 70, 76, 78, 0, 
    
    -- channel=94
    35, 7, 1, 23, 35, 33, 33, 34, 40, 34, 35, 38, 34, 23, 21, 27, 18, 3, 0, 3, 5, 3, 0, 1, 5, 5, 4, 12, 0, 0, 0, 0, 
    130, 107, 89, 109, 127, 136, 141, 144, 147, 137, 133, 136, 133, 123, 109, 113, 102, 74, 56, 61, 69, 66, 59, 50, 50, 51, 61, 80, 76, 55, 52, 0, 
    143, 134, 143, 139, 134, 142, 149, 152, 152, 146, 141, 138, 130, 130, 121, 116, 114, 79, 55, 60, 70, 72, 71, 63, 56, 59, 69, 78, 80, 71, 60, 0, 
    155, 162, 175, 157, 140, 144, 152, 150, 154, 158, 149, 147, 141, 135, 138, 135, 121, 88, 41, 42, 62, 70, 75, 84, 91, 90, 87, 80, 72, 74, 73, 0, 
    157, 161, 178, 162, 143, 152, 163, 158, 162, 165, 162, 163, 156, 143, 147, 157, 138, 108, 52, 26, 49, 59, 58, 71, 89, 100, 99, 89, 72, 74, 84, 3, 
    151, 151, 163, 159, 147, 154, 168, 171, 169, 170, 169, 170, 161, 146, 138, 159, 164, 146, 102, 52, 57, 79, 69, 69, 83, 91, 100, 98, 87, 84, 89, 7, 
    152, 150, 151, 165, 157, 159, 167, 171, 172, 176, 172, 170, 171, 159, 140, 148, 163, 164, 149, 114, 96, 120, 102, 83, 89, 85, 91, 98, 97, 95, 96, 12, 
    152, 131, 153, 166, 163, 166, 169, 178, 178, 180, 180, 177, 176, 171, 158, 150, 154, 167, 168, 155, 126, 128, 107, 83, 85, 79, 72, 82, 92, 94, 98, 13, 
    138, 132, 156, 157, 160, 165, 169, 184, 186, 179, 175, 174, 170, 160, 156, 142, 138, 153, 166, 165, 143, 139, 117, 79, 78, 78, 76, 82, 90, 91, 97, 12, 
    135, 152, 150, 155, 164, 167, 168, 170, 180, 180, 178, 173, 162, 145, 144, 131, 117, 121, 147, 163, 157, 157, 140, 88, 80, 83, 92, 95, 96, 94, 94, 12, 
    134, 152, 150, 163, 179, 179, 172, 170, 177, 189, 190, 170, 141, 127, 152, 156, 121, 104, 123, 142, 146, 149, 134, 93, 74, 81, 83, 87, 93, 95, 96, 13, 
    91, 141, 150, 144, 155, 168, 174, 177, 174, 179, 186, 177, 151, 130, 141, 172, 162, 116, 118, 130, 124, 124, 97, 61, 61, 77, 78, 78, 86, 90, 96, 16, 
    40, 137, 165, 155, 161, 173, 172, 169, 161, 165, 180, 194, 184, 147, 115, 102, 126, 108, 105, 127, 112, 100, 70, 40, 46, 64, 74, 75, 81, 86, 92, 15, 
    24, 115, 178, 189, 193, 183, 178, 162, 144, 156, 178, 189, 184, 161, 128, 76, 77, 96, 101, 111, 106, 83, 53, 33, 31, 47, 63, 65, 76, 79, 85, 13, 
    50, 95, 150, 188, 192, 173, 174, 173, 151, 165, 184, 173, 151, 157, 164, 138, 125, 138, 134, 127, 106, 70, 45, 29, 29, 48, 66, 61, 61, 70, 74, 8, 
    81, 75, 120, 182, 190, 172, 162, 179, 180, 185, 189, 183, 157, 164, 191, 186, 175, 174, 174, 158, 118, 77, 54, 38, 41, 59, 84, 84, 51, 55, 69, 3, 
    99, 81, 107, 166, 185, 170, 141, 165, 199, 191, 200, 210, 185, 172, 198, 209, 192, 179, 185, 180, 155, 106, 62, 41, 36, 65, 105, 117, 70, 37, 59, 5, 
    110, 106, 131, 166, 173, 168, 135, 143, 209, 186, 172, 186, 177, 162, 189, 187, 194, 178, 171, 176, 155, 103, 49, 20, 18, 57, 114, 129, 92, 28, 41, 2, 
    117, 119, 152, 184, 181, 169, 131, 101, 199, 192, 133, 166, 175, 141, 145, 120, 125, 141, 122, 114, 86, 49, 20, 2, 14, 54, 117, 141, 103, 26, 22, 0, 
    119, 109, 130, 181, 190, 175, 134, 60, 134, 208, 170, 180, 174, 129, 148, 145, 95, 86, 69, 54, 27, 13, 22, 14, 25, 69, 126, 160, 128, 29, 2, 0, 
    121, 111, 128, 177, 191, 179, 144, 50, 45, 132, 177, 181, 160, 124, 166, 202, 148, 88, 45, 39, 35, 32, 48, 32, 23, 63, 130, 180, 163, 54, 0, 0, 
    130, 125, 136, 172, 190, 170, 128, 51, 0, 15, 66, 99, 109, 94, 118, 151, 143, 104, 50, 32, 38, 37, 55, 51, 30, 55, 118, 189, 188, 91, 9, 0, 
    137, 133, 124, 152, 179, 155, 104, 50, 17, 10, 5, 14, 32, 49, 65, 85, 79, 68, 46, 22, 15, 7, 27, 53, 58, 69, 95, 165, 198, 117, 19, 0, 
    136, 138, 128, 132, 159, 157, 107, 72, 64, 66, 43, 40, 39, 53, 69, 53, 16, 4, 1, 0, 0, 0, 0, 15, 47, 64, 72, 123, 185, 146, 40, 0, 
    119, 129, 145, 141, 136, 155, 159, 138, 89, 80, 75, 82, 92, 88, 78, 44, 2, 0, 0, 0, 0, 0, 0, 0, 14, 49, 58, 81, 139, 164, 96, 0, 
    116, 132, 147, 147, 123, 126, 166, 192, 127, 108, 125, 104, 107, 103, 87, 65, 34, 9, 0, 0, 0, 0, 0, 0, 0, 40, 43, 41, 76, 104, 127, 16, 
    124, 135, 146, 156, 138, 120, 119, 163, 163, 115, 123, 109, 112, 122, 112, 88, 72, 51, 30, 16, 6, 0, 0, 5, 11, 25, 27, 36, 66, 61, 85, 20, 
    119, 121, 131, 155, 155, 136, 110, 118, 142, 118, 92, 90, 113, 136, 131, 104, 90, 82, 68, 62, 56, 47, 52, 57, 51, 45, 49, 65, 96, 88, 62, 0, 
    128, 117, 107, 129, 145, 129, 112, 110, 110, 104, 102, 107, 117, 134, 136, 120, 105, 103, 98, 95, 90, 89, 100, 103, 93, 89, 88, 86, 92, 90, 86, 0, 
    119, 120, 110, 123, 133, 123, 117, 125, 117, 104, 118, 127, 128, 134, 138, 137, 124, 115, 102, 100, 111, 113, 123, 128, 117, 114, 110, 98, 83, 92, 114, 20, 
    114, 133, 138, 138, 136, 143, 141, 142, 138, 141, 145, 142, 134, 127, 121, 132, 128, 116, 102, 103, 118, 122, 129, 137, 129, 123, 122, 106, 94, 105, 121, 25, 
    145, 176, 180, 163, 140, 142, 156, 163, 157, 154, 161, 159, 155, 142, 118, 118, 130, 135, 133, 131, 139, 147, 151, 160, 158, 148, 145, 142, 135, 136, 142, 62, 
    
    -- channel=95
    52, 0, 7, 32, 36, 33, 36, 41, 39, 31, 33, 39, 33, 26, 26, 31, 23, 5, 4, 18, 25, 22, 17, 19, 18, 16, 21, 31, 19, 7, 13, 0, 
    139, 101, 87, 90, 118, 139, 149, 143, 140, 140, 134, 136, 139, 128, 111, 110, 106, 84, 69, 76, 89, 89, 83, 72, 73, 81, 87, 95, 96, 77, 71, 32, 
    149, 118, 116, 116, 126, 138, 151, 149, 149, 148, 139, 140, 138, 139, 132, 126, 117, 89, 70, 74, 89, 93, 92, 84, 80, 81, 86, 95, 99, 87, 83, 41, 
    157, 133, 140, 134, 128, 136, 145, 146, 151, 153, 147, 150, 143, 140, 145, 137, 131, 103, 66, 62, 82, 91, 98, 104, 107, 107, 105, 97, 92, 97, 94, 41, 
    154, 137, 142, 143, 134, 139, 150, 149, 150, 159, 154, 153, 153, 148, 149, 159, 146, 120, 71, 46, 68, 87, 89, 98, 118, 124, 119, 110, 95, 95, 102, 52, 
    153, 123, 131, 142, 131, 140, 155, 156, 157, 158, 156, 158, 159, 150, 142, 159, 163, 141, 103, 62, 73, 95, 91, 92, 108, 118, 120, 118, 108, 100, 106, 54, 
    149, 114, 129, 139, 136, 144, 151, 159, 158, 158, 156, 160, 165, 158, 143, 143, 160, 157, 142, 112, 99, 116, 115, 103, 113, 113, 113, 119, 118, 113, 113, 58, 
    142, 116, 127, 138, 143, 147, 155, 158, 156, 159, 167, 166, 170, 169, 158, 146, 153, 157, 157, 153, 133, 130, 127, 101, 104, 106, 104, 112, 115, 115, 116, 61, 
    149, 109, 123, 139, 144, 148, 152, 160, 162, 159, 171, 175, 169, 162, 161, 151, 145, 152, 165, 169, 155, 134, 120, 89, 88, 104, 102, 101, 107, 111, 114, 60, 
    135, 114, 135, 141, 143, 148, 147, 152, 164, 166, 167, 162, 157, 149, 150, 140, 122, 126, 154, 170, 163, 148, 133, 89, 81, 101, 106, 107, 110, 111, 114, 61, 
    120, 132, 147, 140, 150, 155, 154, 150, 156, 160, 162, 150, 140, 131, 140, 139, 113, 106, 130, 155, 157, 145, 129, 90, 81, 97, 100, 106, 109, 115, 114, 59, 
    101, 135, 144, 130, 151, 162, 153, 153, 153, 153, 159, 147, 123, 98, 116, 147, 130, 111, 118, 135, 135, 127, 104, 83, 77, 90, 93, 93, 100, 110, 116, 62, 
    69, 126, 151, 136, 141, 142, 143, 147, 144, 141, 147, 140, 126, 107, 92, 104, 130, 125, 111, 126, 121, 107, 90, 60, 61, 80, 90, 92, 100, 106, 112, 62, 
    52, 109, 154, 159, 159, 151, 147, 137, 128, 135, 141, 132, 134, 130, 119, 83, 80, 102, 88, 104, 105, 88, 76, 55, 56, 66, 80, 87, 94, 101, 107, 60, 
    73, 89, 140, 165, 164, 146, 147, 144, 130, 130, 139, 128, 130, 139, 145, 127, 96, 103, 105, 98, 93, 81, 63, 51, 50, 60, 80, 83, 84, 91, 97, 56, 
    103, 99, 125, 158, 163, 145, 134, 146, 146, 140, 147, 146, 134, 136, 152, 149, 131, 134, 129, 123, 108, 80, 59, 50, 50, 66, 95, 95, 74, 75, 88, 49, 
    131, 107, 114, 152, 162, 148, 130, 132, 153, 153, 144, 158, 163, 152, 162, 159, 146, 142, 143, 147, 125, 87, 61, 51, 53, 75, 104, 119, 85, 55, 76, 48, 
    145, 134, 129, 146, 155, 147, 122, 111, 152, 146, 128, 163, 176, 149, 144, 158, 159, 151, 141, 141, 130, 102, 64, 50, 44, 71, 109, 125, 103, 51, 53, 43, 
    153, 138, 145, 166, 157, 142, 120, 92, 140, 158, 121, 142, 152, 125, 137, 138, 132, 143, 123, 114, 100, 81, 63, 43, 39, 65, 110, 128, 106, 50, 35, 32, 
    154, 137, 139, 165, 162, 143, 119, 63, 97, 177, 140, 135, 152, 136, 147, 144, 94, 100, 91, 74, 62, 53, 57, 47, 46, 77, 115, 143, 114, 46, 17, 23, 
    158, 143, 130, 149, 155, 142, 123, 62, 35, 131, 163, 147, 145, 134, 152, 198, 153, 98, 72, 62, 61, 52, 65, 63, 53, 86, 125, 149, 134, 62, 7, 10, 
    162, 144, 140, 157, 157, 136, 115, 72, 26, 42, 85, 112, 125, 121, 134, 175, 167, 124, 76, 51, 59, 61, 74, 79, 63, 75, 114, 153, 151, 87, 19, 7, 
    165, 147, 143, 152, 153, 132, 100, 74, 53, 34, 28, 45, 70, 94, 110, 112, 98, 90, 71, 41, 36, 37, 48, 78, 78, 82, 100, 142, 161, 110, 38, 6, 
    160, 156, 152, 143, 143, 132, 109, 87, 67, 74, 78, 69, 67, 84, 92, 79, 53, 34, 35, 29, 26, 20, 17, 40, 67, 90, 96, 112, 157, 136, 60, 5, 
    153, 156, 168, 149, 130, 142, 140, 113, 88, 95, 109, 111, 117, 115, 111, 83, 39, 14, 8, 11, 14, 15, 10, 11, 40, 73, 80, 86, 134, 154, 103, 11, 
    153, 146, 159, 163, 135, 124, 150, 164, 133, 104, 114, 114, 133, 141, 122, 90, 60, 39, 26, 18, 13, 7, 9, 15, 30, 57, 68, 73, 95, 123, 130, 46, 
    156, 158, 160, 164, 153, 119, 112, 152, 153, 104, 121, 131, 133, 145, 132, 112, 93, 74, 59, 45, 32, 21, 25, 34, 32, 46, 63, 68, 86, 71, 86, 69, 
    155, 149, 146, 165, 167, 145, 118, 113, 146, 115, 100, 120, 129, 152, 155, 133, 113, 104, 92, 79, 74, 70, 72, 75, 69, 66, 70, 79, 99, 97, 77, 49, 
    151, 139, 132, 154, 161, 146, 140, 126, 118, 127, 129, 127, 128, 151, 160, 149, 127, 119, 115, 115, 117, 113, 114, 118, 112, 105, 103, 100, 98, 118, 115, 46, 
    149, 151, 140, 143, 153, 150, 142, 142, 130, 117, 132, 148, 146, 151, 154, 154, 140, 130, 129, 134, 139, 136, 138, 144, 136, 131, 127, 117, 107, 110, 124, 67, 
    144, 153, 152, 154, 152, 157, 157, 153, 153, 142, 147, 154, 152, 145, 139, 146, 147, 140, 134, 130, 140, 145, 146, 152, 148, 141, 137, 130, 117, 119, 134, 76, 
    143, 160, 159, 152, 139, 148, 161, 158, 144, 144, 154, 158, 153, 136, 117, 121, 137, 137, 132, 128, 135, 141, 142, 147, 148, 139, 140, 136, 126, 124, 132, 74, 
    
    -- channel=96
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=97
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 34, 39, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 56, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 71, 33, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 70, 63, 17, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 35, 67, 67, 61, 35, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 23, 28, 33, 49, 74, 74, 56, 31, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 37, 51, 56, 64, 75, 74, 60, 38, 7, 0, 0, 0, 0, 0, 7, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 61, 57, 61, 65, 65, 68, 53, 0, 0, 0, 0, 0, 7, 22, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 53, 61, 60, 60, 57, 56, 66, 64, 29, 0, 0, 14, 27, 33, 21, 5, 0, 
    0, 0, 0, 0, 18, 23, 0, 0, 0, 0, 0, 0, 0, 0, 26, 58, 62, 60, 50, 27, 7, 9, 37, 56, 49, 46, 48, 42, 32, 13, 0, 0, 
    0, 0, 0, 0, 47, 34, 1, 0, 0, 0, 0, 0, 0, 0, 26, 58, 61, 51, 32, 5, 0, 0, 0, 28, 62, 61, 48, 37, 18, 0, 0, 0, 
    0, 0, 0, 0, 11, 25, 6, 0, 0, 0, 0, 0, 0, 7, 34, 59, 58, 45, 23, 0, 0, 0, 0, 0, 30, 48, 42, 21, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 16, 7, 0, 0, 0, 0, 0, 7, 26, 52, 65, 59, 47, 3, 0, 0, 0, 0, 0, 2, 38, 32, 12, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 18, 13, 0, 0, 0, 0, 0, 13, 25, 50, 63, 61, 44, 0, 0, 0, 0, 0, 0, 0, 22, 31, 11, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 13, 0, 0, 0, 0, 16, 16, 22, 50, 57, 59, 37, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 17, 22, 0, 0, 5, 32, 51, 47, 50, 60, 59, 61, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 10, 0, 0, 0, 7, 17, 20, 25, 23, 22, 30, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 12, 10, 9, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=98
    271, 210, 210, 218, 242, 246, 240, 249, 249, 231, 221, 221, 226, 224, 206, 194, 198, 203, 211, 176, 135, 156, 156, 140, 119, 111, 114, 128, 133, 127, 135, 79, 
    351, 289, 288, 292, 320, 328, 322, 329, 329, 310, 293, 286, 289, 289, 273, 257, 253, 249, 238, 216, 215, 213, 198, 189, 153, 103, 119, 176, 173, 155, 162, 98, 
    376, 315, 307, 296, 296, 298, 294, 290, 286, 272, 258, 249, 253, 255, 244, 233, 228, 222, 208, 193, 203, 207, 186, 169, 136, 86, 103, 166, 175, 159, 163, 95, 
    347, 301, 290, 272, 259, 253, 258, 248, 243, 236, 226, 219, 223, 224, 218, 212, 208, 204, 200, 193, 192, 191, 153, 129, 122, 97, 114, 154, 166, 155, 158, 90, 
    315, 263, 260, 244, 234, 228, 227, 215, 214, 213, 205, 199, 200, 201, 202, 200, 196, 193, 192, 193, 202, 175, 109, 80, 103, 113, 140, 161, 157, 150, 146, 84, 
    294, 236, 221, 212, 210, 210, 203, 193, 197, 200, 195, 186, 184, 185, 193, 196, 192, 191, 189, 197, 214, 170, 90, 99, 109, 120, 164, 173, 168, 159, 146, 86, 
    252, 208, 194, 191, 188, 186, 184, 180, 188, 192, 192, 183, 181, 181, 188, 193, 192, 193, 187, 194, 196, 129, 82, 149, 166, 146, 176, 178, 182, 172, 160, 94, 
    217, 185, 176, 180, 180, 178, 176, 174, 183, 187, 190, 184, 187, 184, 185, 184, 185, 193, 187, 183, 154, 82, 70, 161, 198, 171, 171, 175, 178, 175, 169, 96, 
    207, 174, 170, 176, 177, 178, 177, 173, 181, 187, 192, 184, 187, 188, 187, 189, 187, 199, 193, 170, 122, 62, 62, 137, 178, 165, 174, 176, 175, 175, 168, 92, 
    207, 170, 169, 174, 175, 176, 179, 175, 180, 189, 200, 194, 202, 200, 184, 188, 176, 163, 138, 64, 35, 37, 40, 116, 159, 142, 159, 172, 171, 174, 165, 88, 
    212, 170, 167, 171, 174, 173, 177, 175, 181, 185, 198, 196, 198, 175, 121, 125, 136, 144, 136, 52, 8, 0, 0, 37, 169, 172, 141, 134, 158, 170, 161, 88, 
    217, 173, 169, 170, 173, 171, 174, 175, 180, 187, 184, 178, 189, 181, 145, 162, 187, 195, 200, 190, 211, 106, 0, 0, 93, 200, 194, 103, 120, 159, 157, 89, 
    220, 176, 172, 170, 174, 167, 173, 176, 184, 187, 178, 184, 198, 165, 136, 171, 200, 175, 161, 240, 340, 230, 0, 0, 0, 141, 215, 138, 94, 147, 154, 90, 
    220, 176, 173, 170, 174, 161, 168, 181, 188, 182, 154, 157, 166, 111, 53, 85, 152, 128, 103, 225, 303, 204, 40, 0, 0, 39, 162, 155, 109, 137, 155, 93, 
    221, 177, 175, 167, 172, 163, 143, 158, 161, 145, 120, 136, 137, 73, 35, 54, 118, 135, 114, 191, 210, 132, 86, 0, 0, 0, 84, 120, 134, 120, 104, 71, 
    221, 175, 175, 164, 168, 183, 150, 110, 116, 82, 109, 147, 134, 83, 77, 58, 51, 87, 114, 137, 119, 100, 60, 0, 0, 10, 27, 113, 170, 118, 13, 2, 
    220, 170, 172, 163, 158, 184, 189, 132, 108, 76, 83, 159, 150, 176, 219, 146, 84, 108, 121, 113, 107, 82, 7, 0, 88, 109, 34, 116, 193, 129, 0, 0, 
    219, 164, 169, 172, 118, 95, 139, 153, 120, 67, 78, 144, 123, 219, 342, 219, 121, 140, 144, 137, 126, 42, 0, 0, 85, 105, 64, 101, 155, 128, 0, 0, 
    218, 164, 191, 188, 63, 0, 74, 135, 91, 49, 98, 148, 130, 210, 317, 192, 112, 127, 135, 136, 141, 78, 0, 0, 25, 82, 84, 91, 101, 112, 7, 0, 
    213, 184, 245, 199, 7, 0, 19, 110, 67, 40, 102, 153, 173, 248, 278, 147, 100, 115, 98, 109, 188, 238, 137, 4, 20, 67, 73, 79, 84, 76, 18, 0, 
    206, 222, 303, 216, 19, 0, 0, 80, 59, 52, 108, 130, 154, 264, 272, 127, 106, 87, 24, 50, 160, 271, 325, 211, 81, 55, 74, 88, 70, 48, 42, 46, 
    208, 228, 258, 211, 152, 5, 0, 52, 42, 74, 129, 127, 107, 202, 236, 120, 105, 21, 0, 31, 105, 135, 274, 340, 179, 68, 74, 76, 47, 38, 89, 87, 
    213, 197, 135, 125, 219, 74, 0, 33, 49, 93, 154, 167, 129, 188, 190, 105, 72, 0, 0, 80, 98, 84, 148, 298, 246, 88, 56, 24, 7, 67, 124, 83, 
    207, 176, 108, 87, 188, 103, 0, 6, 71, 111, 149, 152, 150, 215, 181, 103, 46, 0, 0, 96, 68, 72, 92, 212, 276, 137, 23, 0, 13, 106, 136, 77, 
    188, 166, 141, 106, 165, 118, 0, 2, 96, 136, 131, 100, 140, 217, 163, 113, 39, 0, 0, 116, 62, 44, 50, 145, 274, 196, 17, 0, 52, 132, 146, 87, 
    168, 152, 147, 114, 156, 123, 0, 0, 97, 131, 109, 58, 83, 143, 114, 99, 25, 0, 0, 141, 82, 8, 11, 81, 228, 215, 37, 0, 79, 131, 141, 93, 
    161, 141, 149, 116, 138, 124, 21, 38, 129, 170, 175, 149, 145, 163, 158, 154, 94, 0, 16, 147, 132, 48, 18, 60, 160, 196, 83, 49, 92, 118, 134, 92, 
    167, 129, 140, 140, 139, 132, 81, 105, 153, 175, 190, 190, 193, 196, 189, 185, 160, 83, 108, 151, 96, 72, 29, 50, 107, 136, 101, 94, 104, 109, 127, 90, 
    175, 125, 106, 106, 116, 108, 86, 85, 97, 109, 115, 114, 118, 121, 119, 117, 117, 103, 151, 194, 110, 58, 37, 39, 92, 105, 100, 104, 110, 114, 123, 84, 
    183, 127, 99, 73, 64, 66, 65, 37, 39, 71, 77, 70, 69, 70, 72, 70, 74, 78, 110, 162, 160, 97, 53, 67, 97, 101, 99, 103, 111, 120, 123, 77, 
    178, 123, 108, 84, 55, 45, 48, 18, 21, 62, 68, 63, 60, 56, 56, 52, 52, 57, 70, 94, 101, 67, 54, 85, 98, 95, 92, 98, 108, 116, 116, 70, 
    180, 156, 171, 178, 165, 142, 127, 99, 98, 126, 127, 127, 129, 127, 126, 119, 111, 108, 110, 119, 120, 95, 83, 102, 115, 114, 109, 112, 123, 130, 128, 98, 
    
    -- channel=99
    15, 14, 16, 18, 20, 24, 25, 25, 24, 23, 20, 17, 15, 16, 17, 13, 10, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=100
    20, 218, 241, 247, 235, 249, 264, 257, 253, 261, 253, 234, 220, 219, 231, 225, 204, 171, 122, 166, 148, 151, 140, 136, 135, 95, 82, 60, 76, 105, 108, 123, 
    0, 280, 303, 299, 268, 279, 301, 287, 280, 293, 290, 269, 247, 243, 263, 263, 238, 199, 142, 172, 169, 175, 171, 153, 140, 104, 46, 11, 66, 136, 146, 178, 
    0, 295, 312, 307, 278, 283, 293, 281, 272, 278, 274, 257, 233, 227, 243, 242, 223, 205, 203, 191, 164, 175, 175, 132, 117, 102, 30, 0, 57, 147, 157, 191, 
    0, 295, 297, 294, 282, 276, 275, 268, 256, 252, 248, 234, 214, 212, 222, 219, 208, 195, 193, 189, 173, 167, 180, 155, 115, 82, 38, 4, 83, 165, 172, 204, 
    0, 254, 243, 240, 248, 245, 248, 247, 231, 222, 221, 213, 200, 201, 206, 203, 198, 190, 190, 188, 167, 145, 184, 174, 120, 88, 51, 52, 126, 185, 184, 210, 
    0, 190, 191, 208, 218, 215, 220, 224, 210, 201, 202, 201, 198, 201, 199, 197, 196, 190, 193, 181, 110, 87, 118, 97, 81, 96, 61, 84, 136, 178, 180, 208, 
    0, 170, 187, 196, 197, 195, 202, 208, 197, 191, 192, 199, 202, 207, 203, 200, 200, 196, 206, 174, 83, 79, 56, 0, 14, 74, 68, 103, 138, 172, 178, 207, 
    0, 173, 185, 184, 186, 190, 194, 200, 192, 191, 194, 203, 205, 214, 220, 222, 219, 204, 209, 163, 112, 127, 55, 0, 0, 86, 120, 151, 161, 177, 176, 208, 
    0, 170, 185, 185, 188, 191, 192, 199, 192, 192, 199, 211, 205, 210, 206, 207, 199, 175, 177, 152, 153, 155, 80, 0, 22, 133, 172, 175, 169, 167, 170, 211, 
    0, 171, 189, 191, 194, 194, 192, 200, 192, 186, 180, 184, 160, 154, 168, 191, 219, 233, 261, 282, 270, 180, 98, 21, 35, 149, 174, 170, 165, 158, 162, 210, 
    0, 179, 195, 197, 198, 199, 193, 199, 191, 176, 153, 156, 141, 180, 241, 252, 241, 211, 190, 264, 253, 207, 220, 83, 0, 61, 118, 172, 165, 149, 152, 205, 
    0, 188, 200, 200, 199, 201, 194, 197, 185, 172, 158, 158, 109, 92, 87, 27, 0, 0, 0, 0, 0, 90, 355, 234, 9, 0, 15, 140, 176, 147, 147, 197, 
    0, 195, 201, 200, 197, 202, 194, 190, 176, 148, 121, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 359, 393, 162, 0, 0, 67, 145, 129, 136, 189, 
    0, 200, 200, 202, 197, 205, 192, 173, 133, 86, 46, 0, 0, 0, 39, 0, 0, 0, 18, 0, 0, 0, 214, 420, 325, 35, 0, 0, 70, 82, 110, 175, 
    0, 197, 198, 204, 196, 210, 206, 166, 93, 66, 52, 27, 4, 77, 109, 55, 0, 30, 62, 0, 0, 0, 65, 316, 378, 144, 0, 0, 9, 59, 129, 189, 
    0, 193, 197, 208, 186, 165, 175, 139, 112, 90, 79, 0, 0, 80, 99, 131, 132, 131, 80, 0, 0, 0, 21, 183, 222, 125, 74, 0, 0, 56, 206, 233, 
    0, 194, 196, 198, 156, 60, 33, 51, 54, 73, 13, 0, 0, 0, 0, 56, 115, 46, 0, 0, 5, 10, 92, 150, 48, 77, 125, 18, 0, 30, 270, 295, 
    0, 196, 191, 180, 168, 92, 0, 0, 0, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 103, 291, 283, 84, 86, 160, 34, 0, 0, 271, 335, 
    0, 198, 177, 144, 234, 206, 11, 0, 0, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 137, 370, 353, 172, 97, 83, 9, 0, 0, 223, 310, 
    0, 186, 92, 71, 269, 258, 57, 0, 24, 59, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 83, 204, 128, 48, 18, 15, 19, 8, 170, 219, 
    4, 103, 0, 0, 179, 244, 96, 0, 42, 43, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 19, 30, 12, 0, 1, 47, 113, 120, 
    0, 0, 0, 0, 0, 142, 106, 6, 61, 26, 0, 0, 0, 0, 0, 0, 0, 42, 164, 57, 0, 0, 0, 0, 0, 4, 0, 0, 32, 72, 58, 69, 
    0, 2, 0, 0, 0, 62, 119, 60, 57, 1, 0, 0, 0, 0, 0, 0, 2, 198, 227, 29, 0, 0, 0, 0, 0, 0, 14, 48, 103, 73, 15, 62, 
    0, 62, 113, 0, 0, 0, 144, 93, 36, 0, 0, 0, 0, 0, 0, 0, 51, 285, 179, 0, 13, 32, 0, 0, 0, 0, 50, 143, 120, 20, 0, 77, 
    0, 66, 55, 0, 0, 0, 156, 104, 0, 0, 0, 0, 0, 0, 0, 0, 87, 292, 128, 0, 40, 51, 29, 0, 0, 0, 75, 164, 62, 0, 0, 76, 
    0, 49, 2, 0, 0, 0, 157, 120, 0, 0, 0, 44, 0, 0, 0, 0, 124, 292, 107, 0, 31, 105, 105, 0, 0, 0, 68, 125, 13, 0, 0, 67, 
    0, 45, 0, 0, 0, 0, 102, 44, 0, 0, 0, 0, 0, 0, 0, 0, 2, 190, 63, 0, 0, 55, 79, 0, 0, 0, 20, 56, 0, 0, 0, 50, 
    0, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 0, 0, 0, 44, 70, 52, 0, 0, 0, 10, 0, 0, 0, 35, 
    0, 79, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 84, 55, 0, 0, 0, 0, 0, 0, 0, 35, 
    0, 68, 83, 66, 38, 38, 50, 62, 45, 1, 0, 5, 8, 8, 9, 11, 10, 13, 0, 0, 0, 0, 41, 38, 0, 0, 0, 0, 0, 0, 0, 42, 
    0, 53, 69, 75, 68, 43, 27, 61, 48, 0, 0, 5, 17, 30, 38, 45, 47, 43, 15, 0, 0, 17, 58, 25, 0, 0, 1, 0, 0, 0, 0, 48, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    
    -- channel=101
    79, 90, 89, 90, 99, 102, 100, 102, 102, 94, 88, 84, 84, 84, 77, 69, 66, 71, 81, 65, 59, 53, 48, 46, 45, 23, 10, 23, 23, 22, 24, 0, 
    79, 61, 49, 39, 41, 35, 26, 27, 24, 18, 15, 15, 18, 18, 11, 9, 11, 14, 11, 0, 0, 0, 0, 7, 5, 0, 0, 0, 0, 2, 5, 0, 
    62, 39, 32, 29, 25, 16, 14, 15, 15, 12, 10, 10, 14, 13, 8, 7, 8, 10, 10, 4, 5, 8, 11, 11, 0, 0, 0, 0, 1, 2, 5, 0, 
    51, 27, 26, 22, 16, 11, 10, 10, 11, 9, 8, 8, 11, 11, 8, 7, 8, 8, 10, 10, 19, 28, 9, 0, 0, 0, 0, 13, 11, 6, 3, 0, 
    52, 22, 13, 9, 4, 4, 7, 6, 8, 9, 8, 7, 9, 9, 10, 11, 12, 12, 12, 15, 44, 52, 5, 0, 0, 0, 13, 21, 19, 7, 0, 0, 
    34, 5, 0, 0, 0, 0, 4, 4, 7, 10, 13, 12, 13, 14, 16, 16, 16, 18, 15, 25, 58, 32, 0, 0, 0, 1, 22, 22, 18, 7, 3, 0, 
    15, 0, 0, 0, 6, 8, 8, 8, 11, 15, 18, 16, 19, 21, 23, 21, 20, 24, 18, 27, 40, 0, 0, 0, 0, 12, 18, 13, 2, 0, 0, 0, 
    15, 2, 6, 12, 14, 14, 14, 13, 15, 18, 21, 20, 26, 27, 28, 28, 24, 28, 25, 31, 16, 0, 0, 0, 4, 1, 10, 2, 0, 0, 2, 0, 
    21, 12, 13, 16, 15, 14, 16, 15, 16, 21, 30, 32, 36, 31, 28, 29, 24, 26, 25, 20, 0, 0, 0, 2, 9, 0, 1, 4, 4, 7, 5, 0, 
    23, 13, 12, 15, 15, 13, 15, 14, 15, 22, 33, 30, 34, 30, 21, 31, 39, 54, 59, 20, 0, 0, 0, 1, 19, 0, 0, 0, 3, 5, 4, 0, 
    24, 14, 14, 14, 15, 12, 14, 12, 15, 20, 26, 35, 60, 61, 50, 64, 77, 94, 104, 73, 73, 47, 0, 0, 0, 9, 6, 0, 0, 3, 2, 0, 
    25, 16, 15, 15, 16, 13, 14, 12, 15, 32, 54, 64, 75, 74, 61, 62, 53, 32, 5, 3, 84, 99, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 
    26, 17, 15, 15, 17, 12, 13, 13, 32, 57, 50, 44, 48, 4, 0, 0, 0, 0, 0, 0, 68, 67, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    27, 17, 16, 14, 16, 8, 8, 24, 48, 38, 9, 0, 0, 0, 0, 0, 0, 0, 0, 70, 132, 68, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28, 17, 16, 12, 18, 24, 19, 25, 25, 0, 0, 0, 0, 0, 0, 0, 11, 38, 83, 146, 130, 63, 9, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    27, 14, 15, 14, 23, 44, 41, 27, 16, 0, 0, 12, 16, 0, 28, 66, 90, 113, 131, 140, 100, 40, 0, 0, 0, 0, 0, 11, 67, 55, 0, 0, 
    27, 13, 14, 16, 17, 22, 19, 19, 13, 0, 0, 0, 0, 28, 140, 157, 149, 157, 132, 90, 49, 0, 0, 0, 0, 0, 0, 57, 104, 76, 0, 0, 
    27, 12, 19, 43, 28, 0, 0, 0, 0, 0, 0, 0, 0, 49, 153, 121, 62, 39, 27, 22, 24, 0, 0, 0, 0, 33, 42, 83, 90, 56, 0, 0, 
    24, 16, 60, 103, 33, 0, 0, 0, 0, 0, 0, 10, 19, 92, 141, 50, 0, 0, 9, 10, 20, 12, 0, 0, 54, 83, 78, 73, 51, 10, 0, 0, 
    20, 46, 140, 137, 19, 0, 0, 0, 0, 0, 0, 1, 21, 101, 128, 34, 2, 17, 0, 0, 0, 15, 41, 56, 76, 73, 49, 18, 0, 0, 0, 0, 
    22, 81, 150, 94, 0, 0, 0, 0, 0, 0, 0, 4, 16, 83, 104, 28, 17, 0, 0, 0, 0, 0, 2, 49, 43, 15, 0, 0, 0, 0, 0, 0, 
    29, 75, 51, 0, 0, 0, 0, 0, 0, 0, 15, 50, 50, 96, 92, 25, 11, 0, 0, 0, 0, 0, 0, 28, 14, 0, 0, 0, 0, 0, 0, 0, 
    32, 48, 0, 0, 0, 0, 0, 0, 0, 0, 43, 65, 65, 118, 100, 28, 0, 0, 0, 0, 0, 0, 2, 34, 17, 0, 0, 0, 0, 0, 0, 0, 
    24, 31, 3, 0, 55, 1, 0, 0, 0, 13, 48, 38, 43, 93, 71, 28, 0, 0, 0, 0, 0, 0, 0, 31, 52, 14, 0, 0, 0, 0, 7, 0, 
    13, 22, 16, 13, 58, 8, 0, 0, 0, 41, 56, 32, 45, 81, 48, 12, 0, 0, 0, 17, 0, 0, 0, 1, 59, 24, 0, 0, 0, 0, 0, 0, 
    9, 17, 19, 8, 37, 11, 0, 0, 32, 72, 78, 60, 65, 68, 29, 8, 0, 0, 0, 31, 20, 0, 0, 0, 34, 7, 0, 0, 0, 0, 0, 0, 
    12, 14, 27, 20, 28, 6, 0, 0, 42, 60, 58, 46, 46, 39, 8, 0, 0, 0, 0, 22, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 11, 12, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 10, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 8, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 6, 18, 29, 32, 31, 22, 0, 0, 7, 8, 8, 6, 4, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=102
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=103
    0, 8, 10, 13, 13, 13, 17, 20, 18, 18, 17, 14, 12, 11, 11, 12, 10, 8, 3, 0, 2, 1, 2, 1, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 19, 20, 24, 18, 13, 15, 14, 9, 10, 12, 11, 10, 8, 10, 12, 12, 1, 0, 5, 4, 2, 13, 6, 6, 0, 0, 0, 0, 0, 4, 0, 
    0, 16, 16, 20, 15, 11, 12, 11, 7, 8, 9, 9, 7, 5, 7, 10, 9, 3, 0, 10, 5, 4, 10, 2, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 15, 10, 12, 8, 8, 8, 8, 7, 7, 7, 7, 5, 3, 5, 7, 6, 5, 4, 7, 10, 8, 2, 0, 0, 0, 0, 0, 0, 1, 3, 0, 
    0, 11, 2, 2, 3, 7, 5, 6, 6, 6, 6, 6, 4, 3, 5, 6, 7, 5, 6, 6, 14, 10, 0, 0, 0, 0, 2, 0, 0, 4, 3, 0, 
    0, 1, 0, 1, 7, 6, 4, 6, 6, 6, 5, 4, 3, 3, 5, 5, 7, 5, 5, 8, 8, 0, 0, 1, 0, 0, 2, 0, 0, 0, 6, 0, 
    0, 0, 1, 4, 6, 4, 3, 6, 5, 3, 2, 1, 1, 1, 3, 4, 7, 6, 8, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 
    0, 1, 1, 2, 1, 2, 1, 4, 3, 2, 1, 4, 8, 4, 4, 5, 6, 6, 10, 4, 0, 0, 1, 0, 0, 0, 0, 0, 3, 3, 6, 0, 
    0, 0, 0, 1, 0, 2, 0, 3, 1, 1, 3, 7, 12, 6, 4, 0, 1, 0, 2, 0, 0, 2, 5, 0, 0, 0, 0, 3, 5, 3, 4, 0, 
    0, 0, 0, 2, 0, 2, 0, 2, 2, 2, 4, 1, 1, 0, 1, 2, 9, 10, 9, 0, 0, 2, 0, 0, 0, 0, 1, 0, 4, 2, 2, 0, 
    0, 1, 1, 2, 1, 3, 1, 3, 3, 2, 0, 0, 7, 6, 9, 10, 8, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 
    0, 3, 1, 2, 1, 4, 2, 4, 5, 5, 5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 2, 2, 0, 3, 2, 4, 8, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 1, 2, 0, 1, 2, 5, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 1, 0, 0, 0, 
    0, 2, 0, 3, 5, 6, 7, 4, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 12, 0, 0, 0, 0, 0, 5, 0, 0, 0, 5, 2, 0, 0, 
    0, 1, 0, 4, 8, 11, 5, 0, 0, 0, 0, 0, 0, 0, 7, 9, 4, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 3, 0, 0, 0, 
    0, 1, 0, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 1, 2, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 1, 0, 0, 0, 0, 4, 
    0, 4, 12, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 13, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 11, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 11, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 4, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=104
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 17, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 58, 32, 8, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 49, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 55, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 83, 102, 104, 78, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 42, 58, 89, 116, 147, 189, 180, 190, 177, 47, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 102, 136, 129, 125, 124, 126, 131, 154, 232, 275, 143, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 43, 62, 93, 103, 65, 38, 52, 47, 19, 69, 205, 314, 262, 75, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 20, 42, 86, 85, 35, 0, 18, 15, 0, 72, 190, 290, 320, 190, 24, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 19, 27, 55, 89, 83, 39, 0, 8, 50, 93, 155, 222, 273, 321, 251, 87, 5, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 18, 26, 53, 53, 29, 49, 72, 69, 87, 103, 129, 190, 215, 225, 265, 295, 268, 178, 106, 34, 0, 0, 52, 69, 39, 
    0, 0, 0, 0, 0, 0, 4, 44, 67, 104, 50, 19, 37, 29, 72, 187, 242, 243, 250, 253, 270, 295, 271, 162, 70, 43, 36, 11, 49, 113, 151, 94, 
    0, 0, 0, 0, 3, 30, 18, 47, 87, 74, 47, 9, 31, 9, 71, 204, 261, 253, 249, 262, 275, 286, 253, 150, 36, 11, 81, 100, 110, 135, 190, 144, 
    0, 0, 0, 0, 115, 126, 53, 32, 66, 57, 28, 0, 38, 27, 63, 197, 261, 246, 249, 260, 256, 268, 297, 217, 110, 111, 150, 160, 150, 161, 188, 150, 
    0, 0, 0, 92, 211, 196, 85, 36, 64, 46, 0, 0, 15, 23, 86, 216, 257, 250, 265, 232, 173, 162, 233, 264, 220, 197, 198, 197, 190, 184, 147, 107, 
    0, 0, 3, 134, 223, 237, 118, 51, 50, 25, 0, 0, 4, 17, 108, 227, 247, 264, 246, 142, 68, 47, 78, 195, 254, 245, 224, 201, 195, 155, 74, 54, 
    0, 0, 26, 68, 147, 210, 136, 65, 37, 14, 0, 15, 62, 59, 125, 229, 247, 270, 188, 91, 48, 22, 0, 64, 200, 234, 200, 189, 156, 79, 20, 22, 
    0, 0, 17, 41, 68, 167, 158, 70, 31, 5, 0, 50, 96, 92, 153, 241, 263, 264, 159, 74, 36, 29, 0, 0, 103, 196, 199, 175, 98, 34, 0, 10, 
    0, 0, 30, 73, 39, 135, 171, 73, 25, 12, 22, 59, 82, 117, 194, 251, 269, 256, 142, 42, 40, 46, 32, 0, 26, 164, 204, 155, 71, 4, 0, 13, 
    0, 0, 23, 69, 49, 121, 173, 82, 21, 25, 58, 91, 105, 134, 192, 237, 260, 255, 128, 39, 75, 62, 40, 0, 0, 114, 187, 132, 39, 0, 0, 8, 
    0, 0, 9, 57, 63, 110, 171, 101, 49, 68, 118, 165, 175, 171, 214, 244, 265, 263, 124, 33, 86, 109, 77, 23, 0, 54, 140, 96, 9, 0, 0, 0, 
    0, 0, 0, 52, 71, 107, 158, 115, 77, 90, 122, 158, 169, 161, 184, 190, 201, 211, 108, 42, 80, 112, 75, 33, 0, 3, 62, 44, 0, 0, 0, 0, 
    0, 0, 0, 34, 56, 72, 89, 63, 31, 30, 38, 53, 66, 68, 74, 75, 80, 102, 53, 31, 62, 75, 80, 39, 0, 0, 6, 7, 0, 0, 0, 3, 
    0, 0, 3, 17, 30, 22, 32, 28, 13, 7, 7, 9, 12, 13, 16, 14, 9, 17, 6, 0, 54, 75, 79, 25, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 14, 32, 41, 45, 62, 71, 49, 28, 28, 33, 32, 29, 25, 21, 12, 6, 0, 0, 26, 53, 31, 16, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 26, 68, 102, 115, 115, 113, 83, 61, 66, 72, 71, 67, 61, 58, 49, 39, 26, 8, 11, 37, 36, 12, 0, 0, 0, 0, 0, 0, 4, 21, 
    0, 0, 0, 29, 54, 64, 61, 62, 54, 38, 37, 41, 40, 39, 35, 33, 28, 22, 16, 11, 11, 16, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=105
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 33, 40, 25, 1, 0, 0, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 13, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 20, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 2, 6, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 1, 13, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 17, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 79, 45, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 76, 110, 135, 127, 55, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 50, 78, 98, 117, 137, 165, 210, 254, 195, 60, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 76, 64, 39, 9, 0, 0, 0, 60, 211, 217, 124, 30, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 19, 2, 0, 0, 0, 0, 0, 0, 42, 145, 156, 156, 121, 50, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 0, 0, 6, 48, 126, 210, 187, 131, 162, 167, 117, 52, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 49, 68, 72, 87, 96, 128, 202, 291, 298, 205, 141, 132, 142, 136, 103, 50, 27, 27, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 15, 46, 44, 39, 51, 74, 91, 147, 238, 300, 321, 329, 334, 261, 180, 122, 27, 0, 56, 84, 84, 126, 150, 79, 26, 
    0, 0, 0, 0, 0, 0, 0, 23, 64, 80, 55, 28, 24, 64, 184, 299, 322, 300, 260, 208, 162, 122, 40, 0, 0, 0, 69, 144, 205, 198, 96, 38, 
    0, 0, 0, 0, 0, 36, 36, 38, 64, 55, 34, 56, 69, 96, 176, 207, 157, 121, 104, 107, 126, 126, 55, 1, 50, 108, 163, 229, 228, 154, 58, 29, 
    0, 0, 0, 10, 119, 127, 102, 91, 78, 38, 41, 85, 124, 169, 202, 145, 98, 106, 116, 119, 114, 121, 147, 191, 222, 228, 228, 219, 176, 106, 27, 0, 
    0, 0, 0, 141, 192, 148, 125, 109, 84, 52, 56, 74, 97, 147, 196, 156, 135, 146, 122, 42, 0, 0, 71, 187, 248, 243, 204, 161, 125, 78, 0, 0, 
    0, 0, 31, 122, 111, 115, 136, 114, 73, 45, 72, 104, 123, 153, 188, 162, 150, 135, 55, 0, 0, 0, 0, 64, 168, 178, 144, 117, 74, 10, 0, 0, 
    0, 0, 0, 0, 0, 90, 127, 110, 65, 55, 108, 174, 225, 235, 213, 164, 147, 104, 10, 0, 51, 60, 10, 15, 73, 107, 101, 68, 12, 0, 0, 16, 
    0, 0, 8, 2, 52, 114, 120, 94, 63, 88, 135, 182, 211, 230, 227, 183, 155, 87, 9, 54, 102, 103, 91, 61, 60, 96, 105, 68, 0, 0, 23, 57, 
    0, 0, 29, 111, 164, 151, 123, 92, 79, 125, 168, 178, 163, 187, 205, 170, 140, 72, 48, 115, 116, 96, 97, 87, 87, 115, 127, 66, 14, 34, 48, 51, 
    0, 0, 37, 120, 161, 149, 108, 92, 106, 158, 202, 203, 182, 195, 171, 132, 118, 73, 76, 126, 134, 129, 106, 90, 92, 98, 88, 38, 21, 33, 19, 24, 
    0, 0, 51, 105, 143, 155, 132, 146, 189, 240, 274, 279, 268, 244, 186, 161, 147, 105, 98, 131, 155, 156, 129, 104, 89, 67, 34, 16, 29, 32, 16, 26, 
    0, 0, 53, 105, 142, 139, 112, 133, 164, 165, 144, 122, 117, 100, 65, 54, 48, 47, 82, 114, 104, 97, 88, 82, 69, 31, 0, 13, 49, 49, 39, 47, 
    5, 0, 29, 62, 77, 60, 20, 31, 48, 26, 0, 0, 0, 0, 0, 0, 0, 0, 25, 110, 96, 69, 67, 71, 64, 45, 15, 37, 66, 67, 60, 60, 
    14, 4, 33, 45, 45, 42, 42, 71, 80, 69, 59, 47, 38, 31, 21, 16, 6, 1, 24, 69, 94, 99, 86, 67, 66, 70, 64, 69, 74, 78, 78, 72, 
    20, 3, 39, 90, 130, 151, 171, 182, 165, 151, 154, 156, 151, 141, 129, 121, 110, 98, 94, 69, 42, 52, 45, 45, 73, 82, 82, 81, 83, 86, 86, 75, 
    36, 25, 73, 148, 215, 238, 227, 199, 179, 183, 191, 191, 186, 179, 173, 169, 159, 145, 140, 139, 120, 86, 66, 76, 94, 99, 98, 96, 97, 98, 90, 71, 
    9, 0, 0, 15, 29, 32, 28, 25, 38, 62, 63, 55, 46, 40, 42, 45, 46, 49, 54, 62, 64, 57, 56, 61, 61, 63, 64, 61, 58, 52, 42, 38, 
    
    -- channel=106
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 24, 50, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 24, 39, 47, 53, 121, 84, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 25, 8, 7, 13, 0, 0, 51, 137, 122, 17, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 76, 145, 137, 83, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 106, 154, 149, 124, 20, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 13, 31, 86, 144, 153, 149, 95, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 71, 66, 93, 119, 148, 149, 148, 111, 33, 0, 0, 0, 0, 0, 35, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 135, 136, 140, 145, 148, 143, 152, 95, 0, 0, 0, 0, 0, 38, 69, 53, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 93, 157, 141, 138, 140, 138, 134, 145, 106, 12, 0, 18, 40, 63, 81, 74, 55, 0, 
    0, 0, 0, 0, 50, 22, 0, 0, 4, 0, 0, 0, 0, 4, 122, 152, 135, 138, 140, 107, 89, 101, 122, 100, 75, 87, 100, 98, 83, 68, 25, 0, 
    0, 0, 0, 57, 104, 58, 0, 0, 0, 0, 0, 0, 0, 8, 126, 146, 131, 146, 115, 56, 34, 27, 63, 129, 137, 125, 106, 96, 80, 36, 0, 0, 
    0, 0, 0, 45, 84, 81, 2, 0, 0, 0, 0, 0, 11, 26, 127, 140, 131, 143, 57, 0, 0, 0, 0, 75, 142, 124, 101, 87, 43, 0, 0, 0, 
    0, 0, 0, 0, 30, 84, 12, 0, 0, 0, 0, 4, 34, 61, 147, 137, 137, 120, 0, 0, 0, 0, 0, 16, 107, 114, 88, 63, 0, 0, 0, 0, 
    0, 0, 0, 0, 18, 90, 27, 0, 0, 0, 0, 33, 45, 82, 144, 138, 144, 93, 0, 0, 0, 0, 0, 0, 57, 101, 89, 37, 0, 0, 0, 0, 
    0, 0, 0, 0, 19, 89, 36, 0, 0, 0, 15, 53, 43, 92, 142, 134, 141, 72, 0, 0, 0, 0, 0, 0, 9, 85, 82, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 17, 84, 51, 0, 0, 20, 59, 85, 75, 112, 137, 128, 134, 69, 0, 0, 23, 7, 0, 0, 0, 55, 50, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 14, 69, 42, 0, 9, 37, 69, 88, 90, 108, 110, 106, 112, 69, 0, 3, 14, 20, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 33, 14, 0, 3, 20, 34, 41, 39, 45, 48, 46, 42, 16, 0, 12, 19, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 21, 26, 25, 1, 0, 3, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 13, 16, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=107
    98, 166, 178, 177, 175, 187, 196, 193, 191, 189, 176, 163, 156, 158, 159, 150, 138, 128, 130, 133, 139, 119, 112, 105, 100, 112, 108, 85, 88, 91, 81, 87, 
    17, 59, 52, 38, 18, 19, 21, 13, 8, 11, 9, 3, 0, 0, 11, 12, 7, 0, 0, 0, 5, 14, 22, 24, 27, 27, 13, 0, 10, 22, 18, 54, 
    0, 16, 21, 24, 16, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 14, 17, 17, 20, 22, 37, 28, 10, 11, 17, 10, 50, 
    0, 1, 16, 28, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 10, 11, 18, 47, 57, 43, 55, 45, 24, 21, 15, 12, 48, 
    0, 6, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 5, 7, 11, 17, 48, 97, 92, 78, 70, 43, 37, 40, 31, 22, 49, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 12, 13, 15, 16, 19, 44, 80, 67, 71, 79, 54, 49, 36, 27, 17, 49, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 16, 21, 22, 30, 32, 15, 29, 39, 10, 31, 61, 47, 23, 6, 8, 9, 51, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 23, 35, 44, 44, 47, 39, 29, 52, 49, 7, 16, 27, 15, 5, 1, 5, 6, 52, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 26, 36, 40, 35, 36, 29, 27, 33, 49, 85, 101, 65, 37, 22, 7, 6, 7, 4, 5, 50, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 25, 25, 30, 30, 55, 90, 132, 179, 192, 168, 158, 90, 38, 37, 25, 12, 8, 4, 3, 46, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 85, 152, 182, 214, 234, 241, 256, 250, 253, 259, 139, 17, 10, 30, 50, 20, 1, 0, 42, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 56, 117, 163, 172, 137, 96, 49, 10, 29, 81, 215, 330, 226, 53, 0, 10, 54, 47, 5, 0, 41, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 64, 79, 34, 6, 0, 0, 0, 0, 0, 0, 0, 128, 309, 310, 170, 15, 0, 23, 42, 10, 2, 42, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 32, 23, 0, 0, 0, 13, 0, 0, 0, 18, 0, 12, 127, 239, 316, 275, 105, 0, 0, 10, 8, 6, 44, 
    0, 0, 0, 0, 0, 0, 9, 30, 22, 15, 5, 22, 46, 91, 106, 81, 58, 79, 141, 157, 156, 154, 188, 285, 281, 162, 58, 17, 14, 40, 71, 83, 
    0, 0, 0, 0, 0, 12, 50, 73, 46, 67, 93, 64, 67, 92, 116, 177, 239, 287, 314, 263, 207, 176, 179, 191, 136, 96, 95, 40, 48, 128, 176, 142, 
    0, 0, 0, 0, 0, 2, 14, 29, 73, 109, 84, 25, 32, 51, 112, 282, 361, 320, 256, 204, 183, 179, 145, 64, 0, 25, 67, 82, 111, 175, 217, 184, 
    0, 0, 0, 0, 30, 45, 14, 25, 51, 73, 39, 13, 31, 38, 48, 162, 190, 145, 123, 137, 158, 168, 191, 150, 52, 64, 137, 168, 146, 139, 194, 198, 
    0, 0, 0, 39, 165, 179, 74, 21, 40, 69, 40, 30, 68, 39, 4, 88, 120, 110, 121, 142, 143, 187, 279, 287, 207, 180, 193, 164, 129, 113, 167, 171, 
    0, 0, 1, 125, 252, 215, 109, 38, 67, 74, 32, 14, 26, 0, 6, 113, 141, 139, 142, 100, 11, 13, 130, 236, 242, 198, 165, 148, 136, 114, 125, 104, 
    0, 0, 0, 87, 173, 197, 143, 63, 73, 58, 29, 10, 10, 0, 21, 130, 145, 140, 110, 0, 0, 0, 0, 33, 151, 178, 152, 127, 117, 83, 47, 51, 
    0, 0, 0, 0, 3, 129, 149, 77, 78, 52, 41, 64, 105, 64, 66, 136, 144, 142, 101, 8, 0, 0, 0, 0, 30, 111, 98, 93, 71, 24, 16, 55, 
    0, 0, 0, 0, 0, 103, 158, 101, 75, 55, 55, 86, 123, 69, 93, 164, 162, 184, 143, 65, 77, 50, 0, 0, 0, 68, 108, 97, 64, 35, 40, 76, 
    0, 0, 20, 51, 30, 102, 161, 113, 74, 65, 56, 57, 64, 53, 122, 166, 168, 218, 143, 59, 77, 88, 42, 0, 0, 59, 131, 130, 84, 52, 50, 79, 
    0, 0, 22, 59, 32, 86, 161, 119, 69, 72, 77, 97, 92, 66, 107, 122, 161, 224, 140, 74, 106, 108, 79, 0, 0, 18, 114, 123, 66, 34, 28, 59, 
    0, 0, 0, 39, 27, 74, 156, 142, 103, 120, 153, 196, 178, 137, 142, 148, 195, 241, 141, 56, 100, 147, 134, 48, 0, 0, 73, 84, 36, 17, 16, 51, 
    0, 0, 1, 35, 40, 75, 142, 129, 97, 87, 86, 100, 82, 63, 64, 56, 88, 144, 96, 42, 80, 102, 102, 52, 0, 0, 18, 40, 31, 25, 20, 53, 
    4, 12, 14, 21, 12, 18, 36, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 9, 0, 41, 58, 77, 79, 4, 0, 15, 37, 38, 33, 27, 57, 
    9, 30, 21, 16, 0, 0, 5, 14, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 92, 106, 79, 38, 34, 43, 46, 46, 45, 42, 70, 
    4, 31, 40, 51, 67, 95, 125, 143, 126, 91, 87, 94, 95, 92, 83, 75, 72, 70, 27, 0, 13, 29, 50, 53, 54, 55, 55, 55, 55, 57, 57, 81, 
    0, 29, 52, 98, 152, 178, 173, 160, 130, 105, 114, 122, 128, 131, 128, 126, 123, 117, 93, 47, 24, 45, 70, 70, 67, 68, 70, 67, 64, 65, 66, 84, 
    0, 0, 0, 0, 5, 2, 0, 15, 24, 21, 20, 20, 24, 28, 30, 32, 35, 38, 40, 32, 26, 35, 42, 42, 43, 43, 42, 39, 36, 29, 26, 42, 
    
    -- channel=108
    92, 113, 127, 132, 142, 157, 158, 155, 156, 149, 134, 124, 121, 124, 118, 101, 88, 91, 109, 126, 111, 70, 59, 56, 35, 30, 31, 30, 30, 17, 5, 0, 
    157, 138, 134, 120, 120, 128, 121, 112, 111, 102, 88, 80, 78, 82, 77, 63, 55, 48, 36, 23, 29, 26, 19, 30, 20, 1, 0, 0, 17, 13, 0, 0, 
    165, 125, 117, 105, 105, 104, 94, 83, 82, 75, 65, 59, 59, 62, 57, 48, 41, 36, 33, 20, 28, 33, 25, 17, 0, 0, 0, 0, 20, 14, 0, 0, 
    149, 103, 108, 104, 101, 87, 72, 61, 57, 54, 48, 43, 44, 48, 42, 36, 33, 29, 30, 28, 27, 41, 42, 15, 0, 0, 0, 1, 32, 21, 6, 0, 
    135, 96, 102, 90, 75, 60, 52, 43, 38, 36, 34, 31, 33, 36, 32, 31, 31, 29, 29, 33, 41, 72, 86, 42, 0, 0, 0, 27, 47, 32, 17, 0, 
    104, 66, 60, 39, 31, 31, 35, 28, 24, 26, 29, 30, 32, 34, 30, 33, 36, 37, 35, 44, 60, 84, 84, 45, 26, 14, 20, 56, 58, 40, 20, 0, 
    57, 19, 19, 18, 22, 24, 27, 21, 23, 27, 32, 36, 40, 42, 40, 45, 46, 49, 47, 54, 57, 42, 0, 0, 30, 37, 42, 52, 39, 24, 7, 0, 
    38, 12, 16, 19, 26, 26, 31, 25, 31, 34, 38, 42, 48, 59, 64, 67, 65, 72, 71, 70, 49, 0, 0, 0, 22, 37, 37, 24, 20, 18, 5, 0, 
    38, 22, 24, 23, 28, 26, 35, 30, 35, 41, 48, 57, 66, 86, 96, 94, 85, 84, 81, 72, 42, 0, 0, 0, 43, 43, 29, 20, 17, 19, 10, 0, 
    42, 26, 26, 25, 29, 26, 35, 30, 35, 44, 58, 76, 83, 97, 103, 101, 104, 124, 145, 137, 90, 53, 39, 37, 67, 54, 34, 23, 13, 16, 12, 0, 
    47, 27, 29, 26, 30, 27, 34, 28, 33, 42, 52, 71, 91, 133, 169, 194, 232, 281, 326, 318, 248, 196, 120, 28, 29, 49, 56, 40, 14, 11, 10, 0, 
    52, 28, 31, 29, 33, 29, 33, 29, 32, 44, 65, 105, 164, 245, 287, 293, 290, 275, 257, 244, 264, 335, 259, 62, 0, 0, 60, 73, 27, 8, 7, 0, 
    57, 28, 34, 32, 36, 32, 31, 32, 39, 69, 112, 157, 184, 183, 130, 76, 50, 22, 0, 16, 153, 338, 337, 155, 0, 0, 18, 64, 39, 10, 5, 0, 
    62, 30, 36, 33, 38, 32, 24, 35, 56, 92, 105, 86, 68, 49, 0, 0, 0, 0, 0, 21, 197, 351, 362, 257, 71, 0, 0, 12, 9, 4, 2, 0, 
    66, 33, 40, 34, 36, 40, 37, 53, 66, 72, 46, 30, 53, 56, 15, 0, 0, 27, 71, 168, 312, 370, 361, 315, 156, 20, 0, 0, 0, 20, 21, 0, 
    65, 33, 40, 35, 36, 59, 92, 101, 81, 56, 38, 61, 85, 70, 60, 88, 126, 195, 271, 355, 394, 371, 341, 260, 131, 50, 0, 0, 28, 113, 106, 10, 
    65, 33, 39, 37, 33, 46, 90, 103, 93, 72, 47, 35, 48, 65, 172, 318, 395, 433, 442, 430, 396, 362, 276, 116, 6, 22, 10, 14, 115, 225, 195, 40, 
    65, 32, 36, 47, 47, 20, 23, 44, 60, 48, 0, 0, 0, 44, 227, 399, 417, 395, 380, 374, 375, 347, 216, 45, 3, 64, 90, 138, 214, 264, 222, 59, 
    62, 30, 49, 110, 139, 75, 29, 30, 34, 0, 0, 0, 30, 85, 249, 350, 333, 323, 331, 349, 366, 372, 301, 191, 157, 191, 229, 250, 252, 235, 200, 54, 
    58, 37, 109, 239, 261, 124, 29, 17, 19, 0, 0, 0, 27, 103, 260, 326, 315, 321, 320, 285, 255, 290, 342, 332, 302, 289, 276, 259, 238, 202, 139, 9, 
    55, 55, 163, 303, 282, 138, 50, 21, 3, 0, 0, 0, 0, 79, 252, 317, 313, 306, 236, 104, 22, 49, 175, 290, 326, 303, 267, 246, 210, 134, 40, 0, 
    53, 50, 111, 167, 163, 133, 64, 18, 0, 0, 0, 2, 52, 126, 265, 310, 305, 262, 117, 0, 0, 0, 16, 159, 266, 265, 223, 185, 118, 20, 0, 0, 
    46, 28, 23, 0, 54, 124, 70, 14, 0, 0, 0, 72, 142, 199, 298, 319, 302, 218, 43, 0, 6, 0, 0, 57, 170, 203, 176, 123, 25, 0, 0, 0, 
    34, 15, 11, 8, 80, 148, 84, 6, 0, 0, 19, 85, 130, 205, 315, 335, 304, 190, 22, 8, 7, 0, 0, 2, 115, 188, 175, 89, 0, 0, 0, 0, 
    20, 1, 12, 44, 89, 149, 90, 4, 0, 19, 70, 112, 138, 227, 311, 307, 280, 162, 27, 43, 46, 23, 0, 0, 64, 160, 151, 46, 0, 0, 0, 0, 
    6, 0, 3, 40, 73, 139, 98, 24, 26, 90, 159, 203, 215, 266, 296, 290, 277, 163, 37, 56, 85, 63, 12, 0, 11, 95, 82, 0, 0, 0, 0, 0, 
    0, 0, 6, 41, 70, 127, 109, 68, 89, 149, 210, 250, 256, 270, 268, 263, 249, 152, 38, 55, 99, 91, 35, 0, 0, 9, 0, 0, 0, 0, 0, 0, 
    4, 0, 3, 28, 47, 66, 39, 2, 6, 16, 26, 34, 37, 46, 49, 45, 47, 21, 0, 39, 52, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 15, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 50, 43, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 29, 20, 0, 0, 0, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 29, 37, 51, 78, 94, 103, 83, 36, 19, 28, 36, 39, 35, 27, 19, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 34, 63, 68, 54, 27, 0, 0, 10, 13, 17, 19, 16, 13, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=109
    178, 151, 149, 149, 166, 169, 158, 156, 154, 140, 129, 126, 131, 132, 116, 100, 96, 106, 120, 113, 107, 68, 67, 64, 46, 33, 21, 42, 49, 33, 25, 0, 
    252, 183, 165, 153, 168, 168, 150, 147, 145, 131, 119, 117, 123, 125, 108, 93, 92, 97, 90, 69, 54, 61, 52, 57, 41, 0, 0, 32, 61, 45, 37, 0, 
    252, 166, 149, 141, 147, 141, 131, 128, 130, 120, 109, 105, 111, 111, 98, 86, 83, 85, 79, 64, 65, 67, 59, 46, 11, 0, 0, 39, 69, 50, 42, 0, 
    230, 151, 150, 139, 133, 125, 118, 114, 114, 108, 99, 95, 101, 101, 90, 81, 78, 78, 79, 69, 69, 89, 69, 18, 0, 0, 0, 61, 79, 59, 48, 0, 
    209, 141, 139, 127, 115, 110, 107, 99, 97, 94, 89, 87, 92, 92, 84, 79, 79, 79, 78, 77, 98, 123, 80, 29, 0, 0, 37, 82, 86, 64, 53, 0, 
    170, 109, 105, 90, 85, 89, 93, 86, 84, 84, 86, 88, 92, 90, 87, 85, 84, 84, 82, 92, 123, 108, 52, 37, 36, 31, 69, 96, 90, 68, 54, 0, 
    124, 73, 71, 77, 81, 86, 85, 80, 82, 86, 92, 96, 102, 100, 97, 95, 94, 96, 91, 100, 101, 38, 0, 15, 58, 66, 82, 86, 76, 59, 44, 0, 
    104, 71, 75, 82, 85, 87, 87, 83, 89, 95, 101, 103, 114, 122, 119, 114, 109, 111, 106, 103, 63, 0, 0, 14, 78, 75, 75, 64, 62, 56, 47, 0, 
    105, 83, 84, 88, 88, 90, 93, 89, 95, 105, 117, 121, 127, 135, 139, 133, 119, 120, 117, 96, 40, 0, 0, 39, 93, 80, 67, 61, 59, 61, 54, 0, 
    112, 88, 88, 90, 90, 92, 96, 92, 97, 110, 129, 126, 127, 139, 141, 150, 155, 175, 188, 130, 52, 24, 6, 53, 105, 79, 66, 61, 55, 59, 56, 0, 
    118, 91, 91, 92, 91, 91, 95, 90, 96, 107, 120, 130, 163, 194, 199, 221, 248, 286, 316, 258, 211, 161, 26, 0, 49, 82, 93, 61, 49, 56, 54, 0, 
    124, 93, 94, 94, 94, 91, 93, 88, 92, 113, 147, 175, 215, 254, 260, 271, 272, 264, 245, 227, 302, 319, 108, 0, 0, 38, 105, 88, 45, 50, 49, 0, 
    129, 94, 96, 96, 99, 89, 88, 86, 106, 147, 163, 181, 213, 190, 111, 81, 81, 49, 14, 100, 301, 362, 191, 0, 0, 0, 80, 76, 48, 50, 47, 0, 
    134, 96, 98, 97, 102, 84, 78, 97, 132, 141, 121, 121, 117, 54, 0, 0, 0, 0, 0, 154, 352, 381, 277, 90, 0, 0, 25, 33, 25, 42, 42, 0, 
    136, 99, 102, 96, 99, 99, 96, 108, 114, 94, 71, 69, 82, 33, 0, 0, 22, 64, 128, 278, 379, 378, 328, 169, 0, 0, 0, 0, 23, 62, 38, 0, 
    136, 99, 104, 94, 97, 124, 139, 124, 100, 67, 36, 92, 99, 58, 77, 120, 162, 226, 295, 374, 395, 361, 283, 115, 29, 15, 0, 2, 108, 148, 65, 0, 
    137, 99, 103, 93, 79, 96, 123, 120, 108, 41, 29, 58, 51, 102, 270, 345, 366, 411, 425, 410, 377, 314, 154, 12, 6, 27, 16, 80, 202, 239, 106, 0, 
    139, 97, 102, 117, 85, 36, 52, 72, 65, 9, 0, 11, 14, 137, 367, 425, 386, 374, 369, 365, 363, 282, 86, 0, 38, 119, 120, 187, 259, 274, 121, 0, 
    137, 93, 144, 210, 123, 12, 27, 69, 31, 0, 0, 24, 54, 196, 390, 374, 309, 316, 333, 340, 354, 322, 190, 113, 169, 222, 240, 261, 263, 237, 97, 0, 
    130, 117, 254, 319, 175, 22, 7, 49, 0, 0, 0, 10, 66, 227, 383, 335, 295, 315, 285, 229, 243, 309, 315, 279, 278, 282, 271, 247, 220, 167, 39, 0, 
    125, 164, 312, 334, 201, 33, 5, 32, 0, 0, 0, 0, 53, 216, 357, 314, 303, 275, 138, 47, 53, 125, 253, 324, 310, 268, 234, 220, 165, 57, 0, 0, 
    128, 165, 204, 192, 164, 63, 9, 4, 0, 0, 0, 59, 100, 238, 344, 305, 295, 173, 0, 0, 0, 9, 127, 265, 286, 226, 199, 148, 42, 0, 0, 0, 
    128, 121, 71, 47, 126, 92, 2, 0, 0, 0, 47, 124, 166, 292, 361, 309, 267, 74, 0, 0, 6, 0, 49, 187, 242, 196, 148, 54, 0, 0, 0, 0, 
    111, 82, 41, 40, 163, 138, 2, 0, 0, 3, 81, 130, 178, 303, 347, 317, 239, 28, 0, 24, 11, 0, 0, 107, 221, 210, 123, 0, 0, 0, 16, 0, 
    83, 61, 55, 67, 163, 150, 0, 0, 0, 62, 122, 139, 192, 305, 327, 296, 208, 8, 0, 64, 39, 5, 0, 33, 182, 203, 79, 0, 0, 0, 15, 0, 
    62, 49, 61, 71, 139, 150, 23, 0, 62, 146, 202, 212, 246, 306, 299, 280, 200, 11, 0, 100, 95, 33, 0, 0, 110, 146, 17, 0, 0, 0, 0, 0, 
    54, 44, 68, 81, 125, 139, 46, 42, 113, 183, 232, 245, 258, 276, 257, 250, 192, 37, 12, 101, 104, 52, 0, 0, 27, 48, 0, 0, 0, 0, 0, 0, 
    59, 44, 55, 61, 84, 70, 6, 2, 39, 60, 70, 67, 67, 74, 72, 69, 46, 0, 14, 96, 69, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    74, 53, 38, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 67, 74, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    82, 62, 39, 15, 1, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 32, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    80, 63, 67, 73, 80, 85, 82, 40, 12, 25, 31, 34, 33, 26, 19, 10, 0, 0, 0, 3, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 22, 37, 58, 71, 68, 50, 11, 0, 10, 19, 19, 19, 17, 16, 12, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=110
    48, 70, 77, 86, 99, 103, 104, 107, 104, 96, 89, 86, 87, 85, 75, 67, 66, 61, 68, 66, 36, 33, 37, 12, 5, 3, 5, 4, 2, 5, 8, 0, 
    142, 201, 208, 215, 232, 240, 239, 241, 237, 225, 210, 201, 200, 200, 187, 172, 164, 157, 164, 147, 124, 116, 105, 86, 71, 49, 45, 51, 52, 60, 62, 13, 
    174, 236, 226, 215, 215, 221, 215, 211, 207, 195, 182, 172, 171, 171, 163, 150, 142, 132, 124, 110, 106, 105, 93, 82, 67, 21, 1, 27, 50, 65, 65, 16, 
    161, 224, 210, 197, 191, 188, 182, 176, 172, 164, 154, 144, 143, 143, 139, 129, 123, 115, 113, 104, 96, 93, 73, 66, 45, 0, 0, 18, 54, 66, 67, 20, 
    136, 194, 190, 182, 172, 159, 152, 147, 144, 138, 129, 121, 120, 123, 122, 114, 110, 104, 106, 102, 96, 83, 64, 46, 20, 6, 15, 33, 61, 67, 69, 20, 
    124, 167, 158, 149, 140, 132, 128, 125, 120, 117, 111, 105, 105, 108, 112, 107, 104, 102, 103, 102, 109, 99, 70, 44, 16, 21, 40, 62, 80, 79, 74, 20, 
    97, 126, 116, 112, 107, 108, 107, 107, 104, 104, 104, 101, 102, 103, 109, 108, 107, 107, 104, 103, 116, 95, 49, 42, 38, 41, 65, 86, 96, 88, 77, 21, 
    62, 92, 91, 95, 96, 96, 95, 96, 97, 101, 106, 106, 109, 108, 110, 108, 110, 113, 109, 107, 99, 52, 1, 24, 51, 62, 81, 90, 91, 87, 78, 23, 
    49, 84, 87, 93, 96, 97, 97, 97, 99, 105, 110, 108, 114, 118, 122, 124, 124, 125, 118, 105, 75, 11, 0, 6, 50, 75, 90, 88, 86, 84, 77, 23, 
    49, 85, 89, 95, 97, 99, 101, 101, 102, 108, 119, 121, 133, 127, 125, 128, 115, 100, 85, 54, 35, 0, 0, 16, 51, 70, 84, 86, 83, 80, 75, 23, 
    53, 87, 91, 97, 98, 98, 101, 102, 103, 107, 124, 129, 124, 98, 82, 94, 102, 112, 121, 88, 43, 0, 0, 11, 63, 73, 56, 67, 76, 75, 73, 22, 
    57, 92, 94, 97, 98, 97, 100, 100, 101, 105, 108, 103, 112, 127, 134, 159, 183, 200, 216, 197, 155, 74, 0, 0, 27, 66, 64, 42, 60, 68, 68, 20, 
    60, 98, 97, 99, 99, 96, 101, 98, 100, 98, 106, 131, 160, 166, 164, 174, 175, 152, 146, 166, 199, 177, 33, 0, 0, 23, 70, 48, 45, 60, 62, 18, 
    63, 101, 98, 100, 101, 96, 98, 95, 98, 109, 124, 132, 128, 94, 53, 41, 56, 32, 19, 71, 157, 199, 114, 0, 0, 0, 33, 49, 35, 47, 56, 15, 
    66, 102, 100, 100, 102, 95, 76, 83, 99, 112, 83, 67, 59, 32, 0, 0, 0, 1, 0, 51, 151, 184, 157, 48, 0, 0, 0, 14, 17, 13, 24, 7, 
    66, 102, 101, 99, 98, 101, 76, 73, 86, 51, 44, 54, 58, 32, 0, 0, 0, 0, 35, 110, 166, 172, 160, 117, 34, 0, 0, 0, 11, 2, 0, 0, 
    64, 99, 102, 98, 93, 111, 111, 86, 63, 30, 37, 65, 67, 69, 55, 39, 62, 107, 156, 184, 186, 172, 148, 94, 50, 15, 0, 0, 39, 54, 0, 0, 
    64, 97, 100, 98, 65, 65, 77, 73, 56, 34, 13, 34, 24, 81, 158, 185, 197, 216, 222, 209, 199, 156, 64, 1, 9, 17, 0, 21, 88, 115, 28, 0, 
    64, 98, 105, 91, 39, 10, 22, 44, 29, 4, 0, 12, 0, 76, 191, 216, 200, 197, 194, 200, 208, 155, 25, 0, 0, 36, 59, 83, 114, 129, 57, 0, 
    62, 103, 122, 116, 66, 0, 0, 22, 0, 0, 0, 15, 36, 105, 177, 182, 166, 164, 167, 197, 231, 227, 138, 51, 58, 91, 108, 112, 114, 111, 67, 0, 
    56, 119, 174, 194, 106, 0, 0, 5, 0, 0, 0, 0, 27, 116, 170, 163, 159, 150, 143, 142, 152, 204, 235, 172, 126, 120, 123, 120, 108, 95, 49, 0, 
    55, 133, 198, 220, 136, 12, 0, 0, 0, 0, 0, 0, 0, 91, 162, 156, 155, 119, 76, 27, 20, 60, 168, 220, 166, 132, 123, 107, 90, 50, 11, 0, 
    57, 121, 120, 105, 115, 31, 0, 0, 0, 0, 0, 15, 36, 104, 148, 149, 139, 68, 5, 0, 0, 0, 50, 170, 168, 114, 90, 66, 33, 0, 0, 0, 
    55, 100, 50, 13, 80, 43, 0, 0, 0, 0, 10, 48, 80, 127, 157, 157, 127, 27, 0, 0, 0, 0, 0, 91, 145, 101, 60, 19, 0, 0, 0, 0, 
    44, 82, 52, 22, 75, 56, 0, 0, 0, 0, 17, 33, 75, 141, 171, 166, 115, 7, 0, 5, 0, 0, 0, 35, 127, 117, 51, 0, 0, 0, 17, 0, 
    28, 61, 54, 34, 70, 60, 0, 0, 0, 7, 24, 23, 62, 130, 147, 145, 95, 0, 0, 28, 2, 0, 0, 0, 95, 114, 40, 0, 0, 0, 13, 0, 
    17, 45, 49, 30, 61, 62, 6, 0, 23, 70, 105, 114, 132, 162, 169, 171, 129, 19, 0, 38, 48, 6, 0, 0, 47, 84, 27, 0, 0, 0, 2, 0, 
    16, 34, 47, 50, 64, 70, 40, 32, 61, 95, 126, 141, 151, 157, 157, 156, 131, 50, 24, 36, 42, 24, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 
    20, 31, 34, 40, 42, 35, 4, 0, 0, 9, 18, 24, 31, 35, 35, 35, 32, 8, 22, 51, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 39, 26, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 41, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 39, 27, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    39, 52, 63, 70, 67, 61, 53, 26, 6, 12, 18, 21, 22, 20, 18, 13, 6, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    
    -- channel=111
    78, 93, 95, 100, 108, 107, 105, 106, 104, 99, 96, 96, 97, 95, 88, 84, 85, 89, 97, 55, 41, 58, 49, 46, 52, 40, 21, 22, 32, 41, 43, 23, 
    201, 253, 260, 268, 284, 291, 289, 289, 288, 278, 266, 259, 259, 257, 246, 231, 225, 212, 192, 205, 169, 163, 161, 149, 126, 86, 69, 88, 112, 119, 123, 72, 
    241, 290, 283, 272, 277, 283, 282, 280, 279, 269, 255, 244, 242, 240, 231, 218, 210, 199, 182, 173, 165, 163, 158, 139, 96, 52, 32, 69, 116, 131, 133, 79, 
    244, 290, 278, 263, 256, 260, 263, 260, 256, 247, 235, 224, 221, 220, 212, 201, 192, 185, 178, 169, 162, 158, 146, 105, 63, 32, 29, 73, 121, 140, 143, 84, 
    220, 260, 253, 244, 242, 239, 242, 235, 229, 220, 211, 203, 202, 202, 196, 186, 180, 176, 172, 169, 166, 151, 110, 68, 55, 39, 57, 97, 131, 143, 141, 86, 
    192, 222, 223, 223, 225, 220, 218, 210, 204, 198, 192, 188, 189, 189, 185, 177, 174, 173, 168, 169, 168, 134, 81, 55, 50, 54, 85, 117, 138, 143, 135, 85, 
    162, 198, 198, 196, 195, 194, 195, 189, 185, 184, 184, 183, 186, 187, 183, 176, 174, 173, 170, 171, 149, 98, 49, 58, 67, 71, 102, 132, 148, 152, 142, 86, 
    139, 175, 177, 180, 179, 179, 179, 178, 179, 182, 185, 187, 190, 189, 189, 184, 176, 175, 174, 160, 119, 57, 13, 40, 91, 111, 135, 151, 157, 157, 149, 86, 
    130, 168, 173, 178, 180, 181, 181, 180, 182, 186, 191, 192, 192, 188, 189, 188, 176, 172, 173, 149, 95, 37, 1, 36, 104, 145, 159, 159, 153, 154, 150, 86, 
    131, 170, 178, 183, 184, 185, 188, 185, 186, 192, 200, 192, 176, 173, 174, 182, 174, 166, 161, 123, 70, 30, 6, 41, 105, 138, 153, 155, 150, 148, 148, 86, 
    135, 175, 183, 185, 185, 185, 188, 187, 187, 193, 196, 181, 164, 160, 152, 161, 158, 147, 137, 80, 29, 11, 0, 39, 94, 109, 120, 135, 142, 143, 144, 87, 
    142, 181, 186, 186, 186, 184, 184, 183, 183, 181, 178, 172, 160, 149, 124, 122, 125, 128, 137, 125, 90, 46, 0, 0, 49, 93, 102, 106, 125, 138, 139, 85, 
    149, 185, 188, 187, 187, 184, 179, 179, 177, 178, 167, 143, 122, 119, 109, 112, 123, 119, 114, 132, 158, 136, 35, 0, 0, 38, 102, 102, 102, 125, 132, 82, 
    152, 187, 187, 187, 189, 184, 177, 176, 177, 159, 124, 111, 111, 86, 54, 55, 71, 58, 38, 74, 124, 142, 100, 0, 0, 0, 58, 90, 84, 107, 121, 75, 
    152, 187, 188, 187, 189, 177, 167, 169, 151, 112, 91, 88, 79, 47, 10, 0, 22, 31, 21, 53, 90, 110, 119, 52, 0, 0, 7, 44, 60, 79, 97, 61, 
    152, 188, 191, 187, 183, 174, 150, 127, 103, 82, 65, 64, 60, 36, 12, 4, 8, 38, 42, 45, 80, 104, 107, 75, 23, 0, 0, 16, 47, 59, 53, 33, 
    152, 188, 192, 186, 167, 151, 135, 90, 81, 40, 31, 57, 59, 52, 61, 51, 29, 45, 61, 83, 102, 106, 72, 55, 74, 63, 21, 30, 58, 65, 42, 11, 
    154, 187, 189, 176, 135, 90, 93, 82, 51, 26, 17, 34, 33, 68, 121, 113, 100, 117, 129, 131, 123, 91, 57, 46, 60, 89, 62, 44, 61, 88, 67, 1, 
    155, 187, 182, 171, 101, 25, 25, 41, 31, 18, 11, 20, 17, 42, 126, 141, 121, 124, 131, 131, 127, 112, 53, 19, 53, 78, 68, 52, 69, 98, 83, 2, 
    154, 189, 194, 161, 65, 0, 2, 30, 23, 0, 8, 26, 38, 55, 117, 118, 102, 105, 106, 109, 129, 150, 111, 51, 48, 59, 65, 74, 78, 79, 69, 12, 
    152, 196, 201, 143, 67, 0, 0, 17, 13, 0, 5, 10, 35, 77, 119, 102, 94, 95, 72, 69, 103, 150, 173, 125, 75, 68, 69, 72, 71, 54, 51, 22, 
    150, 184, 168, 141, 98, 21, 0, 4, 5, 0, 6, 5, 7, 53, 109, 95, 92, 68, 34, 37, 35, 46, 123, 161, 116, 76, 70, 73, 51, 40, 47, 21, 
    143, 153, 110, 95, 105, 47, 0, 0, 0, 0, 17, 25, 14, 40, 96, 91, 82, 40, 12, 18, 7, 0, 26, 119, 129, 85, 67, 42, 28, 30, 33, 17, 
    132, 138, 83, 26, 56, 50, 0, 0, 0, 1, 16, 33, 47, 82, 102, 88, 71, 24, 0, 12, 13, 13, 0, 57, 116, 83, 41, 16, 9, 19, 33, 18, 
    118, 128, 81, 25, 42, 54, 0, 0, 0, 9, 13, 26, 52, 87, 101, 94, 74, 16, 0, 24, 8, 0, 0, 23, 95, 91, 35, 5, 5, 26, 43, 28, 
    100, 107, 78, 42, 44, 54, 0, 0, 4, 17, 23, 23, 36, 76, 93, 92, 71, 6, 0, 35, 22, 2, 0, 2, 63, 88, 38, 2, 9, 31, 47, 31, 
    82, 88, 73, 47, 40, 55, 13, 0, 15, 33, 52, 56, 54, 78, 89, 90, 74, 11, 0, 45, 47, 12, 0, 0, 28, 65, 32, 2, 9, 25, 37, 22, 
    73, 80, 77, 56, 41, 46, 27, 16, 29, 48, 75, 93, 98, 101, 100, 102, 100, 53, 19, 35, 45, 37, 14, 0, 0, 29, 25, 5, 3, 13, 24, 15, 
    76, 82, 65, 55, 37, 32, 20, 11, 14, 20, 29, 36, 40, 45, 45, 45, 50, 41, 38, 51, 28, 29, 0, 0, 0, 1, 0, 0, 0, 4, 14, 8, 
    79, 85, 63, 33, 14, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 47, 55, 22, 7, 0, 0, 0, 0, 0, 0, 3, 9, 2, 
    76, 82, 67, 36, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 25, 28, 12, 0, 0, 0, 0, 0, 0, 3, 8, 0, 
    64, 72, 68, 52, 31, 15, 13, 7, 0, 2, 2, 4, 8, 7, 8, 6, 3, 0, 0, 1, 5, 1, 0, 0, 0, 0, 0, 0, 3, 7, 12, 2, 
    
    -- channel=112
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=113
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 4, 5, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 3, 2, 2, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 8, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 13, 22, 33, 37, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 23, 29, 32, 36, 44, 54, 41, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 41, 43, 46, 41, 26, 21, 21, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 54, 55, 54, 41, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 54, 50, 47, 43, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 37, 25, 19, 20, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 9, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=114
    201, 92, 88, 92, 101, 105, 101, 89, 94, 118, 125, 112, 107, 102, 95, 86, 85, 91, 98, 97, 92, 92, 89, 87, 89, 91, 94, 100, 95, 90, 94, 67, 
    243, 136, 130, 130, 144, 149, 140, 139, 150, 173, 201, 193, 162, 149, 147, 139, 129, 125, 131, 132, 126, 126, 120, 116, 118, 116, 117, 118, 110, 102, 106, 58, 
    241, 134, 131, 126, 143, 149, 123, 150, 183, 178, 206, 231, 200, 164, 162, 164, 147, 135, 134, 132, 129, 133, 126, 122, 121, 117, 114, 113, 108, 103, 108, 43, 
    242, 135, 133, 126, 140, 148, 106, 148, 213, 194, 213, 253, 257, 226, 203, 193, 165, 148, 143, 135, 129, 129, 127, 124, 123, 124, 123, 117, 113, 110, 112, 37, 
    239, 139, 140, 130, 136, 146, 120, 147, 206, 207, 224, 250, 268, 271, 260, 250, 211, 169, 148, 133, 134, 132, 136, 135, 132, 136, 135, 126, 123, 123, 123, 46, 
    235, 139, 144, 138, 126, 130, 149, 181, 197, 216, 240, 255, 265, 277, 285, 283, 263, 230, 190, 150, 145, 152, 155, 149, 138, 143, 143, 132, 129, 130, 130, 54, 
    233, 140, 143, 141, 118, 100, 132, 202, 226, 233, 258, 267, 272, 282, 299, 298, 278, 270, 255, 205, 170, 169, 169, 162, 148, 140, 133, 128, 128, 130, 131, 56, 
    230, 143, 144, 139, 116, 75, 73, 166, 235, 248, 262, 253, 253, 268, 280, 295, 289, 273, 274, 258, 226, 211, 191, 167, 161, 144, 126, 126, 133, 139, 141, 50, 
    232, 141, 140, 135, 126, 76, 32, 125, 231, 258, 279, 254, 238, 243, 240, 264, 293, 289, 280, 276, 271, 259, 237, 196, 173, 158, 136, 136, 141, 146, 152, 45, 
    249, 138, 140, 140, 146, 78, 22, 129, 224, 246, 293, 283, 257, 246, 222, 243, 287, 295, 291, 290, 294, 296, 286, 249, 205, 179, 154, 150, 155, 157, 159, 41, 
    298, 148, 152, 154, 159, 70, 6, 143, 223, 210, 265, 295, 266, 263, 241, 240, 282, 289, 286, 298, 303, 302, 305, 285, 247, 217, 184, 165, 162, 160, 159, 38, 
    336, 158, 157, 159, 163, 85, 0, 114, 230, 205, 226, 271, 248, 240, 262, 253, 275, 278, 265, 284, 301, 291, 295, 301, 264, 238, 212, 178, 163, 156, 151, 38, 
    344, 162, 159, 157, 161, 117, 13, 51, 210, 245, 239, 260, 249, 224, 252, 267, 277, 272, 246, 262, 286, 282, 283, 311, 280, 234, 224, 190, 160, 148, 141, 44, 
    337, 161, 158, 154, 158, 142, 66, 10, 101, 204, 250, 285, 282, 255, 259, 278, 282, 270, 237, 243, 267, 273, 278, 310, 298, 235, 221, 199, 157, 140, 136, 49, 
    324, 159, 158, 156, 158, 151, 122, 74, 44, 69, 155, 263, 270, 244, 263, 286, 289, 270, 239, 231, 248, 266, 278, 298, 304, 248, 210, 203, 166, 142, 137, 41, 
    323, 162, 158, 158, 159, 147, 141, 177, 137, 46, 64, 182, 226, 199, 236, 281, 300, 285, 251, 237, 242, 263, 280, 284, 297, 264, 207, 199, 174, 150, 144, 45, 
    330, 169, 168, 169, 165, 136, 92, 177, 216, 100, 86, 125, 191, 186, 187, 255, 295, 290, 263, 244, 245, 260, 277, 275, 286, 277, 223, 209, 188, 153, 150, 70, 
    344, 172, 170, 167, 157, 131, 52, 86, 236, 173, 118, 102, 155, 219, 171, 225, 286, 285, 268, 251, 250, 260, 269, 270, 278, 284, 242, 217, 198, 157, 146, 84, 
    355, 159, 156, 156, 155, 154, 104, 34, 152, 234, 195, 109, 111, 242, 196, 213, 279, 284, 269, 260, 259, 261, 262, 265, 273, 282, 243, 198, 183, 153, 147, 85, 
    394, 152, 158, 156, 134, 169, 209, 117, 113, 237, 262, 167, 115, 239, 241, 223, 272, 282, 269, 266, 267, 265, 260, 263, 272, 274, 233, 172, 160, 150, 144, 81, 
    458, 154, 157, 145, 72, 117, 256, 228, 186, 244, 270, 221, 191, 248, 265, 252, 275, 280, 271, 270, 267, 263, 264, 267, 272, 269, 235, 164, 136, 145, 143, 75, 
    478, 158, 156, 135, 34, 46, 194, 210, 219, 257, 261, 258, 262, 261, 252, 272, 291, 284, 277, 276, 269, 260, 261, 261, 256, 252, 241, 185, 124, 132, 148, 74, 
    472, 155, 162, 157, 93, 79, 155, 155, 157, 220, 257, 281, 295, 259, 187, 213, 290, 295, 288, 286, 269, 256, 255, 250, 240, 236, 237, 213, 143, 117, 147, 79, 
    454, 170, 161, 156, 144, 138, 156, 156, 123, 139, 211, 269, 296, 263, 163, 129, 215, 267, 270, 281, 270, 251, 245, 234, 213, 218, 232, 227, 182, 123, 129, 76, 
    366, 166, 163, 156, 154, 151, 151, 157, 144, 114, 128, 198, 255, 255, 192, 149, 184, 240, 260, 277, 268, 231, 227, 239, 210, 188, 210, 220, 215, 163, 118, 62, 
    297, 163, 164, 159, 152, 150, 155, 160, 163, 153, 142, 159, 212, 242, 229, 197, 197, 243, 269, 290, 283, 226, 208, 241, 245, 208, 190, 201, 216, 205, 140, 45, 
    274, 158, 158, 161, 162, 161, 162, 165, 169, 176, 183, 162, 159, 212, 249, 227, 207, 241, 268, 291, 301, 251, 220, 242, 260, 238, 203, 194, 204, 216, 179, 49, 
    253, 157, 161, 165, 171, 174, 174, 173, 172, 181, 200, 179, 145, 178, 220, 220, 214, 234, 250, 258, 282, 273, 248, 245, 249, 233, 209, 200, 199, 202, 200, 74, 
    252, 155, 161, 167, 177, 180, 173, 172, 173, 190, 209, 188, 160, 178, 195, 190, 199, 212, 223, 219, 232, 256, 258, 248, 235, 213, 198, 199, 195, 186, 193, 92, 
    258, 160, 162, 167, 177, 178, 168, 164, 167, 190, 214, 195, 177, 179, 179, 179, 182, 185, 197, 194, 195, 220, 231, 227, 218, 198, 184, 189, 189, 176, 175, 96, 
    237, 161, 160, 167, 175, 176, 170, 165, 164, 186, 214, 194, 187, 176, 161, 178, 178, 180, 193, 186, 178, 191, 194, 188, 193, 185, 172, 175, 182, 174, 164, 91, 
    193, 169, 171, 175, 183, 180, 182, 183, 179, 189, 216, 213, 207, 204, 180, 184, 188, 190, 197, 195, 188, 190, 190, 183, 187, 187, 179, 178, 181, 181, 174, 125, 
    
    -- channel=115
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=116
    0, 59, 61, 56, 49, 46, 53, 65, 64, 57, 66, 77, 74, 61, 58, 60, 58, 50, 45, 43, 44, 39, 36, 34, 29, 25, 20, 14, 19, 23, 18, 38, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 23, 17, 3, 2, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 22, 20, 74, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 39, 24, 7, 4, 1, 0, 0, 6, 1, 7, 12, 17, 23, 25, 25, 36, 40, 32, 109, 
    0, 0, 0, 1, 0, 0, 34, 0, 0, 0, 0, 0, 0, 12, 23, 18, 22, 13, 0, 12, 27, 32, 38, 42, 43, 40, 36, 35, 40, 42, 33, 136, 
    0, 0, 0, 0, 0, 0, 46, 0, 0, 0, 0, 0, 0, 0, 0, 6, 30, 31, 25, 36, 47, 48, 45, 43, 43, 32, 28, 32, 33, 32, 28, 140, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 12, 13, 27, 31, 29, 25, 34, 41, 21, 15, 21, 25, 27, 30, 137, 
    0, 0, 0, 0, 11, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 18, 19, 31, 33, 21, 21, 29, 35, 41, 45, 143, 
    0, 0, 0, 0, 45, 100, 84, 0, 0, 0, 0, 0, 13, 4, 0, 0, 11, 0, 0, 0, 0, 0, 18, 39, 40, 34, 41, 41, 40, 46, 52, 162, 
    0, 7, 13, 34, 67, 133, 171, 41, 0, 0, 0, 3, 29, 26, 34, 16, 15, 25, 2, 0, 0, 0, 17, 50, 44, 39, 51, 54, 57, 62, 66, 193, 
    0, 36, 36, 39, 32, 120, 203, 58, 0, 0, 0, 0, 0, 17, 57, 39, 8, 16, 21, 4, 0, 0, 0, 22, 31, 38, 62, 74, 74, 70, 67, 214, 
    0, 20, 13, 9, 2, 143, 222, 50, 0, 0, 0, 0, 0, 0, 33, 36, 8, 12, 21, 16, 4, 0, 0, 0, 9, 21, 51, 73, 74, 72, 70, 225, 
    0, 2, 1, 1, 0, 152, 235, 55, 0, 22, 0, 0, 0, 0, 11, 21, 3, 11, 29, 19, 14, 17, 0, 0, 0, 7, 32, 66, 77, 73, 67, 217, 
    0, 0, 0, 0, 0, 104, 233, 100, 0, 0, 0, 0, 7, 25, 7, 7, 0, 2, 34, 22, 13, 30, 9, 0, 0, 12, 20, 48, 64, 61, 54, 192, 
    0, 0, 0, 2, 0, 51, 197, 195, 41, 0, 0, 0, 0, 7, 0, 0, 0, 0, 36, 31, 16, 31, 19, 0, 0, 16, 8, 20, 46, 49, 44, 166, 
    0, 0, 0, 7, 10, 30, 118, 205, 162, 94, 0, 0, 0, 16, 11, 0, 0, 2, 35, 37, 28, 30, 22, 0, 0, 12, 10, 3, 31, 43, 48, 169, 
    0, 1, 10, 16, 17, 29, 44, 62, 123, 215, 142, 2, 0, 52, 30, 0, 0, 0, 11, 30, 32, 27, 19, 0, 0, 4, 28, 16, 36, 54, 49, 179, 
    0, 6, 10, 10, 20, 67, 104, 22, 46, 207, 206, 61, 35, 68, 76, 14, 0, 0, 0, 20, 33, 26, 17, 15, 0, 0, 30, 19, 27, 45, 41, 161, 
    0, 7, 20, 36, 63, 130, 231, 108, 2, 99, 156, 135, 65, 42, 106, 45, 0, 0, 0, 10, 24, 24, 17, 23, 0, 0, 6, 0, 5, 46, 60, 147, 
    0, 49, 66, 68, 66, 75, 190, 185, 15, 27, 68, 172, 95, 0, 86, 68, 0, 0, 0, 0, 7, 18, 23, 29, 2, 0, 0, 11, 23, 68, 81, 141, 
    0, 61, 50, 33, 27, 0, 2, 148, 64, 0, 0, 135, 112, 0, 49, 69, 0, 0, 0, 0, 0, 9, 25, 28, 7, 0, 18, 59, 64, 74, 73, 137, 
    0, 26, 23, 38, 99, 20, 0, 2, 38, 0, 0, 52, 80, 0, 4, 36, 0, 0, 0, 0, 0, 4, 19, 18, 6, 0, 26, 85, 92, 78, 72, 143, 
    0, 26, 24, 53, 200, 134, 0, 0, 9, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 5, 21, 29, 26, 7, 12, 75, 114, 97, 76, 150, 
    0, 3, 0, 0, 152, 147, 37, 46, 27, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 14, 26, 35, 37, 20, 0, 42, 120, 121, 83, 154, 
    0, 0, 0, 0, 53, 55, 3, 37, 77, 52, 2, 0, 0, 0, 82, 54, 0, 0, 0, 0, 0, 1, 13, 38, 63, 50, 3, 9, 91, 136, 106, 162, 
    0, 0, 0, 0, 0, 0, 0, 18, 83, 113, 77, 14, 0, 0, 60, 90, 13, 0, 0, 0, 0, 6, 18, 36, 85, 84, 44, 9, 43, 113, 128, 180, 
    0, 0, 0, 0, 0, 2, 13, 9, 20, 62, 72, 20, 0, 0, 2, 50, 23, 0, 0, 0, 0, 12, 24, 10, 52, 88, 73, 42, 17, 60, 126, 200, 
    0, 0, 0, 0, 5, 7, 4, 0, 0, 0, 17, 37, 26, 0, 0, 10, 22, 0, 0, 0, 0, 0, 12, 0, 1, 53, 75, 61, 24, 21, 90, 206, 
    0, 3, 3, 0, 0, 0, 0, 6, 19, 17, 3, 51, 83, 27, 0, 6, 18, 0, 0, 0, 0, 0, 0, 0, 0, 27, 56, 57, 44, 22, 44, 188, 
    0, 5, 0, 0, 0, 3, 23, 38, 47, 27, 0, 34, 84, 44, 18, 32, 35, 15, 0, 0, 0, 0, 0, 0, 0, 28, 50, 49, 53, 46, 28, 162, 
    0, 0, 0, 8, 16, 35, 57, 62, 56, 23, 0, 29, 62, 43, 58, 65, 68, 58, 37, 38, 20, 0, 0, 0, 11, 47, 61, 52, 55, 64, 42, 145, 
    0, 8, 25, 37, 38, 46, 59, 60, 61, 26, 0, 33, 51, 59, 84, 72, 75, 71, 50, 55, 57, 33, 27, 39, 44, 64, 76, 63, 55, 63, 59, 138, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 65, 
    
    -- channel=117
    77, 58, 55, 53, 56, 63, 67, 63, 60, 65, 68, 63, 56, 55, 52, 47, 43, 39, 39, 38, 32, 30, 26, 20, 17, 13, 11, 12, 8, 4, 4, 0, 
    59, 0, 0, 0, 0, 5, 0, 0, 0, 0, 1, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    58, 0, 0, 0, 0, 2, 0, 0, 5, 0, 0, 10, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 5, 5, 8, 0, 
    57, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 2, 3, 3, 3, 2, 0, 0, 0, 0, 0, 0, 5, 8, 11, 16, 20, 19, 15, 9, 5, 0, 
    53, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 5, 10, 15, 16, 12, 14, 19, 23, 23, 18, 18, 16, 8, 1, 0, 0, 0, 
    50, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 1, 5, 12, 30, 41, 29, 17, 16, 19, 12, 2, 2, 0, 0, 0, 0, 0, 0, 
    48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 12, 18, 14, 14, 25, 21, 12, 8, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    48, 0, 1, 3, 0, 0, 0, 0, 0, 0, 6, 3, 1, 7, 8, 8, 11, 10, 7, 4, 7, 11, 4, 0, 0, 1, 0, 0, 0, 0, 4, 0, 
    61, 15, 24, 30, 40, 15, 0, 0, 8, 7, 26, 29, 28, 25, 8, 3, 7, 9, 11, 8, 6, 9, 7, 2, 6, 8, 5, 5, 7, 8, 10, 0, 
    97, 44, 52, 56, 59, 3, 0, 0, 8, 0, 22, 33, 31, 27, 5, 0, 11, 9, 6, 10, 10, 10, 12, 10, 13, 17, 12, 12, 14, 16, 15, 0, 
    125, 56, 54, 49, 41, 0, 0, 0, 13, 0, 11, 25, 12, 6, 0, 0, 8, 10, 4, 6, 11, 8, 8, 6, 7, 20, 21, 17, 15, 11, 6, 0, 
    127, 36, 28, 20, 16, 0, 0, 0, 20, 14, 27, 36, 12, 0, 0, 0, 11, 12, 2, 5, 11, 7, 6, 12, 10, 13, 19, 14, 8, 3, 0, 0, 
    118, 15, 11, 8, 7, 0, 0, 0, 3, 24, 37, 43, 22, 2, 0, 0, 15, 16, 2, 3, 8, 3, 3, 19, 18, 11, 14, 10, 0, 0, 0, 0, 
    106, 6, 4, 3, 7, 4, 0, 0, 0, 0, 0, 13, 11, 0, 4, 9, 19, 20, 5, 1, 3, 0, 0, 17, 18, 5, 6, 4, 0, 0, 0, 0, 
    101, 4, 7, 13, 20, 16, 6, 12, 21, 0, 0, 0, 2, 0, 0, 14, 29, 27, 10, 2, 0, 0, 0, 10, 16, 0, 0, 0, 0, 0, 0, 0, 
    106, 18, 22, 26, 26, 10, 0, 14, 32, 13, 8, 27, 26, 4, 1, 18, 30, 28, 13, 0, 0, 0, 2, 5, 14, 4, 0, 2, 1, 0, 2, 0, 
    116, 27, 30, 34, 36, 21, 0, 6, 41, 12, 19, 44, 37, 23, 0, 9, 22, 16, 5, 0, 0, 0, 4, 2, 10, 11, 1, 13, 13, 0, 0, 0, 
    125, 37, 43, 54, 62, 60, 24, 19, 54, 40, 30, 3, 8, 22, 0, 5, 18, 17, 6, 0, 0, 3, 4, 0, 6, 14, 1, 0, 0, 0, 0, 0, 
    158, 63, 73, 81, 82, 83, 65, 21, 20, 10, 29, 0, 0, 19, 0, 0, 15, 17, 9, 4, 7, 9, 3, 0, 2, 9, 0, 0, 0, 0, 0, 0, 
    207, 86, 88, 80, 36, 12, 23, 0, 0, 3, 10, 0, 0, 14, 0, 0, 15, 17, 10, 8, 10, 9, 2, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    221, 75, 63, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 19, 19, 12, 12, 9, 1, 0, 0, 0, 1, 3, 0, 0, 0, 0, 0, 
    210, 38, 30, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 14, 7, 5, 2, 0, 0, 0, 0, 0, 11, 12, 0, 0, 0, 0, 
    191, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 1, 4, 4, 4, 0, 0, 0, 16, 19, 0, 0, 0, 0, 
    123, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 17, 23, 0, 0, 0, 0, 0, 4, 16, 16, 13, 3, 0, 0, 7, 18, 8, 0, 0, 0, 
    70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 19, 0, 0, 12, 21, 18, 31, 38, 19, 2, 1, 0, 0, 0, 10, 12, 5, 0, 0, 
    64, 0, 0, 0, 0, 0, 0, 1, 3, 1, 7, 12, 12, 12, 3, 0, 0, 14, 18, 35, 44, 19, 0, 0, 0, 0, 4, 4, 11, 10, 0, 0, 
    57, 0, 0, 0, 0, 4, 2, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 8, 9, 18, 27, 7, 0, 0, 0, 0, 0, 3, 9, 10, 0, 0, 
    55, 0, 1, 5, 2, 0, 0, 0, 0, 0, 4, 2, 0, 7, 8, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 6, 2, 0, 
    63, 2, 0, 0, 0, 0, 0, 0, 0, 1, 25, 16, 0, 8, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    44, 0, 0, 0, 0, 0, 0, 0, 0, 10, 24, 13, 2, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 6, 21, 9, 1, 0, 0, 0, 0, 1, 6, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=118
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=119
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 10, 7, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 8, 6, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 3, 4, 8, 12, 14, 12, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 11, 10, 9, 10, 14, 14, 12, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 12, 13, 12, 11, 13, 13, 8, 5, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 13, 14, 11, 12, 12, 8, 7, 8, 8, 5, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 6, 3, 11, 10, 7, 9, 8, 6, 9, 12, 15, 10, 8, 9, 8, 9, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 12, 1, 4, 1, 0, 4, 3, 7, 13, 12, 14, 14, 15, 15, 14, 12, 8, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 10, 0, 0, 0, 0, 0, 0, 7, 15, 12, 11, 12, 14, 14, 13, 11, 8, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 5, 0, 1, 5, 0, 0, 3, 9, 14, 11, 8, 8, 10, 10, 11, 12, 8, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 5, 8, 10, 11, 5, 7, 8, 7, 9, 13, 11, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 8, 8, 9, 5, 9, 9, 8, 10, 15, 12, 5, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 7, 6, 7, 4, 7, 8, 9, 12, 16, 11, 5, 4, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 8, 0, 0, 0, 1, 3, 3, 1, 4, 6, 10, 13, 16, 12, 8, 4, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 0, 0, 0, 0, 1, 1, 0, 2, 5, 11, 13, 14, 13, 11, 6, 9, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 3, 2, 2, 5, 10, 11, 12, 13, 13, 7, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 5, 3, 2, 5, 8, 9, 11, 13, 14, 8, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 12, 6, 3, 3, 4, 4, 6, 9, 13, 13, 7, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 18, 7, 1, 8, 3, 2, 4, 3, 0, 1, 7, 12, 12, 6, 2, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 5, 18, 7, 0, 0, 0, 0, 2, 1, 0, 1, 8, 10, 9, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 13, 10, 0, 0, 0, 0, 0, 0, 2, 4, 6, 6, 5, 4, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 1, 0, 0, 1, 0, 0, 4, 6, 5, 2, 0, 1, 3, 3, 0, 0, 0, 4, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 15, 8, 2, 5, 5, 0, 0, 0, 3, 8, 9, 0, 0, 0, 1, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 10, 6, 5, 2, 0, 0, 0, 5, 12, 11, 6, 0, 0, 0, 1, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 5, 0, 0, 0, 0, 3, 6, 9, 10, 7, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 1, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=120
    33, 89, 90, 83, 78, 78, 86, 92, 88, 79, 80, 84, 82, 78, 78, 77, 72, 66, 60, 60, 59, 54, 51, 46, 39, 33, 26, 21, 22, 18, 12, 18, 
    0, 88, 90, 83, 72, 73, 83, 81, 73, 64, 60, 72, 80, 78, 70, 72, 73, 67, 58, 56, 54, 49, 47, 41, 35, 29, 23, 20, 23, 25, 21, 41, 
    0, 88, 87, 85, 70, 75, 84, 53, 51, 65, 53, 54, 73, 78, 67, 63, 65, 60, 53, 50, 47, 40, 36, 34, 33, 32, 33, 34, 38, 41, 36, 62, 
    0, 86, 86, 86, 71, 72, 80, 44, 39, 57, 44, 31, 41, 57, 57, 51, 57, 53, 48, 46, 48, 44, 44, 48, 49, 49, 51, 52, 53, 53, 48, 74, 
    0, 82, 81, 83, 74, 65, 71, 52, 25, 34, 30, 16, 13, 26, 32, 30, 43, 51, 58, 64, 66, 65, 62, 65, 64, 59, 60, 62, 59, 54, 47, 71, 
    0, 76, 74, 76, 76, 62, 44, 28, 18, 25, 20, 12, 9, 3, 4, 12, 27, 45, 64, 84, 80, 73, 68, 73, 72, 64, 59, 58, 51, 43, 36, 64, 
    0, 72, 69, 70, 73, 55, 21, 0, 14, 18, 10, 5, 1, 0, 0, 0, 12, 24, 39, 70, 78, 75, 77, 71, 65, 61, 57, 54, 48, 39, 32, 64, 
    0, 69, 68, 69, 71, 78, 62, 4, 0, 11, 8, 12, 8, 6, 2, 0, 4, 10, 17, 39, 61, 67, 69, 65, 59, 60, 61, 56, 47, 37, 30, 72, 
    0, 72, 81, 92, 104, 135, 115, 26, 0, 8, 11, 29, 35, 35, 31, 7, 2, 12, 14, 17, 30, 41, 54, 67, 60, 57, 58, 51, 44, 38, 35, 87, 
    4, 106, 120, 132, 142, 172, 136, 41, 5, 13, 0, 23, 48, 58, 60, 30, 7, 11, 13, 11, 11, 20, 32, 51, 55, 49, 53, 52, 49, 44, 40, 95, 
    17, 138, 145, 153, 157, 187, 154, 41, 7, 23, 0, 11, 52, 57, 62, 45, 18, 16, 14, 7, 5, 10, 14, 29, 40, 38, 48, 52, 49, 48, 45, 100, 
    9, 150, 155, 160, 162, 185, 176, 49, 3, 35, 27, 25, 61, 61, 55, 51, 27, 27, 27, 10, 6, 14, 11, 13, 28, 28, 35, 49, 54, 55, 52, 98, 
    2, 151, 154, 153, 154, 167, 184, 92, 4, 21, 40, 40, 64, 78, 51, 45, 33, 38, 41, 23, 11, 17, 16, 5, 26, 28, 27, 48, 58, 58, 51, 87, 
    0, 143, 144, 145, 143, 149, 170, 144, 48, 24, 20, 15, 38, 62, 42, 32, 35, 45, 57, 44, 25, 21, 19, 4, 17, 39, 27, 41, 58, 55, 44, 78, 
    0, 137, 137, 139, 141, 149, 158, 160, 127, 79, 21, 0, 20, 44, 35, 25, 36, 56, 73, 64, 42, 27, 19, 9, 8, 41, 36, 32, 46, 46, 43, 85, 
    0, 136, 139, 144, 150, 157, 146, 119, 143, 134, 87, 32, 40, 58, 37, 23, 36, 60, 76, 73, 53, 32, 21, 17, 9, 33, 43, 28, 41, 49, 46, 85, 
    1, 141, 145, 148, 152, 162, 167, 105, 118, 182, 156, 100, 55, 76, 65, 33, 35, 55, 73, 73, 58, 40, 28, 26, 16, 25, 47, 37, 43, 44, 28, 55, 
    2, 144, 150, 160, 181, 208, 241, 190, 124, 179, 165, 160, 83, 77, 90, 50, 40, 54, 69, 71, 62, 50, 38, 34, 25, 21, 45, 36, 23, 17, 0, 34, 
    7, 176, 196, 218, 240, 250, 272, 275, 160, 149, 161, 184, 122, 53, 89, 69, 44, 56, 66, 68, 64, 57, 51, 42, 33, 23, 37, 23, 0, 0, 0, 30, 
    36, 236, 247, 257, 269, 237, 223, 267, 195, 112, 131, 158, 133, 44, 74, 74, 49, 56, 66, 66, 64, 61, 58, 48, 36, 24, 26, 22, 0, 0, 0, 28, 
    43, 263, 264, 276, 292, 207, 137, 159, 155, 97, 92, 102, 110, 52, 50, 59, 47, 55, 64, 64, 61, 59, 52, 43, 31, 19, 18, 28, 7, 0, 0, 32, 
    28, 276, 280, 284, 286, 194, 97, 102, 110, 74, 53, 55, 62, 51, 37, 23, 27, 46, 55, 54, 50, 44, 40, 42, 34, 21, 9, 24, 29, 2, 0, 34, 
    30, 275, 257, 231, 220, 190, 119, 115, 99, 48, 23, 21, 22, 36, 52, 21, 0, 17, 30, 31, 36, 45, 50, 49, 38, 15, 0, 10, 39, 22, 0, 35, 
    7, 208, 183, 165, 166, 162, 120, 107, 104, 68, 29, 4, 1, 35, 73, 48, 0, 8, 23, 28, 43, 57, 56, 54, 46, 14, 0, 0, 24, 38, 9, 39, 
    0, 147, 146, 139, 123, 106, 95, 91, 104, 102, 68, 30, 16, 33, 62, 73, 34, 18, 31, 32, 53, 79, 75, 61, 52, 29, 0, 0, 2, 34, 34, 49, 
    0, 115, 105, 95, 89, 89, 91, 88, 86, 92, 84, 55, 23, 14, 35, 58, 48, 27, 33, 36, 63, 98, 91, 61, 49, 41, 9, 0, 0, 12, 40, 67, 
    0, 77, 76, 79, 84, 85, 80, 70, 57, 44, 39, 46, 31, 13, 19, 40, 45, 29, 30, 32, 47, 83, 89, 61, 39, 34, 20, 0, 0, 0, 23, 82, 
    0, 70, 72, 73, 68, 64, 51, 34, 19, 9, 9, 32, 43, 17, 15, 26, 26, 16, 14, 16, 15, 42, 63, 55, 42, 28, 7, 0, 0, 0, 0, 74, 
    0, 69, 60, 49, 36, 26, 16, 4, 0, 0, 0, 20, 40, 30, 18, 4, 0, 0, 0, 0, 0, 7, 25, 31, 27, 15, 0, 0, 0, 0, 0, 51, 
    0, 45, 29, 12, 1, 0, 0, 0, 0, 0, 0, 12, 28, 28, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 
    0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 15, 20, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=121
    140, 166, 164, 158, 154, 156, 164, 166, 154, 138, 130, 131, 136, 141, 147, 149, 146, 141, 138, 135, 133, 130, 128, 124, 119, 113, 109, 105, 104, 101, 100, 96, 
    103, 79, 78, 74, 70, 71, 70, 57, 42, 22, 8, 19, 39, 46, 48, 54, 63, 68, 66, 62, 59, 59, 61, 60, 61, 64, 68, 73, 78, 81, 87, 85, 
    103, 79, 79, 75, 71, 70, 57, 32, 27, 22, 0, 0, 14, 29, 29, 33, 42, 50, 55, 53, 46, 50, 56, 61, 71, 80, 88, 93, 95, 94, 94, 87, 
    101, 79, 80, 77, 71, 67, 54, 32, 23, 0, 0, 0, 0, 0, 0, 5, 21, 38, 53, 59, 62, 70, 76, 83, 87, 89, 93, 93, 88, 81, 74, 66, 
    97, 71, 74, 73, 65, 55, 46, 42, 20, 0, 0, 0, 0, 0, 0, 0, 0, 43, 79, 85, 83, 82, 80, 78, 73, 68, 67, 62, 52, 43, 37, 38, 
    95, 68, 67, 66, 58, 36, 10, 12, 1, 0, 0, 0, 0, 0, 0, 0, 0, 4, 56, 74, 66, 55, 50, 46, 39, 37, 37, 33, 26, 19, 17, 25, 
    91, 67, 68, 64, 56, 40, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 29, 30, 21, 12, 13, 28, 36, 32, 27, 23, 20, 31, 
    89, 67, 73, 79, 87, 93, 75, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 34, 44, 37, 27, 21, 19, 36, 
    103, 94, 110, 126, 137, 136, 98, 34, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 29, 31, 25, 21, 17, 13, 31, 
    135, 138, 147, 148, 140, 108, 40, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 12, 9, 7, 5, 1, 17, 
    141, 131, 123, 111, 97, 66, 10, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    122, 90, 78, 69, 62, 52, 35, 24, 14, 19, 28, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    109, 61, 56, 52, 51, 49, 57, 49, 13, 0, 9, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    102, 52, 50, 50, 55, 58, 72, 95, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    104, 56, 58, 62, 70, 69, 62, 87, 120, 85, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 18, 35, 
    108, 72, 76, 79, 76, 60, 23, 8, 52, 95, 94, 68, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 20, 18, 28, 
    112, 76, 74, 73, 76, 78, 59, 33, 48, 70, 100, 94, 43, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    114, 81, 88, 105, 129, 149, 158, 119, 72, 52, 62, 59, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    150, 136, 151, 161, 162, 148, 141, 132, 65, 0, 0, 33, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    192, 173, 160, 142, 97, 30, 0, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    179, 135, 115, 94, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    161, 92, 82, 62, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    143, 47, 10, 0, 0, 4, 60, 46, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    70, 0, 0, 0, 0, 12, 36, 25, 23, 5, 0, 0, 0, 0, 24, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    53, 0, 0, 9, 19, 20, 19, 17, 30, 58, 54, 26, 7, 0, 0, 5, 18, 3, 0, 0, 14, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    72, 12, 23, 27, 31, 33, 35, 34, 21, 13, 22, 19, 0, 0, 0, 0, 0, 0, 0, 0, 14, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    70, 27, 30, 35, 39, 38, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    74, 36, 39, 34, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    76, 35, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=122
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 4, 7, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 11, 20, 26, 29, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    46, 28, 32, 32, 32, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    55, 30, 32, 30, 30, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    52, 29, 29, 26, 24, 24, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    47, 22, 22, 20, 21, 21, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    39, 17, 18, 19, 20, 19, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 12, 15, 18, 24, 29, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    43, 19, 25, 33, 45, 48, 44, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    66, 41, 49, 60, 73, 78, 84, 50, 0, 2, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    104, 74, 84, 98, 108, 79, 81, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    136, 112, 117, 123, 114, 34, 25, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    158, 125, 123, 120, 99, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    157, 114, 104, 93, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    119, 85, 76, 57, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    75, 36, 23, 12, 7, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=123
    110, 202, 202, 198, 191, 189, 192, 202, 210, 216, 223, 226, 213, 195, 184, 181, 178, 175, 169, 166, 163, 152, 145, 139, 130, 122, 114, 108, 107, 104, 96, 93, 
    28, 118, 119, 116, 106, 97, 100, 102, 103, 121, 137, 147, 153, 139, 117, 108, 110, 109, 105, 104, 101, 92, 89, 87, 85, 83, 79, 76, 83, 91, 94, 110, 
    27, 116, 117, 117, 108, 100, 103, 88, 92, 141, 153, 153, 165, 171, 155, 130, 112, 99, 92, 99, 100, 93, 91, 94, 100, 104, 107, 109, 115, 118, 116, 132, 
    28, 116, 118, 121, 112, 102, 111, 100, 107, 151, 150, 139, 148, 167, 173, 158, 135, 110, 95, 106, 116, 121, 124, 132, 138, 136, 132, 128, 125, 121, 113, 134, 
    26, 110, 110, 116, 109, 102, 121, 116, 116, 136, 145, 142, 146, 163, 175, 170, 157, 138, 131, 145, 154, 156, 152, 149, 145, 132, 121, 116, 109, 101, 92, 119, 
    27, 107, 105, 108, 105, 98, 94, 86, 117, 155, 168, 174, 174, 175, 178, 184, 182, 160, 151, 157, 157, 146, 137, 135, 129, 110, 97, 91, 85, 80, 77, 110, 
    31, 109, 107, 108, 106, 92, 73, 80, 124, 166, 174, 175, 177, 181, 189, 192, 186, 160, 130, 125, 133, 139, 140, 127, 103, 89, 85, 87, 89, 91, 92, 121, 
    34, 112, 113, 115, 126, 147, 156, 131, 135, 171, 183, 193, 202, 200, 199, 195, 184, 169, 144, 130, 133, 144, 145, 135, 110, 95, 101, 105, 105, 105, 105, 138, 
    39, 129, 143, 163, 191, 230, 234, 169, 153, 184, 194, 212, 230, 230, 226, 207, 197, 199, 184, 164, 151, 152, 164, 163, 137, 112, 109, 112, 115, 118, 121, 156, 
    55, 181, 195, 208, 212, 232, 231, 158, 153, 174, 158, 170, 206, 224, 240, 227, 206, 209, 210, 198, 186, 178, 175, 171, 146, 120, 119, 126, 128, 127, 121, 159, 
    55, 192, 187, 181, 174, 207, 220, 149, 141, 169, 147, 145, 181, 200, 214, 226, 213, 210, 217, 216, 207, 199, 183, 169, 147, 121, 117, 121, 118, 114, 111, 156, 
    19, 157, 153, 151, 149, 197, 225, 160, 130, 179, 188, 183, 199, 208, 211, 219, 212, 209, 219, 216, 212, 213, 200, 177, 156, 126, 102, 105, 110, 107, 101, 144, 
    0, 138, 134, 132, 130, 175, 222, 182, 120, 133, 172, 189, 215, 230, 227, 216, 206, 204, 216, 212, 208, 216, 208, 188, 171, 142, 103, 93, 99, 93, 84, 124, 
    0, 120, 120, 123, 127, 155, 214, 213, 159, 118, 109, 109, 155, 199, 206, 206, 200, 203, 218, 219, 212, 217, 212, 188, 173, 152, 111, 82, 83, 80, 73, 116, 
    0, 124, 127, 131, 141, 159, 203, 231, 222, 188, 117, 75, 120, 187, 197, 202, 203, 216, 233, 233, 227, 223, 218, 193, 172, 158, 129, 88, 77, 81, 90, 138, 
    11, 144, 149, 155, 161, 166, 164, 163, 192, 236, 209, 173, 176, 208, 208, 197, 198, 209, 226, 233, 231, 226, 223, 207, 182, 170, 154, 117, 106, 115, 115, 145, 
    21, 163, 163, 160, 158, 172, 186, 156, 166, 274, 284, 217, 190, 192, 225, 205, 187, 196, 210, 225, 230, 230, 230, 222, 195, 180, 175, 151, 128, 114, 86, 102, 
    18, 162, 164, 175, 201, 253, 305, 278, 218, 227, 256, 222, 189, 168, 224, 218, 195, 199, 211, 224, 233, 236, 237, 234, 209, 186, 176, 141, 93, 63, 46, 82, 
    19, 203, 227, 247, 258, 267, 307, 302, 233, 184, 198, 230, 196, 138, 196, 225, 206, 204, 213, 223, 229, 237, 243, 243, 221, 190, 164, 115, 61, 47, 58, 92, 
    37, 260, 253, 234, 213, 168, 159, 224, 204, 150, 144, 202, 184, 144, 185, 222, 212, 211, 217, 220, 224, 233, 244, 244, 225, 188, 158, 122, 81, 61, 63, 94, 
    1, 218, 200, 194, 196, 125, 33, 96, 139, 133, 123, 163, 176, 158, 175, 196, 203, 216, 222, 218, 216, 220, 225, 224, 214, 180, 155, 137, 107, 74, 62, 94, 
    0, 189, 187, 191, 210, 156, 77, 119, 158, 140, 128, 143, 163, 156, 150, 143, 158, 197, 209, 201, 192, 193, 206, 221, 218, 181, 142, 127, 122, 96, 68, 96, 
    0, 173, 138, 109, 149, 177, 181, 197, 191, 155, 139, 151, 156, 151, 153, 134, 110, 137, 166, 166, 171, 193, 218, 230, 214, 164, 114, 106, 122, 114, 81, 97, 
    0, 70, 44, 54, 109, 143, 146, 155, 168, 183, 179, 163, 153, 166, 185, 157, 127, 140, 170, 181, 188, 203, 214, 218, 207, 159, 99, 82, 102, 121, 106, 110, 
    0, 50, 81, 100, 97, 86, 84, 114, 163, 201, 212, 199, 171, 163, 181, 184, 173, 177, 196, 197, 198, 217, 226, 220, 210, 177, 118, 74, 82, 111, 124, 129, 
    0, 98, 96, 88, 87, 99, 114, 124, 136, 160, 170, 165, 137, 119, 141, 174, 184, 180, 187, 188, 195, 225, 231, 215, 209, 183, 140, 93, 72, 89, 117, 144, 
    5, 85, 87, 103, 121, 129, 122, 105, 83, 71, 79, 99, 112, 111, 122, 159, 179, 173, 172, 159, 151, 181, 209, 204, 192, 177, 143, 99, 68, 71, 98, 144, 
    16, 107, 115, 117, 115, 105, 89, 67, 54, 52, 67, 107, 132, 124, 121, 141, 144, 138, 135, 117, 104, 126, 167, 190, 189, 168, 127, 85, 65, 62, 75, 126, 
    34, 119, 105, 87, 72, 65, 63, 63, 65, 63, 63, 97, 130, 131, 121, 112, 102, 101, 101, 98, 95, 104, 128, 147, 149, 134, 105, 73, 60, 58, 57, 103, 
    20, 81, 60, 48, 48, 61, 75, 78, 70, 55, 50, 80, 110, 114, 108, 90, 85, 83, 85, 98, 100, 90, 88, 90, 90, 95, 88, 66, 53, 54, 52, 91, 
    0, 39, 42, 49, 56, 64, 67, 68, 68, 54, 45, 71, 94, 100, 104, 81, 69, 70, 72, 81, 85, 78, 72, 70, 67, 73, 73, 61, 50, 50, 53, 88, 
    0, 3, 8, 7, 2, 0, 0, 4, 8, 0, 0, 0, 0, 7, 11, 4, 3, 2, 3, 8, 12, 10, 9, 8, 3, 3, 6, 5, 1, 2, 6, 33, 
    
    -- channel=124
    77, 126, 123, 117, 118, 126, 136, 141, 137, 137, 139, 132, 121, 114, 111, 104, 92, 82, 77, 74, 68, 60, 51, 40, 29, 18, 10, 6, 3, 0, 0, 0, 
    72, 98, 95, 87, 88, 93, 99, 99, 96, 94, 99, 103, 97, 81, 74, 72, 68, 62, 56, 51, 42, 32, 24, 15, 6, 0, 0, 0, 0, 0, 0, 0, 
    70, 94, 91, 84, 83, 91, 84, 68, 79, 88, 89, 101, 109, 95, 74, 66, 61, 55, 49, 45, 34, 26, 22, 16, 14, 14, 18, 23, 30, 29, 31, 10, 
    69, 95, 93, 88, 84, 89, 70, 44, 73, 91, 79, 80, 93, 96, 83, 70, 57, 45, 45, 48, 45, 43, 45, 48, 54, 59, 67, 71, 71, 64, 57, 26, 
    63, 87, 88, 87, 79, 79, 67, 47, 67, 66, 51, 48, 54, 62, 65, 67, 67, 62, 69, 80, 87, 92, 95, 98, 96, 92, 93, 90, 82, 71, 58, 23, 
    56, 78, 78, 81, 72, 57, 43, 41, 53, 45, 44, 48, 50, 51, 52, 58, 71, 87, 115, 125, 123, 121, 119, 116, 106, 95, 91, 83, 69, 54, 41, 9, 
    51, 73, 71, 73, 65, 34, 0, 4, 29, 39, 42, 44, 45, 48, 59, 73, 77, 78, 103, 122, 121, 118, 116, 111, 97, 83, 74, 66, 57, 47, 39, 10, 
    49, 72, 75, 79, 78, 60, 20, 2, 18, 28, 40, 46, 48, 54, 65, 76, 78, 69, 70, 86, 102, 115, 115, 99, 84, 82, 78, 71, 65, 61, 56, 25, 
    59, 91, 104, 122, 145, 151, 98, 32, 24, 36, 65, 90, 96, 100, 92, 78, 77, 75, 71, 71, 79, 94, 105, 102, 95, 96, 92, 84, 79, 77, 77, 45, 
    101, 153, 180, 206, 227, 218, 123, 34, 32, 36, 62, 103, 123, 133, 119, 91, 83, 80, 76, 72, 73, 81, 96, 107, 106, 109, 108, 105, 105, 104, 102, 61, 
    161, 225, 241, 250, 253, 223, 104, 26, 41, 35, 41, 83, 112, 124, 119, 97, 88, 87, 82, 77, 76, 75, 77, 89, 99, 116, 127, 126, 121, 115, 107, 62, 
    187, 241, 243, 243, 240, 220, 113, 33, 50, 62, 68, 99, 115, 105, 101, 96, 93, 97, 92, 85, 83, 79, 69, 78, 92, 108, 126, 129, 124, 115, 105, 58, 
    186, 232, 231, 226, 220, 214, 147, 55, 46, 77, 105, 129, 139, 117, 102, 95, 96, 108, 103, 92, 89, 83, 67, 76, 99, 107, 117, 123, 119, 105, 87, 41, 
    172, 212, 210, 207, 205, 208, 189, 109, 54, 46, 67, 94, 119, 114, 99, 94, 97, 113, 111, 100, 92, 84, 66, 70, 98, 102, 102, 106, 98, 80, 61, 23, 
    156, 193, 198, 202, 210, 217, 222, 195, 144, 79, 22, 31, 74, 86, 81, 95, 109, 126, 128, 116, 100, 85, 69, 65, 85, 90, 81, 79, 72, 62, 55, 26, 
    154, 198, 208, 218, 229, 229, 210, 205, 209, 166, 85, 73, 112, 115, 96, 101, 118, 137, 141, 128, 107, 88, 75, 68, 73, 84, 73, 68, 68, 72, 75, 44, 
    166, 218, 231, 242, 250, 244, 200, 171, 218, 227, 190, 168, 162, 151, 121, 102, 108, 124, 130, 124, 108, 92, 83, 75, 69, 83, 82, 85, 96, 90, 69, 24, 
    184, 239, 253, 272, 296, 320, 303, 243, 268, 290, 258, 206, 162, 169, 151, 112, 105, 116, 125, 124, 115, 104, 94, 82, 69, 80, 86, 83, 83, 59, 25, 0, 
    218, 289, 322, 359, 395, 423, 427, 342, 276, 271, 267, 245, 156, 160, 155, 115, 105, 113, 123, 125, 122, 117, 105, 89, 72, 75, 77, 56, 40, 19, 5, 0, 
    296, 391, 420, 434, 420, 386, 384, 348, 252, 225, 228, 236, 145, 136, 145, 120, 107, 113, 120, 124, 127, 125, 114, 94, 75, 69, 68, 42, 24, 18, 14, 0, 
    355, 442, 439, 426, 362, 254, 218, 224, 174, 167, 172, 170, 118, 119, 132, 116, 112, 118, 123, 127, 129, 123, 107, 87, 70, 64, 71, 60, 40, 28, 20, 0, 
    358, 428, 424, 409, 329, 178, 118, 119, 101, 110, 114, 98, 85, 94, 95, 86, 102, 116, 119, 120, 120, 110, 94, 81, 70, 62, 75, 84, 64, 38, 25, 0, 
    345, 396, 368, 332, 274, 182, 166, 158, 109, 69, 54, 49, 62, 81, 69, 42, 56, 80, 87, 93, 100, 102, 103, 101, 87, 69, 72, 90, 84, 51, 29, 1, 
    274, 290, 237, 196, 180, 170, 177, 167, 121, 65, 30, 30, 55, 93, 97, 51, 26, 38, 56, 76, 102, 118, 124, 116, 88, 61, 59, 80, 92, 69, 40, 3, 
    156, 155, 145, 145, 148, 143, 130, 127, 127, 113, 77, 55, 68, 99, 107, 77, 58, 66, 79, 100, 128, 138, 132, 126, 109, 74, 56, 61, 80, 86, 61, 10, 
    108, 124, 129, 123, 116, 112, 117, 127, 137, 137, 118, 99, 84, 85, 83, 78, 65, 69, 84, 111, 149, 161, 139, 121, 114, 96, 74, 56, 63, 84, 76, 20, 
    85, 103, 99, 101, 112, 122, 124, 115, 98, 81, 74, 73, 56, 45, 60, 81, 72, 63, 74, 95, 132, 148, 128, 106, 98, 92, 77, 60, 51, 66, 75, 32, 
    69, 90, 101, 110, 114, 107, 90, 68, 47, 36, 50, 76, 69, 53, 60, 71, 62, 52, 56, 58, 72, 90, 95, 93, 88, 79, 64, 48, 42, 48, 59, 33, 
    78, 102, 100, 89, 74, 58, 40, 26, 22, 31, 58, 84, 78, 68, 70, 61, 41, 30, 32, 32, 32, 44, 64, 78, 77, 60, 43, 34, 36, 35, 37, 18, 
    69, 79, 60, 40, 28, 26, 25, 23, 24, 30, 55, 76, 76, 70, 62, 45, 34, 25, 26, 30, 28, 28, 38, 44, 44, 35, 27, 24, 28, 26, 20, 0, 
    31, 25, 13, 9, 17, 25, 28, 26, 22, 24, 48, 65, 67, 68, 50, 35, 33, 24, 27, 33, 27, 22, 25, 24, 24, 26, 22, 16, 16, 17, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 15, 15, 20, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=125
    114, 99, 92, 90, 96, 108, 118, 117, 110, 110, 105, 91, 83, 86, 86, 78, 67, 58, 56, 53, 45, 40, 33, 22, 13, 6, 2, 2, 0, 0, 0, 0, 
    137, 83, 75, 71, 80, 95, 95, 87, 86, 77, 76, 76, 66, 55, 57, 56, 50, 45, 45, 38, 26, 21, 13, 4, 0, 0, 0, 2, 0, 0, 0, 0, 
    135, 79, 74, 65, 77, 88, 61, 61, 83, 63, 60, 75, 74, 54, 42, 41, 40, 40, 42, 32, 19, 17, 15, 11, 10, 13, 20, 27, 28, 26, 30, 0, 
    132, 79, 77, 67, 76, 80, 37, 43, 75, 52, 39, 51, 57, 50, 38, 34, 25, 26, 40, 41, 35, 35, 40, 42, 46, 53, 63, 68, 65, 57, 52, 0, 
    125, 73, 75, 67, 66, 66, 36, 39, 55, 27, 9, 13, 20, 15, 12, 23, 29, 44, 64, 70, 73, 78, 83, 85, 80, 83, 87, 81, 72, 61, 49, 0, 
    116, 64, 67, 65, 52, 32, 21, 37, 37, 3, 0, 0, 1, 0, 2, 12, 29, 67, 104, 106, 101, 102, 106, 97, 83, 82, 83, 74, 61, 47, 35, 0, 
    109, 59, 60, 59, 38, 5, 0, 8, 7, 0, 0, 0, 0, 0, 9, 25, 33, 51, 89, 103, 102, 101, 93, 82, 77, 76, 71, 60, 51, 42, 34, 0, 
    105, 58, 65, 70, 65, 34, 0, 0, 0, 0, 0, 0, 0, 1, 13, 24, 28, 31, 46, 65, 81, 91, 83, 68, 69, 80, 74, 64, 58, 55, 54, 0, 
    123, 86, 103, 119, 139, 102, 9, 0, 0, 0, 22, 39, 40, 41, 24, 19, 22, 19, 26, 38, 50, 64, 67, 62, 74, 90, 87, 79, 74, 73, 73, 0, 
    185, 150, 173, 193, 212, 138, 4, 0, 0, 0, 33, 71, 75, 72, 37, 16, 22, 17, 13, 17, 25, 36, 52, 61, 80, 103, 104, 98, 96, 96, 94, 0, 
    259, 213, 227, 232, 233, 127, 0, 0, 15, 0, 23, 69, 68, 62, 41, 16, 20, 20, 12, 10, 14, 14, 26, 45, 69, 108, 123, 118, 113, 106, 97, 0, 
    298, 228, 227, 221, 216, 131, 0, 0, 40, 25, 43, 79, 62, 40, 28, 16, 27, 33, 18, 16, 18, 7, 8, 34, 62, 96, 125, 125, 115, 104, 91, 0, 
    299, 215, 211, 205, 199, 155, 36, 0, 33, 62, 78, 98, 78, 40, 26, 19, 37, 48, 31, 24, 25, 8, 0, 33, 63, 84, 113, 120, 108, 91, 73, 0, 
    281, 197, 195, 191, 191, 181, 112, 33, 25, 27, 40, 76, 76, 38, 29, 31, 46, 58, 41, 30, 27, 9, 0, 26, 57, 64, 88, 102, 85, 65, 53, 0, 
    261, 181, 186, 192, 202, 199, 172, 128, 93, 22, 0, 42, 60, 24, 20, 42, 62, 72, 55, 39, 24, 7, 0, 11, 43, 44, 52, 68, 64, 58, 55, 0, 
    258, 186, 197, 208, 214, 197, 164, 174, 163, 86, 40, 71, 90, 55, 38, 53, 72, 80, 68, 45, 23, 7, 0, 2, 28, 36, 31, 54, 65, 66, 68, 0, 
    272, 201, 215, 228, 236, 215, 146, 165, 214, 151, 111, 129, 131, 106, 55, 47, 63, 69, 62, 44, 24, 13, 7, 0, 15, 35, 33, 62, 82, 72, 52, 0, 
    294, 228, 247, 271, 294, 294, 221, 189, 250, 233, 192, 133, 124, 138, 74, 46, 53, 62, 59, 47, 34, 24, 14, 0, 5, 31, 33, 49, 64, 43, 21, 0, 
    353, 288, 318, 349, 373, 389, 346, 240, 227, 223, 226, 149, 96, 144, 87, 37, 46, 55, 57, 52, 47, 39, 21, 1, 0, 21, 19, 17, 29, 18, 10, 0, 
    456, 374, 398, 409, 372, 343, 346, 237, 171, 191, 205, 143, 76, 122, 84, 40, 46, 54, 54, 56, 56, 49, 27, 2, 0, 10, 14, 5, 19, 26, 24, 0, 
    528, 419, 420, 395, 270, 182, 208, 157, 103, 135, 143, 100, 48, 83, 72, 46, 57, 59, 55, 60, 62, 46, 20, 0, 0, 7, 32, 30, 30, 36, 32, 0, 
    545, 403, 395, 354, 198, 91, 108, 74, 37, 65, 68, 40, 22, 35, 31, 40, 66, 59, 51, 54, 54, 42, 22, 1, 0, 9, 52, 67, 45, 32, 35, 0, 
    519, 347, 316, 271, 173, 108, 129, 94, 32, 9, 0, 0, 11, 34, 11, 0, 31, 38, 31, 40, 49, 45, 37, 21, 9, 21, 65, 90, 61, 32, 31, 0, 
    406, 243, 204, 169, 136, 122, 139, 113, 52, 0, 0, 0, 29, 68, 36, 2, 9, 10, 11, 32, 56, 64, 62, 45, 13, 14, 55, 91, 82, 46, 29, 0, 
    271, 134, 120, 120, 125, 125, 119, 109, 85, 46, 11, 8, 52, 77, 53, 15, 20, 32, 32, 61, 90, 81, 64, 57, 38, 24, 40, 73, 89, 71, 36, 0, 
    196, 102, 109, 110, 110, 107, 108, 115, 114, 88, 64, 57, 59, 65, 52, 26, 15, 27, 38, 77, 115, 95, 61, 51, 45, 37, 45, 55, 79, 84, 49, 0, 
    157, 94, 94, 97, 104, 108, 106, 96, 80, 67, 68, 55, 30, 24, 43, 39, 16, 17, 28, 62, 103, 87, 47, 32, 35, 32, 35, 48, 63, 78, 62, 0, 
    141, 85, 94, 101, 99, 85, 66, 51, 39, 43, 70, 68, 38, 39, 49, 32, 13, 13, 19, 31, 53, 51, 33, 26, 24, 20, 24, 41, 51, 61, 63, 0, 
    144, 90, 86, 74, 60, 43, 28, 21, 24, 48, 86, 85, 53, 52, 49, 33, 17, 10, 15, 14, 18, 23, 27, 30, 25, 15, 17, 36, 48, 46, 50, 0, 
    126, 63, 49, 36, 31, 28, 23, 24, 30, 54, 88, 82, 63, 52, 39, 33, 27, 23, 28, 21, 13, 20, 26, 25, 23, 15, 15, 32, 43, 37, 32, 0, 
    80, 24, 16, 18, 29, 35, 34, 33, 28, 48, 83, 75, 63, 52, 31, 31, 35, 31, 36, 32, 20, 25, 28, 24, 27, 26, 20, 24, 31, 30, 22, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 17, 14, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=126
    10, 0, 0, 0, 0, 0, 0, 0, 3, 15, 13, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    75, 61, 57, 56, 61, 65, 69, 76, 79, 90, 97, 86, 70, 64, 62, 53, 43, 39, 40, 39, 33, 29, 22, 17, 12, 6, 3, 3, 0, 0, 0, 0, 
    74, 60, 56, 52, 60, 63, 62, 81, 81, 83, 98, 104, 87, 71, 66, 60, 51, 43, 41, 39, 32, 29, 23, 16, 10, 5, 2, 3, 2, 0, 1, 0, 
    74, 59, 56, 50, 58, 63, 47, 65, 87, 90, 99, 117, 119, 99, 83, 72, 54, 45, 41, 37, 28, 26, 22, 19, 18, 18, 19, 22, 23, 23, 23, 0, 
    73, 60, 59, 52, 57, 62, 44, 52, 89, 94, 94, 105, 118, 118, 109, 95, 67, 47, 39, 38, 37, 37, 42, 43, 44, 47, 48, 48, 48, 46, 42, 0, 
    69, 57, 59, 55, 49, 53, 58, 68, 79, 85, 87, 92, 101, 111, 112, 105, 93, 80, 69, 61, 65, 70, 73, 70, 66, 66, 67, 63, 59, 53, 47, 0, 
    66, 53, 55, 52, 40, 31, 44, 72, 80, 83, 88, 94, 98, 102, 109, 112, 110, 117, 118, 99, 90, 89, 88, 86, 74, 66, 64, 58, 52, 47, 41, 0, 
    63, 52, 52, 48, 33, 4, 2, 54, 79, 79, 79, 79, 84, 91, 105, 121, 121, 120, 126, 124, 113, 107, 97, 83, 73, 63, 56, 52, 50, 49, 45, 0, 
    60, 49, 49, 47, 43, 16, 4, 42, 71, 76, 82, 79, 81, 86, 95, 114, 124, 121, 119, 125, 128, 125, 111, 85, 74, 71, 64, 59, 57, 57, 58, 0, 
    63, 57, 65, 76, 91, 63, 33, 47, 67, 76, 104, 108, 107, 105, 98, 107, 121, 124, 122, 123, 128, 133, 129, 108, 89, 84, 77, 74, 73, 74, 76, 0, 
    99, 96, 111, 124, 137, 86, 31, 53, 66, 61, 98, 120, 123, 130, 113, 106, 117, 120, 121, 125, 126, 130, 136, 123, 107, 102, 95, 93, 92, 90, 87, 2, 
    143, 134, 141, 148, 152, 92, 12, 44, 72, 56, 76, 111, 114, 121, 122, 107, 113, 113, 112, 121, 124, 121, 127, 124, 109, 114, 114, 106, 100, 94, 88, 5, 
    160, 146, 146, 147, 147, 106, 18, 18, 80, 88, 92, 118, 118, 106, 117, 110, 114, 113, 107, 113, 121, 119, 118, 124, 111, 110, 119, 111, 102, 92, 83, 5, 
    159, 142, 140, 138, 137, 117, 51, 0, 38, 86, 118, 140, 140, 123, 117, 115, 117, 117, 105, 107, 116, 117, 113, 124, 122, 105, 115, 110, 95, 82, 70, 0, 
    148, 129, 129, 129, 129, 124, 99, 46, 12, 30, 75, 116, 120, 116, 116, 120, 124, 121, 110, 104, 111, 114, 110, 117, 127, 103, 100, 101, 84, 65, 53, 0, 
    139, 122, 123, 127, 133, 133, 133, 131, 80, 26, 12, 64, 93, 92, 109, 127, 138, 136, 123, 112, 110, 111, 110, 110, 121, 104, 84, 82, 68, 58, 56, 0, 
    139, 127, 133, 140, 145, 131, 106, 145, 137, 70, 46, 62, 108, 93, 99, 127, 141, 143, 131, 118, 111, 109, 111, 105, 113, 107, 82, 78, 72, 70, 75, 9, 
    149, 138, 142, 145, 143, 130, 83, 106, 177, 136, 111, 82, 121, 122, 104, 121, 135, 136, 129, 119, 112, 110, 111, 106, 108, 110, 90, 88, 88, 79, 68, 4, 
    153, 138, 145, 157, 172, 189, 155, 111, 180, 193, 163, 102, 112, 151, 121, 119, 130, 131, 127, 121, 117, 116, 112, 107, 105, 108, 90, 79, 75, 60, 49, 0, 
    174, 167, 188, 207, 218, 253, 252, 176, 165, 196, 195, 143, 108, 150, 137, 120, 127, 129, 125, 123, 123, 123, 118, 110, 104, 101, 79, 52, 49, 45, 44, 0, 
    236, 219, 233, 234, 205, 230, 263, 222, 169, 169, 189, 167, 124, 138, 143, 129, 129, 130, 126, 125, 126, 129, 125, 114, 104, 94, 73, 43, 39, 47, 46, 0, 
    273, 241, 243, 234, 168, 138, 166, 159, 145, 150, 164, 155, 131, 121, 125, 136, 137, 136, 131, 130, 131, 128, 120, 105, 93, 84, 83, 62, 41, 48, 49, 0, 
    275, 244, 249, 239, 162, 92, 100, 95, 96, 120, 129, 127, 119, 96, 74, 103, 137, 140, 135, 129, 122, 116, 112, 102, 90, 83, 91, 90, 58, 45, 52, 0, 
    278, 236, 214, 186, 141, 109, 113, 102, 68, 62, 81, 94, 103, 89, 55, 49, 89, 110, 110, 113, 110, 112, 114, 102, 84, 82, 92, 106, 83, 49, 48, 0, 
    217, 169, 143, 124, 117, 114, 109, 99, 71, 40, 33, 57, 88, 106, 83, 48, 63, 87, 95, 106, 110, 110, 114, 110, 84, 69, 86, 102, 104, 70, 46, 0, 
    134, 113, 109, 104, 97, 92, 89, 92, 93, 79, 56, 57, 91, 115, 102, 76, 77, 95, 104, 119, 126, 117, 113, 119, 107, 80, 76, 89, 105, 97, 59, 0, 
    106, 94, 90, 87, 85, 87, 93, 99, 104, 104, 92, 70, 73, 97, 104, 91, 85, 96, 106, 127, 149, 137, 117, 116, 116, 96, 80, 84, 95, 105, 80, 0, 
    87, 76, 77, 85, 95, 99, 99, 95, 87, 83, 87, 75, 60, 73, 88, 92, 87, 91, 97, 111, 140, 140, 118, 105, 103, 93, 83, 83, 85, 94, 92, 3, 
    78, 75, 84, 93, 98, 92, 81, 72, 65, 72, 87, 87, 73, 73, 80, 81, 78, 81, 83, 83, 99, 112, 109, 101, 96, 81, 73, 77, 79, 80, 87, 12, 
    87, 83, 84, 82, 78, 69, 59, 56, 57, 74, 94, 95, 84, 78, 78, 70, 69, 70, 71, 67, 71, 83, 90, 93, 88, 70, 62, 69, 74, 71, 72, 10, 
    80, 71, 62, 59, 58, 60, 60, 57, 56, 71, 92, 92, 90, 77, 68, 68, 69, 68, 71, 68, 62, 66, 68, 71, 72, 65, 59, 62, 68, 64, 58, 2, 
    51, 50, 49, 52, 59, 64, 66, 63, 59, 67, 90, 98, 96, 88, 71, 69, 70, 71, 73, 72, 64, 64, 65, 63, 66, 68, 62, 58, 60, 60, 55, 12, 
    
    -- channel=127
    23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    62, 33, 30, 29, 35, 42, 48, 46, 43, 45, 45, 36, 31, 32, 34, 34, 29, 24, 24, 22, 18, 20, 17, 13, 11, 9, 10, 12, 11, 7, 6, 0, 
    61, 32, 31, 29, 35, 41, 39, 43, 48, 38, 41, 44, 32, 23, 26, 31, 31, 29, 28, 26, 21, 21, 19, 16, 14, 13, 14, 17, 16, 13, 13, 0, 
    60, 31, 31, 27, 33, 38, 28, 36, 51, 35, 30, 44, 45, 30, 20, 22, 26, 31, 32, 28, 21, 23, 24, 22, 20, 20, 22, 24, 27, 26, 27, 4, 
    60, 32, 32, 29, 30, 38, 28, 23, 40, 35, 28, 32, 43, 41, 30, 24, 22, 26, 33, 32, 28, 28, 31, 32, 31, 35, 41, 43, 43, 42, 41, 13, 
    56, 30, 32, 31, 29, 35, 36, 25, 29, 27, 23, 21, 23, 27, 29, 32, 34, 34, 38, 38, 40, 40, 47, 49, 48, 52, 54, 53, 51, 50, 47, 19, 
    53, 27, 29, 31, 26, 22, 30, 40, 28, 13, 16, 19, 19, 23, 29, 30, 34, 44, 57, 55, 51, 53, 56, 57, 57, 58, 56, 53, 51, 48, 46, 17, 
    52, 28, 27, 28, 25, 17, 11, 21, 22, 6, 8, 13, 18, 23, 32, 40, 38, 39, 55, 63, 57, 52, 47, 52, 59, 59, 53, 47, 47, 47, 46, 16, 
    53, 29, 30, 32, 35, 22, 0, 0, 14, 5, 11, 12, 11, 17, 22, 34, 45, 38, 33, 43, 51, 53, 51, 44, 52, 61, 57, 53, 54, 57, 59, 20, 
    63, 38, 40, 45, 50, 35, 5, 5, 15, 8, 24, 32, 28, 26, 20, 22, 35, 38, 32, 30, 39, 47, 50, 46, 48, 64, 70, 69, 69, 68, 69, 26, 
    88, 54, 61, 68, 73, 51, 14, 16, 19, 3, 24, 45, 42, 39, 28, 21, 31, 34, 32, 31, 31, 38, 42, 47, 54, 73, 84, 83, 83, 82, 82, 33, 
    115, 78, 84, 87, 87, 60, 5, 13, 31, 6, 9, 36, 32, 32, 33, 21, 27, 34, 31, 33, 34, 31, 30, 37, 51, 77, 97, 96, 92, 88, 83, 34, 
    128, 89, 90, 88, 87, 72, 13, 2, 40, 35, 20, 32, 30, 14, 22, 22, 27, 34, 30, 32, 38, 31, 23, 34, 44, 66, 97, 101, 92, 84, 77, 33, 
    125, 87, 89, 86, 83, 79, 41, 0, 24, 56, 50, 50, 48, 24, 17, 25, 30, 36, 31, 30, 34, 30, 21, 33, 48, 55, 81, 94, 85, 74, 65, 28, 
    115, 80, 82, 82, 82, 82, 73, 30, 5, 16, 38, 59, 57, 42, 33, 34, 34, 37, 27, 23, 26, 25, 20, 26, 45, 47, 57, 75, 69, 60, 55, 20, 
    107, 72, 76, 82, 84, 82, 82, 84, 51, 5, 5, 40, 49, 35, 35, 41, 42, 37, 29, 22, 20, 22, 20, 19, 34, 39, 34, 51, 60, 57, 56, 17, 
    109, 75, 80, 84, 87, 80, 68, 89, 100, 57, 19, 29, 54, 46, 36, 41, 43, 42, 34, 26, 22, 21, 19, 15, 23, 35, 29, 42, 56, 61, 64, 32, 
    117, 80, 87, 93, 99, 93, 55, 56, 100, 74, 56, 51, 68, 77, 41, 36, 37, 36, 31, 25, 22, 19, 17, 13, 14, 29, 32, 43, 65, 71, 73, 43, 
    129, 91, 99, 107, 113, 114, 87, 38, 84, 109, 87, 65, 56, 91, 59, 33, 34, 29, 27, 24, 23, 21, 16, 12, 10, 22, 30, 42, 70, 81, 75, 33, 
    154, 106, 114, 121, 127, 140, 150, 88, 55, 103, 111, 83, 40, 83, 71, 36, 30, 27, 23, 25, 27, 26, 18, 10, 8, 16, 30, 41, 65, 76, 71, 31, 
    188, 126, 138, 143, 122, 121, 154, 127, 67, 80, 95, 89, 45, 58, 69, 45, 32, 27, 23, 27, 32, 32, 25, 14, 10, 17, 36, 43, 57, 71, 71, 34, 
    213, 149, 151, 143, 94, 63, 94, 99, 69, 59, 62, 65, 48, 45, 58, 55, 46, 35, 29, 33, 38, 36, 30, 19, 13, 24, 49, 59, 56, 66, 72, 35, 
    213, 145, 143, 135, 102, 52, 49, 39, 26, 34, 36, 38, 36, 33, 35, 50, 58, 45, 34, 35, 43, 43, 32, 20, 16, 29, 59, 80, 65, 60, 72, 37, 
    195, 125, 119, 120, 112, 73, 60, 47, 18, 15, 15, 16, 26, 36, 18, 13, 39, 40, 30, 33, 40, 38, 30, 25, 26, 42, 68, 90, 84, 62, 64, 35, 
    155, 108, 96, 81, 75, 71, 69, 70, 49, 12, 0, 6, 26, 38, 34, 15, 14, 19, 15, 22, 33, 33, 32, 32, 27, 40, 67, 90, 98, 76, 58, 27, 
    108, 70, 62, 57, 60, 66, 66, 64, 64, 50, 22, 16, 31, 45, 44, 29, 18, 20, 20, 29, 39, 30, 22, 34, 42, 37, 58, 80, 96, 94, 64, 21, 
    82, 54, 57, 60, 58, 55, 59, 64, 69, 70, 67, 52, 50, 58, 51, 34, 19, 21, 24, 36, 50, 40, 22, 24, 38, 48, 58, 74, 86, 96, 80, 21, 
    75, 55, 55, 56, 57, 59, 62, 66, 70, 73, 80, 71, 46, 43, 50, 46, 35, 29, 29, 35, 53, 51, 31, 23, 29, 41, 58, 78, 85, 89, 90, 31, 
    71, 50, 56, 61, 65, 65, 66, 69, 73, 76, 82, 78, 57, 48, 49, 54, 56, 50, 46, 40, 45, 50, 44, 36, 33, 40, 57, 79, 88, 85, 87, 42, 
    76, 56, 62, 66, 70, 71, 68, 67, 71, 80, 91, 84, 68, 59, 63, 69, 72, 66, 63, 55, 46, 50, 54, 57, 57, 59, 63, 79, 90, 86, 80, 43, 
    75, 64, 67, 70, 74, 75, 73, 70, 71, 78, 92, 90, 78, 68, 69, 77, 81, 79, 75, 68, 60, 61, 66, 71, 77, 77, 74, 79, 86, 83, 74, 38, 
    60, 62, 62, 66, 73, 76, 79, 74, 69, 72, 88, 88, 83, 78, 68, 76, 83, 81, 79, 77, 71, 70, 72, 72, 77, 79, 76, 74, 75, 75, 69, 34, 
    
    -- channel=128
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=129
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 27, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 32, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 7, 0, 0, 4, 5, 5, 4, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 32, 28, 12, 0, 0, 0, 0, 0, 0, 0, 0, 21, 13, 6, 20, 27, 26, 23, 14, 8, 8, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 26, 25, 22, 10, 0, 0, 0, 0, 0, 0, 0, 18, 9, 1, 20, 30, 24, 20, 7, 0, 6, 20, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 13, 19, 18, 14, 6, 0, 0, 0, 0, 0, 0, 14, 9, 4, 21, 28, 20, 8, 0, 0, 0, 18, 
    0, 0, 0, 0, 5, 2, 0, 0, 0, 0, 12, 16, 14, 10, 0, 0, 0, 0, 0, 0, 0, 7, 4, 10, 24, 25, 19, 3, 0, 0, 0, 4, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 1, 16, 17, 14, 5, 0, 0, 0, 0, 0, 0, 0, 5, 0, 8, 24, 26, 19, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 11, 11, 9, 0, 0, 0, 0, 0, 0, 2, 8, 3, 7, 24, 29, 23, 14, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 0, 0, 1, 7, 6, 0, 4, 7, 5, 12, 23, 26, 26, 26, 12, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 4, 3, 6, 8, 0, 0, 8, 15, 1, 3, 12, 6, 3, 13, 19, 20, 23, 29, 23, 9, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 11, 15, 9, 10, 19, 15, 0, 0, 12, 0, 0, 5, 5, 0, 0, 11, 17, 20, 22, 22, 14, 8, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 12, 11, 16, 12, 8, 15, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 15, 18, 12, 6, 10, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 28, 26, 23, 20, 14, 10, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 21, 27, 36, 38, 28, 22, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 2, 0, 0, 0, 0, 3, 8, 6, 4, 13, 23, 30, 36, 32, 24, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 0, 0, 0, 5, 4, 9, 13, 5, 7, 9, 11, 20, 30, 29, 25, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 4, 0, 0, 7, 10, 7, 9, 14, 12, 6, 0, 2, 10, 12, 19, 19, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 8, 0, 0, 4, 16, 15, 10, 13, 18, 11, 0, 0, 1, 3, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 7, 2, 0, 0, 15, 21, 21, 19, 17, 10, 2, 0, 0, 4, 9, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 2, 0, 0, 0, 11, 20, 22, 19, 5, 0, 0, 3, 1, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 0, 0, 8, 20, 20, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 0, 0, 3, 21, 21, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 19, 21, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 19, 23, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 20, 24, 14, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 16, 22, 15, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 15, 9, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=130
    120, 88, 122, 244, 255, 143, 114, 109, 105, 128, 148, 139, 131, 128, 132, 132, 109, 62, 28, 76, 138, 170, 184, 135, 113, 122, 120, 127, 125, 121, 123, 0, 
    127, 93, 115, 262, 352, 247, 190, 182, 164, 168, 205, 230, 215, 201, 205, 211, 195, 134, 47, 38, 148, 264, 266, 199, 194, 205, 206, 213, 212, 206, 207, 0, 
    128, 96, 101, 222, 355, 273, 189, 191, 166, 135, 141, 201, 218, 193, 191, 197, 196, 165, 77, 12, 110, 268, 258, 186, 193, 203, 208, 216, 215, 208, 207, 0, 
    128, 97, 96, 182, 333, 290, 190, 210, 191, 129, 93, 133, 204, 211, 211, 209, 197, 174, 107, 57, 144, 264, 240, 184, 184, 188, 195, 204, 207, 203, 202, 0, 
    130, 96, 93, 146, 293, 303, 199, 215, 222, 153, 80, 68, 141, 196, 231, 241, 216, 179, 136, 111, 178, 249, 231, 214, 203, 188, 190, 191, 184, 184, 182, 0, 
    132, 100, 98, 122, 251, 309, 209, 189, 221, 183, 93, 36, 68, 142, 194, 215, 213, 183, 165, 183, 197, 196, 192, 219, 210, 187, 184, 188, 178, 177, 179, 0, 
    119, 65, 101, 138, 223, 267, 196, 167, 212, 195, 116, 53, 29, 81, 137, 138, 163, 173, 166, 228, 234, 168, 171, 217, 189, 161, 164, 161, 176, 196, 198, 0, 
    175, 0, 47, 147, 223, 222, 162, 148, 220, 221, 145, 99, 60, 62, 90, 86, 111, 148, 152, 220, 250, 176, 180, 239, 195, 158, 166, 151, 178, 233, 226, 0, 
    323, 58, 66, 161, 211, 187, 142, 121, 199, 237, 176, 140, 117, 94, 78, 72, 113, 143, 146, 200, 238, 196, 198, 237, 198, 167, 158, 149, 189, 256, 267, 0, 
    400, 154, 156, 193, 199, 183, 132, 112, 181, 211, 170, 151, 141, 119, 90, 77, 113, 152, 141, 190, 227, 217, 241, 240, 196, 182, 156, 146, 197, 249, 284, 0, 
    419, 178, 178, 205, 210, 186, 128, 126, 194, 188, 148, 145, 133, 111, 96, 100, 133, 137, 127, 178, 208, 207, 267, 266, 208, 191, 170, 151, 196, 242, 273, 0, 
    430, 195, 183, 201, 220, 196, 146, 142, 198, 193, 151, 147, 138, 97, 80, 109, 152, 122, 108, 160, 180, 186, 256, 276, 219, 197, 182, 155, 177, 229, 255, 0, 
    433, 205, 195, 205, 209, 201, 198, 163, 163, 182, 169, 168, 157, 110, 92, 121, 145, 115, 108, 151, 156, 188, 250, 265, 224, 207, 195, 162, 149, 198, 242, 0, 
    436, 205, 199, 208, 184, 168, 244, 202, 122, 125, 125, 153, 149, 89, 97, 176, 167, 106, 126, 160, 140, 177, 253, 258, 224, 215, 212, 182, 139, 173, 238, 0, 
    437, 207, 203, 207, 163, 115, 244, 246, 130, 124, 113, 132, 144, 93, 64, 144, 198, 129, 122, 183, 168, 159, 240, 287, 246, 222, 220, 197, 159, 184, 233, 0, 
    432, 196, 210, 214, 170, 89, 204, 273, 155, 131, 145, 132, 126, 133, 100, 86, 176, 202, 127, 176, 217, 154, 187, 302, 342, 285, 235, 193, 185, 229, 235, 0, 
    434, 173, 193, 221, 198, 109, 141, 247, 186, 118, 128, 122, 95, 121, 132, 70, 118, 252, 170, 144, 225, 159, 98, 180, 328, 360, 293, 223, 223, 273, 250, 0, 
    441, 160, 159, 205, 206, 147, 122, 181, 205, 160, 146, 127, 78, 88, 109, 62, 70, 224, 216, 148, 221, 177, 98, 111, 180, 281, 294, 241, 255, 310, 286, 0, 
    450, 172, 149, 189, 202, 165, 142, 143, 181, 201, 190, 173, 135, 101, 89, 73, 52, 137, 218, 177, 191, 169, 150, 159, 135, 184, 230, 201, 213, 287, 317, 0, 
    455, 188, 161, 188, 210, 172, 164, 162, 153, 178, 187, 177, 183, 166, 115, 101, 80, 64, 155, 193, 158, 143, 176, 193, 156, 167, 189, 165, 171, 216, 268, 20, 
    459, 198, 166, 174, 215, 192, 161, 175, 171, 159, 150, 138, 181, 208, 163, 156, 147, 87, 114, 165, 141, 150, 182, 193, 172, 170, 164, 149, 162, 184, 198, 10, 
    459, 208, 173, 153, 204, 217, 167, 158, 177, 173, 139, 104, 157, 208, 176, 173, 177, 143, 126, 125, 140, 185, 192, 179, 179, 166, 140, 141, 159, 170, 168, 5, 
    453, 213, 190, 144, 187, 235, 190, 157, 159, 162, 141, 113, 141, 183, 169, 161, 163, 151, 127, 106, 149, 210, 195, 170, 183, 166, 129, 138, 146, 141, 150, 0, 
    449, 212, 208, 160, 178, 235, 202, 168, 163, 150, 133, 156, 180, 176, 163, 164, 162, 144, 116, 108, 166, 211, 186, 167, 196, 183, 136, 140, 144, 134, 144, 0, 
    444, 207, 213, 187, 192, 234, 204, 163, 161, 131, 102, 188, 255, 196, 161, 174, 172, 148, 121, 125, 178, 205, 178, 164, 192, 191, 160, 152, 150, 152, 151, 0, 
    441, 203, 210, 203, 216, 247, 219, 161, 147, 99, 41, 163, 278, 209, 162, 180, 176, 154, 136, 141, 183, 203, 171, 168, 176, 172, 176, 180, 167, 151, 140, 0, 
    438, 199, 206, 205, 223, 263, 247, 176, 140, 96, 38, 118, 218, 187, 165, 180, 176, 161, 142, 154, 196, 199, 166, 167, 165, 146, 167, 198, 193, 159, 142, 0, 
    435, 198, 206, 201, 219, 267, 264, 191, 141, 118, 98, 126, 162, 155, 171, 177, 165, 158, 140, 163, 206, 187, 164, 163, 152, 136, 161, 193, 201, 178, 153, 0, 
    428, 202, 219, 201, 203, 267, 277, 199, 146, 134, 141, 146, 140, 144, 171, 174, 156, 144, 141, 179, 204, 179, 175, 167, 144, 136, 162, 186, 191, 181, 160, 0, 
    410, 209, 237, 213, 179, 245, 289, 212, 153, 146, 149, 137, 131, 153, 185, 186, 154, 132, 149, 188, 187, 173, 184, 171, 149, 144, 162, 174, 179, 179, 166, 0, 
    382, 216, 256, 243, 186, 211, 287, 240, 166, 155, 155, 128, 112, 148, 199, 211, 175, 143, 159, 182, 170, 177, 187, 170, 154, 158, 165, 170, 178, 180, 168, 0, 
    354, 264, 296, 300, 266, 249, 304, 316, 278, 263, 249, 211, 176, 180, 206, 232, 223, 207, 221, 224, 218, 232, 244, 233, 227, 224, 215, 225, 243, 252, 241, 107, 
    
    -- channel=131
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 2, 3, 1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 2, 1, 1, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=132
    0, 10, 0, 0, 0, 142, 187, 177, 164, 142, 145, 163, 175, 176, 169, 168, 184, 213, 204, 109, 48, 24, 51, 157, 193, 194, 197, 191, 194, 197, 195, 340, 
    0, 0, 0, 0, 0, 25, 113, 99, 89, 68, 56, 60, 81, 99, 89, 80, 104, 175, 237, 153, 12, 0, 0, 72, 111, 115, 117, 107, 112, 120, 119, 421, 
    0, 0, 0, 0, 0, 0, 104, 75, 61, 83, 68, 39, 44, 82, 85, 70, 69, 115, 216, 227, 52, 0, 0, 84, 102, 104, 103, 97, 103, 114, 116, 431, 
    0, 0, 0, 0, 0, 0, 91, 35, 11, 73, 109, 55, 5, 17, 26, 36, 44, 72, 167, 223, 51, 0, 0, 84, 103, 109, 107, 101, 103, 109, 111, 436, 
    0, 0, 2, 0, 0, 0, 77, 8, 0, 27, 123, 110, 14, 0, 0, 0, 6, 52, 125, 151, 7, 0, 0, 36, 68, 89, 95, 98, 110, 117, 118, 453, 
    0, 0, 0, 0, 0, 0, 69, 41, 0, 0, 108, 165, 97, 17, 0, 0, 0, 18, 58, 50, 0, 0, 0, 6, 33, 66, 68, 74, 93, 98, 105, 468, 
    0, 63, 14, 0, 0, 0, 79, 74, 0, 0, 79, 179, 183, 108, 33, 22, 1, 12, 11, 0, 0, 12, 32, 0, 36, 77, 67, 64, 64, 47, 55, 474, 
    9, 224, 155, 38, 0, 0, 69, 76, 0, 0, 31, 131, 188, 147, 103, 113, 56, 31, 10, 0, 0, 19, 25, 0, 29, 59, 49, 63, 31, 0, 4, 477, 
    0, 252, 191, 25, 0, 0, 105, 118, 0, 0, 0, 53, 106, 125, 129, 133, 69, 12, 10, 0, 0, 12, 8, 0, 26, 53, 66, 98, 35, 0, 0, 463, 
    0, 142, 110, 5, 0, 47, 137, 156, 0, 0, 0, 23, 47, 87, 118, 125, 48, 8, 12, 0, 0, 0, 0, 0, 38, 64, 109, 129, 55, 0, 0, 436, 
    0, 77, 57, 16, 14, 54, 152, 146, 5, 0, 14, 27, 41, 76, 101, 103, 32, 14, 34, 0, 0, 0, 0, 0, 31, 54, 117, 137, 70, 0, 0, 399, 
    0, 60, 55, 16, 1, 49, 144, 111, 0, 0, 11, 14, 40, 93, 127, 86, 20, 42, 65, 0, 0, 0, 0, 0, 17, 47, 100, 143, 95, 28, 0, 383, 
    0, 51, 55, 25, 6, 43, 83, 76, 21, 0, 0, 0, 15, 98, 124, 64, 10, 67, 63, 0, 0, 0, 0, 0, 6, 37, 75, 137, 130, 71, 17, 402, 
    0, 56, 58, 34, 49, 68, 6, 49, 101, 61, 59, 22, 32, 103, 85, 0, 0, 68, 43, 0, 15, 0, 0, 0, 9, 26, 44, 98, 148, 94, 15, 432, 
    0, 57, 56, 35, 105, 137, 0, 5, 123, 111, 92, 29, 27, 100, 99, 0, 0, 61, 46, 0, 12, 0, 0, 0, 0, 19, 21, 57, 127, 72, 1, 456, 
    0, 57, 43, 15, 107, 183, 0, 0, 69, 73, 51, 28, 31, 71, 105, 33, 0, 4, 60, 0, 0, 13, 0, 0, 0, 0, 0, 47, 83, 21, 0, 476, 
    0, 79, 45, 0, 58, 182, 37, 0, 36, 84, 67, 86, 94, 46, 54, 112, 9, 0, 57, 27, 0, 58, 96, 0, 0, 0, 0, 9, 13, 0, 0, 491, 
    0, 115, 86, 15, 22, 136, 98, 0, 5, 62, 57, 86, 133, 93, 62, 165, 102, 0, 19, 63, 0, 60, 185, 114, 0, 0, 0, 0, 0, 0, 0, 479, 
    0, 122, 120, 41, 12, 71, 99, 45, 0, 0, 0, 20, 84, 91, 94, 162, 169, 7, 9, 46, 0, 57, 118, 120, 96, 0, 0, 19, 0, 0, 0, 413, 
    0, 96, 114, 36, 0, 34, 55, 65, 32, 0, 0, 0, 4, 28, 84, 121, 184, 140, 50, 26, 36, 75, 53, 56, 112, 57, 18, 62, 39, 0, 0, 352, 
    0, 66, 98, 41, 0, 16, 37, 53, 61, 45, 41, 40, 0, 0, 37, 42, 87, 162, 79, 34, 76, 82, 35, 43, 75, 50, 42, 75, 65, 27, 0, 314, 
    0, 45, 89, 72, 0, 0, 49, 55, 51, 51, 82, 108, 16, 0, 11, 3, 11, 97, 87, 83, 90, 44, 22, 36, 39, 43, 75, 92, 60, 37, 30, 285, 
    0, 28, 71, 101, 11, 0, 25, 60, 49, 49, 100, 137, 62, 9, 35, 33, 26, 62, 98, 138, 82, 4, 14, 37, 22, 50, 107, 93, 69, 64, 65, 283, 
    0, 21, 46, 108, 30, 0, 0, 37, 41, 54, 83, 83, 31, 27, 53, 48, 48, 64, 120, 147, 59, 0, 17, 40, 0, 32, 96, 82, 86, 91, 81, 292, 
    0, 27, 30, 88, 33, 0, 0, 24, 31, 65, 95, 0, 0, 16, 59, 42, 42, 73, 124, 118, 31, 0, 32, 43, 0, 8, 59, 67, 74, 76, 62, 284, 
    0, 37, 34, 62, 22, 0, 0, 35, 47, 125, 187, 12, 0, 9, 63, 37, 41, 77, 103, 88, 13, 0, 40, 41, 0, 8, 24, 37, 51, 69, 78, 301, 
    0, 44, 46, 56, 16, 0, 0, 30, 66, 170, 255, 81, 0, 35, 61, 37, 48, 67, 82, 68, 0, 0, 45, 33, 28, 43, 22, 3, 23, 66, 91, 321, 
    0, 47, 48, 61, 27, 0, 0, 9, 71, 143, 195, 94, 30, 64, 59, 47, 62, 66, 87, 47, 0, 13, 51, 40, 55, 73, 35, 0, 0, 43, 68, 323, 
    0, 38, 34, 61, 44, 0, 0, 0, 64, 95, 95, 71, 80, 91, 59, 56, 74, 72, 90, 18, 0, 20, 35, 40, 69, 80, 39, 4, 0, 22, 51, 312, 
    0, 23, 2, 55, 72, 0, 0, 0, 46, 70, 63, 77, 97, 71, 24, 32, 65, 90, 75, 0, 2, 23, 19, 35, 74, 76, 41, 16, 9, 19, 51, 311, 
    0, 1, 0, 9, 75, 0, 0, 0, 20, 46, 46, 80, 92, 44, 0, 0, 34, 81, 41, 2, 20, 20, 6, 34, 61, 51, 29, 18, 18, 25, 49, 314, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 127, 
    
    -- channel=133
    3, 0, 9, 86, 141, 131, 120, 115, 107, 108, 118, 124, 120, 117, 119, 124, 116, 86, 47, 42, 63, 116, 147, 134, 135, 137, 137, 137, 135, 132, 131, 12, 
    0, 0, 0, 53, 91, 46, 21, 23, 21, 12, 12, 27, 32, 27, 31, 37, 39, 28, 0, 0, 0, 70, 87, 47, 36, 40, 39, 40, 37, 34, 33, 0, 
    0, 0, 0, 36, 88, 43, 7, 26, 36, 20, 7, 17, 32, 31, 35, 39, 39, 30, 0, 0, 28, 100, 86, 37, 30, 34, 33, 35, 35, 32, 32, 0, 
    0, 0, 0, 19, 77, 43, 0, 35, 57, 38, 9, 6, 17, 27, 41, 46, 39, 20, 0, 0, 45, 116, 83, 40, 33, 31, 30, 31, 30, 29, 28, 0, 
    1, 0, 0, 3, 59, 47, 6, 38, 67, 54, 12, 0, 0, 0, 6, 21, 16, 0, 0, 0, 59, 89, 56, 37, 40, 38, 38, 40, 35, 30, 29, 0, 
    1, 0, 0, 0, 51, 68, 27, 36, 66, 54, 12, 0, 0, 0, 0, 0, 0, 0, 0, 36, 83, 65, 30, 30, 33, 31, 38, 41, 39, 41, 44, 0, 
    22, 0, 0, 23, 92, 92, 33, 31, 67, 56, 16, 0, 0, 0, 9, 0, 0, 0, 2, 55, 85, 50, 33, 61, 53, 40, 43, 28, 23, 39, 48, 0, 
    104, 15, 12, 73, 120, 99, 32, 0, 39, 57, 29, 13, 14, 25, 21, 1, 3, 10, 19, 58, 71, 29, 31, 70, 59, 46, 37, 13, 13, 39, 52, 0, 
    151, 62, 85, 118, 115, 67, 0, 0, 22, 48, 29, 21, 22, 23, 13, 0, 5, 29, 22, 51, 63, 33, 46, 67, 46, 30, 9, 0, 0, 34, 54, 0, 
    151, 28, 52, 85, 72, 31, 0, 0, 39, 58, 30, 18, 15, 2, 0, 0, 0, 12, 12, 40, 55, 41, 62, 75, 48, 32, 10, 0, 6, 34, 48, 0, 
    156, 26, 27, 41, 44, 25, 0, 0, 55, 68, 36, 24, 10, 0, 0, 0, 12, 21, 9, 39, 50, 36, 58, 70, 48, 35, 14, 0, 10, 30, 40, 0, 
    156, 27, 26, 34, 35, 17, 0, 9, 49, 53, 28, 16, 8, 0, 0, 0, 33, 28, 16, 44, 43, 34, 61, 66, 44, 33, 20, 1, 6, 21, 31, 0, 
    156, 22, 18, 27, 20, 0, 14, 26, 21, 11, 0, 8, 10, 0, 0, 35, 52, 25, 25, 38, 30, 38, 69, 69, 46, 38, 34, 21, 10, 20, 44, 0, 
    156, 22, 17, 26, 4, 0, 29, 44, 21, 11, 0, 14, 19, 0, 0, 38, 62, 19, 14, 37, 30, 33, 65, 71, 46, 39, 41, 35, 12, 27, 57, 0, 
    154, 19, 20, 29, 2, 0, 43, 67, 32, 36, 42, 41, 34, 13, 0, 15, 32, 18, 5, 33, 41, 30, 49, 63, 56, 43, 42, 27, 9, 35, 58, 0, 
    153, 8, 10, 26, 11, 0, 46, 82, 35, 17, 24, 27, 9, 4, 18, 11, 19, 33, 9, 19, 38, 14, 0, 4, 46, 61, 46, 13, 5, 41, 55, 0, 
    156, 0, 0, 12, 18, 1, 39, 69, 39, 21, 25, 15, 4, 15, 15, 0, 0, 31, 10, 9, 41, 7, 0, 0, 0, 20, 28, 4, 15, 53, 52, 0, 
    161, 0, 0, 16, 32, 24, 40, 60, 41, 38, 55, 54, 30, 24, 18, 0, 0, 27, 17, 11, 52, 20, 0, 7, 12, 5, 0, 0, 3, 53, 57, 0, 
    165, 8, 5, 35, 50, 39, 40, 43, 29, 26, 38, 39, 34, 38, 22, 0, 0, 13, 22, 29, 39, 0, 0, 18, 27, 41, 32, 1, 0, 20, 34, 0, 
    169, 17, 10, 35, 53, 38, 31, 33, 29, 20, 15, 4, 10, 27, 23, 27, 23, 15, 33, 35, 18, 0, 0, 19, 18, 41, 45, 16, 8, 16, 13, 0, 
    172, 25, 11, 17, 37, 35, 26, 25, 31, 40, 21, 0, 7, 22, 15, 32, 42, 25, 38, 22, 0, 0, 17, 29, 30, 36, 25, 2, 4, 16, 11, 0, 
    169, 28, 14, 3, 28, 45, 36, 33, 33, 38, 22, 0, 10, 29, 17, 20, 20, 5, 6, 0, 0, 15, 36, 35, 34, 29, 6, 0, 4, 5, 0, 0, 
    167, 27, 19, 0, 22, 54, 46, 40, 41, 30, 9, 2, 28, 41, 25, 26, 21, 4, 0, 0, 0, 35, 38, 26, 35, 26, 3, 8, 6, 0, 0, 0, 
    164, 25, 20, 0, 22, 56, 44, 30, 32, 18, 0, 3, 49, 49, 29, 31, 28, 10, 0, 0, 13, 45, 29, 13, 32, 29, 10, 7, 5, 6, 9, 0, 
    162, 21, 17, 3, 22, 54, 43, 22, 16, 0, 0, 0, 54, 42, 19, 21, 18, 0, 0, 0, 21, 39, 16, 8, 21, 15, 1, 3, 6, 4, 8, 0, 
    160, 18, 13, 2, 15, 51, 49, 27, 15, 0, 0, 0, 61, 32, 4, 12, 5, 0, 0, 0, 20, 28, 8, 7, 13, 0, 0, 7, 14, 10, 5, 0, 
    158, 15, 9, 0, 9, 42, 54, 34, 15, 0, 0, 39, 68, 17, 0, 1, 0, 0, 0, 0, 21, 23, 4, 7, 3, 0, 0, 11, 25, 24, 16, 0, 
    153, 11, 9, 0, 4, 43, 60, 36, 13, 0, 11, 53, 52, 7, 0, 1, 0, 0, 0, 0, 26, 19, 7, 9, 2, 0, 5, 27, 31, 22, 14, 0, 
    139, 3, 12, 2, 0, 38, 65, 39, 13, 8, 17, 26, 12, 0, 0, 4, 0, 0, 0, 12, 28, 15, 14, 17, 4, 0, 17, 30, 27, 16, 4, 0, 
    119, 0, 17, 10, 0, 21, 61, 43, 16, 13, 17, 0, 0, 0, 1, 8, 0, 0, 0, 21, 20, 11, 18, 15, 5, 11, 21, 21, 17, 13, 8, 0, 
    99, 0, 16, 14, 0, 6, 52, 45, 17, 10, 3, 0, 0, 0, 0, 0, 0, 0, 10, 20, 13, 14, 24, 14, 7, 8, 11, 13, 16, 19, 15, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=134
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=135
    0, 0, 0, 0, 0, 0, 6, 4, 1, 1, 3, 6, 6, 6, 7, 7, 5, 2, 1, 1, 0, 0, 0, 0, 2, 3, 4, 5, 4, 4, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 10, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=136
    0, 4, 0, 0, 29, 104, 121, 123, 116, 99, 93, 100, 106, 107, 105, 108, 118, 127, 115, 72, 48, 40, 83, 130, 131, 128, 129, 128, 129, 127, 122, 193, 
    0, 4, 0, 0, 0, 74, 110, 110, 111, 101, 80, 78, 91, 95, 94, 100, 117, 141, 159, 118, 32, 12, 69, 118, 126, 119, 120, 118, 117, 116, 110, 216, 
    0, 4, 0, 0, 0, 52, 109, 107, 128, 139, 121, 91, 97, 114, 119, 125, 135, 158, 185, 157, 56, 23, 90, 146, 144, 133, 130, 125, 125, 124, 119, 226, 
    0, 4, 2, 0, 0, 24, 97, 93, 129, 167, 176, 132, 104, 112, 117, 128, 139, 150, 165, 154, 84, 59, 119, 170, 167, 157, 148, 142, 136, 133, 128, 232, 
    0, 5, 6, 0, 0, 0, 81, 84, 114, 175, 211, 182, 113, 90, 85, 99, 122, 133, 136, 133, 103, 103, 142, 175, 180, 180, 170, 164, 163, 157, 152, 254, 
    0, 4, 5, 0, 0, 0, 80, 100, 109, 172, 219, 213, 147, 85, 66, 78, 87, 103, 106, 109, 127, 148, 164, 174, 187, 197, 193, 193, 195, 189, 184, 291, 
    3, 30, 5, 0, 0, 26, 121, 130, 115, 161, 208, 223, 188, 123, 96, 91, 73, 83, 90, 86, 135, 184, 181, 174, 204, 217, 222, 225, 209, 199, 201, 319, 
    36, 114, 62, 32, 65, 103, 148, 150, 110, 135, 193, 218, 212, 176, 141, 125, 99, 86, 95, 81, 117, 185, 182, 180, 220, 234, 236, 231, 197, 181, 199, 330, 
    37, 189, 143, 113, 118, 142, 177, 160, 99, 114, 176, 199, 205, 201, 177, 158, 115, 91, 101, 86, 107, 167, 184, 190, 219, 237, 238, 222, 187, 160, 178, 327, 
    3, 193, 181, 152, 151, 179, 193, 159, 109, 116, 165, 186, 194, 196, 186, 156, 109, 99, 105, 91, 111, 150, 174, 197, 228, 241, 244, 222, 180, 152, 154, 308, 
    0, 187, 181, 165, 174, 190, 194, 159, 124, 139, 177, 188, 194, 186, 169, 136, 111, 106, 116, 99, 116, 143, 151, 194, 238, 243, 247, 233, 182, 155, 147, 274, 
    0, 188, 186, 171, 172, 184, 187, 167, 134, 150, 183, 182, 178, 178, 161, 128, 111, 136, 134, 119, 131, 146, 141, 185, 236, 246, 248, 244, 199, 163, 150, 258, 
    0, 183, 184, 169, 169, 167, 155, 170, 151, 145, 156, 147, 159, 180, 158, 134, 135, 161, 153, 144, 144, 141, 145, 181, 231, 247, 251, 253, 234, 182, 159, 277, 
    0, 182, 180, 165, 171, 147, 106, 157, 173, 160, 156, 151, 169, 188, 163, 120, 140, 172, 166, 147, 156, 153, 147, 182, 227, 242, 246, 258, 260, 207, 181, 305, 
    0, 185, 177, 162, 170, 151, 75, 133, 202, 196, 191, 181, 171, 186, 173, 123, 129, 176, 173, 137, 169, 171, 139, 158, 207, 233, 239, 255, 254, 222, 203, 322, 
    0, 191, 172, 155, 158, 165, 80, 105, 206, 207, 191, 185, 177, 180, 187, 167, 104, 135, 176, 134, 138, 168, 145, 97, 123, 183, 224, 244, 231, 214, 213, 334, 
    2, 202, 165, 138, 136, 161, 120, 103, 190, 213, 197, 211, 208, 178, 179, 186, 112, 81, 157, 135, 103, 165, 156, 84, 55, 103, 166, 199, 191, 182, 211, 342, 
    2, 213, 176, 133, 131, 159, 166, 135, 173, 217, 221, 224, 237, 215, 190, 192, 155, 60, 111, 138, 104, 154, 162, 124, 68, 52, 98, 146, 147, 138, 182, 335, 
    2, 217, 197, 152, 150, 167, 181, 183, 175, 191, 204, 216, 237, 233, 220, 202, 184, 102, 80, 130, 126, 138, 137, 128, 114, 71, 81, 125, 124, 106, 127, 288, 
    3, 217, 213, 173, 162, 180, 186, 194, 190, 179, 187, 197, 197, 213, 223, 209, 210, 182, 108, 135, 145, 127, 106, 101, 118, 111, 110, 130, 119, 92, 92, 226, 
    3, 216, 217, 189, 162, 181, 192, 188, 197, 195, 201, 196, 162, 170, 200, 204, 207, 215, 161, 141, 138, 115, 98, 99, 120, 130, 127, 126, 114, 105, 102, 181, 
    0, 211, 220, 207, 160, 168, 200, 198, 196, 207, 213, 201, 159, 146, 174, 182, 183, 198, 188, 150, 118, 96, 105, 114, 126, 135, 138, 128, 118, 109, 101, 158, 
    0, 206, 214, 218, 168, 157, 198, 214, 206, 210, 212, 204, 172, 152, 172, 176, 176, 182, 183, 148, 103, 88, 110, 125, 121, 141, 152, 134, 125, 107, 92, 158, 
    1, 201, 203, 216, 177, 154, 193, 215, 213, 215, 206, 170, 158, 166, 176, 177, 179, 181, 171, 140, 103, 88, 113, 125, 116, 137, 152, 141, 122, 112, 104, 167, 
    1, 200, 194, 200, 181, 156, 189, 212, 208, 215, 184, 100, 106, 164, 178, 170, 168, 171, 157, 135, 95, 89, 114, 120, 111, 119, 137, 129, 115, 118, 107, 160, 
    2, 199, 190, 185, 171, 150, 182, 213, 209, 210, 170, 71, 68, 151, 172, 153, 151, 150, 143, 119, 85, 90, 113, 112, 108, 106, 105, 101, 112, 112, 106, 170, 
    2, 198, 187, 176, 156, 140, 169, 211, 217, 207, 180, 103, 87, 142, 153, 137, 131, 127, 125, 95, 75, 87, 106, 103, 104, 99, 84, 81, 95, 113, 121, 187, 
    1, 193, 179, 170, 149, 128, 154, 204, 221, 207, 188, 153, 127, 137, 134, 121, 115, 114, 106, 73, 68, 85, 101, 102, 101, 101, 80, 68, 85, 114, 125, 188, 
    0, 178, 162, 165, 148, 118, 140, 194, 219, 209, 187, 169, 152, 142, 116, 111, 111, 103, 84, 63, 67, 83, 92, 99, 105, 98, 78, 78, 91, 104, 114, 181, 
    0, 155, 141, 156, 157, 116, 116, 177, 212, 206, 189, 182, 162, 123, 91, 89, 98, 95, 70, 63, 67, 79, 83, 98, 104, 98, 92, 89, 88, 91, 103, 182, 
    0, 132, 117, 131, 154, 118, 87, 149, 197, 198, 188, 177, 139, 89, 53, 50, 76, 78, 69, 67, 70, 75, 80, 95, 99, 102, 91, 80, 79, 91, 106, 185, 
    0, 39, 27, 32, 49, 40, 11, 36, 70, 71, 64, 60, 47, 17, 0, 0, 4, 14, 12, 5, 13, 12, 11, 19, 25, 21, 16, 15, 16, 19, 24, 63, 
    
    -- channel=137
    93, 98, 79, 69, 104, 127, 130, 138, 138, 121, 113, 115, 119, 118, 120, 129, 145, 155, 143, 117, 111, 129, 156, 163, 147, 142, 141, 140, 139, 133, 129, 147, 
    87, 81, 62, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 64, 65, 36, 29, 43, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    86, 81, 68, 35, 0, 0, 0, 0, 38, 56, 25, 0, 0, 0, 2, 12, 15, 21, 42, 63, 71, 80, 64, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    85, 79, 73, 49, 0, 0, 0, 0, 62, 93, 79, 39, 0, 0, 0, 0, 4, 0, 0, 13, 67, 108, 74, 19, 4, 0, 0, 0, 0, 0, 0, 0, 
    84, 80, 80, 62, 8, 0, 0, 0, 60, 97, 98, 68, 17, 0, 0, 0, 0, 0, 0, 17, 79, 100, 43, 1, 6, 10, 8, 8, 5, 0, 0, 0, 
    80, 73, 76, 69, 30, 0, 0, 27, 69, 90, 93, 75, 44, 6, 0, 0, 0, 0, 0, 32, 105, 110, 46, 15, 19, 29, 32, 36, 35, 32, 34, 30, 
    115, 91, 71, 88, 110, 89, 40, 35, 65, 85, 80, 82, 89, 77, 58, 31, 0, 0, 10, 45, 91, 88, 51, 55, 73, 76, 75, 61, 34, 27, 37, 32, 
    180, 190, 165, 164, 181, 137, 41, 0, 22, 59, 68, 78, 101, 115, 103, 74, 56, 54, 53, 63, 67, 48, 34, 57, 75, 67, 57, 33, 1, 4, 29, 25, 
    133, 149, 179, 188, 165, 84, 10, 0, 18, 49, 57, 61, 69, 86, 85, 60, 56, 62, 61, 65, 61, 42, 43, 68, 61, 45, 30, 0, 0, 0, 12, 13, 
    90, 43, 71, 103, 84, 39, 5, 0, 49, 87, 73, 60, 55, 48, 37, 36, 40, 54, 55, 59, 61, 37, 36, 64, 57, 43, 28, 1, 0, 0, 0, 0, 
    87, 29, 36, 42, 39, 26, 1, 4, 67, 108, 92, 74, 59, 30, 7, 14, 52, 79, 71, 72, 74, 40, 21, 37, 48, 38, 20, 5, 0, 0, 0, 0, 
    79, 17, 25, 26, 18, 3, 0, 16, 59, 74, 65, 53, 44, 34, 30, 46, 86, 106, 96, 95, 89, 54, 34, 39, 42, 37, 26, 19, 10, 1, 0, 0, 
    76, 4, 6, 11, 0, 0, 0, 18, 45, 26, 10, 17, 31, 40, 55, 93, 120, 112, 95, 100, 83, 52, 49, 50, 39, 35, 37, 40, 35, 24, 21, 19, 
    75, 3, 2, 4, 0, 0, 0, 18, 63, 74, 69, 73, 85, 71, 44, 62, 97, 89, 71, 88, 85, 66, 54, 46, 35, 29, 35, 42, 44, 40, 45, 41, 
    73, 0, 2, 5, 0, 0, 0, 27, 63, 98, 114, 110, 93, 83, 87, 73, 61, 59, 60, 62, 75, 69, 27, 3, 8, 24, 31, 27, 22, 33, 56, 33, 
    78, 0, 0, 0, 0, 0, 0, 31, 51, 66, 66, 76, 65, 59, 89, 92, 38, 16, 40, 34, 34, 25, 0, 0, 0, 0, 11, 9, 0, 15, 45, 18, 
    82, 1, 0, 0, 0, 4, 36, 49, 51, 80, 90, 97, 97, 88, 78, 66, 17, 0, 8, 22, 26, 25, 9, 0, 0, 0, 0, 0, 0, 0, 24, 8, 
    84, 12, 7, 9, 16, 28, 64, 73, 51, 68, 104, 125, 126, 125, 106, 68, 34, 8, 0, 7, 33, 25, 9, 25, 16, 0, 0, 0, 0, 0, 0, 0, 
    86, 17, 28, 48, 59, 53, 61, 75, 53, 35, 46, 58, 78, 108, 111, 84, 73, 48, 11, 17, 44, 3, 0, 0, 31, 32, 8, 0, 0, 0, 0, 0, 
    90, 20, 29, 46, 60, 52, 41, 52, 57, 48, 36, 27, 22, 47, 80, 89, 104, 106, 67, 39, 32, 0, 0, 0, 7, 38, 44, 13, 0, 0, 0, 0, 
    92, 24, 31, 35, 40, 43, 44, 38, 49, 72, 67, 39, 15, 19, 35, 53, 72, 81, 72, 39, 0, 0, 0, 12, 22, 38, 28, 0, 0, 0, 0, 0, 
    90, 22, 30, 33, 35, 43, 58, 60, 54, 59, 61, 43, 33, 35, 31, 36, 33, 20, 23, 3, 0, 0, 22, 32, 29, 32, 15, 0, 0, 0, 0, 0, 
    91, 20, 23, 29, 35, 48, 59, 69, 69, 56, 38, 35, 56, 60, 48, 50, 45, 24, 2, 0, 0, 13, 33, 28, 27, 31, 23, 17, 19, 6, 0, 0, 
    92, 17, 12, 17, 34, 55, 55, 53, 52, 39, 3, 0, 26, 54, 45, 41, 42, 26, 0, 0, 1, 30, 23, 9, 13, 23, 18, 14, 13, 12, 20, 32, 
    92, 16, 4, 0, 20, 51, 57, 52, 40, 9, 0, 0, 0, 24, 22, 15, 11, 0, 0, 0, 8, 19, 10, 4, 9, 1, 0, 0, 0, 6, 12, 14, 
    91, 13, 0, 0, 0, 28, 52, 62, 50, 19, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 7, 1, 1, 8, 0, 0, 0, 4, 19, 18, 18, 
    90, 9, 0, 0, 0, 7, 43, 62, 55, 32, 28, 60, 65, 10, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 6, 0, 0, 0, 6, 22, 30, 38, 
    82, 0, 0, 0, 0, 5, 44, 61, 53, 36, 43, 74, 62, 0, 0, 0, 0, 0, 0, 0, 3, 13, 4, 10, 13, 2, 4, 12, 14, 16, 18, 18, 
    67, 0, 0, 0, 0, 0, 46, 60, 50, 41, 38, 37, 14, 0, 0, 0, 0, 0, 0, 0, 16, 7, 3, 15, 16, 11, 18, 26, 21, 7, 0, 1, 
    52, 0, 0, 0, 0, 0, 36, 53, 49, 45, 43, 21, 0, 0, 0, 0, 0, 0, 0, 11, 21, 4, 7, 13, 14, 18, 29, 25, 8, 0, 1, 13, 
    42, 0, 0, 0, 0, 0, 24, 38, 37, 31, 18, 0, 0, 0, 0, 0, 0, 0, 6, 26, 14, 6, 14, 13, 7, 8, 10, 2, 1, 12, 19, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=138
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 21, 42, 25, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 30, 11, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 22, 66, 63, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 30, 20, 14, 9, 0, 0, 0, 0, 0, 35, 
    0, 0, 0, 0, 0, 0, 0, 0, 17, 73, 82, 45, 2, 0, 0, 0, 0, 0, 0, 0, 11, 39, 29, 25, 29, 29, 26, 26, 23, 16, 13, 63, 
    0, 0, 0, 0, 0, 0, 0, 0, 13, 76, 85, 61, 22, 0, 0, 0, 0, 0, 0, 0, 36, 58, 28, 38, 56, 52, 54, 53, 35, 35, 36, 88, 
    11, 0, 0, 0, 0, 1, 4, 0, 0, 67, 83, 66, 41, 15, 3, 0, 0, 0, 0, 0, 44, 62, 28, 47, 74, 71, 71, 62, 35, 32, 47, 102, 
    32, 0, 0, 0, 8, 28, 12, 0, 0, 47, 71, 68, 54, 40, 26, 6, 0, 0, 0, 2, 43, 52, 31, 55, 76, 75, 69, 40, 12, 12, 36, 110, 
    56, 1, 0, 3, 29, 23, 10, 0, 0, 40, 64, 65, 59, 49, 31, 10, 0, 0, 3, 2, 37, 37, 29, 62, 70, 64, 55, 16, 0, 0, 16, 98, 
    63, 14, 8, 13, 24, 24, 10, 0, 0, 45, 62, 61, 61, 44, 24, 1, 0, 13, 5, 5, 38, 32, 25, 61, 67, 62, 48, 11, 0, 0, 0, 75, 
    63, 15, 15, 14, 20, 20, 6, 0, 0, 42, 61, 56, 57, 45, 17, 0, 3, 30, 11, 18, 41, 31, 27, 59, 68, 65, 50, 20, 0, 0, 0, 56, 
    61, 9, 11, 5, 14, 0, 0, 1, 4, 29, 41, 44, 53, 38, 14, 10, 26, 40, 23, 35, 42, 30, 34, 59, 66, 65, 58, 39, 8, 0, 0, 58, 
    60, 2, 5, 0, 10, 0, 0, 19, 16, 32, 32, 30, 49, 46, 13, 7, 53, 52, 23, 41, 49, 29, 30, 60, 60, 61, 62, 58, 36, 0, 3, 73, 
    63, 0, 4, 0, 12, 0, 0, 29, 28, 34, 41, 40, 52, 60, 39, 15, 35, 50, 23, 21, 47, 30, 22, 39, 57, 58, 61, 66, 48, 20, 28, 91, 
    68, 0, 0, 0, 14, 0, 0, 30, 53, 47, 45, 60, 56, 46, 47, 35, 6, 30, 29, 0, 30, 36, 4, 0, 19, 53, 62, 63, 37, 25, 44, 96, 
    71, 5, 0, 0, 9, 5, 0, 21, 63, 67, 57, 64, 53, 48, 52, 44, 0, 0, 25, 0, 12, 32, 0, 0, 0, 1, 39, 42, 16, 21, 44, 93, 
    73, 11, 0, 0, 11, 18, 8, 29, 54, 68, 66, 81, 77, 59, 61, 49, 0, 0, 12, 0, 0, 24, 0, 0, 0, 0, 0, 6, 0, 2, 34, 93, 
    74, 16, 0, 0, 21, 34, 33, 43, 46, 57, 69, 82, 83, 81, 75, 48, 15, 0, 0, 0, 1, 11, 0, 0, 0, 0, 0, 0, 0, 0, 3, 82, 
    78, 21, 6, 0, 30, 46, 40, 44, 47, 48, 57, 68, 65, 79, 80, 58, 44, 6, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 
    80, 27, 22, 9, 26, 49, 47, 38, 40, 46, 53, 48, 36, 60, 65, 53, 58, 39, 3, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 
    82, 31, 32, 17, 16, 46, 54, 44, 42, 46, 54, 40, 14, 38, 50, 46, 57, 46, 18, 7, 0, 0, 0, 0, 0, 8, 4, 0, 0, 0, 0, 6, 
    82, 30, 34, 25, 6, 42, 62, 58, 57, 56, 50, 31, 12, 28, 37, 39, 48, 39, 20, 0, 0, 0, 0, 0, 0, 18, 2, 0, 0, 0, 0, 0, 
    81, 27, 27, 24, 3, 37, 68, 68, 65, 63, 43, 12, 20, 34, 32, 32, 38, 33, 14, 0, 0, 0, 0, 0, 0, 17, 6, 0, 0, 0, 0, 0, 
    80, 23, 18, 13, 0, 30, 68, 72, 65, 63, 22, 0, 14, 39, 27, 22, 27, 22, 3, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 3, 
    79, 19, 10, 0, 0, 16, 61, 71, 62, 57, 7, 0, 0, 31, 16, 9, 13, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    78, 15, 3, 0, 0, 0, 48, 70, 61, 48, 4, 0, 2, 17, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    75, 8, 0, 0, 0, 0, 41, 70, 64, 44, 13, 0, 15, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    66, 0, 0, 0, 0, 0, 37, 72, 66, 46, 27, 19, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    53, 0, 0, 0, 0, 0, 23, 73, 67, 47, 38, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    36, 0, 0, 0, 0, 0, 2, 64, 64, 46, 35, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 4, 14, 7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=139
    53, 73, 76, 88, 166, 282, 309, 293, 285, 282, 282, 289, 298, 299, 296, 294, 298, 293, 263, 207, 164, 172, 235, 315, 331, 325, 328, 329, 329, 326, 320, 311, 
    29, 50, 34, 0, 0, 110, 155, 134, 129, 135, 137, 128, 140, 152, 150, 152, 165, 191, 210, 166, 85, 41, 96, 171, 174, 172, 174, 172, 171, 169, 165, 255, 
    30, 50, 44, 0, 0, 74, 134, 111, 118, 152, 157, 132, 124, 151, 165, 167, 171, 189, 217, 197, 119, 64, 123, 183, 177, 170, 168, 168, 169, 169, 166, 262, 
    31, 50, 49, 0, 0, 46, 117, 91, 97, 158, 187, 160, 122, 118, 131, 146, 155, 155, 170, 182, 134, 99, 155, 195, 194, 188, 182, 177, 174, 169, 165, 262, 
    31, 51, 53, 16, 0, 25, 103, 83, 75, 132, 195, 180, 112, 66, 58, 75, 101, 114, 129, 149, 137, 126, 160, 177, 189, 197, 195, 190, 191, 187, 180, 284, 
    32, 51, 49, 28, 0, 24, 125, 123, 83, 109, 177, 191, 143, 79, 44, 50, 55, 63, 90, 112, 132, 162, 170, 161, 175, 190, 192, 199, 208, 208, 207, 316, 
    62, 112, 64, 41, 33, 114, 198, 167, 91, 90, 154, 195, 194, 158, 114, 94, 67, 61, 78, 86, 115, 180, 186, 163, 185, 207, 204, 212, 205, 189, 200, 328, 
    118, 255, 203, 164, 165, 194, 205, 165, 76, 56, 127, 188, 218, 209, 180, 154, 117, 104, 98, 72, 81, 150, 174, 160, 187, 203, 198, 195, 173, 155, 175, 330, 
    122, 319, 300, 246, 200, 190, 205, 172, 73, 49, 103, 148, 180, 194, 191, 178, 131, 101, 104, 67, 67, 139, 171, 166, 181, 186, 195, 200, 170, 150, 155, 317, 
    38, 253, 248, 204, 188, 201, 221, 191, 101, 81, 108, 129, 146, 162, 164, 142, 106, 92, 98, 72, 73, 137, 162, 177, 205, 217, 236, 243, 206, 165, 152, 300, 
    12, 207, 199, 181, 183, 203, 222, 196, 132, 123, 140, 142, 142, 144, 129, 117, 95, 107, 116, 84, 84, 123, 135, 165, 209, 228, 255, 267, 237, 192, 162, 286, 
    10, 201, 194, 178, 174, 190, 213, 192, 144, 125, 132, 129, 123, 134, 140, 124, 113, 138, 148, 107, 110, 125, 124, 155, 202, 226, 256, 278, 261, 222, 185, 290, 
    10, 200, 193, 175, 169, 173, 168, 168, 150, 105, 85, 74, 99, 146, 154, 137, 143, 167, 158, 127, 123, 119, 122, 159, 199, 222, 247, 280, 286, 256, 218, 323, 
    17, 209, 198, 180, 172, 159, 113, 137, 174, 142, 131, 123, 137, 166, 150, 104, 105, 163, 152, 123, 130, 139, 132, 159, 202, 216, 228, 260, 286, 266, 236, 349, 
    20, 213, 199, 178, 179, 166, 89, 112, 203, 209, 200, 177, 154, 152, 142, 105, 96, 143, 158, 133, 143, 160, 129, 127, 170, 203, 213, 233, 256, 242, 230, 354, 
    21, 216, 190, 155, 163, 168, 87, 79, 164, 190, 162, 137, 138, 146, 159, 143, 104, 99, 153, 138, 108, 132, 112, 58, 46, 115, 179, 210, 222, 210, 222, 356, 
    26, 225, 188, 131, 128, 153, 109, 87, 132, 170, 170, 182, 181, 152, 149, 152, 103, 71, 128, 131, 92, 137, 147, 67, 12, 24, 86, 149, 167, 174, 213, 361, 
    28, 242, 211, 148, 126, 161, 146, 120, 135, 176, 193, 206, 220, 196, 165, 184, 151, 81, 98, 132, 111, 154, 200, 158, 93, 37, 40, 101, 122, 122, 169, 339, 
    26, 255, 243, 192, 155, 164, 164, 152, 147, 138, 137, 158, 184, 189, 191, 206, 193, 134, 106, 120, 127, 144, 157, 165, 156, 105, 91, 125, 122, 91, 99, 265, 
    20, 251, 251, 206, 161, 158, 165, 163, 158, 143, 123, 120, 123, 134, 168, 194, 228, 215, 169, 140, 141, 131, 108, 116, 148, 143, 142, 154, 129, 85, 72, 214, 
    15, 235, 240, 202, 155, 147, 160, 171, 175, 180, 174, 152, 104, 94, 139, 158, 195, 225, 191, 150, 133, 115, 106, 122, 143, 144, 139, 131, 121, 113, 100, 200, 
    6, 219, 233, 213, 156, 139, 169, 183, 185, 189, 191, 183, 133, 105, 125, 123, 131, 170, 166, 149, 120, 102, 118, 135, 132, 129, 137, 134, 126, 122, 103, 176, 
    3, 209, 223, 225, 170, 131, 164, 184, 180, 179, 188, 193, 164, 147, 151, 138, 134, 153, 158, 151, 118, 106, 127, 132, 118, 132, 159, 151, 136, 121, 105, 181, 
    4, 205, 215, 229, 185, 132, 144, 165, 165, 166, 166, 144, 127, 154, 167, 154, 152, 158, 160, 155, 128, 113, 124, 123, 106, 123, 155, 150, 139, 133, 138, 206, 
    7, 208, 210, 225, 191, 145, 138, 151, 150, 150, 123, 48, 42, 127, 163, 145, 139, 143, 152, 148, 120, 104, 119, 117, 95, 103, 121, 122, 128, 137, 133, 191, 
    9, 213, 211, 220, 191, 146, 139, 160, 164, 160, 133, 41, 24, 115, 151, 129, 121, 130, 136, 127, 101, 98, 120, 114, 92, 91, 85, 93, 115, 129, 127, 201, 
    11, 216, 216, 217, 191, 146, 135, 167, 183, 194, 190, 121, 93, 129, 133, 118, 113, 115, 119, 109, 83, 97, 115, 107, 99, 95, 84, 85, 103, 133, 153, 225, 
    11, 210, 209, 217, 199, 144, 125, 161, 186, 202, 208, 169, 135, 131, 121, 110, 113, 114, 113, 95, 81, 104, 116, 113, 116, 118, 99, 85, 101, 128, 142, 216, 
    6, 192, 189, 211, 208, 141, 107, 145, 179, 187, 180, 154, 144, 138, 120, 115, 120, 112, 109, 89, 91, 107, 108, 115, 128, 126, 109, 104, 108, 112, 115, 198, 
    1, 167, 167, 203, 218, 146, 84, 117, 167, 177, 169, 167, 155, 119, 89, 88, 102, 110, 106, 90, 100, 100, 100, 115, 129, 128, 126, 117, 100, 95, 110, 204, 
    5, 151, 141, 178, 206, 145, 65, 84, 144, 162, 159, 150, 122, 77, 41, 41, 71, 100, 103, 101, 104, 99, 100, 113, 124, 125, 114, 94, 90, 105, 129, 213, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 
    
    -- channel=140
    0, 0, 0, 60, 199, 268, 268, 259, 248, 244, 255, 260, 260, 257, 256, 259, 257, 229, 166, 113, 119, 167, 241, 297, 305, 302, 299, 301, 302, 299, 293, 207, 
    0, 0, 0, 19, 163, 239, 234, 221, 213, 207, 211, 221, 232, 231, 228, 233, 246, 242, 187, 99, 71, 131, 243, 291, 284, 282, 277, 276, 275, 270, 263, 188, 
    0, 0, 0, 0, 130, 224, 218, 209, 222, 230, 219, 212, 230, 243, 245, 250, 263, 272, 244, 156, 101, 164, 278, 307, 298, 295, 287, 285, 285, 281, 274, 196, 
    0, 0, 0, 0, 94, 199, 194, 194, 235, 266, 253, 221, 224, 244, 260, 271, 276, 272, 238, 168, 140, 224, 316, 326, 317, 308, 300, 296, 295, 291, 285, 205, 
    0, 0, 0, 0, 57, 167, 176, 181, 237, 289, 291, 234, 193, 183, 199, 230, 249, 245, 215, 178, 182, 261, 320, 330, 335, 332, 325, 321, 316, 306, 298, 214, 
    0, 0, 0, 0, 29, 147, 188, 193, 238, 293, 310, 251, 179, 141, 141, 164, 181, 184, 175, 192, 237, 290, 301, 310, 328, 336, 338, 344, 345, 339, 335, 247, 
    0, 0, 0, 0, 56, 183, 239, 231, 246, 293, 311, 275, 211, 164, 152, 148, 132, 139, 146, 195, 277, 322, 311, 329, 354, 361, 359, 358, 348, 346, 355, 271, 
    109, 89, 38, 67, 170, 277, 286, 229, 219, 275, 306, 303, 276, 236, 209, 176, 139, 146, 154, 196, 274, 312, 305, 343, 386, 389, 380, 358, 324, 326, 354, 280, 
    231, 259, 219, 227, 285, 309, 275, 205, 179, 239, 288, 306, 303, 284, 252, 202, 163, 168, 171, 194, 256, 297, 308, 352, 384, 375, 356, 317, 280, 296, 341, 284, 
    253, 297, 284, 297, 313, 307, 278, 210, 182, 237, 276, 289, 293, 285, 248, 193, 152, 157, 167, 185, 242, 291, 326, 376, 391, 386, 365, 313, 275, 280, 315, 270, 
    260, 303, 290, 296, 311, 315, 282, 218, 215, 268, 288, 292, 289, 264, 214, 169, 150, 170, 170, 185, 238, 274, 315, 376, 399, 398, 378, 326, 286, 277, 292, 244, 
    263, 311, 300, 296, 306, 309, 283, 236, 243, 281, 291, 286, 277, 244, 192, 157, 173, 202, 195, 204, 245, 266, 302, 365, 397, 399, 386, 345, 298, 277, 277, 219, 
    262, 306, 296, 289, 291, 280, 271, 257, 245, 244, 241, 239, 249, 239, 212, 198, 222, 241, 225, 230, 250, 262, 303, 365, 393, 401, 400, 379, 331, 296, 293, 227, 
    267, 307, 296, 288, 281, 242, 237, 272, 259, 231, 211, 217, 248, 244, 207, 216, 256, 257, 229, 242, 247, 256, 305, 366, 389, 397, 406, 406, 370, 327, 328, 263, 
    270, 307, 299, 292, 287, 225, 213, 286, 298, 293, 283, 278, 286, 266, 211, 196, 238, 253, 228, 240, 266, 274, 297, 349, 384, 392, 401, 405, 379, 344, 355, 283, 
    270, 299, 287, 285, 291, 236, 208, 287, 314, 309, 294, 281, 263, 254, 250, 227, 224, 243, 239, 227, 259, 263, 238, 253, 310, 364, 388, 384, 354, 344, 370, 286, 
    275, 294, 261, 253, 274, 257, 220, 273, 312, 310, 291, 289, 271, 256, 261, 237, 182, 204, 237, 210, 232, 246, 200, 140, 163, 254, 325, 336, 315, 336, 374, 287, 
    281, 301, 252, 236, 261, 285, 268, 280, 308, 334, 345, 355, 329, 293, 279, 250, 174, 178, 224, 208, 234, 269, 238, 175, 145, 164, 215, 245, 254, 306, 363, 286, 
    285, 319, 276, 260, 283, 309, 308, 294, 296, 316, 336, 357, 356, 338, 313, 280, 220, 179, 206, 215, 239, 254, 225, 216, 195, 179, 200, 217, 214, 242, 299, 254, 
    289, 333, 303, 286, 303, 317, 317, 310, 296, 290, 294, 302, 311, 325, 325, 306, 287, 240, 226, 238, 250, 226, 193, 207, 207, 207, 234, 238, 213, 204, 221, 187, 
    293, 342, 318, 287, 293, 310, 312, 309, 309, 312, 302, 279, 260, 284, 308, 312, 335, 315, 271, 256, 227, 193, 186, 212, 226, 236, 245, 225, 199, 197, 199, 148, 
    289, 343, 329, 290, 279, 307, 325, 323, 326, 334, 324, 282, 239, 261, 284, 285, 303, 306, 274, 241, 187, 176, 203, 229, 238, 246, 234, 206, 191, 192, 183, 118, 
    284, 338, 333, 297, 270, 304, 341, 348, 347, 341, 326, 293, 261, 274, 288, 284, 286, 285, 260, 211, 162, 180, 221, 232, 237, 250, 237, 214, 199, 178, 155, 95, 
    280, 330, 328, 303, 270, 300, 337, 349, 350, 341, 311, 284, 281, 297, 303, 295, 294, 286, 251, 196, 169, 200, 226, 221, 229, 255, 247, 222, 206, 182, 168, 116, 
    278, 323, 317, 300, 272, 298, 328, 334, 330, 312, 250, 209, 246, 294, 299, 288, 284, 269, 234, 189, 179, 204, 214, 204, 208, 233, 228, 212, 198, 186, 180, 124, 
    276, 319, 306, 287, 266, 288, 322, 332, 322, 290, 200, 140, 212, 279, 281, 267, 256, 239, 208, 178, 172, 193, 201, 192, 193, 195, 185, 188, 191, 190, 175, 112, 
    275, 315, 298, 273, 251, 266, 313, 338, 328, 300, 232, 187, 236, 267, 253, 238, 226, 208, 181, 155, 158, 184, 187, 178, 177, 163, 149, 163, 191, 205, 199, 137, 
    271, 306, 289, 263, 238, 249, 301, 338, 333, 308, 282, 268, 277, 251, 222, 212, 199, 178, 154, 130, 149, 177, 178, 172, 171, 153, 142, 158, 188, 209, 211, 145, 
    257, 286, 275, 257, 227, 229, 288, 332, 332, 309, 297, 286, 266, 223, 203, 200, 186, 161, 133, 120, 154, 172, 174, 179, 175, 154, 149, 165, 190, 203, 196, 130, 
    227, 250, 251, 255, 223, 203, 261, 316, 325, 310, 297, 277, 237, 196, 180, 181, 170, 141, 117, 123, 154, 157, 165, 178, 176, 163, 163, 175, 181, 182, 181, 125, 
    191, 210, 222, 243, 219, 181, 221, 289, 311, 303, 290, 256, 190, 132, 115, 131, 138, 128, 118, 136, 150, 150, 166, 178, 175, 168, 168, 165, 163, 173, 188, 137, 
    84, 90, 97, 113, 107, 74, 91, 140, 160, 156, 142, 113, 63, 26, 14, 25, 41, 46, 51, 66, 63, 66, 79, 87, 82, 78, 69, 62, 72, 93, 103, 72, 
    
    -- channel=141
    0, 0, 7, 140, 252, 245, 218, 210, 204, 210, 221, 224, 220, 215, 215, 221, 211, 163, 92, 75, 112, 197, 267, 265, 261, 260, 256, 258, 257, 253, 249, 41, 
    0, 0, 0, 132, 273, 249, 203, 198, 198, 194, 197, 213, 220, 211, 212, 222, 227, 202, 118, 49, 87, 220, 301, 279, 264, 264, 257, 257, 254, 247, 243, 0, 
    0, 0, 0, 92, 256, 249, 188, 202, 224, 213, 194, 205, 230, 231, 232, 240, 250, 241, 168, 78, 118, 265, 322, 285, 273, 272, 265, 264, 263, 257, 252, 1, 
    0, 0, 0, 55, 220, 238, 171, 209, 261, 256, 210, 195, 218, 237, 255, 265, 264, 246, 176, 98, 161, 307, 337, 298, 286, 279, 274, 272, 271, 266, 261, 5, 
    0, 0, 0, 25, 173, 223, 166, 209, 284, 300, 242, 179, 176, 185, 211, 240, 241, 218, 173, 145, 212, 307, 316, 302, 302, 296, 294, 295, 287, 278, 272, 6, 
    0, 0, 0, 5, 133, 227, 192, 207, 287, 319, 269, 182, 137, 138, 166, 177, 182, 173, 162, 203, 276, 299, 282, 291, 303, 301, 308, 313, 307, 304, 303, 20, 
    32, 0, 0, 33, 170, 255, 217, 212, 286, 326, 288, 216, 154, 143, 155, 140, 138, 145, 159, 243, 318, 303, 283, 327, 340, 332, 333, 318, 305, 316, 326, 27, 
    168, 43, 27, 120, 242, 292, 236, 181, 248, 320, 306, 263, 220, 201, 182, 144, 137, 152, 170, 253, 324, 293, 288, 356, 371, 361, 346, 303, 285, 313, 339, 28, 
    307, 176, 177, 243, 301, 293, 207, 139, 206, 293, 301, 288, 270, 244, 206, 150, 145, 178, 179, 243, 310, 293, 308, 362, 367, 350, 310, 249, 240, 288, 338, 35, 
    367, 228, 235, 285, 304, 270, 194, 139, 209, 285, 290, 285, 277, 247, 195, 142, 147, 167, 172, 226, 289, 298, 333, 374, 365, 346, 294, 230, 222, 263, 316, 26, 
    387, 257, 252, 276, 292, 269, 193, 161, 237, 296, 290, 285, 268, 221, 163, 134, 159, 179, 167, 222, 274, 284, 333, 376, 365, 349, 296, 230, 217, 241, 280, 11, 
    395, 268, 261, 273, 283, 261, 206, 193, 252, 291, 282, 273, 258, 208, 147, 143, 194, 200, 184, 233, 265, 272, 331, 372, 363, 348, 310, 246, 217, 223, 245, 0, 
    393, 262, 251, 260, 258, 228, 229, 228, 229, 238, 229, 244, 248, 201, 175, 203, 242, 219, 212, 241, 251, 273, 336, 374, 364, 353, 336, 290, 237, 225, 254, 0, 
    392, 257, 246, 257, 233, 187, 242, 265, 229, 218, 203, 230, 247, 200, 170, 234, 281, 231, 212, 246, 249, 266, 333, 376, 359, 354, 356, 334, 269, 253, 292, 16, 
    391, 252, 249, 265, 232, 166, 250, 308, 262, 258, 257, 265, 269, 230, 187, 221, 262, 234, 203, 244, 265, 261, 312, 360, 367, 356, 364, 343, 289, 288, 321, 22, 
    389, 237, 236, 262, 249, 177, 250, 337, 293, 268, 267, 266, 246, 231, 228, 214, 234, 250, 207, 223, 265, 240, 215, 259, 332, 368, 364, 321, 284, 308, 333, 15, 
    393, 219, 204, 235, 260, 219, 249, 323, 310, 281, 280, 264, 235, 244, 248, 187, 178, 239, 212, 197, 260, 226, 145, 138, 204, 289, 321, 284, 275, 324, 338, 11, 
    401, 215, 186, 220, 269, 269, 269, 309, 314, 313, 329, 328, 285, 264, 260, 190, 135, 212, 218, 193, 264, 242, 169, 142, 160, 204, 236, 220, 236, 314, 344, 18, 
    410, 233, 201, 237, 287, 301, 296, 291, 292, 306, 329, 339, 320, 308, 277, 224, 163, 182, 213, 220, 253, 221, 185, 181, 167, 198, 226, 201, 201, 253, 303, 20, 
    418, 257, 224, 251, 297, 305, 300, 287, 279, 281, 290, 290, 299, 314, 293, 273, 237, 197, 224, 242, 230, 191, 183, 202, 187, 212, 239, 210, 191, 211, 240, 0, 
    425, 278, 244, 241, 282, 300, 292, 286, 286, 294, 278, 242, 261, 297, 288, 297, 303, 253, 249, 238, 189, 170, 192, 215, 221, 234, 231, 197, 183, 193, 197, 0, 
    427, 290, 259, 227, 264, 309, 306, 301, 305, 308, 281, 226, 232, 277, 278, 283, 293, 264, 237, 194, 152, 180, 213, 229, 239, 242, 210, 181, 179, 177, 163, 0, 
    422, 292, 271, 222, 247, 318, 330, 324, 328, 314, 279, 239, 247, 279, 276, 278, 280, 259, 211, 150, 147, 201, 226, 224, 245, 245, 204, 191, 178, 156, 141, 0, 
    416, 286, 274, 224, 239, 314, 334, 328, 330, 308, 260, 250, 286, 295, 282, 282, 281, 255, 195, 145, 165, 220, 222, 209, 242, 251, 217, 195, 178, 162, 154, 0, 
    411, 275, 264, 227, 236, 303, 326, 317, 312, 264, 183, 217, 298, 298, 273, 272, 267, 233, 183, 149, 179, 219, 205, 194, 222, 230, 206, 190, 181, 166, 160, 0, 
    407, 266, 249, 218, 222, 287, 323, 312, 298, 228, 129, 179, 293, 285, 249, 251, 239, 205, 167, 147, 179, 204, 187, 183, 198, 187, 176, 186, 187, 176, 161, 0, 
    403, 257, 234, 203, 202, 261, 319, 318, 292, 235, 169, 222, 293, 256, 224, 220, 205, 183, 146, 134, 174, 192, 173, 174, 171, 151, 150, 175, 198, 197, 180, 0, 
    395, 246, 226, 191, 181, 243, 316, 323, 290, 255, 238, 271, 280, 228, 199, 197, 180, 155, 118, 127, 172, 180, 168, 168, 158, 133, 142, 180, 205, 204, 190, 0, 
    372, 227, 223, 190, 160, 222, 313, 326, 292, 268, 266, 265, 238, 190, 186, 185, 163, 133, 104, 133, 170, 170, 172, 175, 156, 134, 153, 182, 199, 197, 179, 0, 
    332, 201, 218, 196, 146, 188, 295, 325, 294, 275, 269, 235, 181, 159, 173, 176, 153, 111, 105, 143, 160, 158, 173, 175, 157, 152, 164, 176, 181, 184, 175, 0, 
    283, 168, 200, 195, 137, 150, 264, 315, 290, 270, 252, 196, 129, 102, 119, 145, 133, 109, 122, 144, 148, 154, 177, 172, 161, 156, 158, 162, 171, 182, 182, 0, 
    117, 65, 81, 82, 48, 54, 124, 160, 152, 142, 124, 80, 32, 15, 26, 43, 43, 41, 54, 68, 61, 71, 84, 82, 76, 73, 65, 62, 77, 96, 99, 0, 
    
    -- channel=142
    0, 0, 0, 49, 64, 45, 40, 34, 35, 45, 51, 48, 45, 44, 47, 44, 30, 6, 0, 1, 19, 37, 46, 46, 46, 48, 50, 52, 50, 50, 50, 0, 
    0, 0, 0, 105, 190, 182, 169, 158, 147, 149, 170, 181, 175, 171, 171, 172, 160, 118, 57, 42, 86, 139, 171, 182, 186, 193, 196, 197, 195, 192, 191, 32, 
    0, 0, 0, 78, 188, 191, 171, 159, 142, 130, 136, 169, 174, 166, 167, 172, 171, 149, 91, 37, 64, 143, 186, 191, 196, 204, 205, 205, 203, 198, 197, 31, 
    0, 0, 0, 48, 169, 187, 163, 162, 153, 133, 112, 138, 171, 178, 184, 185, 182, 174, 131, 72, 85, 159, 199, 197, 196, 200, 202, 203, 205, 202, 200, 33, 
    0, 0, 0, 23, 140, 178, 151, 161, 175, 154, 118, 112, 146, 172, 194, 201, 193, 179, 145, 99, 118, 181, 216, 215, 208, 202, 203, 201, 199, 197, 194, 26, 
    0, 0, 0, 6, 107, 163, 138, 147, 181, 177, 141, 100, 100, 126, 151, 172, 182, 163, 145, 130, 140, 177, 203, 213, 211, 206, 205, 205, 202, 199, 195, 15, 
    0, 0, 0, 6, 67, 134, 141, 147, 181, 190, 161, 108, 71, 80, 101, 115, 134, 128, 126, 155, 174, 178, 190, 201, 199, 200, 200, 205, 215, 214, 212, 18, 
    0, 0, 0, 14, 79, 149, 155, 149, 186, 198, 174, 138, 95, 79, 88, 82, 87, 99, 108, 160, 203, 193, 196, 214, 216, 215, 218, 214, 220, 230, 227, 23, 
    103, 32, 21, 72, 144, 177, 155, 132, 165, 193, 185, 170, 146, 120, 104, 86, 93, 98, 108, 154, 199, 200, 200, 226, 236, 230, 224, 211, 209, 233, 244, 29, 
    190, 143, 129, 156, 184, 186, 151, 121, 136, 171, 180, 177, 170, 154, 127, 101, 99, 106, 110, 147, 185, 206, 221, 233, 237, 235, 214, 194, 195, 219, 251, 41, 
    211, 180, 177, 192, 201, 192, 152, 125, 140, 160, 166, 171, 168, 157, 132, 105, 97, 99, 103, 136, 170, 202, 241, 249, 244, 242, 219, 189, 193, 207, 238, 49, 
    221, 195, 186, 199, 212, 200, 158, 134, 161, 177, 171, 175, 167, 138, 109, 97, 103, 94, 100, 126, 158, 187, 232, 255, 252, 245, 225, 192, 187, 200, 218, 36, 
    226, 205, 195, 201, 205, 203, 180, 147, 164, 182, 180, 177, 161, 130, 104, 97, 112, 112, 111, 129, 155, 182, 220, 251, 254, 247, 231, 201, 178, 190, 202, 14, 
    226, 205, 194, 199, 185, 182, 200, 167, 147, 140, 138, 145, 143, 122, 116, 140, 140, 128, 132, 143, 143, 173, 224, 248, 253, 251, 245, 221, 186, 189, 203, 13, 
    228, 206, 193, 196, 169, 143, 199, 193, 152, 135, 124, 139, 154, 123, 97, 138, 171, 140, 135, 158, 148, 168, 226, 263, 258, 253, 254, 242, 214, 202, 218, 23, 
    226, 201, 197, 198, 170, 119, 185, 220, 177, 166, 166, 156, 155, 143, 107, 110, 178, 170, 130, 165, 182, 167, 202, 274, 291, 270, 259, 246, 231, 228, 232, 26, 
    226, 188, 189, 195, 179, 126, 154, 222, 196, 165, 162, 147, 135, 144, 139, 111, 145, 192, 143, 152, 186, 154, 138, 182, 258, 288, 275, 248, 236, 247, 243, 25, 
    231, 177, 163, 174, 175, 149, 147, 198, 209, 179, 172, 162, 133, 133, 142, 109, 100, 177, 163, 141, 176, 161, 118, 98, 148, 225, 246, 226, 231, 260, 259, 31, 
    237, 181, 150, 161, 172, 174, 171, 179, 204, 210, 211, 205, 177, 153, 142, 120, 83, 129, 166, 144, 168, 172, 149, 121, 109, 147, 177, 175, 193, 243, 273, 52, 
    241, 194, 163, 172, 188, 186, 193, 189, 183, 196, 208, 211, 213, 192, 163, 143, 102, 92, 143, 154, 162, 158, 157, 151, 128, 130, 151, 153, 160, 189, 231, 60, 
    244, 206, 178, 179, 200, 193, 191, 197, 182, 177, 180, 181, 203, 207, 187, 179, 162, 123, 136, 163, 159, 143, 143, 151, 144, 147, 158, 153, 147, 150, 171, 41, 
    246, 215, 188, 172, 195, 200, 186, 188, 194, 193, 177, 154, 172, 194, 187, 195, 199, 172, 155, 154, 147, 139, 140, 150, 158, 158, 150, 142, 137, 143, 147, 24, 
    243, 221, 201, 166, 184, 207, 199, 191, 198, 202, 184, 151, 156, 176, 176, 183, 186, 179, 159, 138, 130, 143, 149, 153, 165, 156, 141, 134, 129, 130, 124, 5, 
    240, 221, 213, 173, 175, 207, 210, 206, 206, 200, 186, 182, 177, 177, 179, 182, 181, 171, 151, 123, 125, 149, 155, 155, 169, 165, 146, 137, 133, 115, 107, 0, 
    236, 216, 215, 188, 179, 206, 209, 205, 209, 189, 172, 198, 209, 193, 186, 190, 189, 174, 145, 121, 136, 154, 152, 148, 165, 173, 158, 145, 134, 122, 119, 9, 
    234, 212, 210, 195, 191, 210, 207, 196, 196, 160, 116, 157, 210, 201, 187, 191, 186, 168, 142, 127, 140, 151, 145, 143, 149, 159, 158, 148, 134, 126, 118, 2, 
    232, 209, 203, 193, 192, 210, 213, 199, 188, 145, 83, 112, 183, 197, 181, 179, 175, 158, 134, 129, 137, 145, 138, 136, 135, 131, 134, 144, 143, 128, 116, 0, 
    231, 206, 198, 185, 183, 202, 214, 206, 188, 156, 119, 133, 177, 180, 169, 163, 155, 143, 123, 121, 130, 138, 130, 127, 122, 110, 116, 134, 145, 141, 133, 9, 
    228, 204, 198, 178, 171, 194, 214, 208, 189, 170, 163, 170, 172, 160, 155, 149, 139, 126, 111, 112, 127, 133, 130, 125, 115, 106, 110, 125, 143, 150, 140, 13, 
    218, 197, 196, 178, 154, 179, 214, 207, 189, 179, 174, 167, 160, 153, 152, 148, 130, 110, 101, 108, 123, 126, 130, 127, 118, 106, 111, 127, 141, 144, 133, 5, 
    196, 183, 194, 189, 149, 154, 206, 209, 191, 185, 179, 161, 141, 135, 144, 146, 125, 102, 95, 109, 116, 120, 128, 128, 121, 116, 124, 130, 132, 131, 128, 5, 
    190, 183, 200, 209, 178, 156, 205, 243, 238, 230, 217, 181, 135, 112, 118, 134, 132, 119, 124, 133, 134, 142, 156, 157, 152, 149, 145, 144, 153, 165, 168, 65, 
    
    -- channel=143
    5, 0, 7, 49, 54, 25, 17, 18, 16, 19, 23, 23, 22, 22, 22, 20, 14, 2, 0, 6, 15, 24, 37, 22, 18, 25, 23, 23, 23, 23, 24, 0, 
    13, 10, 20, 86, 161, 148, 129, 126, 122, 120, 131, 139, 136, 131, 132, 134, 124, 100, 61, 42, 72, 113, 137, 138, 143, 149, 146, 145, 146, 147, 148, 62, 
    14, 10, 15, 66, 153, 158, 130, 127, 121, 103, 104, 126, 133, 127, 124, 122, 123, 116, 76, 28, 51, 114, 145, 140, 146, 151, 150, 148, 148, 149, 148, 63, 
    15, 11, 12, 47, 134, 156, 125, 128, 124, 105, 84, 100, 127, 128, 124, 121, 121, 124, 105, 66, 65, 113, 140, 134, 139, 145, 147, 149, 151, 151, 152, 63, 
    16, 11, 12, 32, 109, 150, 121, 127, 137, 120, 91, 76, 103, 128, 139, 142, 135, 130, 113, 86, 86, 118, 136, 136, 135, 135, 138, 141, 144, 146, 147, 60, 
    19, 13, 12, 23, 84, 139, 118, 112, 140, 138, 105, 72, 75, 98, 121, 138, 136, 128, 117, 101, 94, 109, 122, 136, 140, 135, 136, 138, 133, 133, 133, 42, 
    18, 9, 13, 22, 69, 125, 111, 96, 127, 142, 120, 84, 61, 73, 88, 95, 108, 110, 103, 118, 118, 107, 105, 126, 135, 131, 131, 131, 128, 130, 133, 39, 
    26, 0, 2, 37, 71, 95, 95, 93, 122, 144, 131, 107, 75, 63, 71, 69, 76, 90, 88, 115, 140, 123, 114, 139, 142, 135, 132, 121, 124, 136, 138, 45, 
    98, 8, 4, 40, 75, 100, 98, 82, 110, 148, 137, 122, 108, 87, 77, 73, 68, 82, 85, 106, 140, 132, 119, 140, 151, 142, 135, 122, 119, 137, 144, 48, 
    152, 88, 69, 75, 101, 110, 96, 74, 93, 129, 132, 127, 124, 113, 94, 75, 80, 90, 87, 104, 130, 135, 126, 135, 144, 139, 121, 104, 102, 119, 144, 54, 
    163, 107, 104, 112, 117, 111, 94, 82, 95, 114, 120, 121, 120, 113, 98, 85, 77, 84, 82, 99, 122, 130, 141, 148, 141, 136, 119, 94, 91, 102, 125, 54, 
    168, 113, 107, 115, 123, 115, 99, 88, 107, 119, 117, 118, 115, 103, 89, 84, 86, 81, 75, 93, 114, 118, 138, 154, 144, 134, 122, 95, 84, 93, 105, 45, 
    167, 117, 112, 114, 122, 120, 114, 98, 104, 123, 121, 119, 124, 104, 81, 79, 91, 83, 77, 92, 106, 117, 133, 148, 143, 135, 126, 104, 82, 85, 97, 29, 
    166, 111, 111, 116, 114, 113, 137, 121, 91, 98, 106, 115, 115, 99, 92, 99, 99, 90, 85, 93, 100, 117, 134, 145, 142, 139, 136, 123, 92, 85, 103, 20, 
    168, 109, 109, 117, 116, 104, 143, 151, 104, 90, 85, 92, 102, 87, 75, 110, 127, 97, 84, 104, 103, 101, 134, 153, 147, 141, 143, 138, 111, 98, 110, 27, 
    166, 107, 111, 121, 129, 106, 136, 169, 122, 109, 104, 97, 109, 109, 83, 79, 120, 117, 84, 104, 119, 105, 122, 163, 170, 155, 145, 136, 125, 116, 117, 31, 
    165, 95, 103, 121, 140, 119, 125, 169, 136, 106, 113, 110, 93, 104, 110, 79, 98, 140, 105, 90, 130, 113, 83, 121, 179, 184, 159, 135, 125, 131, 127, 32, 
    167, 87, 84, 109, 139, 140, 117, 142, 145, 120, 110, 105, 90, 91, 104, 91, 72, 124, 128, 94, 125, 119, 80, 63, 98, 152, 162, 144, 132, 144, 142, 37, 
    170, 92, 75, 95, 124, 138, 129, 121, 133, 136, 135, 135, 114, 97, 100, 92, 63, 91, 131, 109, 118, 125, 112, 95, 71, 94, 128, 122, 120, 147, 161, 56, 
    171, 101, 83, 93, 118, 129, 135, 120, 110, 126, 137, 142, 143, 129, 110, 103, 82, 63, 109, 120, 108, 114, 118, 123, 104, 99, 113, 109, 100, 118, 151, 76, 
    174, 107, 93, 94, 120, 127, 125, 130, 116, 110, 114, 115, 130, 143, 131, 123, 115, 80, 88, 114, 109, 108, 115, 123, 117, 111, 114, 112, 108, 110, 115, 63, 
    177, 114, 100, 87, 112, 133, 122, 123, 130, 121, 106, 97, 110, 131, 132, 133, 139, 124, 102, 106, 106, 112, 111, 116, 117, 116, 113, 110, 108, 108, 101, 48, 
    175, 118, 108, 86, 101, 136, 135, 124, 129, 130, 122, 103, 100, 120, 123, 124, 130, 129, 115, 99, 100, 113, 112, 110, 118, 121, 107, 102, 99, 96, 98, 44, 
    172, 116, 114, 90, 92, 132, 143, 138, 135, 130, 130, 125, 119, 119, 120, 124, 124, 119, 109, 96, 95, 109, 112, 111, 123, 124, 108, 102, 97, 91, 91, 31, 
    171, 112, 112, 98, 90, 122, 138, 137, 138, 131, 123, 145, 158, 135, 123, 129, 131, 120, 109, 96, 97, 111, 111, 108, 121, 130, 117, 105, 105, 98, 90, 34, 
    169, 109, 106, 100, 93, 116, 134, 129, 128, 115, 104, 138, 174, 148, 124, 129, 131, 122, 110, 96, 102, 113, 108, 105, 110, 120, 117, 114, 105, 97, 93, 40, 
    168, 106, 102, 93, 92, 113, 134, 129, 120, 109, 89, 110, 154, 142, 123, 127, 126, 117, 105, 96, 103, 111, 103, 103, 103, 100, 107, 115, 110, 102, 94, 29, 
    168, 106, 100, 90, 84, 104, 134, 132, 119, 117, 108, 110, 127, 128, 121, 120, 119, 111, 95, 92, 104, 105, 100, 97, 97, 91, 92, 104, 116, 110, 100, 35, 
    165, 106, 103, 89, 78, 97, 131, 133, 121, 118, 121, 120, 124, 117, 116, 117, 109, 98, 88, 89, 100, 100, 100, 96, 92, 84, 89, 100, 109, 110, 104, 42, 
    157, 104, 107, 92, 69, 87, 130, 135, 122, 116, 116, 118, 113, 108, 113, 114, 104, 90, 85, 87, 95, 96, 103, 101, 92, 86, 90, 96, 102, 108, 105, 40, 
    142, 96, 104, 98, 66, 69, 125, 141, 125, 120, 118, 105, 95, 103, 113, 118, 104, 85, 83, 85, 89, 93, 101, 99, 96, 93, 90, 94, 101, 106, 104, 36, 
    125, 95, 106, 111, 90, 73, 116, 150, 142, 133, 128, 113, 94, 86, 96, 109, 104, 94, 87, 90, 92, 99, 105, 106, 103, 99, 99, 105, 108, 110, 108, 51, 
    
    -- channel=144
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=145
    0, 42, 38, 28, 30, 42, 36, 22, 16, 20, 23, 29, 35, 37, 41, 38, 36, 36, 40, 47, 45, 36, 35, 40, 45, 43, 29, 21, 24, 23, 17, 15, 
    0, 40, 39, 38, 39, 40, 35, 15, 4, 5, 18, 25, 22, 30, 36, 40, 44, 45, 43, 39, 33, 28, 26, 27, 36, 41, 35, 24, 18, 19, 18, 23, 
    3, 52, 51, 49, 48, 50, 41, 23, 16, 13, 20, 25, 22, 20, 20, 28, 35, 35, 42, 37, 19, 16, 21, 25, 31, 33, 35, 23, 11, 11, 23, 30, 
    4, 54, 54, 54, 53, 50, 34, 15, 13, 27, 26, 28, 38, 23, 21, 26, 17, 21, 29, 27, 16, 5, 15, 30, 30, 29, 31, 16, 0, 0, 19, 32, 
    5, 54, 54, 54, 54, 55, 49, 14, 5, 38, 47, 52, 59, 53, 54, 50, 36, 39, 32, 22, 20, 17, 17, 33, 36, 26, 21, 9, 0, 0, 9, 29, 
    5, 54, 54, 54, 50, 49, 53, 35, 27, 54, 74, 80, 75, 78, 87, 84, 79, 73, 68, 58, 37, 24, 24, 33, 38, 30, 17, 4, 0, 0, 0, 24, 
    5, 54, 54, 52, 48, 43, 40, 42, 49, 67, 84, 90, 84, 78, 85, 92, 93, 90, 85, 88, 77, 42, 17, 25, 32, 33, 25, 14, 3, 0, 0, 17, 
    5, 54, 53, 54, 53, 43, 36, 47, 46, 46, 57, 71, 75, 77, 85, 88, 90, 90, 85, 82, 85, 78, 37, 15, 27, 34, 29, 21, 4, 0, 0, 8, 
    4, 53, 53, 54, 48, 33, 39, 53, 45, 55, 66, 64, 65, 76, 82, 86, 87, 87, 84, 84, 87, 82, 61, 39, 37, 38, 41, 41, 26, 12, 11, 22, 
    1, 51, 53, 53, 39, 28, 41, 48, 44, 57, 71, 64, 65, 70, 75, 80, 80, 77, 77, 80, 83, 87, 73, 47, 40, 48, 54, 55, 49, 39, 40, 49, 
    0, 45, 51, 52, 52, 47, 39, 45, 32, 32, 51, 58, 61, 61, 65, 70, 70, 66, 66, 65, 69, 76, 72, 53, 43, 49, 53, 53, 50, 52, 54, 60, 
    0, 35, 44, 45, 43, 35, 43, 54, 33, 16, 29, 53, 67, 65, 57, 55, 56, 55, 57, 61, 56, 48, 49, 47, 41, 42, 51, 55, 54, 54, 54, 60, 
    0, 26, 32, 34, 23, 10, 26, 48, 46, 38, 48, 57, 72, 87, 73, 56, 55, 60, 66, 76, 68, 40, 23, 16, 14, 22, 30, 41, 52, 54, 54, 59, 
    0, 29, 26, 22, 12, 3, 17, 22, 21, 55, 76, 65, 57, 69, 70, 53, 45, 46, 50, 58, 54, 31, 17, 14, 18, 21, 19, 21, 39, 55, 54, 59, 
    0, 25, 15, 0, 0, 5, 22, 14, 15, 51, 57, 34, 21, 23, 26, 24, 24, 26, 27, 24, 15, 10, 12, 13, 11, 13, 23, 28, 35, 51, 55, 60, 
    0, 11, 9, 0, 0, 0, 3, 15, 28, 46, 54, 39, 27, 20, 18, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 37, 41, 48, 54, 60, 
    0, 19, 17, 8, 0, 0, 0, 0, 13, 39, 31, 29, 42, 46, 46, 37, 19, 9, 9, 8, 24, 33, 15, 1, 0, 4, 40, 54, 43, 44, 52, 60, 
    0, 25, 24, 10, 0, 0, 0, 0, 0, 23, 21, 0, 14, 33, 38, 42, 39, 34, 37, 36, 42, 57, 49, 38, 35, 42, 45, 37, 31, 37, 48, 60, 
    0, 36, 31, 5, 0, 0, 4, 0, 0, 2, 21, 6, 0, 0, 6, 21, 24, 28, 26, 24, 35, 34, 23, 27, 33, 45, 41, 22, 16, 26, 44, 60, 
    0, 39, 35, 9, 0, 0, 0, 0, 0, 0, 6, 11, 6, 0, 0, 0, 17, 47, 39, 28, 34, 37, 31, 31, 25, 29, 42, 26, 9, 20, 44, 60, 
    0, 36, 40, 25, 0, 0, 0, 0, 0, 0, 0, 0, 7, 12, 15, 1, 0, 7, 21, 20, 21, 19, 18, 23, 17, 15, 24, 32, 29, 23, 40, 59, 
    0, 35, 39, 21, 7, 0, 0, 0, 0, 0, 0, 0, 0, 22, 36, 12, 0, 5, 24, 21, 19, 23, 23, 37, 36, 1, 0, 24, 35, 25, 33, 58, 
    0, 45, 45, 14, 0, 0, 8, 8, 10, 0, 0, 0, 0, 0, 8, 11, 0, 0, 14, 27, 22, 29, 26, 26, 34, 9, 0, 0, 14, 10, 30, 63, 
    0, 55, 54, 21, 0, 0, 5, 27, 26, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 10, 25, 23, 8, 14, 0, 0, 0, 0, 0, 31, 71, 
    3, 60, 69, 49, 8, 0, 0, 27, 35, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 44, 48, 46, 43, 15, 0, 0, 0, 0, 0, 37, 78, 
    1, 57, 68, 64, 45, 27, 22, 29, 25, 15, 6, 0, 0, 0, 0, 0, 0, 0, 0, 9, 40, 48, 47, 46, 22, 0, 0, 0, 0, 13, 47, 80, 
    4, 53, 51, 52, 55, 47, 32, 26, 18, 14, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 28, 33, 39, 10, 0, 0, 0, 0, 20, 48, 81, 
    6, 54, 54, 56, 51, 42, 22, 17, 14, 10, 12, 0, 0, 0, 0, 0, 0, 0, 0, 4, 10, 19, 34, 45, 8, 0, 0, 0, 0, 19, 48, 82, 
    1, 58, 62, 58, 51, 42, 23, 11, 6, 7, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 20, 37, 13, 0, 0, 0, 0, 15, 51, 83, 
    4, 60, 60, 61, 59, 53, 34, 9, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 15, 4, 0, 0, 0, 0, 22, 61, 88, 
    10, 68, 71, 68, 62, 62, 51, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 9, 12, 14, 14, 14, 10, 0, 0, 0, 13, 38, 73, 85, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=146
    335, 59, 59, 76, 87, 51, 28, 54, 81, 55, 49, 57, 55, 50, 42, 68, 87, 92, 85, 62, 56, 75, 88, 72, 41, 28, 66, 104, 70, 51, 80, 0, 
    434, 147, 146, 150, 158, 128, 74, 109, 177, 157, 128, 137, 152, 156, 157, 157, 169, 170, 169, 171, 165, 168, 188, 190, 155, 129, 142, 172, 168, 147, 168, 0, 
    449, 146, 146, 147, 151, 124, 42, 63, 150, 143, 137, 139, 136, 173, 195, 184, 200, 189, 176, 191, 194, 189, 197, 203, 182, 161, 152, 165, 193, 188, 166, 0, 
    462, 147, 149, 150, 151, 122, 29, 33, 127, 105, 104, 118, 78, 122, 150, 147, 194, 192, 184, 225, 212, 208, 217, 195, 179, 181, 159, 164, 220, 241, 184, 0, 
    465, 148, 149, 151, 145, 108, 0, 0, 78, 62, 37, 45, 9, 26, 35, 30, 81, 101, 114, 195, 246, 228, 219, 184, 155, 175, 167, 163, 231, 276, 233, 0, 
    464, 148, 150, 149, 135, 113, 7, 0, 6, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 175, 263, 229, 176, 140, 142, 155, 156, 204, 280, 282, 0, 
    464, 148, 152, 141, 113, 122, 53, 0, 0, 77, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 175, 268, 220, 153, 129, 137, 142, 149, 229, 296, 0, 
    463, 148, 153, 132, 88, 114, 53, 0, 17, 122, 80, 88, 20, 0, 0, 0, 0, 0, 0, 8, 8, 34, 198, 252, 180, 148, 143, 125, 129, 175, 263, 0, 
    464, 150, 153, 129, 82, 99, 43, 0, 28, 87, 32, 93, 77, 0, 0, 0, 0, 13, 0, 12, 29, 0, 105, 216, 177, 156, 145, 97, 97, 142, 187, 0, 
    465, 156, 154, 124, 56, 68, 37, 0, 37, 72, 0, 24, 46, 3, 0, 0, 4, 14, 5, 17, 44, 1, 53, 185, 201, 173, 146, 99, 82, 117, 138, 0, 
    465, 174, 161, 119, 23, 5, 0, 0, 27, 96, 37, 7, 10, 9, 1, 0, 6, 10, 14, 32, 54, 35, 35, 132, 218, 211, 167, 133, 131, 135, 140, 0, 
    446, 193, 168, 114, 56, 46, 0, 0, 0, 82, 73, 16, 0, 0, 0, 3, 6, 9, 19, 23, 29, 61, 66, 104, 198, 224, 176, 146, 149, 149, 149, 0, 
    414, 189, 161, 105, 85, 116, 26, 0, 0, 17, 29, 9, 0, 0, 0, 0, 0, 0, 7, 0, 0, 30, 91, 133, 205, 230, 209, 190, 170, 152, 149, 0, 
    390, 151, 122, 90, 86, 111, 77, 3, 0, 0, 0, 0, 10, 0, 0, 0, 14, 27, 40, 30, 0, 33, 93, 137, 181, 198, 196, 226, 235, 177, 149, 0, 
    392, 123, 65, 83, 132, 128, 96, 20, 0, 0, 0, 3, 45, 43, 15, 17, 33, 39, 39, 39, 37, 58, 78, 98, 128, 148, 144, 174, 265, 231, 156, 0, 
    398, 129, 26, 42, 160, 200, 146, 21, 0, 1, 0, 0, 0, 7, 16, 5, 31, 64, 59, 64, 53, 43, 73, 90, 110, 122, 92, 89, 210, 257, 175, 0, 
    366, 100, 4, 0, 134, 193, 127, 44, 34, 35, 21, 32, 0, 0, 0, 0, 0, 29, 13, 39, 33, 0, 0, 29, 48, 90, 55, 28, 125, 234, 199, 0, 
    365, 82, 3, 0, 142, 150, 30, 33, 124, 79, 48, 94, 88, 47, 11, 0, 14, 20, 5, 39, 61, 0, 0, 5, 21, 45, 23, 34, 110, 229, 237, 0, 
    384, 75, 0, 0, 159, 149, 0, 7, 139, 107, 44, 62, 105, 125, 102, 98, 102, 44, 63, 109, 101, 63, 68, 76, 107, 77, 0, 34, 117, 237, 268, 0, 
    394, 85, 0, 0, 124, 165, 21, 12, 91, 96, 56, 27, 43, 73, 93, 155, 143, 24, 29, 75, 69, 48, 61, 65, 103, 102, 0, 6, 106, 228, 269, 0, 
    396, 106, 0, 0, 37, 123, 71, 27, 41, 76, 97, 64, 36, 34, 33, 73, 134, 89, 41, 46, 51, 44, 63, 60, 53, 78, 43, 9, 47, 196, 275, 0, 
    386, 110, 0, 0, 28, 48, 61, 39, 11, 46, 91, 108, 95, 63, 0, 0, 87, 133, 40, 0, 25, 21, 55, 68, 0, 3, 123, 63, 6, 167, 289, 0, 
    373, 92, 0, 0, 99, 83, 27, 35, 0, 7, 66, 108, 146, 152, 67, 0, 75, 204, 104, 0, 36, 26, 65, 119, 0, 0, 149, 138, 44, 186, 297, 0, 
    358, 70, 0, 0, 94, 171, 94, 27, 0, 0, 44, 80, 108, 144, 122, 40, 89, 204, 192, 101, 103, 74, 75, 114, 17, 0, 105, 109, 89, 227, 287, 0, 
    332, 53, 0, 0, 6, 119, 148, 51, 0, 0, 18, 51, 75, 90, 91, 83, 84, 131, 191, 140, 63, 27, 24, 0, 0, 33, 85, 83, 97, 212, 254, 0, 
    315, 57, 3, 0, 0, 29, 110, 51, 0, 0, 0, 16, 63, 83, 84, 89, 73, 102, 234, 233, 110, 59, 50, 0, 0, 14, 98, 107, 107, 178, 213, 0, 
    310, 68, 53, 7, 0, 0, 82, 46, 0, 28, 0, 0, 44, 81, 83, 91, 84, 89, 190, 236, 169, 134, 106, 0, 0, 22, 104, 130, 112, 159, 194, 0, 
    305, 66, 54, 33, 3, 0, 60, 60, 5, 45, 14, 0, 38, 77, 82, 89, 106, 114, 131, 144, 133, 133, 104, 0, 0, 43, 105, 128, 112, 159, 185, 0, 
    305, 47, 35, 29, 25, 0, 14, 51, 45, 52, 26, 16, 40, 75, 83, 82, 89, 98, 104, 103, 106, 114, 104, 0, 0, 41, 110, 120, 117, 173, 173, 0, 
    293, 33, 29, 23, 22, 0, 0, 21, 74, 58, 33, 39, 50, 64, 74, 68, 66, 74, 79, 78, 85, 93, 94, 31, 0, 19, 103, 115, 125, 171, 137, 0, 
    278, 28, 22, 13, 12, 0, 0, 0, 80, 74, 54, 55, 59, 57, 58, 50, 51, 63, 64, 49, 48, 56, 59, 34, 0, 1, 69, 108, 132, 149, 94, 0, 
    311, 174, 177, 169, 159, 134, 72, 58, 122, 126, 128, 134, 131, 130, 128, 120, 122, 140, 151, 142, 135, 140, 140, 127, 103, 102, 126, 173, 231, 242, 216, 29, 
    
    -- channel=147
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=148
    0, 199, 200, 174, 174, 194, 212, 180, 156, 176, 173, 175, 169, 189, 194, 172, 167, 166, 184, 205, 209, 187, 181, 194, 225, 228, 181, 158, 192, 200, 164, 327, 
    0, 63, 70, 48, 37, 80, 132, 77, 8, 33, 43, 28, 21, 29, 31, 16, 1, 0, 9, 29, 45, 29, 11, 16, 79, 106, 73, 27, 75, 83, 47, 416, 
    0, 54, 57, 58, 40, 86, 171, 108, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 20, 0, 0, 34, 57, 65, 43, 49, 46, 37, 451, 
    0, 39, 38, 36, 30, 70, 174, 102, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 25, 57, 67, 10, 0, 34, 472, 
    0, 30, 30, 28, 32, 84, 219, 160, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 37, 27, 61, 66, 0, 0, 0, 479, 
    0, 30, 28, 25, 38, 87, 245, 248, 36, 0, 0, 21, 60, 30, 45, 65, 23, 13, 0, 0, 0, 0, 0, 20, 64, 54, 69, 69, 0, 0, 0, 461, 
    0, 30, 28, 30, 57, 53, 168, 266, 47, 0, 10, 69, 96, 53, 19, 27, 35, 36, 34, 16, 0, 0, 0, 0, 45, 86, 84, 111, 66, 0, 0, 415, 
    0, 32, 24, 49, 99, 49, 116, 242, 0, 0, 0, 0, 21, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 75, 88, 115, 102, 0, 0, 376, 
    0, 29, 22, 62, 112, 39, 100, 190, 0, 0, 0, 0, 0, 51, 0, 0, 0, 0, 0, 0, 0, 39, 0, 0, 14, 53, 77, 129, 145, 84, 0, 413, 
    0, 20, 25, 63, 110, 43, 61, 128, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 51, 155, 170, 122, 69, 482, 
    0, 0, 16, 68, 174, 125, 105, 114, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 87, 89, 58, 46, 518, 
    0, 0, 0, 65, 174, 122, 140, 159, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 29, 29, 29, 528, 
    0, 0, 0, 64, 87, 27, 114, 195, 72, 0, 0, 0, 0, 24, 12, 0, 0, 0, 0, 1, 20, 0, 0, 0, 0, 0, 0, 0, 0, 24, 30, 527, 
    0, 0, 28, 91, 70, 13, 86, 143, 74, 0, 0, 0, 0, 4, 15, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 527, 
    0, 35, 96, 76, 28, 15, 84, 112, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 529, 
    0, 50, 153, 98, 0, 0, 16, 124, 86, 0, 1, 38, 17, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 530, 
    0, 102, 239, 188, 0, 0, 0, 110, 45, 0, 27, 66, 98, 93, 64, 110, 74, 42, 73, 57, 70, 139, 98, 43, 8, 0, 0, 0, 0, 0, 0, 528, 
    0, 110, 222, 169, 0, 0, 91, 87, 0, 0, 0, 0, 0, 0, 47, 134, 108, 118, 151, 62, 68, 205, 183, 147, 96, 12, 19, 0, 0, 0, 0, 515, 
    0, 98, 214, 151, 0, 0, 204, 93, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 23, 13, 0, 0, 0, 29, 0, 0, 0, 0, 498, 
    0, 103, 240, 190, 0, 0, 167, 87, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 78, 24, 0, 0, 0, 481, 
    0, 75, 241, 257, 0, 0, 75, 66, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 41, 0, 0, 0, 466, 
    0, 52, 214, 254, 75, 6, 48, 52, 58, 0, 0, 0, 0, 0, 65, 57, 0, 0, 12, 63, 26, 22, 0, 8, 98, 51, 0, 0, 20, 0, 0, 451, 
    0, 40, 199, 197, 15, 12, 57, 68, 112, 67, 0, 0, 0, 0, 5, 114, 0, 0, 3, 114, 53, 62, 0, 0, 194, 112, 0, 0, 0, 0, 0, 441, 
    0, 28, 208, 212, 0, 0, 10, 58, 155, 107, 30, 0, 0, 0, 0, 69, 0, 0, 0, 0, 0, 8, 0, 0, 137, 94, 0, 0, 0, 0, 0, 426, 
    0, 21, 213, 277, 55, 0, 0, 31, 156, 121, 61, 17, 0, 0, 0, 3, 0, 0, 0, 0, 56, 110, 85, 92, 192, 79, 0, 0, 0, 0, 0, 407, 
    0, 11, 157, 259, 165, 15, 0, 26, 141, 104, 92, 65, 12, 0, 0, 0, 0, 0, 0, 0, 3, 65, 62, 192, 226, 44, 0, 0, 0, 0, 0, 395, 
    0, 0, 48, 127, 127, 60, 0, 40, 115, 51, 92, 95, 32, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 153, 234, 59, 0, 0, 0, 0, 0, 384, 
    0, 0, 0, 38, 90, 92, 0, 32, 71, 4, 68, 104, 53, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 159, 220, 54, 0, 0, 0, 0, 0, 383, 
    0, 0, 11, 33, 54, 90, 5, 25, 25, 0, 48, 81, 49, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 140, 192, 45, 0, 0, 0, 0, 0, 386, 
    0, 2, 13, 23, 31, 88, 90, 40, 0, 0, 32, 48, 36, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 85, 170, 58, 0, 0, 0, 0, 0, 393, 
    0, 10, 18, 33, 39, 99, 160, 78, 0, 0, 15, 21, 34, 24, 14, 19, 18, 3, 1, 12, 3, 0, 0, 55, 148, 94, 0, 0, 0, 0, 0, 402, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 156, 
    
    -- channel=149
    218, 171, 166, 169, 175, 168, 138, 136, 148, 141, 133, 138, 148, 142, 146, 158, 168, 179, 184, 183, 176, 179, 184, 186, 168, 152, 153, 163, 148, 135, 144, 4, 
    191, 40, 41, 45, 50, 26, 0, 0, 19, 26, 33, 45, 49, 62, 80, 86, 85, 73, 50, 40, 35, 31, 35, 40, 36, 36, 41, 43, 28, 30, 45, 0, 
    203, 44, 44, 45, 52, 35, 0, 0, 11, 0, 4, 14, 0, 9, 21, 15, 30, 25, 17, 19, 13, 18, 33, 39, 36, 36, 29, 21, 30, 44, 46, 0, 
    205, 42, 43, 43, 42, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 13, 15, 41, 43, 30, 30, 14, 0, 27, 51, 47, 0, 
    204, 34, 34, 36, 32, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 42, 52, 41, 25, 20, 5, 0, 17, 50, 52, 0, 
    203, 34, 35, 34, 19, 6, 0, 0, 0, 21, 21, 21, 5, 21, 24, 8, 3, 0, 0, 0, 0, 46, 75, 49, 25, 9, 0, 0, 3, 38, 57, 0, 
    203, 33, 36, 27, 0, 3, 0, 0, 15, 81, 70, 63, 40, 22, 24, 26, 29, 30, 27, 36, 29, 13, 42, 57, 26, 12, 13, 2, 3, 20, 51, 0, 
    202, 33, 37, 23, 0, 10, 0, 0, 2, 61, 36, 51, 35, 2, 0, 0, 2, 11, 12, 27, 29, 12, 18, 31, 23, 27, 30, 14, 3, 21, 45, 0, 
    202, 35, 36, 21, 0, 0, 0, 0, 3, 36, 0, 0, 0, 0, 0, 0, 2, 8, 0, 14, 18, 0, 27, 59, 45, 41, 39, 9, 0, 21, 50, 0, 
    199, 37, 37, 18, 0, 0, 0, 0, 7, 32, 0, 0, 0, 0, 0, 0, 2, 2, 0, 10, 22, 0, 17, 54, 62, 63, 51, 28, 39, 62, 78, 0, 
    188, 43, 39, 14, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 1, 0, 16, 40, 56, 44, 37, 51, 71, 69, 0, 
    175, 41, 33, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 51, 58, 45, 34, 35, 35, 35, 0, 
    163, 33, 15, 0, 0, 0, 0, 0, 0, 18, 11, 10, 15, 0, 0, 0, 0, 4, 22, 12, 0, 0, 0, 22, 59, 60, 39, 41, 46, 37, 34, 0, 
    163, 29, 0, 0, 0, 0, 0, 0, 15, 37, 24, 1, 0, 0, 0, 0, 1, 11, 19, 4, 0, 0, 0, 8, 17, 3, 0, 5, 48, 50, 35, 0, 
    170, 24, 0, 0, 0, 29, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 56, 40, 0, 
    153, 7, 0, 0, 0, 46, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 52, 67, 43, 0, 
    149, 0, 0, 0, 23, 49, 0, 0, 0, 4, 11, 41, 41, 32, 17, 0, 0, 0, 0, 13, 32, 0, 0, 0, 0, 25, 31, 29, 57, 77, 56, 0, 
    163, 17, 0, 0, 49, 46, 0, 0, 0, 22, 0, 10, 19, 38, 22, 20, 63, 71, 68, 95, 95, 60, 64, 71, 83, 86, 41, 18, 38, 81, 72, 0, 
    166, 10, 0, 0, 21, 17, 0, 0, 13, 11, 0, 0, 0, 0, 0, 38, 57, 27, 25, 46, 35, 0, 13, 37, 64, 60, 0, 0, 0, 61, 79, 0, 
    165, 11, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 1, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 79, 102, 0, 
    162, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 80, 112, 0, 
    161, 16, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 22, 45, 8, 0, 0, 21, 0, 0, 0, 0, 6, 34, 0, 0, 15, 34, 3, 72, 118, 0, 
    160, 13, 0, 0, 0, 23, 10, 0, 0, 0, 0, 0, 5, 32, 1, 0, 0, 71, 53, 21, 41, 31, 53, 77, 0, 0, 22, 5, 0, 74, 121, 0, 
    151, 4, 0, 0, 0, 12, 44, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 14, 6, 27, 23, 22, 0, 0, 0, 0, 0, 0, 70, 122, 0, 
    140, 0, 0, 0, 0, 20, 34, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 39, 44, 37, 16, 11, 0, 0, 0, 0, 0, 10, 92, 112, 0, 
    134, 9, 2, 0, 17, 30, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 93, 123, 92, 66, 54, 0, 0, 0, 0, 16, 37, 91, 103, 0, 
    135, 21, 18, 7, 8, 5, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 28, 63, 43, 0, 0, 0, 0, 0, 0, 0, 26, 35, 78, 95, 0, 
    143, 17, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 12, 23, 35, 7, 0, 0, 0, 0, 0, 0, 8, 29, 29, 73, 91, 0, 
    139, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 7, 0, 0, 0, 6, 20, 27, 82, 87, 0, 
    123, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 19, 49, 97, 73, 0, 
    124, 7, 12, 9, 5, 0, 0, 0, 0, 0, 0, 0, 0, 4, 8, 2, 2, 13, 19, 12, 7, 3, 0, 0, 0, 0, 10, 40, 82, 98, 62, 0, 
    17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 13, 8, 0, 0, 
    
    -- channel=150
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=151
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=152
    103, 235, 232, 223, 225, 237, 234, 199, 182, 189, 183, 179, 186, 198, 197, 198, 213, 231, 247, 254, 251, 241, 240, 245, 252, 232, 209, 203, 226, 208, 185, 245, 
    26, 251, 247, 241, 231, 254, 254, 205, 171, 192, 191, 186, 204, 203, 220, 233, 230, 241, 245, 249, 252, 244, 226, 233, 251, 256, 239, 214, 221, 221, 204, 298, 
    31, 264, 264, 263, 260, 267, 286, 226, 165, 178, 174, 182, 184, 171, 188, 202, 199, 228, 230, 226, 234, 230, 215, 223, 240, 254, 247, 228, 206, 222, 223, 314, 
    32, 273, 273, 271, 272, 280, 297, 227, 153, 161, 150, 161, 168, 145, 148, 152, 151, 173, 179, 173, 191, 202, 202, 221, 232, 237, 243, 226, 194, 202, 228, 333, 
    28, 275, 274, 273, 276, 281, 294, 235, 140, 147, 154, 154, 174, 157, 154, 159, 139, 139, 144, 125, 131, 165, 197, 227, 235, 228, 232, 219, 178, 166, 208, 347, 
    28, 275, 273, 274, 280, 272, 297, 273, 152, 149, 187, 196, 215, 207, 208, 215, 195, 180, 172, 147, 120, 133, 187, 230, 250, 237, 215, 207, 166, 140, 177, 339, 
    27, 274, 272, 280, 278, 248, 281, 297, 168, 152, 218, 244, 272, 263, 246, 247, 237, 231, 223, 202, 182, 140, 149, 205, 247, 236, 213, 207, 190, 151, 145, 306, 
    28, 273, 272, 281, 277, 244, 277, 283, 178, 160, 215, 213, 266, 272, 232, 235, 234, 237, 243, 224, 233, 188, 127, 171, 221, 230, 240, 235, 209, 155, 124, 268, 
    26, 272, 272, 280, 289, 258, 259, 252, 163, 148, 194, 181, 225, 258, 231, 221, 223, 222, 244, 221, 228, 245, 162, 147, 213, 246, 251, 252, 215, 179, 162, 279, 
    22, 266, 270, 282, 301, 237, 220, 227, 154, 159, 210, 188, 189, 224, 217, 207, 211, 213, 226, 216, 214, 244, 205, 162, 206, 238, 257, 274, 260, 237, 227, 335, 
    8, 249, 265, 283, 290, 236, 237, 216, 138, 121, 177, 182, 176, 190, 195, 194, 195, 194, 192, 195, 192, 217, 216, 164, 160, 210, 263, 282, 284, 267, 263, 374, 
    0, 225, 255, 275, 269, 246, 250, 224, 130, 83, 136, 172, 186, 185, 174, 171, 167, 163, 163, 174, 175, 172, 176, 151, 146, 203, 257, 276, 274, 273, 274, 383, 
    0, 200, 232, 244, 226, 198, 223, 217, 160, 128, 145, 170, 198, 209, 182, 161, 156, 164, 175, 196, 193, 155, 144, 148, 146, 172, 216, 242, 259, 272, 274, 382, 
    0, 195, 219, 210, 189, 153, 170, 196, 205, 174, 166, 174, 177, 203, 187, 158, 150, 158, 166, 176, 177, 145, 117, 114, 112, 135, 170, 177, 201, 254, 274, 382, 
    1, 212, 224, 177, 132, 122, 155, 216, 200, 173, 163, 149, 120, 125, 141, 132, 119, 120, 122, 121, 125, 110, 95, 93, 96, 108, 129, 126, 127, 211, 268, 383, 
    0, 192, 211, 149, 79, 99, 164, 221, 185, 150, 141, 134, 130, 115, 119, 120, 92, 72, 72, 64, 77, 86, 68, 61, 53, 68, 111, 127, 100, 166, 258, 384, 
    0, 186, 227, 168, 78, 91, 157, 164, 155, 122, 138, 151, 173, 155, 147, 139, 90, 70, 89, 77, 111, 144, 95, 76, 73, 90, 136, 159, 139, 146, 236, 383, 
    23, 219, 241, 180, 82, 105, 160, 112, 93, 115, 135, 131, 146, 155, 175, 150, 142, 157, 165, 156, 172, 208, 185, 155, 151, 158, 185, 185, 148, 112, 197, 378, 
    26, 233, 247, 186, 72, 109, 165, 109, 49, 91, 117, 97, 85, 108, 113, 123, 176, 191, 165, 157, 161, 192, 192, 168, 153, 184, 204, 150, 109, 89, 163, 370, 
    20, 237, 263, 203, 66, 69, 141, 117, 50, 53, 95, 106, 83, 66, 76, 90, 115, 163, 155, 140, 148, 153, 142, 138, 135, 160, 186, 136, 95, 75, 140, 362, 
    14, 229, 267, 220, 96, 53, 107, 111, 66, 42, 60, 84, 89, 89, 98, 74, 69, 134, 146, 128, 121, 129, 114, 126, 133, 103, 140, 150, 121, 74, 127, 355, 
    14, 224, 266, 221, 118, 90, 93, 98, 84, 53, 33, 40, 77, 102, 149, 131, 42, 56, 136, 147, 122, 127, 108, 127, 188, 122, 86, 154, 165, 77, 112, 347, 
    25, 226, 261, 207, 86, 102, 105, 111, 121, 79, 38, 28, 45, 71, 132, 132, 43, 33, 140, 170, 144, 157, 134, 147, 230, 141, 53, 105, 126, 62, 103, 339, 
    29, 229, 258, 198, 56, 51, 110, 148, 161, 106, 54, 33, 14, 23, 50, 90, 50, 13, 67, 129, 133, 149, 150, 143, 166, 133, 43, 47, 80, 51, 104, 331, 
    31, 226, 247, 219, 102, 52, 105, 170, 171, 129, 74, 43, 25, 16, 17, 45, 41, 0, 0, 115, 176, 203, 199, 195, 167, 109, 46, 43, 62, 45, 108, 323, 
    29, 214, 235, 259, 197, 128, 96, 160, 176, 135, 104, 68, 32, 20, 19, 20, 30, 20, 16, 121, 213, 229, 224, 248, 191, 71, 27, 40, 68, 63, 119, 317, 
    25, 207, 230, 254, 233, 174, 117, 163, 171, 128, 123, 87, 37, 19, 21, 21, 34, 50, 37, 77, 153, 176, 197, 223, 182, 66, 16, 34, 73, 77, 132, 311, 
    36, 216, 217, 215, 217, 202, 143, 150, 152, 117, 117, 99, 54, 27, 30, 32, 40, 56, 49, 55, 104, 133, 163, 209, 160, 58, 19, 33, 68, 80, 139, 310, 
    44, 214, 213, 211, 204, 200, 159, 122, 128, 106, 108, 95, 64, 38, 37, 40, 39, 44, 59, 72, 90, 106, 129, 181, 155, 52, 19, 34, 59, 80, 152, 308, 
    39, 211, 214, 208, 203, 206, 181, 111, 97, 98, 99, 82, 69, 52, 49, 54, 57, 56, 62, 72, 80, 88, 103, 138, 154, 61, 20, 37, 56, 98, 175, 311, 
    40, 212, 216, 221, 220, 219, 209, 127, 77, 80, 82, 75, 76, 73, 72, 78, 76, 73, 82, 99, 102, 103, 111, 125, 136, 91, 50, 48, 82, 140, 199, 319, 
    0, 100, 102, 104, 102, 101, 106, 68, 21, 22, 28, 29, 25, 29, 30, 33, 33, 32, 36, 44, 47, 47, 47, 51, 57, 49, 23, 16, 33, 54, 88, 146, 
    
    -- channel=153
    229, 288, 284, 275, 283, 284, 265, 236, 234, 250, 257, 266, 279, 295, 304, 311, 315, 312, 310, 306, 297, 285, 283, 288, 294, 285, 269, 263, 263, 252, 250, 232, 
    154, 100, 101, 109, 111, 103, 79, 49, 44, 69, 91, 100, 106, 114, 133, 151, 143, 124, 97, 73, 67, 64, 57, 59, 77, 94, 105, 84, 66, 71, 96, 80, 
    165, 111, 110, 112, 116, 112, 91, 73, 72, 71, 72, 78, 68, 47, 46, 47, 41, 49, 49, 34, 24, 28, 41, 56, 64, 71, 69, 46, 34, 63, 95, 59, 
    163, 102, 103, 103, 103, 87, 60, 48, 66, 83, 83, 90, 81, 62, 49, 24, 10, 13, 3, 0, 1, 15, 46, 67, 58, 51, 39, 16, 10, 41, 72, 46, 
    162, 95, 95, 96, 95, 88, 73, 69, 102, 138, 164, 180, 171, 180, 178, 150, 126, 97, 55, 17, 3, 38, 75, 81, 63, 43, 23, 0, 0, 10, 38, 40, 
    161, 95, 95, 94, 87, 76, 94, 142, 201, 239, 275, 291, 279, 291, 303, 299, 289, 260, 229, 179, 93, 63, 85, 87, 73, 54, 17, 0, 0, 0, 18, 25, 
    161, 93, 95, 93, 78, 63, 85, 141, 218, 280, 304, 312, 311, 298, 287, 287, 298, 305, 298, 289, 234, 113, 42, 44, 55, 54, 42, 46, 42, 21, 11, 1, 
    161, 95, 96, 95, 86, 84, 108, 132, 183, 226, 204, 187, 216, 240, 240, 241, 247, 259, 268, 259, 253, 185, 75, 32, 44, 56, 75, 68, 42, 25, 13, 0, 
    159, 92, 94, 92, 88, 88, 108, 127, 190, 228, 185, 141, 147, 187, 231, 250, 248, 241, 248, 247, 238, 204, 150, 108, 90, 98, 103, 83, 61, 71, 96, 54, 
    152, 86, 93, 90, 75, 63, 82, 127, 196, 230, 221, 206, 179, 184, 228, 243, 239, 227, 223, 230, 237, 220, 178, 127, 96, 103, 105, 108, 127, 157, 168, 111, 
    133, 70, 87, 89, 94, 110, 153, 164, 167, 165, 172, 203, 199, 196, 219, 227, 217, 203, 192, 197, 205, 199, 175, 120, 70, 74, 95, 98, 115, 136, 132, 80, 
    120, 59, 72, 62, 61, 120, 203, 194, 171, 155, 172, 218, 239, 231, 213, 202, 194, 188, 198, 209, 189, 155, 138, 127, 110, 104, 100, 95, 96, 96, 95, 50, 
    122, 56, 47, 27, 16, 50, 115, 169, 226, 259, 262, 250, 271, 276, 249, 225, 227, 245, 271, 274, 231, 171, 133, 120, 109, 73, 40, 52, 81, 94, 95, 50, 
    137, 74, 49, 20, 20, 41, 75, 133, 225, 277, 273, 236, 223, 223, 221, 216, 214, 216, 211, 187, 152, 137, 128, 112, 87, 46, 11, 8, 43, 82, 95, 50, 
    139, 78, 38, 0, 4, 66, 122, 162, 202, 206, 181, 140, 121, 115, 128, 151, 159, 152, 135, 103, 77, 93, 112, 106, 83, 62, 56, 49, 46, 70, 91, 52, 
    108, 36, 16, 1, 14, 56, 99, 126, 152, 188, 195, 187, 199, 189, 174, 153, 115, 89, 83, 93, 109, 109, 90, 71, 71, 97, 133, 144, 119, 93, 89, 51, 
    129, 59, 62, 80, 97, 88, 43, 13, 92, 180, 192, 215, 258, 269, 248, 210, 178, 186, 198, 216, 255, 255, 208, 182, 185, 216, 250, 238, 193, 128, 90, 49, 
    148, 95, 90, 84, 109, 103, 42, 0, 92, 173, 159, 124, 131, 166, 197, 198, 235, 279, 283, 282, 283, 270, 273, 284, 292, 302, 257, 192, 147, 101, 83, 46, 
    150, 97, 87, 65, 71, 69, 50, 61, 133, 146, 118, 92, 64, 58, 88, 125, 186, 180, 135, 139, 138, 103, 118, 143, 160, 191, 158, 99, 84, 88, 98, 48, 
    145, 91, 98, 84, 63, 37, 40, 101, 150, 122, 105, 127, 137, 123, 99, 99, 128, 121, 123, 128, 120, 106, 107, 113, 108, 109, 101, 107, 128, 139, 129, 55, 
    139, 84, 100, 110, 111, 70, 62, 113, 130, 101, 94, 121, 159, 185, 182, 136, 78, 76, 125, 139, 123, 114, 127, 142, 134, 97, 102, 177, 208, 172, 135, 57, 
    145, 92, 88, 88, 135, 138, 114, 124, 129, 116, 103, 104, 149, 212, 224, 166, 112, 126, 168, 176, 169, 174, 183, 214, 200, 129, 126, 192, 204, 156, 129, 59, 
    162, 111, 92, 54, 71, 125, 155, 168, 164, 136, 115, 101, 102, 106, 118, 105, 106, 139, 178, 191, 205, 216, 208, 201, 176, 128, 111, 106, 96, 112, 140, 69, 
    173, 123, 101, 65, 52, 71, 143, 207, 186, 138, 116, 108, 91, 52, 22, 29, 87, 91, 57, 67, 126, 153, 144, 102, 34, 46, 108, 78, 57, 121, 167, 80, 
    186, 141, 142, 144, 170, 152, 151, 179, 154, 132, 129, 111, 101, 95, 73, 68, 98, 102, 102, 164, 234, 233, 218, 181, 80, 58, 105, 111, 134, 181, 187, 84, 
    188, 152, 171, 215, 254, 231, 185, 149, 123, 142, 151, 124, 100, 94, 99, 104, 111, 117, 144, 189, 201, 192, 178, 166, 120, 91, 90, 120, 170, 207, 203, 102, 
    193, 166, 168, 179, 200, 189, 162, 144, 128, 145, 146, 125, 105, 101, 107, 118, 137, 161, 160, 100, 38, 45, 80, 76, 50, 73, 101, 133, 173, 196, 205, 115, 
    206, 175, 162, 142, 144, 154, 138, 120, 114, 141, 130, 111, 109, 115, 120, 123, 120, 128, 134, 98, 59, 77, 112, 99, 61, 80, 114, 142, 163, 186, 210, 122, 
    205, 170, 157, 152, 156, 160, 136, 100, 98, 135, 122, 108, 111, 117, 120, 123, 120, 109, 105, 107, 111, 119, 118, 106, 87, 97, 110, 133, 154, 190, 222, 127, 
    201, 168, 173, 180, 184, 174, 143, 107, 106, 130, 117, 107, 115, 128, 132, 135, 136, 135, 137, 136, 132, 124, 110, 89, 90, 110, 116, 139, 175, 226, 245, 130, 
    214, 199, 214, 215, 207, 196, 163, 125, 113, 111, 111, 118, 133, 148, 160, 160, 159, 164, 176, 182, 180, 170, 158, 136, 129, 148, 164, 181, 221, 264, 244, 126, 
    30, 0, 0, 0, 0, 0, 0, 0, 19, 11, 4, 11, 16, 20, 26, 24, 21, 18, 13, 9, 6, 1, 0, 0, 0, 13, 37, 26, 8, 0, 0, 0, 
    
    -- channel=154
    53, 44, 39, 31, 41, 52, 39, 14, 20, 29, 22, 22, 26, 29, 25, 24, 29, 36, 48, 54, 48, 39, 42, 49, 52, 33, 19, 14, 31, 10, 12, 50, 
    129, 85, 81, 80, 88, 97, 82, 39, 40, 60, 60, 66, 64, 67, 72, 80, 83, 98, 95, 89, 85, 76, 73, 81, 86, 72, 58, 46, 53, 38, 42, 85, 
    142, 102, 101, 98, 101, 111, 103, 48, 54, 78, 68, 93, 84, 78, 94, 96, 96, 111, 91, 84, 71, 66, 67, 79, 85, 83, 73, 51, 42, 49, 64, 101, 
    153, 117, 117, 115, 116, 119, 109, 54, 71, 101, 84, 114, 105, 87, 104, 96, 90, 109, 83, 74, 65, 53, 62, 84, 78, 81, 74, 40, 23, 44, 72, 111, 
    159, 124, 123, 122, 125, 124, 121, 57, 71, 123, 113, 139, 128, 120, 129, 114, 106, 117, 91, 65, 48, 57, 66, 89, 80, 70, 60, 30, 4, 30, 64, 118, 
    159, 123, 124, 124, 126, 114, 123, 80, 72, 139, 148, 166, 156, 156, 170, 159, 154, 147, 130, 107, 58, 53, 85, 98, 90, 73, 47, 28, 0, 7, 46, 119, 
    159, 123, 123, 127, 123, 102, 127, 101, 73, 154, 170, 176, 184, 175, 187, 195, 187, 188, 174, 159, 134, 72, 67, 99, 94, 74, 53, 32, 9, 0, 24, 114, 
    159, 122, 122, 129, 121, 95, 141, 114, 86, 159, 169, 169, 202, 188, 193, 202, 194, 196, 194, 178, 177, 126, 69, 78, 89, 77, 66, 47, 16, 6, 15, 95, 
    157, 121, 123, 128, 120, 96, 145, 121, 96, 173, 169, 150, 183, 178, 182, 198, 194, 192, 197, 180, 200, 156, 90, 92, 94, 85, 87, 77, 36, 21, 29, 95, 
    152, 120, 123, 127, 124, 89, 143, 112, 105, 172, 172, 158, 180, 171, 179, 190, 189, 187, 190, 178, 199, 186, 125, 105, 105, 109, 116, 101, 73, 62, 69, 126, 
    137, 115, 123, 128, 127, 95, 133, 103, 98, 139, 158, 160, 167, 162, 172, 178, 178, 175, 175, 169, 186, 190, 157, 124, 110, 124, 127, 114, 104, 107, 112, 150, 
    120, 105, 119, 121, 103, 87, 147, 110, 85, 100, 131, 150, 163, 153, 151, 154, 156, 152, 151, 157, 153, 146, 141, 119, 107, 117, 129, 124, 124, 124, 124, 157, 
    110, 92, 112, 103, 79, 67, 127, 97, 101, 97, 129, 145, 173, 176, 150, 139, 143, 146, 150, 161, 139, 108, 100, 87, 89, 110, 116, 116, 128, 125, 123, 157, 
    108, 92, 98, 75, 61, 50, 84, 75, 106, 121, 159, 153, 166, 175, 151, 131, 128, 137, 146, 153, 128, 89, 77, 76, 88, 100, 99, 90, 116, 136, 123, 157, 
    105, 88, 81, 35, 37, 47, 70, 79, 105, 140, 152, 122, 123, 128, 123, 111, 109, 121, 125, 120, 94, 70, 70, 70, 75, 83, 97, 91, 96, 137, 129, 156, 
    96, 75, 76, 12, 12, 28, 65, 89, 100, 118, 137, 102, 95, 80, 86, 77, 54, 58, 60, 56, 66, 52, 38, 50, 54, 84, 111, 103, 96, 132, 133, 156, 
    107, 69, 71, 2, 8, 34, 68, 54, 77, 92, 97, 75, 95, 77, 87, 63, 31, 31, 32, 21, 59, 59, 19, 27, 28, 61, 113, 121, 106, 121, 139, 158, 
    116, 74, 84, 13, 18, 58, 62, 4, 46, 89, 87, 65, 97, 99, 115, 71, 62, 54, 52, 54, 83, 89, 55, 47, 49, 90, 115, 113, 106, 106, 143, 161, 
    129, 92, 100, 18, 12, 62, 49, 0, 27, 74, 84, 59, 63, 62, 86, 75, 101, 94, 86, 95, 124, 108, 83, 92, 86, 135, 126, 89, 93, 82, 136, 165, 
    132, 94, 104, 23, 2, 45, 37, 0, 25, 50, 71, 52, 43, 49, 61, 48, 117, 129, 98, 101, 113, 109, 99, 102, 93, 117, 112, 67, 67, 68, 138, 169, 
    127, 95, 112, 36, 12, 19, 25, 9, 20, 16, 35, 44, 52, 53, 60, 49, 75, 88, 91, 93, 96, 93, 83, 98, 87, 91, 94, 80, 80, 60, 134, 174, 
    128, 99, 116, 30, 22, 34, 14, 25, 19, 0, 6, 16, 50, 66, 94, 42, 24, 69, 98, 75, 70, 82, 62, 94, 105, 30, 56, 103, 92, 52, 129, 175, 
    135, 111, 124, 28, 2, 49, 37, 39, 31, 0, 0, 0, 20, 45, 89, 43, 0, 26, 89, 67, 65, 83, 57, 91, 107, 16, 30, 84, 84, 49, 130, 176, 
    145, 130, 132, 28, 0, 23, 51, 79, 51, 6, 0, 0, 4, 14, 40, 11, 0, 9, 59, 65, 66, 89, 73, 89, 78, 11, 20, 51, 39, 31, 138, 181, 
    152, 145, 143, 57, 4, 24, 46, 103, 71, 26, 0, 0, 0, 0, 0, 0, 0, 2, 39, 81, 89, 100, 85, 111, 41, 0, 6, 16, 25, 42, 147, 185, 
    143, 143, 144, 102, 60, 48, 65, 115, 64, 41, 19, 0, 0, 0, 0, 0, 0, 0, 1, 86, 110, 116, 109, 118, 35, 0, 0, 6, 37, 62, 156, 187, 
    133, 140, 141, 129, 116, 92, 69, 113, 55, 55, 38, 0, 0, 0, 0, 0, 0, 0, 14, 84, 105, 109, 112, 115, 17, 0, 0, 6, 53, 76, 160, 187, 
    136, 137, 142, 141, 127, 104, 64, 95, 53, 62, 49, 8, 0, 0, 0, 0, 0, 5, 33, 74, 79, 88, 107, 112, 2, 0, 0, 11, 56, 80, 163, 185, 
    141, 148, 147, 134, 122, 107, 73, 71, 45, 59, 45, 12, 0, 0, 0, 0, 1, 13, 27, 45, 59, 80, 100, 105, 17, 0, 0, 14, 47, 82, 169, 180, 
    146, 150, 148, 139, 133, 120, 78, 45, 38, 52, 35, 12, 0, 0, 0, 1, 5, 11, 25, 37, 49, 66, 79, 81, 25, 0, 0, 12, 42, 98, 175, 178, 
    146, 150, 156, 150, 142, 133, 99, 27, 26, 36, 27, 16, 8, 6, 15, 18, 19, 23, 35, 46, 50, 59, 65, 66, 35, 0, 0, 15, 60, 120, 177, 175, 
    46, 79, 83, 83, 84, 76, 54, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 12, 16, 18, 20, 20, 5, 0, 0, 0, 17, 68, 99, 95, 
    
    -- channel=155
    187, 406, 406, 400, 388, 389, 391, 362, 330, 329, 328, 324, 336, 357, 368, 379, 401, 420, 429, 433, 432, 424, 416, 416, 419, 411, 394, 391, 398, 389, 354, 352, 
    0, 216, 223, 209, 198, 202, 211, 175, 139, 147, 149, 157, 175, 197, 216, 233, 229, 210, 208, 205, 211, 202, 186, 182, 213, 240, 244, 232, 229, 227, 222, 323, 
    0, 214, 218, 219, 209, 214, 226, 179, 104, 96, 86, 73, 88, 70, 73, 91, 94, 117, 148, 164, 187, 177, 163, 167, 192, 209, 224, 216, 210, 205, 211, 325, 
    0, 198, 198, 198, 194, 206, 211, 135, 33, 26, 17, 0, 18, 0, 0, 0, 0, 8, 45, 76, 130, 154, 145, 162, 180, 177, 202, 216, 197, 187, 198, 329, 
    0, 182, 183, 182, 183, 188, 204, 136, 5, 0, 0, 0, 19, 6, 5, 4, 0, 0, 0, 7, 58, 116, 153, 170, 182, 180, 196, 208, 178, 153, 174, 332, 
    0, 182, 180, 179, 180, 185, 218, 194, 70, 23, 58, 82, 100, 87, 98, 105, 77, 61, 41, 38, 62, 88, 132, 178, 190, 189, 187, 182, 163, 135, 147, 321, 
    0, 181, 180, 180, 175, 154, 185, 202, 94, 48, 121, 159, 168, 143, 107, 101, 103, 102, 101, 89, 87, 97, 83, 118, 172, 186, 190, 212, 206, 164, 122, 283, 
    0, 182, 181, 182, 182, 154, 159, 167, 52, 19, 64, 75, 102, 101, 48, 36, 55, 69, 77, 86, 90, 89, 70, 83, 140, 180, 211, 244, 221, 151, 100, 252, 
    0, 180, 179, 189, 198, 158, 125, 115, 15, 0, 4, 0, 24, 59, 37, 29, 35, 49, 62, 48, 65, 112, 94, 89, 154, 199, 218, 229, 219, 181, 155, 297, 
    0, 170, 176, 190, 189, 107, 54, 71, 8, 0, 35, 2, 2, 24, 21, 20, 23, 30, 42, 28, 36, 85, 92, 94, 129, 163, 196, 238, 257, 256, 237, 354, 
    0, 142, 168, 187, 182, 127, 96, 87, 0, 0, 0, 0, 0, 1, 2, 3, 3, 0, 0, 0, 0, 26, 41, 30, 36, 93, 169, 222, 230, 223, 213, 352, 
    0, 113, 146, 170, 188, 155, 139, 116, 10, 0, 0, 6, 24, 31, 11, 0, 0, 0, 0, 0, 6, 2, 4, 10, 36, 100, 162, 182, 181, 180, 181, 341, 
    0, 93, 108, 126, 121, 90, 100, 108, 67, 48, 41, 40, 36, 54, 47, 17, 9, 26, 47, 76, 87, 52, 39, 51, 53, 70, 101, 123, 150, 177, 182, 341, 
    0, 96, 109, 110, 84, 59, 72, 114, 108, 72, 41, 23, 7, 21, 33, 24, 18, 18, 11, 23, 45, 37, 24, 4, 0, 0, 18, 36, 65, 137, 182, 341, 
    0, 125, 133, 90, 40, 48, 110, 155, 94, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 75, 167, 343, 
    0, 104, 112, 69, 14, 42, 115, 139, 64, 0, 0, 20, 22, 23, 17, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 148, 343, 
    0, 124, 163, 138, 55, 44, 70, 65, 0, 20, 74, 116, 145, 144, 116, 115, 72, 54, 82, 90, 108, 149, 115, 63, 53, 31, 48, 61, 34, 50, 120, 339, 
    0, 166, 188, 153, 59, 48, 81, 33, 0, 17, 68, 57, 47, 63, 96, 133, 150, 212, 231, 203, 211, 245, 240, 234, 205, 159, 142, 93, 21, 0, 70, 329, 
    0, 153, 174, 130, 27, 34, 116, 62, 0, 0, 8, 0, 0, 0, 0, 37, 101, 139, 96, 41, 47, 94, 99, 98, 81, 79, 93, 18, 0, 0, 42, 318, 
    0, 157, 195, 152, 13, 0, 90, 81, 7, 0, 0, 21, 10, 0, 0, 0, 0, 4, 10, 0, 0, 0, 0, 0, 0, 10, 41, 23, 0, 0, 32, 311, 
    0, 142, 195, 177, 53, 20, 58, 70, 34, 0, 0, 12, 30, 40, 36, 0, 0, 0, 14, 3, 0, 0, 0, 7, 1, 0, 10, 52, 54, 1, 22, 303, 
    0, 130, 187, 186, 87, 72, 77, 59, 67, 36, 2, 0, 15, 57, 106, 93, 0, 0, 36, 75, 42, 42, 47, 60, 117, 80, 4, 59, 95, 5, 2, 293, 
    0, 120, 164, 150, 58, 47, 86, 90, 119, 97, 43, 10, 0, 0, 48, 81, 18, 5, 96, 154, 123, 130, 119, 124, 190, 122, 0, 0, 10, 0, 0, 287, 
    0, 96, 152, 130, 15, 4, 49, 117, 159, 117, 70, 17, 0, 0, 0, 20, 6, 0, 0, 32, 56, 79, 67, 44, 83, 44, 0, 0, 0, 0, 0, 273, 
    0, 72, 138, 172, 92, 48, 54, 92, 136, 108, 89, 57, 26, 0, 0, 21, 6, 0, 0, 37, 144, 179, 149, 120, 136, 60, 8, 13, 11, 0, 0, 248, 
    0, 65, 138, 212, 209, 130, 51, 67, 112, 97, 109, 97, 58, 34, 30, 24, 27, 18, 13, 90, 183, 191, 175, 199, 174, 63, 12, 16, 22, 0, 0, 238, 
    0, 76, 121, 161, 151, 109, 52, 77, 105, 77, 105, 104, 66, 42, 39, 38, 53, 55, 3, 0, 0, 22, 45, 125, 137, 54, 18, 8, 13, 0, 0, 233, 
    0, 90, 80, 78, 90, 97, 65, 69, 73, 48, 79, 97, 82, 62, 56, 52, 54, 40, 0, 0, 0, 0, 19, 111, 137, 60, 26, 5, 1, 0, 0, 234, 
    0, 69, 63, 74, 90, 104, 69, 52, 37, 37, 65, 83, 81, 65, 55, 45, 24, 9, 0, 0, 0, 0, 4, 85, 124, 72, 20, 1, 0, 0, 4, 239, 
    0, 58, 62, 72, 82, 111, 101, 58, 22, 38, 59, 66, 68, 66, 58, 56, 52, 39, 27, 20, 5, 0, 0, 58, 107, 81, 26, 10, 9, 0, 38, 242, 
    0, 68, 81, 98, 105, 117, 132, 92, 28, 30, 43, 60, 76, 76, 74, 76, 72, 64, 66, 72, 64, 51, 43, 73, 112, 105, 72, 50, 46, 48, 74, 244, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 
    
    -- channel=156
    309, 418, 407, 403, 418, 420, 392, 355, 342, 334, 319, 315, 316, 320, 317, 328, 363, 405, 440, 451, 442, 434, 442, 447, 429, 388, 362, 370, 375, 343, 325, 233, 
    316, 379, 377, 369, 374, 370, 334, 276, 269, 290, 295, 304, 317, 342, 363, 385, 402, 408, 401, 395, 388, 372, 369, 375, 384, 369, 355, 348, 344, 316, 316, 247, 
    338, 405, 403, 402, 405, 403, 354, 272, 248, 258, 259, 271, 273, 279, 309, 330, 346, 365, 362, 360, 360, 352, 350, 364, 382, 385, 377, 349, 338, 336, 348, 266, 
    350, 419, 418, 418, 416, 405, 343, 241, 206, 206, 196, 211, 202, 189, 205, 210, 229, 268, 282, 298, 315, 318, 336, 365, 372, 374, 364, 331, 318, 344, 366, 272, 
    349, 413, 414, 414, 414, 393, 309, 172, 125, 142, 136, 159, 153, 143, 149, 136, 138, 159, 165, 197, 245, 296, 338, 374, 368, 359, 350, 315, 292, 324, 361, 283, 
    349, 413, 413, 413, 407, 388, 331, 196, 123, 151, 174, 199, 197, 198, 212, 199, 179, 171, 159, 167, 197, 275, 356, 388, 377, 354, 329, 290, 260, 283, 339, 289, 
    348, 412, 413, 410, 388, 358, 338, 234, 160, 211, 266, 294, 285, 261, 262, 260, 250, 242, 231, 233, 233, 250, 317, 373, 378, 355, 321, 295, 264, 262, 306, 275, 
    348, 412, 413, 408, 374, 336, 321, 225, 154, 230, 291, 324, 329, 278, 238, 231, 236, 246, 244, 256, 277, 257, 258, 314, 352, 354, 349, 339, 296, 261, 269, 240, 
    347, 412, 412, 407, 374, 335, 303, 200, 141, 203, 212, 220, 257, 233, 208, 215, 225, 240, 242, 238, 272, 267, 260, 313, 353, 372, 388, 360, 300, 264, 279, 234, 
    342, 408, 411, 405, 357, 282, 234, 155, 138, 199, 202, 194, 214, 198, 195, 205, 214, 227, 232, 226, 260, 274, 268, 320, 374, 403, 415, 398, 367, 360, 379, 295, 
    325, 394, 409, 402, 338, 238, 190, 130, 104, 149, 165, 166, 168, 161, 168, 176, 182, 185, 185, 186, 219, 246, 248, 271, 317, 372, 411, 423, 422, 430, 431, 326, 
    295, 367, 394, 384, 332, 274, 247, 143, 66, 75, 115, 150, 156, 148, 144, 142, 140, 137, 139, 150, 162, 176, 192, 212, 267, 351, 408, 414, 414, 414, 414, 318, 
    272, 340, 358, 333, 280, 251, 238, 157, 102, 98, 139, 168, 189, 176, 140, 121, 124, 139, 165, 190, 171, 143, 152, 193, 267, 343, 379, 393, 409, 413, 414, 318, 
    264, 317, 313, 275, 228, 202, 188, 164, 169, 178, 188, 168, 179, 182, 154, 133, 138, 162, 190, 209, 185, 144, 142, 163, 205, 245, 268, 304, 365, 408, 414, 318, 
    270, 322, 287, 214, 193, 201, 217, 200, 177, 147, 137, 105, 88, 93, 90, 87, 86, 89, 83, 82, 73, 71, 85, 99, 125, 155, 178, 203, 280, 378, 413, 319, 
    265, 310, 246, 134, 129, 197, 268, 247, 151, 103, 98, 66, 44, 41, 49, 44, 27, 19, 13, 14, 18, 17, 19, 25, 40, 73, 116, 151, 225, 344, 405, 319, 
    254, 283, 230, 132, 130, 197, 226, 174, 95, 108, 139, 163, 179, 160, 139, 98, 41, 24, 25, 40, 83, 76, 27, 9, 21, 70, 144, 182, 230, 329, 398, 318, 
    283, 316, 270, 168, 167, 210, 165, 51, 49, 119, 151, 164, 189, 193, 195, 171, 163, 192, 210, 219, 267, 265, 212, 199, 195, 215, 233, 223, 236, 295, 379, 317, 
    294, 319, 257, 139, 141, 191, 138, 11, 41, 111, 118, 78, 72, 91, 138, 167, 233, 260, 241, 234, 259, 250, 236, 247, 250, 271, 228, 155, 148, 215, 350, 314, 
    293, 325, 267, 132, 93, 138, 111, 31, 39, 65, 72, 57, 42, 39, 58, 103, 193, 179, 130, 130, 147, 138, 128, 130, 145, 188, 155, 85, 98, 192, 344, 313, 
    286, 328, 283, 147, 68, 79, 77, 48, 31, 15, 34, 58, 67, 70, 71, 64, 98, 121, 132, 128, 121, 110, 113, 128, 123, 131, 121, 110, 128, 194, 336, 314, 
    277, 323, 285, 166, 107, 94, 75, 60, 34, 0, 0, 23, 70, 116, 132, 65, 31, 71, 105, 93, 79, 81, 94, 140, 127, 65, 95, 160, 170, 190, 322, 310, 
    276, 321, 271, 135, 100, 122, 106, 91, 70, 24, 2, 3, 51, 113, 156, 82, 23, 102, 196, 187, 169, 176, 183, 246, 230, 97, 79, 141, 142, 154, 306, 306, 
    266, 308, 253, 97, 37, 92, 134, 161, 128, 52, 12, 0, 0, 1, 36, 11, 1, 70, 153, 163, 175, 197, 187, 204, 167, 46, 26, 46, 41, 115, 302, 301, 
    244, 285, 250, 124, 49, 81, 142, 197, 154, 68, 24, 0, 0, 0, 0, 0, 0, 4, 64, 137, 198, 223, 209, 177, 78, 1, 17, 30, 45, 131, 295, 284, 
    223, 268, 275, 229, 182, 158, 171, 189, 134, 89, 56, 11, 0, 0, 0, 0, 0, 0, 96, 263, 345, 346, 316, 263, 119, 13, 3, 32, 76, 152, 285, 268, 
    210, 266, 289, 289, 252, 195, 170, 185, 127, 107, 87, 33, 0, 0, 0, 0, 16, 35, 97, 204, 241, 248, 245, 212, 77, 0, 0, 33, 91, 158, 276, 263, 
    219, 275, 276, 255, 221, 180, 158, 171, 116, 102, 90, 42, 1, 0, 0, 12, 40, 69, 93, 119, 126, 156, 195, 172, 48, 0, 0, 38, 89, 150, 269, 257, 
    225, 272, 254, 232, 217, 193, 148, 127, 85, 89, 80, 47, 19, 10, 15, 19, 24, 34, 48, 73, 99, 136, 175, 166, 53, 0, 2, 34, 78, 150, 275, 254, 
    207, 244, 236, 233, 227, 204, 139, 88, 66, 79, 68, 48, 32, 25, 28, 32, 34, 38, 49, 61, 75, 95, 114, 126, 55, 4, 2, 33, 84, 173, 290, 248, 
    198, 239, 244, 246, 245, 228, 156, 69, 53, 63, 58, 50, 50, 52, 58, 61, 61, 66, 82, 92, 97, 103, 109, 114, 78, 35, 30, 65, 133, 229, 312, 245, 
    97, 129, 142, 145, 138, 124, 86, 18, 0, 0, 0, 8, 17, 18, 24, 25, 22, 28, 46, 58, 59, 60, 60, 56, 42, 21, 20, 37, 85, 146, 172, 142, 
    
    -- channel=157
    391, 349, 334, 340, 357, 353, 306, 284, 290, 282, 274, 274, 279, 270, 272, 294, 323, 355, 376, 376, 363, 364, 372, 374, 341, 304, 298, 314, 291, 258, 268, 56, 
    478, 341, 336, 341, 359, 334, 263, 228, 258, 270, 280, 298, 300, 321, 343, 360, 377, 383, 369, 358, 343, 331, 340, 351, 338, 317, 308, 309, 280, 263, 286, 23, 
    508, 372, 369, 369, 381, 359, 262, 206, 246, 248, 256, 280, 264, 288, 317, 320, 349, 351, 338, 337, 314, 308, 330, 352, 354, 345, 325, 296, 292, 303, 318, 25, 
    528, 391, 390, 390, 390, 354, 229, 164, 214, 209, 214, 230, 203, 214, 229, 226, 261, 279, 281, 301, 291, 286, 331, 356, 347, 345, 313, 266, 284, 325, 333, 24, 
    533, 390, 390, 392, 387, 342, 201, 93, 145, 175, 184, 200, 174, 185, 184, 164, 182, 192, 191, 222, 266, 309, 347, 359, 340, 330, 291, 243, 257, 318, 341, 28, 
    533, 390, 391, 391, 371, 338, 227, 100, 142, 214, 232, 243, 219, 236, 244, 216, 211, 201, 193, 202, 241, 323, 380, 371, 342, 310, 270, 223, 223, 285, 342, 36, 
    532, 389, 392, 381, 339, 327, 260, 124, 189, 307, 325, 324, 289, 267, 276, 274, 270, 264, 254, 263, 267, 288, 348, 379, 345, 307, 281, 240, 214, 244, 322, 42, 
    531, 389, 393, 372, 322, 320, 260, 125, 196, 314, 321, 357, 326, 261, 261, 263, 270, 276, 267, 290, 288, 269, 305, 342, 335, 326, 310, 270, 220, 230, 294, 30, 
    530, 390, 392, 369, 313, 297, 238, 132, 199, 284, 246, 280, 278, 227, 239, 258, 267, 281, 263, 284, 302, 252, 298, 364, 357, 353, 347, 289, 233, 243, 295, 25, 
    525, 391, 391, 364, 272, 229, 201, 123, 204, 267, 229, 245, 251, 220, 233, 251, 259, 268, 254, 274, 309, 277, 294, 365, 389, 399, 389, 338, 317, 335, 363, 53, 
    506, 392, 395, 357, 253, 208, 165, 103, 158, 217, 212, 211, 210, 203, 213, 222, 226, 224, 222, 239, 279, 277, 271, 315, 369, 407, 399, 381, 383, 403, 406, 59, 
    478, 381, 383, 333, 260, 252, 206, 98, 95, 156, 184, 198, 199, 184, 182, 187, 187, 184, 199, 212, 214, 224, 234, 273, 352, 401, 402, 391, 392, 392, 392, 45, 
    447, 359, 350, 286, 237, 246, 202, 115, 122, 161, 195, 216, 229, 201, 166, 162, 174, 194, 227, 229, 185, 173, 192, 242, 328, 381, 381, 389, 402, 394, 391, 45, 
    432, 339, 295, 238, 209, 212, 188, 154, 167, 214, 233, 217, 227, 203, 174, 168, 184, 210, 239, 231, 178, 154, 168, 205, 258, 283, 286, 329, 399, 410, 391, 45, 
    442, 323, 233, 176, 200, 240, 245, 184, 160, 189, 173, 138, 150, 146, 133, 132, 144, 151, 145, 125, 96, 103, 130, 150, 176, 202, 219, 265, 369, 419, 399, 45, 
    426, 294, 177, 102, 173, 265, 287, 189, 139, 149, 142, 105, 86, 83, 89, 67, 53, 62, 58, 64, 71, 53, 56, 77, 102, 158, 189, 224, 347, 424, 404, 45, 
    413, 273, 154, 90, 188, 267, 215, 113, 119, 168, 174, 190, 185, 168, 156, 84, 59, 70, 56, 94, 133, 72, 39, 45, 73, 155, 215, 245, 324, 413, 417, 46, 
    430, 291, 183, 120, 223, 257, 105, 27, 115, 186, 177, 186, 205, 224, 198, 164, 194, 205, 199, 247, 277, 219, 189, 191, 215, 263, 251, 238, 286, 394, 432, 51, 
    446, 293, 170, 86, 199, 218, 52, 3, 121, 164, 136, 109, 113, 137, 165, 225, 267, 237, 231, 265, 278, 228, 220, 241, 282, 296, 198, 158, 210, 343, 433, 57, 
    451, 300, 170, 54, 137, 168, 57, 23, 97, 118, 103, 78, 75, 91, 113, 183, 248, 194, 158, 177, 179, 163, 162, 166, 206, 208, 127, 100, 168, 331, 448, 65, 
    447, 313, 189, 57, 85, 111, 68, 44, 52, 62, 79, 90, 101, 114, 110, 124, 158, 152, 159, 162, 156, 140, 157, 174, 161, 165, 140, 143, 184, 319, 449, 71, 
    441, 314, 193, 74, 109, 114, 77, 66, 33, 22, 41, 77, 128, 177, 142, 48, 92, 170, 155, 108, 117, 119, 157, 208, 116, 64, 166, 206, 179, 300, 446, 74, 
    436, 314, 180, 50, 115, 143, 119, 104, 50, 12, 21, 56, 108, 181, 149, 37, 75, 211, 223, 169, 187, 184, 224, 288, 141, 56, 157, 181, 149, 283, 443, 76, 
    427, 307, 162, 9, 71, 139, 181, 176, 79, 24, 12, 21, 46, 72, 57, 0, 47, 161, 194, 181, 207, 211, 220, 217, 86, 24, 91, 91, 81, 260, 438, 81, 
    406, 294, 184, 48, 65, 145, 205, 201, 102, 39, 15, 1, 5, 13, 12, 0, 19, 83, 183, 229, 241, 227, 217, 150, 6, 0, 53, 68, 105, 277, 425, 78, 
    385, 294, 256, 174, 152, 176, 237, 192, 94, 74, 39, 0, 0, 0, 7, 19, 18, 58, 224, 344, 345, 317, 298, 175, 21, 4, 37, 83, 143, 285, 411, 75, 
    374, 301, 295, 255, 215, 189, 225, 182, 98, 111, 65, 6, 0, 0, 5, 27, 50, 88, 202, 277, 262, 260, 254, 132, 0, 0, 34, 99, 159, 279, 397, 77, 
    379, 297, 286, 256, 210, 166, 187, 160, 106, 120, 77, 15, 0, 11, 22, 42, 72, 105, 161, 187, 178, 209, 229, 106, 0, 0, 45, 107, 157, 274, 388, 72, 
    377, 285, 265, 239, 219, 175, 148, 120, 98, 112, 76, 32, 16, 25, 36, 46, 61, 78, 97, 124, 157, 199, 223, 118, 0, 0, 46, 97, 149, 281, 383, 67, 
    357, 262, 253, 247, 239, 187, 106, 83, 96, 102, 69, 46, 37, 40, 51, 55, 58, 72, 91, 106, 127, 152, 170, 110, 3, 0, 46, 92, 170, 306, 372, 59, 
    348, 268, 273, 266, 254, 209, 103, 52, 82, 85, 72, 66, 60, 69, 80, 79, 81, 99, 119, 123, 130, 141, 145, 115, 44, 28, 62, 127, 232, 335, 369, 55, 
    187, 166, 173, 171, 161, 132, 57, 22, 27, 22, 19, 27, 35, 40, 48, 47, 46, 59, 76, 82, 85, 88, 87, 71, 38, 24, 45, 88, 155, 213, 215, 25, 
    
    -- channel=158
    74, 37, 33, 38, 44, 32, 24, 34, 31, 13, 11, 14, 10, 3, 0, 10, 24, 38, 45, 42, 40, 46, 53, 45, 29, 21, 28, 44, 27, 24, 21, 0, 
    231, 199, 193, 192, 201, 188, 161, 165, 175, 156, 151, 156, 159, 161, 157, 167, 192, 205, 221, 225, 216, 216, 227, 222, 201, 177, 175, 196, 186, 162, 158, 0, 
    242, 210, 207, 205, 209, 198, 145, 141, 163, 155, 168, 165, 177, 201, 211, 224, 236, 227, 236, 238, 233, 224, 225, 229, 224, 211, 206, 210, 208, 187, 183, 10, 
    258, 224, 223, 223, 225, 209, 145, 127, 139, 125, 138, 136, 132, 154, 173, 189, 210, 213, 228, 239, 226, 218, 220, 222, 230, 230, 219, 213, 219, 221, 206, 10, 
    266, 231, 231, 231, 228, 207, 121, 77, 93, 74, 68, 75, 61, 62, 73, 79, 109, 132, 152, 197, 214, 203, 214, 217, 218, 227, 220, 204, 223, 245, 228, 12, 
    266, 231, 231, 231, 224, 206, 110, 17, 38, 34, 24, 23, 16, 19, 16, 6, 15, 30, 46, 89, 165, 210, 218, 219, 207, 210, 211, 187, 203, 240, 245, 26, 
    266, 231, 232, 226, 213, 209, 129, 24, 39, 55, 50, 48, 29, 41, 50, 36, 27, 17, 23, 38, 83, 187, 245, 234, 214, 203, 187, 168, 164, 207, 249, 41, 
    265, 230, 232, 220, 194, 193, 130, 48, 61, 102, 122, 141, 95, 72, 77, 70, 69, 60, 52, 70, 71, 119, 207, 238, 221, 200, 181, 169, 162, 178, 227, 46, 
    266, 231, 232, 218, 181, 181, 128, 47, 63, 95, 110, 153, 131, 80, 66, 65, 71, 79, 64, 89, 91, 81, 147, 207, 205, 202, 199, 171, 154, 146, 178, 18, 
    267, 233, 232, 214, 169, 171, 110, 41, 59, 76, 59, 88, 100, 73, 58, 62, 69, 80, 74, 86, 98, 83, 122, 194, 220, 223, 212, 177, 145, 146, 169, 0, 
    269, 238, 234, 210, 146, 110, 56, 25, 56, 91, 63, 57, 64, 59, 52, 56, 64, 72, 74, 83, 102, 97, 110, 178, 235, 240, 227, 210, 196, 201, 210, 11, 
    257, 240, 235, 209, 152, 105, 38, 2, 23, 61, 56, 40, 27, 33, 43, 48, 51, 51, 53, 58, 80, 104, 108, 137, 196, 232, 235, 230, 231, 232, 232, 21, 
    232, 233, 226, 199, 165, 151, 79, 12, 0, 0, 28, 35, 24, 6, 14, 24, 23, 19, 27, 33, 42, 73, 95, 121, 186, 239, 251, 246, 236, 231, 232, 21, 
    212, 203, 196, 174, 142, 144, 103, 38, 0, 12, 26, 40, 50, 27, 9, 15, 26, 39, 62, 73, 54, 54, 81, 118, 171, 209, 225, 251, 256, 235, 231, 21, 
    205, 179, 161, 155, 139, 123, 97, 50, 39, 44, 42, 51, 66, 62, 33, 27, 40, 52, 65, 70, 53, 47, 57, 81, 114, 142, 153, 190, 253, 248, 231, 21, 
    214, 187, 123, 110, 130, 141, 131, 81, 41, 41, 16, 1, 0, 9, 9, 9, 27, 35, 32, 30, 14, 16, 39, 49, 70, 77, 74, 104, 202, 247, 234, 21, 
    196, 162, 84, 58, 93, 145, 150, 109, 44, 33, 15, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 36, 54, 143, 235, 238, 20, 
    184, 149, 86, 58, 98, 125, 100, 73, 53, 43, 49, 84, 76, 52, 27, 6, 0, 0, 0, 8, 32, 0, 0, 0, 0, 24, 53, 78, 138, 230, 245, 21, 
    202, 157, 87, 60, 118, 120, 43, 10, 44, 65, 55, 72, 90, 97, 85, 71, 66, 78, 92, 109, 123, 102, 84, 84, 100, 91, 78, 97, 123, 206, 246, 23, 
    212, 160, 74, 36, 102, 118, 29, 0, 26, 58, 32, 12, 23, 45, 58, 105, 124, 85, 79, 95, 102, 93, 92, 91, 114, 119, 62, 45, 76, 176, 238, 24, 
    215, 172, 81, 14, 40, 79, 33, 0, 5, 28, 32, 14, 0, 0, 9, 63, 105, 75, 49, 58, 63, 54, 58, 51, 70, 94, 45, 6, 37, 161, 236, 24, 
    208, 176, 93, 30, 18, 21, 30, 5, 0, 0, 19, 29, 16, 13, 0, 0, 57, 68, 29, 22, 28, 18, 39, 40, 1, 41, 61, 29, 37, 153, 235, 26, 
    197, 167, 92, 44, 63, 30, 14, 2, 0, 0, 0, 19, 53, 80, 45, 0, 22, 78, 50, 22, 25, 16, 51, 82, 11, 7, 78, 92, 67, 145, 226, 26, 
    192, 154, 75, 20, 62, 78, 37, 9, 0, 0, 0, 2, 35, 77, 72, 5, 12, 101, 128, 85, 81, 71, 87, 127, 74, 10, 51, 74, 55, 134, 215, 24, 
    178, 136, 61, 0, 0, 51, 79, 51, 10, 0, 0, 0, 0, 9, 16, 0, 2, 58, 101, 70, 61, 58, 66, 48, 22, 7, 16, 18, 20, 118, 202, 20, 
    165, 127, 73, 0, 0, 26, 91, 68, 23, 0, 0, 0, 0, 0, 0, 0, 0, 9, 88, 120, 114, 107, 99, 36, 0, 0, 11, 11, 21, 109, 181, 12, 
    155, 122, 109, 72, 37, 41, 89, 59, 28, 14, 0, 0, 0, 0, 0, 0, 0, 0, 95, 181, 187, 168, 146, 72, 0, 0, 2, 20, 37, 107, 166, 6, 
    146, 123, 129, 115, 77, 47, 82, 66, 35, 30, 7, 0, 0, 0, 0, 0, 9, 27, 73, 119, 128, 128, 120, 44, 0, 0, 0, 25, 47, 106, 157, 2, 
    149, 120, 113, 100, 81, 52, 60, 63, 39, 30, 14, 0, 0, 0, 0, 0, 14, 31, 45, 58, 71, 93, 104, 37, 0, 0, 4, 25, 49, 103, 149, 0, 
    146, 106, 95, 87, 78, 51, 32, 40, 37, 26, 14, 2, 0, 0, 0, 0, 0, 9, 19, 30, 49, 70, 86, 47, 0, 0, 3, 20, 45, 96, 141, 0, 
    132, 91, 85, 79, 75, 53, 6, 11, 33, 30, 16, 4, 0, 0, 0, 0, 0, 4, 8, 11, 22, 34, 47, 33, 0, 0, 0, 19, 46, 102, 138, 0, 
    181, 160, 164, 161, 155, 131, 70, 30, 44, 45, 42, 42, 41, 41, 44, 43, 43, 54, 67, 69, 72, 78, 82, 74, 46, 24, 33, 70, 129, 188, 210, 80, 
    
    -- channel=159
    77, 0, 0, 1, 6, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 6, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    186, 121, 115, 109, 126, 125, 106, 105, 116, 110, 105, 109, 101, 94, 87, 86, 93, 106, 122, 124, 121, 118, 129, 135, 123, 103, 93, 100, 96, 84, 92, 15, 
    195, 126, 126, 123, 127, 126, 101, 92, 110, 116, 119, 122, 124, 133, 141, 136, 140, 140, 136, 133, 127, 124, 131, 140, 138, 126, 114, 104, 111, 107, 108, 31, 
    206, 136, 136, 136, 136, 135, 101, 82, 105, 101, 108, 119, 106, 119, 134, 136, 148, 150, 140, 136, 121, 124, 134, 139, 138, 137, 127, 110, 116, 123, 117, 36, 
    211, 144, 144, 144, 142, 129, 89, 62, 95, 92, 80, 95, 79, 79, 90, 91, 108, 122, 124, 142, 125, 115, 135, 139, 134, 139, 126, 108, 111, 129, 132, 39, 
    211, 144, 144, 145, 143, 134, 85, 25, 53, 76, 55, 60, 59, 54, 53, 44, 49, 67, 71, 92, 125, 125, 128, 142, 133, 129, 124, 108, 105, 128, 141, 46, 
    211, 144, 145, 142, 136, 137, 114, 38, 34, 72, 65, 59, 53, 61, 63, 52, 45, 45, 53, 52, 77, 128, 141, 149, 138, 121, 116, 103, 90, 112, 141, 56, 
    211, 143, 145, 139, 125, 129, 115, 57, 54, 102, 99, 101, 76, 60, 77, 77, 76, 67, 64, 81, 67, 78, 136, 158, 143, 133, 120, 104, 83, 90, 134, 65, 
    211, 144, 144, 139, 123, 121, 100, 57, 61, 101, 107, 135, 121, 77, 72, 76, 78, 82, 70, 81, 96, 76, 97, 139, 145, 137, 124, 103, 93, 97, 116, 59, 
    212, 146, 145, 139, 118, 108, 104, 61, 64, 87, 68, 87, 105, 79, 68, 74, 76, 85, 78, 77, 96, 88, 95, 136, 144, 135, 136, 116, 100, 103, 106, 32, 
    214, 152, 148, 135, 96, 89, 87, 55, 60, 89, 73, 68, 81, 77, 70, 73, 76, 79, 82, 83, 96, 98, 94, 127, 156, 159, 149, 140, 124, 121, 127, 35, 
    210, 162, 153, 137, 109, 77, 56, 31, 34, 78, 86, 68, 65, 62, 64, 65, 67, 67, 71, 74, 82, 94, 92, 104, 149, 163, 152, 143, 145, 145, 145, 51, 
    197, 162, 155, 136, 123, 113, 83, 28, 23, 48, 65, 68, 60, 45, 45, 53, 58, 60, 64, 59, 47, 63, 88, 100, 127, 151, 156, 150, 148, 145, 144, 51, 
    183, 151, 147, 130, 115, 118, 101, 65, 47, 40, 46, 59, 77, 61, 40, 48, 61, 66, 71, 70, 50, 49, 73, 90, 119, 146, 159, 166, 164, 150, 144, 51, 
    185, 139, 126, 119, 114, 107, 101, 70, 55, 68, 63, 56, 71, 79, 64, 54, 58, 66, 75, 87, 82, 67, 68, 81, 102, 118, 123, 145, 180, 166, 145, 51, 
    189, 138, 108, 96, 124, 132, 121, 64, 48, 59, 51, 45, 46, 59, 58, 46, 44, 52, 51, 52, 55, 50, 51, 58, 68, 91, 105, 104, 157, 179, 151, 50, 
    181, 145, 103, 60, 95, 129, 130, 89, 57, 59, 58, 45, 24, 18, 27, 11, 14, 32, 29, 36, 36, 7, 15, 31, 46, 72, 75, 75, 120, 170, 158, 51, 
    181, 127, 88, 50, 82, 109, 90, 71, 77, 73, 65, 79, 71, 52, 47, 31, 29, 27, 17, 27, 44, 9, 0, 11, 12, 38, 61, 74, 98, 157, 169, 53, 
    185, 117, 88, 59, 102, 109, 57, 27, 69, 82, 61, 66, 97, 95, 85, 85, 83, 64, 70, 75, 96, 92, 67, 65, 65, 68, 63, 77, 108, 158, 180, 57, 
    191, 121, 79, 39, 86, 110, 59, 15, 37, 71, 69, 42, 45, 60, 91, 102, 106, 86, 89, 105, 105, 97, 96, 99, 116, 113, 67, 61, 91, 136, 176, 60, 
    193, 131, 82, 22, 50, 91, 66, 25, 23, 48, 64, 43, 33, 37, 41, 63, 113, 92, 62, 63, 72, 69, 67, 72, 68, 91, 74, 44, 61, 118, 172, 63, 
    189, 136, 95, 33, 29, 52, 52, 34, 22, 20, 43, 55, 55, 44, 32, 18, 57, 85, 68, 53, 60, 58, 64, 68, 44, 59, 89, 67, 48, 103, 174, 68, 
    185, 130, 91, 44, 62, 47, 38, 42, 21, 6, 20, 42, 66, 77, 52, 3, 35, 88, 66, 31, 43, 44, 53, 84, 24, 5, 80, 87, 59, 107, 176, 69, 
    184, 124, 85, 23, 65, 88, 58, 48, 18, 2, 14, 17, 44, 76, 89, 40, 34, 92, 108, 74, 71, 71, 73, 104, 73, 18, 49, 81, 81, 116, 172, 68, 
    177, 121, 80, 14, 20, 81, 93, 65, 30, 12, 10, 12, 18, 27, 50, 41, 25, 50, 105, 96, 75, 79, 66, 64, 63, 35, 33, 43, 54, 101, 163, 69, 
    162, 115, 96, 34, 12, 34, 75, 82, 49, 27, 9, 5, 11, 16, 17, 21, 19, 35, 91, 105, 73, 65, 71, 38, 0, 14, 36, 43, 51, 88, 150, 68, 
    152, 112, 115, 81, 43, 44, 73, 78, 47, 47, 21, 0, 5, 15, 17, 21, 23, 26, 78, 136, 130, 123, 112, 77, 10, 9, 33, 49, 58, 89, 142, 63, 
    152, 108, 106, 103, 83, 65, 77, 76, 45, 53, 37, 12, 4, 12, 15, 23, 37, 36, 52, 100, 120, 123, 111, 71, 13, 13, 26, 45, 62, 92, 139, 61, 
    150, 104, 102, 97, 86, 63, 60, 74, 51, 52, 44, 23, 11, 16, 20, 23, 34, 50, 61, 72, 82, 94, 103, 63, 4, 12, 28, 44, 61, 94, 135, 55, 
    148, 101, 98, 90, 83, 69, 44, 52, 54, 48, 41, 31, 20, 20, 25, 26, 28, 34, 43, 53, 65, 78, 92, 81, 14, 5, 28, 41, 60, 97, 127, 50, 
    142, 90, 89, 86, 85, 67, 34, 29, 49, 47, 37, 36, 29, 24, 28, 28, 27, 32, 38, 41, 47, 57, 65, 67, 28, 5, 22, 41, 66, 94, 114, 44, 
    132, 107, 106, 100, 97, 92, 53, 25, 41, 49, 49, 43, 41, 40, 41, 40, 42, 49, 55, 54, 55, 60, 62, 61, 48, 26, 28, 57, 83, 108, 128, 62, 
    
    
    others => 0);
end gold_package;
