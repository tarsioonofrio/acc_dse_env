LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
	PACKAGE inmem_package is
		type padroes is array(0 to 4000000) of integer;

		constant input_mem: padroes := ( 
					-- bias

					-- weights

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			90, 65, 72, 94, 62, 25, 71, 
			36, 94, 52, 18, 45, 3, 58, 
			0, 38, 0, 0, 0, 0, 25, 
			0, 14, 0, 7, 14, 11, 59, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 14, 0, 0, 0, 3, 0, 
			0, 0, 0, 23, 0, 28, 75, 
			108, 0, 0, 147, 0, 103, 87, 
			156, 48, 0, 17, 0, 110, 0, 
			116, 0, 0, 71, 0, 0, 0, 
			0, 0, 0, 0, 12, 0, 0, 
			74, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 63, 
			0, 9, 0, 0, 0, 45, 34, 
			0, 0, 0, 0, 0, 61, 0, 
			0, 0, 23, 3, 0, 96, 26, 
			0, 0, 0, 0, 50, 42, 39, 
			0, 14, 0, 7, 0, 0, 0, 
			

			57, 34, 30, 86, 84, 110, 63, 
			87, 59, 38, 110, 79, 78, 54, 
			81, 45, 0, 87, 68, 103, 85, 
			98, 129, 67, 84, 0, 59, 51, 
			35, 98, 49, 49, 124, 55, 60, 
			69, 0, 79, 45, 89, 74, 90, 
			70, 105, 99, 82, 68, 74, 58, 
			

			0, 0, 0, 108, 104, 117, 51, 
			106, 1, 84, 0, 0, 0, 84, 
			0, 99, 0, 0, 0, 0, 0, 
			0, 51, 0, 0, 0, 0, 0, 
			0, 0, 110, 0, 101, 99, 59, 
			14, 0, 208, 105, 20, 0, 0, 
			64, 55, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 23, 0, 0, 
			49, 0, 0, 3, 149, 58, 0, 
			117, 0, 0, 2, 31, 47, 0, 
			31, 220, 112, 51, 60, 0, 0, 
			142, 152, 169, 54, 103, 102, 131, 
			100, 163, 111, 77, 67, 98, 99, 
			

			123, 154, 13, 39, 0, 0, 56, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 6, 0, 0, 39, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 4, 0, 0, 0, 
			

			19, 0, 0, 161, 0, 58, 65, 
			117, 9, 5, 58, 0, 162, 32, 
			246, 0, 0, 169, 0, 200, 0, 
			154, 84, 0, 225, 0, 131, 9, 
			46, 139, 68, 0, 202, 40, 0, 
			38, 0, 271, 42, 0, 0, 0, 
			0, 28, 5, 0, 0, 0, 0, 
			

			0, 0, 9, 0, 27, 0, 0, 
			0, 24, 13, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 56, 
			65, 38, 98, 0, 0, 0, 0, 
			0, 0, 0, 63, 25, 13, 46, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 134, 0, 0, 0, 0, 0, 
			

			0, 23, 7, 78, 29, 86, 21, 
			84, 4, 96, 112, 36, 140, 102, 
			107, 118, 0, 163, 24, 129, 84, 
			62, 115, 12, 124, 95, 62, 52, 
			20, 38, 93, 0, 114, 50, 3, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 52, 0, 0, 0, 0, 0, 
			0, 0, 46, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			101, 90, 82, 78, 13, 0, 100, 
			121, 121, 65, 0, 72, 4, 15, 
			1, 166, 32, 0, 108, 0, 0, 
			0, 16, 74, 11, 73, 0, 39, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 155, 0, 0, 
			0, 0, 164, 0, 12, 0, 0, 
			20, 0, 0, 134, 5, 0, 5, 
			0, 347, 0, 0, 0, 0, 0, 
			0, 123, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 18, 0, 
			0, 0, 0, 51, 0, 4, 31, 
			13, 0, 0, 0, 0, 0, 0, 
			0, 120, 49, 0, 0, 0, 0, 
			0, 0, 0, 0, 32, 34, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 20, 0, 
			26, 0, 0, 0, 0, 52, 0, 
			0, 0, 29, 24, 55, 118, 0, 
			68, 0, 202, 212, 223, 200, 209, 
			153, 363, 221, 150, 174, 163, 216, 
			

			6, 22, 29, 0, 78, 0, 0, 
			0, 82, 0, 0, 163, 0, 0, 
			0, 101, 84, 0, 169, 0, 0, 
			0, 0, 141, 0, 61, 0, 24, 
			0, 0, 0, 0, 0, 0, 46, 
			64, 85, 0, 0, 0, 89, 39, 
			39, 0, 0, 12, 102, 89, 85, 
			

			0, 0, 0, 0, 0, 12, 0, 
			0, 0, 0, 15, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 16, 33, 55, 87, 26, 
			63, 0, 184, 132, 208, 230, 246, 
			191, 69, 197, 171, 180, 190, 181, 
			

			67, 87, 0, 62, 0, 5, 50, 
			0, 0, 0, 56, 0, 44, 187, 
			15, 253, 0, 26, 2, 176, 5, 
			0, 89, 0, 23, 104, 200, 7, 
			0, 0, 0, 0, 35, 0, 0, 
			22, 0, 0, 0, 0, 0, 0, 
			115, 0, 0, 1, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			101, 0, 0, 28, 0, 0, 25, 
			73, 0, 0, 0, 19, 38, 0, 
			

			85, 70, 33, 168, 0, 32, 47, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 20, 0, 0, 
			0, 0, 120, 111, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			107, 45, 106, 147, 23, 0, 79, 
			0, 55, 0, 0, 28, 0, 0, 
			0, 8, 46, 0, 0, 4, 0, 
			0, 0, 83, 19, 0, 29, 38, 
			0, 0, 0, 0, 84, 0, 36, 
			90, 0, 136, 14, 0, 0, 0, 
			0, 89, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 53, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			39, 44, 0, 0, 47, 23, 51, 
			0, 0, 0, 0, 0, 0, 10, 
			0, 0, 0, 0, 0, 0, 22, 
			0, 0, 0, 0, 0, 0, 26, 
			0, 0, 0, 0, 0, 0, 49, 
			0, 0, 0, 0, 80, 201, 201, 
			196, 0, 53, 167, 208, 198, 145, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 33, 0, 0, 10, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 132, 0, 0, 2, 0, 
			0, 0, 0, 0, 0, 36, 55, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 21, 0, 0, 0, 0, 
			0, 0, 8, 11, 0, 0, 0, 
			53, 0, 0, 0, 0, 0, 0, 
			110, 138, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 6, 2, 52, 
			

			3, 0, 84, 43, 137, 19, 66, 
			278, 113, 84, 0, 293, 49, 0, 
			145, 0, 0, 0, 582, 0, 0, 
			0, 0, 191, 41, 400, 0, 54, 
			227, 417, 0, 0, 0, 0, 74, 
			39, 447, 0, 0, 0, 0, 0, 
			0, 0, 119, 0, 0, 0, 0, 
			

			117, 145, 38, 0, 34, 0, 72, 
			162, 199, 0, 0, 38, 0, 0, 
			0, 0, 0, 0, 100, 0, 0, 
			0, 18, 0, 0, 0, 0, 17, 
			0, 105, 0, 0, 0, 0, 34, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			33, 15, 41, 46, 31, 19, 28, 
			25, 52, 96, 61, 14, 21, 8, 
			0, 18, 64, 17, 0, 39, 0, 
			0, 58, 8, 0, 0, 24, 0, 
			0, 0, 63, 0, 26, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 77, 0, 
			53, 0, 92, 121, 0, 106, 21, 
			113, 0, 0, 285, 0, 135, 53, 
			252, 95, 0, 0, 0, 38, 0, 
			157, 112, 130, 51, 28, 0, 0, 
			0, 0, 107, 0, 26, 0, 14, 
			0, 0, 11, 39, 25, 0, 50, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 33, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 53, 0, 0, 0, 81, 0, 
			0, 0, 0, 0, 36, 50, 0, 
			0, 0, 39, 53, 47, 62, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 131, 0, 0, 0, 0, 
			125, 0, 0, 0, 0, 0, 0, 
			

			58, 48, 67, 86, 65, 63, 63, 
			92, 107, 103, 125, 126, 117, 58, 
			61, 138, 84, 155, 236, 112, 46, 
			63, 122, 141, 114, 127, 74, 37, 
			110, 174, 86, 52, 102, 43, 35, 
			0, 192, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 30, 
			68, 0, 0, 73, 92, 0, 123, 
			0, 133, 0, 0, 312, 97, 0, 
			0, 120, 0, 0, 78, 14, 0, 
			0, 32, 93, 0, 5, 59, 0, 
			0, 0, 40, 0, 110, 59, 47, 
			206, 0, 83, 24, 28, 45, 4, 
			

			0, 45, 0, 0, 0, 0, 0, 
			0, 0, 0, 19, 0, 42, 0, 
			8, 0, 0, 75, 0, 25, 0, 
			59, 0, 0, 0, 0, 0, 0, 
			0, 50, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 124, 64, 88, 
			0, 0, 86, 140, 121, 86, 59, 
			

			133, 114, 126, 117, 92, 69, 120, 
			156, 172, 131, 99, 148, 118, 65, 
			127, 92, 143, 118, 193, 118, 90, 
			69, 133, 78, 98, 111, 57, 102, 
			61, 208, 120, 21, 59, 11, 57, 
			21, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 52, 40, 0, 
			61, 0, 0, 56, 169, 18, 78, 
			161, 49, 30, 19, 50, 0, 5, 
			169, 146, 62, 83, 51, 20, 37, 
			102, 197, 0, 15, 51, 84, 101, 
			118, 0, 24, 94, 114, 139, 190, 
			

			29, 0, 58, 0, 0, 0, 1, 
			224, 77, 23, 0, 164, 0, 0, 
			149, 89, 0, 0, 411, 0, 0, 
			0, 0, 66, 0, 244, 0, 0, 
			132, 402, 61, 0, 0, 0, 0, 
			0, 421, 0, 0, 0, 0, 0, 
			0, 0, 89, 0, 0, 0, 0, 
			

			0, 0, 18, 115, 113, 102, 62, 
			20, 45, 82, 86, 74, 51, 7, 
			84, 129, 128, 0, 11, 24, 25, 
			4, 55, 62, 43, 11, 18, 22, 
			0, 15, 135, 57, 187, 105, 154, 
			25, 141, 223, 68, 126, 103, 106, 
			0, 0, 0, 0, 0, 0, 0, 
			

			53, 77, 22, 0, 0, 0, 37, 
			53, 72, 0, 3, 40, 40, 29, 
			75, 0, 54, 56, 77, 97, 68, 
			91, 84, 0, 19, 0, 0, 57, 
			30, 153, 42, 74, 0, 0, 1, 
			6, 0, 0, 0, 0, 76, 2, 
			0, 0, 0, 42, 51, 40, 10, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 81, 0, 0, 0, 0, 
			0, 0, 92, 73, 0, 0, 36, 
			154, 0, 0, 0, 0, 0, 0, 
			39, 18, 0, 225, 0, 43, 50, 
			0, 329, 65, 114, 102, 124, 92, 
			

			65, 0, 32, 160, 135, 133, 164, 
			43, 34, 0, 0, 0, 0, 37, 
			53, 31, 0, 0, 0, 0, 0, 
			0, 138, 43, 0, 0, 0, 0, 
			0, 0, 0, 4, 73, 48, 217, 
			192, 0, 86, 123, 61, 28, 74, 
			129, 60, 28, 0, 0, 0, 0, 
			

			24, 39, 0, 0, 0, 0, 4, 
			0, 0, 0, 59, 0, 93, 36, 
			0, 0, 0, 101, 0, 100, 24, 
			24, 0, 0, 126, 0, 145, 0, 
			81, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 25, 37, 0, 0, 
			0, 0, 152, 81, 67, 27, 32, 
			

			68, 70, 0, 167, 112, 0, 47, 
			0, 156, 29, 0, 56, 27, 0, 
			0, 0, 55, 0, 0, 147, 34, 
			0, 59, 0, 120, 0, 29, 33, 
			0, 0, 69, 0, 149, 146, 0, 
			150, 0, 126, 166, 0, 0, 33, 
			0, 328, 0, 21, 0, 92, 0, 
			

			0, 0, 0, 0, 118, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 64, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 47, 0, 192, 0, 
			0, 137, 0, 0, 142, 0, 0, 
			0, 0, 63, 0, 0, 0, 80, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			173, 190, 121, 0, 0, 0, 55, 
			0, 149, 0, 0, 40, 0, 0, 
			0, 21, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 31, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 25, 
			0, 0, 0, 0, 0, 0, 0, 
			78, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 82, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 20, 0, 0, 
			0, 0, 0, 0, 34, 0, 0, 
			0, 0, 109, 14, 0, 8, 61, 
			117, 113, 0, 99, 72, 158, 143, 
			164, 0, 55, 72, 117, 106, 140, 
			

			167, 190, 183, 219, 204, 128, 122, 
			96, 212, 181, 2, 17, 0, 0, 
			0, 0, 27, 0, 14, 0, 22, 
			54, 91, 0, 0, 0, 0, 0, 
			0, 51, 92, 45, 119, 173, 239, 
			0, 0, 32, 113, 73, 94, 114, 
			34, 0, 0, 12, 29, 0, 1, 
			

			101, 121, 133, 115, 80, 41, 67, 
			0, 113, 100, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 21, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			16, 0, 64, 0, 60, 0, 0, 
			0, 54, 0, 12, 0, 0, 0, 
			65, 0, 287, 178, 0, 0, 145, 
			159, 23, 0, 0, 0, 111, 14, 
			146, 152, 0, 209, 0, 0, 0, 
			0, 0, 270, 0, 195, 66, 129, 
			79, 9, 178, 107, 71, 9, 0, 
			

			65, 60, 104, 48, 70, 86, 66, 
			105, 137, 114, 108, 102, 33, 51, 
			7, 0, 0, 120, 120, 48, 120, 
			74, 164, 21, 0, 0, 12, 33, 
			0, 140, 71, 95, 125, 49, 60, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			72, 0, 0, 0, 0, 0, 0, 
			0, 30, 0, 47, 71, 179, 162, 
			73, 0, 75, 169, 209, 219, 275, 
			

			26, 0, 32, 100, 90, 100, 65, 
			88, 4, 136, 28, 18, 0, 58, 
			0, 72, 2, 0, 0, 0, 0, 
			2, 102, 49, 37, 93, 60, 16, 
			0, 0, 61, 0, 75, 78, 53, 
			47, 0, 95, 123, 0, 0, 0, 
			70, 100, 0, 0, 0, 0, 0, 
			

			49, 151, 0, 0, 0, 0, 0, 
			0, 8, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 107, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 35, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			

			0, 0, 23, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 0, 
			0, 0, 0, 0, 0, 0, 52, 
			0, 0, 0, 62, 0, 0, 78, 
			0, 159, 0, 0, 0, 118, 31, 
			0, 0, 0, 0, 73, 0, 81, 
			
