library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    0, 0, 0, 
    0, 314, 59, 
    0, 0, 0, 
    
    -- channel=1
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=2
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 1299, 
    
    -- channel=3
    0, 256, 87, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=4
    0, 0, 516, 
    0, 0, 551, 
    0, 0, 0, 
    
    -- channel=5
    0, 0, 0, 
    0, 0, 0, 
    64, 0, 0, 
    
    -- channel=6
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 339, 
    
    -- channel=7
    0, 0, 0, 
    0, 0, 350, 
    1101, 0, 1304, 
    
    -- channel=8
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=9
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=10
    0, 0, 280, 
    0, 0, 0, 
    422, 273, 119, 
    
    -- channel=11
    0, 0, 213, 
    0, 0, 0, 
    1359, 0, 0, 
    
    -- channel=12
    1048, 48, 1075, 
    1994, 0, 0, 
    0, 240, 573, 
    
    -- channel=13
    1374, 0, 788, 
    702, 0, 0, 
    1924, 1226, 1128, 
    
    -- channel=14
    0, 141, 0, 
    0, 0, 0, 
    0, 0, 177, 
    
    -- channel=15
    1696, 687, 620, 
    1330, 193, 0, 
    509, 724, 1213, 
    
    -- channel=16
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=17
    0, 0, 0, 
    25, 0, 0, 
    8, 0, 522, 
    
    -- channel=18
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=19
    93, 64, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=20
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=21
    0, 0, 111, 
    0, 617, 431, 
    807, 1137, 823, 
    
    -- channel=22
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=23
    0, 0, 0, 
    0, 0, 0, 
    478, 0, 0, 
    
    -- channel=24
    0, 585, 0, 
    111, 0, 0, 
    0, 0, 0, 
    
    -- channel=25
    0, 0, 0, 
    0, 48, 795, 
    0, 0, 0, 
    
    -- channel=26
    0, 0, 0, 
    40, 0, 0, 
    0, 0, 0, 
    
    -- channel=27
    0, 0, 0, 
    0, 0, 0, 
    0, 47, 924, 
    
    -- channel=28
    440, 0, 755, 
    0, 0, 248, 
    1737, 1071, 1744, 
    
    -- channel=29
    376, 815, 0, 
    2137, 289, 584, 
    0, 84, 0, 
    
    -- channel=30
    0, 452, 751, 
    1026, 51, 155, 
    0, 1088, 0, 
    
    -- channel=31
    0, 0, 0, 
    0, 0, 0, 
    566, 0, 190, 
    
    -- channel=32
    43, 262, 0, 
    0, 0, 0, 
    0, 1084, 0, 
    
    -- channel=33
    0, 0, 0, 
    0, 0, 0, 
    197, 0, 0, 
    
    -- channel=34
    405, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=35
    0, 0, 0, 
    0, 0, 0, 
    0, 41, 283, 
    
    -- channel=36
    0, 0, 584, 
    0, 622, 415, 
    1106, 0, 64, 
    
    -- channel=37
    0, 0, 0, 
    0, 0, 0, 
    0, 569, 433, 
    
    -- channel=38
    75, 90, 244, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=39
    0, 245, 0, 
    0, 256, 0, 
    377, 0, 690, 
    
    -- channel=40
    0, 160, 0, 
    0, 0, 0, 
    0, 0, 580, 
    
    -- channel=41
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=42
    0, 728, 158, 
    0, 967, 0, 
    0, 0, 0, 
    
    -- channel=43
    0, 0, 842, 
    0, 0, 910, 
    1006, 1360, 560, 
    
    -- channel=44
    0, 0, 0, 
    0, 0, 0, 
    318, 0, 0, 
    
    -- channel=45
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=46
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=47
    0, 1072, 0, 
    0, 743, 0, 
    8, 207, 0, 
    
    -- channel=48
    0, 0, 0, 
    0, 0, 0, 
    33, 354, 414, 
    
    -- channel=49
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=50
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=51
    0, 0, 0, 
    252, 620, 0, 
    198, 0, 893, 
    
    -- channel=52
    60, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=53
    613, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=54
    0, 0, 0, 
    0, 160, 0, 
    0, 0, 0, 
    
    -- channel=55
    0, 83, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=56
    0, 118, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=57
    0, 0, 0, 
    0, 602, 392, 
    0, 0, 0, 
    
    -- channel=58
    0, 0, 0, 
    0, 0, 793, 
    0, 0, 0, 
    
    -- channel=59
    138, 0, 760, 
    1072, 0, 1201, 
    0, 0, 0, 
    
    -- channel=60
    0, 25, 0, 
    0, 186, 0, 
    0, 0, 0, 
    
    -- channel=61
    0, 0, 230, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=62
    0, 344, 295, 
    0, 0, 0, 
    1036, 1624, 2233, 
    
    -- channel=63
    0, 0, 0, 
    0, 0, 40, 
    0, 0, 232, 
    
    -- channel=64
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=65
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 751, 
    
    -- channel=66
    0, 26, 0, 
    0, 147, 0, 
    0, 0, 0, 
    
    -- channel=67
    1211, 435, 828, 
    1019, 0, 0, 
    0, 0, 0, 
    
    -- channel=68
    0, 0, 0, 
    0, 0, 0, 
    0, 39, 405, 
    
    -- channel=69
    662, 433, 549, 
    606, 0, 0, 
    272, 0, 520, 
    
    -- channel=70
    0, 60, 45, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=71
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=72
    0, 2036, 0, 
    1254, 0, 0, 
    0, 861, 0, 
    
    -- channel=73
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 54, 
    
    -- channel=74
    0, 0, 0, 
    0, 0, 427, 
    0, 0, 0, 
    
    -- channel=75
    137, 152, 0, 
    0, 328, 232, 
    0, 0, 0, 
    
    -- channel=76
    0, 0, 0, 
    0, 0, 0, 
    61, 0, 134, 
    
    -- channel=77
    309, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=78
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=79
    1484, 0, 0, 
    1450, 0, 0, 
    0, 0, 0, 
    
    -- channel=80
    644, 1231, 0, 
    107, 382, 43, 
    0, 121, 0, 
    
    -- channel=81
    0, 0, 0, 
    0, 0, 0, 
    0, 659, 1097, 
    
    -- channel=82
    0, 1045, 821, 
    829, 206, 501, 
    1363, 1493, 1700, 
    
    -- channel=83
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=84
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=85
    0, 0, 0, 
    0, 0, 0, 
    43, 375, 430, 
    
    -- channel=86
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 22, 
    
    -- channel=87
    0, 0, 0, 
    0, 0, 90, 
    1128, 1276, 2430, 
    
    -- channel=88
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=89
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=90
    0, 0, 0, 
    0, 0, 315, 
    0, 0, 0, 
    
    -- channel=91
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=92
    470, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=93
    996, 790, 335, 
    88, 927, 80, 
    642, 0, 0, 
    
    -- channel=94
    0, 21, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=95
    0, 0, 0, 
    0, 790, 4, 
    0, 1751, 0, 
    
    -- channel=96
    474, 243, 0, 
    287, 0, 0, 
    0, 0, 0, 
    
    -- channel=97
    0, 0, 0, 
    0, 0, 0, 
    396, 0, 0, 
    
    -- channel=98
    655, 342, 0, 
    524, 0, 0, 
    0, 0, 0, 
    
    -- channel=99
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 485, 
    
    -- channel=100
    0, 0, 0, 
    0, 0, 0, 
    883, 0, 0, 
    
    -- channel=101
    0, 0, 0, 
    0, 0, 0, 
    0, 1615, 3059, 
    
    -- channel=102
    0, 0, 0, 
    0, 0, 0, 
    75, 232, 0, 
    
    -- channel=103
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=104
    0, 0, 0, 
    0, 0, 0, 
    26, 208, 0, 
    
    -- channel=105
    97, 0, 1, 
    0, 354, 836, 
    1534, 1196, 1070, 
    
    -- channel=106
    10, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=107
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=108
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=109
    286, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=110
    0, 2124, 314, 
    123, 1575, 2794, 
    0, 664, 0, 
    
    -- channel=111
    0, 1595, 718, 
    623, 0, 1287, 
    0, 0, 0, 
    
    -- channel=112
    1011, 0, 0, 
    80, 0, 28, 
    0, 0, 0, 
    
    -- channel=113
    0, 0, 36, 
    0, 361, 319, 
    0, 0, 0, 
    
    -- channel=114
    0, 0, 0, 
    0, 0, 0, 
    0, 461, 502, 
    
    -- channel=115
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=116
    1185, 1064, 0, 
    0, 0, 0, 
    0, 207, 0, 
    
    -- channel=117
    0, 0, 133, 
    0, 0, 0, 
    1669, 2058, 1237, 
    
    -- channel=118
    1417, 1193, 1285, 
    869, 0, 0, 
    2130, 1705, 4234, 
    
    -- channel=119
    0, 0, 0, 
    0, 0, 0, 
    194, 95, 206, 
    
    -- channel=120
    0, 130, 0, 
    0, 0, 97, 
    0, 603, 291, 
    
    -- channel=121
    137, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=122
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=123
    297, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=124
    1199, 947, 371, 
    0, 155, 0, 
    0, 0, 0, 
    
    -- channel=125
    0, 12, 118, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=126
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=127
    369, 1547, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=128
    0, 398, 322, 
    0, 63, 143, 
    0, 0, 0, 
    
    -- channel=129
    0, 0, 0, 
    0, 1042, 685, 
    1633, 830, 341, 
    
    -- channel=130
    0, 0, 0, 
    0, 0, 0, 
    85, 1247, 1433, 
    
    -- channel=131
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=132
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=133
    0, 0, 0, 
    0, 0, 0, 
    876, 0, 0, 
    
    -- channel=134
    684, 798, 404, 
    813, 301, 607, 
    1355, 1492, 1195, 
    
    -- channel=135
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=136
    0, 440, 245, 
    0, 0, 67, 
    0, 0, 0, 
    
    -- channel=137
    0, 258, 1234, 
    0, 0, 161, 
    953, 421, 0, 
    
    -- channel=138
    0, 0, 0, 
    0, 0, 432, 
    0, 0, 0, 
    
    -- channel=139
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=140
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=141
    172, 750, 0, 
    307, 0, 0, 
    0, 0, 0, 
    
    -- channel=142
    0, 0, 198, 
    0, 0, 127, 
    0, 0, 0, 
    
    -- channel=143
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=144
    587, 727, 710, 
    657, 0, 0, 
    132, 840, 1133, 
    
    -- channel=145
    1205, 0, 109, 
    170, 9, 0, 
    0, 0, 0, 
    
    -- channel=146
    1363, 466, 442, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=147
    1413, 1606, 0, 
    426, 0, 0, 
    251, 809, 1917, 
    
    -- channel=148
    0, 1531, 888, 
    0, 59, 0, 
    0, 343, 0, 
    
    -- channel=149
    3, 0, 423, 
    0, 0, 0, 
    1091, 0, 140, 
    
    -- channel=150
    0, 0, 0, 
    143, 0, 0, 
    305, 1082, 994, 
    
    -- channel=151
    0, 0, 772, 
    1367, 303, 187, 
    2551, 3112, 4033, 
    
    -- channel=152
    0, 81, 0, 
    0, 0, 0, 
    966, 1422, 855, 
    
    -- channel=153
    0, 0, 0, 
    0, 0, 0, 
    0, 826, 1220, 
    
    -- channel=154
    0, 0, 0, 
    0, 247, 0, 
    0, 39, 0, 
    
    -- channel=155
    109, 0, 115, 
    0, 0, 0, 
    0, 282, 1270, 
    
    -- channel=156
    0, 880, 288, 
    0, 679, 919, 
    0, 0, 0, 
    
    -- channel=157
    0, 0, 245, 
    0, 0, 0, 
    0, 0, 177, 
    
    -- channel=158
    705, 0, 644, 
    93, 0, 17, 
    0, 0, 0, 
    
    -- channel=159
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=160
    509, 18, 0, 
    1226, 196, 140, 
    0, 0, 42, 
    
    -- channel=161
    223, 275, 0, 
    0, 0, 0, 
    62, 649, 492, 
    
    -- channel=162
    0, 0, 970, 
    1063, 0, 692, 
    0, 0, 0, 
    
    -- channel=163
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=164
    431, 180, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=165
    59, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=166
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=167
    1155, 0, 301, 
    0, 0, 0, 
    1875, 1168, 2630, 
    
    -- channel=168
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=169
    0, 0, 0, 
    98, 0, 0, 
    847, 0, 13, 
    
    -- channel=170
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=171
    1026, 10, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=172
    2149, 3442, 1490, 
    2624, 908, 167, 
    1607, 3260, 3876, 
    
    -- channel=173
    546, 47, 296, 
    1312, 459, 240, 
    2321, 1356, 883, 
    
    -- channel=174
    40, 123, 4, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=175
    0, 0, 0, 
    0, 0, 0, 
    1141, 953, 1354, 
    
    -- channel=176
    1371, 0, 435, 
    2256, 0, 0, 
    1777, 1663, 1451, 
    
    -- channel=177
    415, 745, 0, 
    963, 1005, 205, 
    0, 0, 0, 
    
    -- channel=178
    278, 0, 0, 
    110, 0, 0, 
    609, 0, 0, 
    
    -- channel=179
    0, 0, 0, 
    0, 0, 0, 
    0, 193, 274, 
    
    -- channel=180
    0, 0, 0, 
    0, 49, 135, 
    0, 0, 0, 
    
    -- channel=181
    438, 96, 226, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=182
    0, 612, 93, 
    0, 0, 647, 
    242, 1103, 0, 
    
    -- channel=183
    0, 0, 0, 
    0, 0, 217, 
    0, 604, 1368, 
    
    -- channel=184
    433, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=185
    262, 140, 0, 
    730, 0, 0, 
    0, 0, 493, 
    
    -- channel=186
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=187
    0, 0, 0, 
    0, 0, 0, 
    280, 902, 1025, 
    
    -- channel=188
    567, 0, 0, 
    0, 0, 0, 
    2384, 132, 0, 
    
    -- channel=189
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=190
    36, 0, 0, 
    0, 0, 0, 
    0, 371, 818, 
    
    -- channel=191
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 644, 
    
    -- channel=192
    0, 0, 0, 
    0, 32, 0, 
    772, 633, 943, 
    
    -- channel=193
    0, 177, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=194
    0, 0, 0, 
    0, 0, 98, 
    0, 203, 179, 
    
    -- channel=195
    0, 0, 0, 
    0, 0, 0, 
    0, 542, 321, 
    
    -- channel=196
    1414, 0, 0, 
    203, 0, 0, 
    16, 311, 492, 
    
    -- channel=197
    0, 160, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=198
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 72, 
    
    -- channel=199
    1542, 11, 232, 
    344, 0, 0, 
    0, 0, 0, 
    
    -- channel=200
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=201
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=202
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=203
    0, 0, 0, 
    0, 0, 0, 
    284, 33, 0, 
    
    -- channel=204
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=205
    0, 0, 0, 
    0, 0, 327, 
    0, 0, 0, 
    
    -- channel=206
    0, 0, 0, 
    0, 0, 0, 
    375, 286, 566, 
    
    -- channel=207
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=208
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 115, 
    
    -- channel=209
    0, 0, 0, 
    0, 0, 0, 
    1606, 1054, 99, 
    
    -- channel=210
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=211
    0, 0, 1052, 
    371, 1326, 0, 
    533, 0, 780, 
    
    -- channel=212
    0, 1673, 708, 
    0, 591, 814, 
    0, 0, 456, 
    
    -- channel=213
    508, 0, 1044, 
    0, 0, 353, 
    0, 0, 0, 
    
    -- channel=214
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=215
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=216
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=217
    0, 0, 0, 
    0, 0, 0, 
    2115, 0, 1158, 
    
    -- channel=218
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=219
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=220
    0, 0, 0, 
    0, 259, 0, 
    0, 0, 0, 
    
    -- channel=221
    0, 0, 246, 
    0, 0, 0, 
    993, 0, 0, 
    
    -- channel=222
    373, 0, 5, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=223
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 121, 
    
    -- channel=224
    0, 0, 368, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=225
    576, 499, 673, 
    855, 32, 314, 
    807, 756, 1267, 
    
    -- channel=226
    0, 0, 0, 
    0, 0, 99, 
    0, 0, 0, 
    
    -- channel=227
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=228
    0, 0, 0, 
    509, 0, 0, 
    696, 1266, 649, 
    
    -- channel=229
    1822, 1556, 236, 
    795, 307, 575, 
    64, 1500, 2053, 
    
    -- channel=230
    124, 0, 0, 
    0, 0, 0, 
    516, 0, 0, 
    
    -- channel=231
    182, 0, 25, 
    0, 0, 0, 
    808, 0, 0, 
    
    -- channel=232
    0, 0, 0, 
    0, 0, 0, 
    0, 232, 609, 
    
    -- channel=233
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=234
    0, 0, 0, 
    0, 0, 0, 
    0, 2, 0, 
    
    -- channel=235
    602, 0, 171, 
    56, 0, 32, 
    0, 0, 0, 
    
    -- channel=236
    144, 0, 359, 
    602, 0, 0, 
    0, 0, 0, 
    
    -- channel=237
    1471, 0, 0, 
    977, 152, 97, 
    0, 0, 0, 
    
    -- channel=238
    0, 0, 0, 
    0, 0, 0, 
    0, 651, 2035, 
    
    -- channel=239
    190, 581, 516, 
    2246, 315, 0, 
    0, 0, 0, 
    
    -- channel=240
    815, 0, 0, 
    0, 0, 0, 
    1161, 350, 0, 
    
    -- channel=241
    0, 0, 0, 
    0, 0, 0, 
    57, 129, 664, 
    
    -- channel=242
    0, 0, 0, 
    553, 0, 0, 
    1222, 3164, 3730, 
    
    -- channel=243
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=244
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 46, 
    
    -- channel=245
    346, 0, 0, 
    1050, 0, 0, 
    791, 624, 1366, 
    
    -- channel=246
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=247
    0, 615, 0, 
    0, 378, 0, 
    0, 0, 0, 
    
    -- channel=248
    0, 145, 0, 
    569, 0, 1016, 
    0, 0, 0, 
    
    -- channel=249
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=250
    0, 0, 0, 
    0, 0, 0, 
    1083, 1598, 2535, 
    
    -- channel=251
    529, 0, 0, 
    39, 0, 0, 
    0, 0, 0, 
    
    -- channel=252
    0, 42, 0, 
    0, 0, 289, 
    0, 0, 0, 
    
    -- channel=253
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=254
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    -- channel=255
    0, 0, 0, 
    0, 0, 0, 
    0, 0, 0, 
    
    
    others => 0);
end gold_package;
