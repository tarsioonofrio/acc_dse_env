library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 4000000) of integer;

  constant input_wght : mem := (
    -- bias
    -- layer=3
    -10672, -3316, -981, 5515, 10964, -10702, 14608, -9602, 7586, -3873,

    -- weights
    -- layer=3 channel=0
    -28, -27, 34, -13, 0, 19, 0, 14, -24, 10, 25, 29, -89, 42, -48, 44, -21, -17, 4, -18, 40, -44, -12, 30, -15, -56, 11, -18, 22, -19, -29, 5, -28, -9, -78, 36, -30, -118, -9, -9, -11, -37, -13, 23, -33, -21, -6, 47, -4, -3, 17, 8, 20, 7, -15, -8, 23, 37, -22, -31, -16, 39, -35, 33, -26, 15, -26, -25, 0, 22, 4, 13, 12, 26, -9, 36, -34, -16, 10, -8, 3, -2, -67, 13, 23, -31, -37, -14, 0, -16, 2, 16, -20, 0, -26, 46, -37, 32, -67, 37, -32, -57, -3, -23, 24, 23, 13, 9, 4, -15, 19, 54, -15, 21, 43, -2, 32, 60, 10, -20, 23, -25, -52, -14, -23, 32, 24, -20, 11, 9, -3, -27, 33, 35, -9, 10, 8, 6, 15, 0, -34, -6, 5, 5, 5, -8, 28, 53, 34, -11, -32, 9, -23, -20, -23, -28, -11, -39, -7, 57, 23, 40, -7, -17, -37, -61, -38, -48, 22, 73, 40, -2, -19, -46, 18, 7, -64, 0, -8, 2, -6, -2, -63, 27, 14, -7, 5, -8, -54, -90, 3, 43, -2, -19, -8, 10, -19, -28, -68, 8, 60, 63, -30, -57, 25, -3, -8, 12, 23, -67, -41, 30, -5, -46, 56, 7, -28, -83, -16, -10, 10, 6, -16, 8, -28, -40, -32, 17, 18, -60, 5, 24, 20, 4, -34, -18, 20, -33, 2, -25, 3, 3, 2, 11, -25, 52, -8, 3, 26, 45, -32, -10, -20, 8, -6, -6, 21, 16, -30, -5, 19, 17, -25, 2, 7, -18, -18, -60, 25, 30, 21, 0, 5, -83, -22, 16, -31, -21, 21, 51, -4, -70, -16, -27, -5, -73, 0, -20, 5, -29, 42, -27, 7, -12, -24, 10, 19, 2, 7, 49, 14, -24, 34, -11, -38, 2, 27, -23, -27, -2, -11, -17, 3, 34, -26, -6, -33, 8, 16, -10, 40, -10, -30, 21, 12, 8, -62, -10, 40, -34, 8, -58, 40, -27, 5, 13, 76, -95, 6, 52, 10, -19, 16, -44, 3, -71, -49, 10, 3, -38, 14, 32, -10, -74, -39, 9, -40, 3, -7, 15, -7, 42, 67, -11, -52, -14, 39, -26, -62, 7, -38, -18, -30, 26, -56, 46, 21, 22, 72, -10, -23, -25, 34, 13, -14, -53, -2, 19, 17, -11, 32, 23, 9, 34, -79, -28, -10, -12, -77, -48, -17, 9, 29, 53, -40, -24, -40, 24, 22, -9, -2, 8, -17, 21, -7, 92, -45, 4, 6, 3, -34, 4, -43, -5, 61, 47, 2, -17, 0, -7, -60, 3, 15, 38, -11, 14, -73, 24, 44, -45, -19, -27, -12, -5, 2, -13, 36, 37, -40, 3, -31, 8, -5, -21, 36, -25, 14, 13, -35, 39, 17, 18, 3, 24, -37, -16, 67, 9, -25, 0, -10, -9, -4, -38, 7, 12, 16, 17, 9, 8, -22, 35, 0, 35, -64, 24, 7, 4, 75, 3, -29, 53, 45, -44, -6, 38, -11, -22, -21, -8, -17, 1, 3, -6, 27, 23, 0, 80, 32, 39, -17, -13, 33, -71, -35, 20, 29, 22, 14, 19, -62, -1, -55, -11, -41, 78, -5, 0, 19, -67, 30, 14, -11, -44, 6, -44, -23, -9, 12, 17, -13, 29, -24, -12, 8, 10, -18, 52, -55, -7, 14, -16, -28, -6, 10, -25, -40, -11, -31, -21, -1, -59, -3, 14, -6, 10, -38, 21, 68, 52, 2, 47, -12, -34, 33, -20,
    -- layer=3 channel=1
    16, -18, 7, -16, -40, -59, -17, -3, -18, 13, -6, -11, 3, -35, 32, -37, 18, 44, -5, 6, -6, -23, -12, 12, 0, -7, -28, 10, -14, -12, -33, 23, -25, -26, 11, 3, 20, 16, 2, 6, 4, 2, -9, 37, -19, -23, -10, -9, -19, -28, 18, 1, 0, -9, 3, -6, -72, -11, -30, 23, -4, -89, 2, 2, -45, -17, -30, -12, -53, -34, -42, 14, 8, -16, -49, -17, 23, 35, 51, -9, 2, -7, -17, 17, -18, 34, 24, -42, 2, 7, -28, 15, 6, 2, -4, -34, 2, -51, 23, -21, -18, 33, -26, 49, 20, -41, 59, 8, 22, -6, 2, -35, -24, -13, -1, 16, -61, 5, 19, 14, -7, 3, 4, -8, -34, -47, 29, 48, 19, -25, 6, 15, -45, -1, 14, -20, -15, -24, -13, -28, -23, 21, -16, 13, -19, 32, -41, 8, 37, 49, 34, 5, 19, -4, -1, -17, -9, 17, -4, -50, -27, -43, -25, -29, -2, 46, -59, 25, 8, -19, 27, 1, 37, 2, -4, -33, -125, -43, -26, 7, 30, -7, 13, 30, -39, 2, 0, -2, -16, 35, 48, -24, -10, 5, 5, 6, 66, -34, -13, -20, -29, -10, -108, -30, -33, 6, -37, 16, -25, 33, 22, 46, 22, 14, 14, -25, 24, 7, 1, -15, 6, 21, 20, -47, 50, -63, 11, -36, 17, -28, 35, -24, 36, -42, -46, 52, -62, 2, 15, -50, 75, -48, 28, 3, -65, -9, 9, -21, 2, 48, 13, -8, -33, -39, 14, 24, 8, 1, 28, -5, 47, 48, -32, -1, 14, -29, -107, -58, 7, 41, -27, 8, 0, -2, 4, 11, 42, 5, -10, 56, 21, -77, 34, 20, -6, -81, 25, -59, 44, -48, 10, -44, -11, -5, -6, 43, 0, 9, -59, -12, -13, -29, 0, -61, 2, -25, -36, -6, -76, 24, -27, -35, 36, 25, 17, 10, -23, 19, 0, 41, -52, 44, -22, 23, 37, 50, -27, -20, -45, -54, -28, -61, -106, 59, -10, 11, -2, -24, -45, 21, 40, 70, -14, 11, -18, -50, 22, 20, 0, -51, -17, 18, 25, -104, -27, 14, -32, 8, -13, 38, -29, 35, -21, 0, -10, -5, -8, -76, -25, 12, -15, 12, -47, -18, 33, -22, 12, -20, 40, 74, -28, -68, -3, -16, 6, 69, -41, -9, 26, -19, -28, 0, -60, -8, -58, 4, 54, 23, -2, 64, 22, 21, -5, -4, -66, -14, 29, -8, 5, -66, -24, -6, 25, -52, -6, -14, -26, 51, 12, 22, -65, -81, 43, -92, -49, -83, -25, 42, 19, -13, -10, -47, 60, -63, 23, -23, -18, 40, 53, 42, -45, 64, -15, -23, -1, 75, -93, 35, 27, 77, 18, 2, 13, 31, -78, -29, -38, -69, 57, -52, 14, -3, 74, 7, -22, -12, -31, 41, -36, 34, 0, 29, 25, -30, 2, 11, 3, 18, 27, -5, -18, -99, 106, -9, 0, 6, -31, -40, -43, -13, 74, 54, 39, 16, 14, 0, 11, 21, -41, -25, 10, 47, 13, 9, 11, 50, -25, 29, -45, 11, -20, 30, -9, 110, -2, 0, 11, -55, -24, -20, -61, -65, -23, 33, 43, -27, -6, 15, -63, 47, 56, 8, -6, 71, 10, 26, 1, -67, -8, -8, 4, -33, -9, 86, 10, -6, -32, -64, -51, -25, -61, -59, -26, 72, 9, 67, 28, 6, -16, -23, -50, 0, -4, 2, -47, 20, 36, -32, 5, -40, -27, 11, -22, -17, -53, 24,
    -- layer=3 channel=2
    -18, -33, -59, 9, 6, 19, 27, 17, 17, 42, -15, 3, -13, -11, -25, 10, -12, 39, -52, 9, 11, -21, 9, -56, -22, 8, -37, 3, 19, 0, 4, -14, -62, 16, 30, 40, -12, -28, 41, -4, 31, 6, -7, -25, 2, -23, 20, 25, 9, 8, -2, 9, -28, -18, -31, -48, 17, -8, 23, -1, 31, 12, 10, -4, -14, -10, 19, 4, -43, -3, -35, -9, -37, 43, 3, -16, -14, 20, 4, 11, 25, 12, -17, -13, 3, 21, 0, 61, 11, -21, -6, 3, 0, -19, 0, 36, -3, -13, -14, 7, -39, -5, 78, 20, 8, 18, -27, -61, -5, -37, -21, 48, 9, 19, 14, -6, 10, -67, -17, 29, -6, -15, 22, -10, -39, -7, 11, -11, -25, -13, -1, 7, 33, 36, -4, -18, -14, 27, 21, -24, 25, -3, -2, -33, 15, 52, 12, -48, 25, 29, -13, -5, 22, 17, -13, 2, -5, -12, 9, -8, -11, -15, 46, -6, -29, -10, 8, -17, -11, 30, -19, -54, 13, -10, -12, 30, -33, -27, 42, -26, 22, 14, -1, -40, -25, -22, 11, 25, 14, -23, -1, -37, -25, -12, -19, 14, -34, 50, -13, 21, 47, -14, 2, 28, 15, -18, 6, -24, -28, 7, -60, 31, -12, -57, -9, -12, -28, 23, -18, 7, -18, -17, 7, -13, -49, 43, 54, 44, -58, -37, 26, 0, 30, 15, 11, -30, 17, 9, 3, 14, -47, -57, 72, -18, -16, 21, -32, -16, -6, -54, -36, 5, 33, 35, 44, 22, -37, 10, 38, 3, -27, -29, -61, -3, -15, -27, -11, -10, 18, -28, 41, -56, -4, -6, 10, 19, -5, 27, -18, 17, -10, 2, -39, 14, -24, -7, -16, 41, 61, -27, -14, 48, -81, -15, 45, 32, -25, 7, 4, -25, 41, -25, -56, -21, -22, -30, 52, 0, -3, -73, -39, 89, 11, -14, 12, -45, -21, 53, -32, 19, -36, 0, 20, 11, -50, 41, -4, -13, -5, 2, 13, 8, 37, -3, 12, -48, -34, 40, 27, -32, 3, 2, -40, -45, -13, -32, -7, 18, -2, -5, 8, 17, 37, 5, -9, 27, -51, 12, 43, -33, 27, 8, 65, -25, -35, 0, 19, 39, -19, 44, 81, 16, 26, 9, -23, -12, -16, 46, -21, 21, -4, -17, 58, -27, -29, -34, 36, 15, -39, 50, -7, -18, 105, -23, -2, 4, -51, -15, -19, -40, -14, -40, 28, 25, 53, -28, -30, 31, -21, 19, 27, 9, -3, 30, -23, 6, 1, 12, 6, -24, 53, -13, -12, 55, 9, 14, 21, -65, -60, 14, 9, -1, -44, 0, -1, -8, -11, 23, -25, -62, 38, 15, -74, 4, 50, -40, -5, -18, 21, -37, 26, -7, 13, -18, -12, 4, 52, 36, -28, -3, 2, 6, -10, -24, -9, -30, -26, -22, 72, 32, -1, 15, 4, 15, -3, 19, -9, -33, -2, -14, -6, 55, -48, -9, -26, -16, 40, 38, -44, 2, -26, -27, -32, -4, -17, 37, -8, 11, -5, -9, 11, -70, -6, -21, -15, 19, 10, -10, 16, 3, -63, -20, -46, -65, 0, 9, -30, 40, 15, 19, 17, 17, -5, 1, -44, 45, -5, -25, 15, 27, -7, -22, 11, -35, -13, -61, -15, 23, -21, -16, 14, -18, -3, -57, -49, 23, 22, 12, -4, 6, 74, 16, 0, -17, -5, -81, -79, 6, 13, 55, 42, 53, 31, -23, 12, 40, 0, -49, 0, 61, 27, 8, 28, -46, 0, 16,
    -- layer=3 channel=3
    2, 16, 27, -4, 4, -10, -11, -24, -28, -5, 30, 0, 48, 16, 13, -18, -19, -15, -52, -17, -16, 7, -4, 12, 14, -16, -2, -23, -26, -1, 10, 24, 1, 13, -39, -3, 7, 24, 17, 10, 9, -3, -19, 0, 11, -8, -21, 55, -46, -52, -10, 2, 7, 10, 17, 21, -8, -37, -22, -42, -5, 35, -27, -43, 26, 38, 18, 20, 14, -10, -17, -11, 6, -9, -11, 14, 7, -28, 16, -17, -10, 12, 19, -5, -21, 5, -18, -12, 20, 25, -44, -9, 9, 0, 19, 24, 1, 27, 1, 21, 1, -15, 13, -29, -9, -52, -57, 18, 16, -10, -19, -8, -2, -16, 16, -20, 40, 0, 4, -15, 3, -8, 10, 12, 28, 40, 9, -44, 14, 5, -9, 6, 15, -38, 20, 12, -25, 0, 18, -2, 9, -13, 18, -5, 2, 10, -22, 21, -16, 20, -9, -18, 22, 28, -4, -4, 7, 5, -41, -11, -9, -35, -6, 14, 13, -11, 14, -34, 0, -17, -12, 19, 14, -14, -12, 4, -14, 0, -46, 6, -5, -9, -12, -1, -36, -13, 21, 12, -30, 28, -1, -35, -30, -27, 1, -6, 20, 10, -2, 6, -14, 19, -18, 39, -9, -23, 28, -10, -2, -21, -15, -50, 27, 34, -11, -51, 3, 35, -10, -9, 23, -12, 29, 58, -17, 6, -4, -3, -26, 0, 11, -15, -14, -18, 9, -23, -16, -24, -58, 49, -70, 28, -5, 7, 16, -63, 24, -11, -59, -22, 26, 5, -9, -5, 17, -27, -21, -60, 10, -12, 1, -80, 21, -7, 14, 32, 30, 50, -35, -20, 17, -67, 26, 48, -3, -11, 5, -73, -12, -21, -17, 44, 1, -27, 14, 0, 15, 1, -48, 3, 18, -2, 3, 26, -40, 17, -1, 23, -30, -38, -11, -18, -42, 23, 12, 89, 5, 9, 13, -60, 27, -15, -23, -37, -18, 2, 51, -42, -22, 3, -13, -37, 10, 5, 4, -42, 31, 17, 11, 19, 11, 23, -17, -22, -14, 5, 16, 29, -6, 14, 18, -50, -17, -19, 0, 16, 51, -11, 18, -5, 9, -46, -30, 21, 27, 31, -8, -1, 9, 3, 16, -12, -36, 0, 9, 2, -34, 0, 31, 19, 21, -16, 19, -46, -16, 0, -26, -43, -9, -24, 0, 7, -21, -5, -20, -1, 14, -13, -16, 9, -14, 10, 1, -5, 15, -3, -30, 3, 1, 11, 0, -27, -15, -56, 54, -11, 2, -4, 14, -19, 39, -23, -16, -27, -9, 6, 12, 21, -43, 27, 13, -5, -6, 30, 0, 40, 24, -47, -10, 1, -7, 43, -7, 16, 8, 4, 10, -17, 0, 10, -5, -36, -12, -17, -44, -20, 8, 9, -23, -56, -10, -20, -19, -33, -15, -7, -14, -16, -4, 0, 6, 0, -23, -27, 26, 17, -19, 25, 10, -25, -2, -15, 22, 18, -4, 5, -6, 12, -16, -23, -40, -11, -14, 13, -14, 45, -5, 8, 33, 49, 36, -21, 22, 10, -1, -25, -82, -43, -6, 17, -31, 44, -34, -17, -38, -43, 1, -51, -19, -7, 25, -6, -2, -55, 30, -11, -20, 16, 6, -15, 6, 29, 19, 6, 8, -1, -19, -17, 73, -22, -35, -11, 35, -25, -16, 17, -19, -13, 14, 14, 3, 9, 9, -51, -36, -6, 27, 31, -8, -2, -13, 21, 30, 7, 22, -30, -12, 9, -24, -8, 35, 1, 4, -1, -2, 16, -37, -18, -15, -24, 10, -61, -16, -13, 26, -28,
    -- layer=3 channel=4
    -45, -16, -23, -17, 48, -32, -12, 3, 43, -6, -2, 19, -17, -36, 32, 17, 13, 13, -17, 1, 14, 19, -36, 26, 0, -11, -28, -9, 1, -21, -12, -58, -24, -5, 0, -8, 31, 61, -94, -35, -57, -53, 29, -28, -29, 14, 17, 16, -12, 7, -18, -7, 0, 22, 34, -24, 42, 24, -40, -7, 16, -7, -8, -9, -42, 2, -56, -12, 24, 20, 35, -8, -5, -27, 52, 47, 3, -38, -23, 19, -47, 49, -45, -20, -65, -65, -33, -34, 25, -3, -12, -17, -25, 18, -8, -4, -56, -14, 8, 39, 11, -2, -71, -73, -62, -45, 5, -41, -22, 3, -6, -14, -43, 21, -45, -8, 13, -7, -5, -56, 57, 11, -37, 62, 35, -40, -22, -11, 19, 7, -77, 0, 13, -3, -23, -11, -59, 20, -12, 42, 2, -38, -41, -18, -1, 20, 4, 22, -28, -64, -59, -12, -19, 23, 22, 11, 6, -24, 0, 37, -11, 5, 20, -35, 1, 4, -83, -35, -34, 13, 46, -52, -11, 22, -3, -20, 38, 64, -77, 5, -27, 3, -7, -53, 3, -5, 11, 21, 33, -125, -26, 4, -13, 5, -52, -21, 10, 46, 5, 25, 24, -74, 19, 13, -19, 0, -45, 20, -25, -13, 16, -33, 28, 17, 12, 47, 23, -3, 39, 5, 18, -28, -22, -10, -34, 12, -2, 31, -32, 14, -43, -3, -39, 18, 3, -18, 23, 9, 17, -26, -74, -24, 18, -5, -12, 45, -50, 6, 65, 27, 16, -14, -23, 36, 7, -66, 27, 11, 56, 7, -80, 10, 19, -4, -90, 45, -10, -4, 32, -40, 9, -35, -23, 0, 60, -38, 19, -26, 22, 63, 24, 23, 4, -19, -16, 6, 0, 8, 1, 10, -46, -40, 8, -20, -39, -35, -20, -29, -22, 7, -14, 24, -37, -19, -43, -28, -12, -16, 24, -22, 11, 40, -40, -15, 11, -10, -16, 18, -39, -56, -9, 18, 44, -12, 0, 32, 32, 19, -56, 23, -40, -25, 17, -2, 37, -21, 25, 6, 17, -15, -10, -21, -57, 84, -13, 13, 9, 19, 13, 29, 16, -41, 51, 31, -17, -1, -21, -38, -15, -49, -18, -17, -24, -1, 0, -2, 20, -28, -24, -43, 8, 21, -43, 49, 35, 13, 12, 27, 28, -7, 31, -56, 28, 3, 40, -2, -45, 19, 37, 36, 19, 17, -28, -16, 18, 33, -25, 49, -10, 14, 0, 23, 15, -17, 28, 21, -42, 34, -10, 9, 22, 4, -1, 39, -13, -32, 24, -24, -64, 15, 28, 26, -2, 5, -45, 25, 7, -89, 9, -1, 46, -27, -37, 23, 21, 10, -15, -11, -7, -44, -47, 33, -39, 3, 46, -65, 15, -28, 49, 23, 14, -12, -65, -15, 40, 21, -18, -24, 23, 47, 22, 19, 30, -37, -30, 52, -54, -61, -7, -10, 2, 28, -19, 21, 3, 11, 10, -4, 27, -67, -18, 40, -37, 12, 13, -25, -3, 37, -4, 24, -47, -81, 62, -31, 60, 33, -26, -31, -15, 9, 20, -13, -10, -40, -24, -77, -12, -8, 29, -4, 16, -21, 26, -68, -17, -16, 5, 10, 5, -18, -5, -50, 14, 45, -36, 24, 26, 22, 22, 26, 32, -24, -14, -50, 14, 55, -18, 22, -33, -13, 9, 38, 21, -102, -8, 48, -31, -19, -27, -21, 2, 41, -18, 2, -40, -54, -5, -6, 58, -10, 40, -46, 3, -8, 14, 17, 62, -20, 12, -18, 5, 26, 3, -12, 19, -25,
    -- layer=3 channel=5
    26, 17, 24, -3, -38, 27, -31, 6, -33, 2, -2, -18, -19, -12, -34, -52, 12, -14, 4, -51, -19, -21, 9, -10, 16, 22, -58, 6, 0, -69, -13, 11, 28, -38, 34, -35, -22, -21, 58, -9, 25, 25, -17, 19, 0, -15, -13, 41, -68, -69, 0, 9, 17, -37, 62, -19, -23, -8, 56, 10, 18, 42, 16, -38, 31, 45, 36, 10, -5, 25, -1, 4, -6, 36, -27, -54, -35, 0, 6, -51, 4, -40, 5, -59, -17, 8, 23, 61, -16, 15, -17, -22, 22, -2, 13, -39, 36, -48, 57, 12, 1, 12, 14, 1, 37, -24, 2, -11, 9, 7, -66, 11, 61, -8, -36, -3, 27, -6, 40, -24, 0, 18, 16, 11, -11, 33, 23, -57, 0, 19, 29, 4, 59, -21, -36, -7, 0, 29, 23, -45, 28, -2, -3, -55, 32, -12, 1, -11, -1, 34, -25, 63, 11, 4, 2, 0, -13, 21, -15, -33, 12, -11, -47, 22, -30, 20, 12, 36, 5, -17, -26, -3, 17, -5, -26, -1, 8, 54, 3, -18, 7, -20, 22, -3, -22, -4, 1, -47, 6, 63, -65, -10, 0, 10, -40, 19, -7, 6, -4, 8, -30, -23, -8, 11, -2, 4, -3, -16, -40, 12, -24, -74, -6, -54, -19, -31, -24, 14, -1, -17, 23, -11, -7, -6, -14, 32, -12, -12, -33, -23, 20, -34, 23, 26, -41, 7, 32, -26, 24, 58, -59, -2, 33, -24, 12, -53, -9, -27, -39, -79, 8, -28, -13, -11, 38, -84, -2, -9, -29, 6, -21, -71, -23, 15, 1, 32, -13, 25, 21, -42, 52, -46, -39, -14, 2, -36, 10, -21, 55, -5, -17, 47, 32, 13, 17, 44, -26, -14, -73, 5, 16, 6, 7, 24, -7, -5, -31, 29, -11, 39, 16, -4, -79, -20, 15, 43, -33, -23, -13, 40, -14, -16, -75, -66, -4, -36, 0, 15, -6, -15, -23, -7, 18, 7, -3, -46, -2, -13, -4, -17, 24, 29, 13, -23, 44, -24, -9, -11, -12, -37, 24, -3, -42, -12, -18, 29, 33, -2, 16, 22, 6, -96, -70, 34, -8, 26, 34, -21, 25, -21, -33, -4, -59, 17, 6, -30, -19, 19, 37, -2, -13, 19, 36, -18, -13, 13, -34, -3, -66, -61, 11, 43, -18, -19, 3, -57, 11, -6, -12, -11, 8, 5, -13, -10, 27, -6, -23, -6, 26, -28, -12, 6, -14, -30, 19, -14, -41, -32, -22, -6, -40, 18, 13, -44, 9, -18, 18, -3, -33, 12, -28, -11, 38, 16, 13, 35, 45, -23, 8, 0, 39, 36, -51, -6, 19, -16, -12, -20, -63, 34, -3, -56, 6, -15, -15, -9, 3, -51, -9, -8, -21, 21, 12, -17, 7, -5, -31, 9, 5, 32, 23, 27, 13, 9, -29, 11, -17, -68, -8, -26, -35, 8, 16, 6, 25, 7, -18, 2, -19, -13, -40, -11, -65, -17, -11, -6, 3, 27, 50, -35, -6, -24, 8, -25, 5, -1, 4, -36, 12, 1, -20, -13, 12, -10, -49, -62, -28, -78, 2, -6, 5, -38, -14, -98, 16, 8, 4, 0, 22, 5, -19, 39, 5, -1, 2, 3, 20, -27, 17, 3, -31, -43, 16, -42, -43, -32, -3, -17, 40, -8, 0, 39, -2, -64, -2, -7, -29, 41, -1, 15, 11, 24, 29, -13, 1, -13, 1, -33, 13, -1, -19, -44, 12, -8, 9, -68, -25, 8, -47, -21, -14, -29, -21, -6, 14, -16,
    -- layer=3 channel=6
    0, -18, -71, -19, 46, 16, -35, 0, -1, -5, -4, 12, 7, -27, -10, -47, -22, -19, -28, -79, -26, 8, 39, -93, -5, 16, -43, 17, -26, -10, -24, 10, 19, 23, -26, -4, 40, 24, -24, -1, 6, 34, -74, -28, 2, -2, -25, -45, -70, 52, -124, 20, 23, -12, 0, -14, 45, -22, 12, 22, 40, -56, -60, -5, -47, -1, -71, 0, 96, -1, 18, -5, -33, -63, -20, 32, 23, -36, -52, 23, 57, 45, 4, 42, 18, -1, -17, -20, 9, 18, -30, -6, -14, 6, -8, 44, -27, 5, -46, -4, 40, -14, -85, 11, -24, -3, -101, 52, -39, 10, 54, -35, -51, -40, 26, 12, -8, -6, -18, -2, -5, -1, -4, -3, 21, -36, -37, -8, -25, -11, -6, -22, 0, -14, 2, 19, -38, 30, 28, 30, -27, 7, -67, -59, 36, -2, 24, -51, -35, -15, 38, 0, -17, -5, -49, -15, 20, 15, 27, -17, -33, 7, 28, 19, -3, 10, -12, -32, -25, -81, -90, -26, -19, 12, 39, -37, 40, 0, 75, -24, 8, -14, 20, 2, 3, -26, -60, -9, 27, 27, -31, -41, -49, -77, 37, 6, -19, 3, -44, -20, -6, 49, -15, -30, 16, -8, 25, 20, -29, -7, -57, -72, -83, 8, 17, -97, 26, -2, -19, -10, -25, 42, -6, -5, -8, 14, 38, 18, 8, 23, 24, 33, -52, 16, -14, -23, -41, -11, -24, 11, 84, 34, -41, -13, 41, -40, 40, -15, 16, -3, 63, 7, 41, 30, -53, 21, -43, 12, 2, 11, -32, 98, 2, 17, -52, -22, 39, 52, -91, -45, -88, 50, 114, 75, -23, -31, -1, -14, -21, -73, -26, 53, -81, 4, 12, 0, 6, -18, -36, 52, 76, 51, -65, 9, -30, 3, 6, -12, -42, -42, -129, -22, 21, 23, -15, -1, -34, -19, 26, -48, -29, 26, -3, 37, -27, 59, 63, -71, -12, 1, 0, -62, 15, -25, -12, -44, -12, -24, -56, 44, 8, 7, 0, -41, -14, -14, 26, -27, -13, -35, -32, -51, 32, -65, -12, 22, -54, 25, -12, -6, 0, 71, -25, 16, 31, -6, 8, 1, 27, 24, -11, 10, -27, -9, -29, -18, 27, -20, -40, -49, 85, 9, -9, -70, 26, 18, 52, -58, 5, 16, 20, 19, 25, 0, -4, -52, -29, 11, -49, 1, -50, 18, -1, 6, -29, 11, 3, -60, -36, 7, -61, 31, -48, -56, -30, -26, 4, -124, -13, 19, -46, -15, -24, 4, -19, -92, -49, 9, 65, 46, 10, -11, -5, 30, -11, -1, -54, 1, -8, 23, 3, -8, 48, -26, -26, 18, 43, 11, 20, -1, 41, -32, -8, -15, -24, 19, 19, -37, 1, 0, 3, -21, -34, 0, -65, -22, -90, 28, 40, -42, 11, -30, 22, 32, -21, -45, 3, -48, -53, -29, 54, -80, -16, 3, -36, 14, -1, -29, 14, -40, -34, -50, -8, -5, -7, 23, -43, 18, 33, 52, -37, -10, 12, -5, -38, -35, 20, 34, 4, -21, 21, -44, 34, -18, 27, -36, 8, 15, -14, 25, 1, -50, 24, 13, -25, -26, -16, -33, -43, 22, -60, 31, 9, -39, 40, -66, -23, -45, -44, 17, -3, -41, -32, -11, -1, -88, -22, 27, -21, -19, -15, -9, 8, -18, 13, 3, 19, 5, 30, 38, -52, 18, 10, 50, -23, -9, 6, 8, 14, -38, -55, 16, 18, -24, -18, -19, -13, -34, 56, -50, 22, 4, 26, -23, -4, -54,
    -- layer=3 channel=7
    -5, -2, 12, 16, 3, -3, -27, -7, 0, -2, -62, 14, 30, 58, 6, 12, -3, -87, 37, 16, 37, -18, 6, 38, -2, -3, 33, 17, -3, 9, 9, -63, 2, -19, 15, -57, -61, 17, -64, 51, -21, -7, 13, -7, 5, 11, 25, -76, 87, 15, 1, -24, -14, 8, -22, 21, -6, 44, 0, -7, -21, -29, -5, -10, 30, -18, 44, 16, -10, -5, -39, 0, -71, 19, -44, 0, 63, -12, -14, 39, -15, -53, -5, -6, 35, -36, 2, -7, -23, -1, 5, 23, 15, -34, 8, -47, -43, -2, -9, -32, -4, 2, -24, -32, -5, 34, 53, -23, 37, -23, -127, -2, -56, -7, -70, -8, 34, -42, 34, 31, -25, -27, -27, -46, -51, 60, -12, -28, -35, 0, 1, -26, 8, 21, 21, -4, 35, -13, -56, -47, -8, 17, 19, 60, 8, -45, 70, -16, 41, -44, -12, 48, 12, -3, 27, 0, 2, -4, -43, 11, 35, -1, -56, -24, -14, -38, 21, 4, -25, -12, -20, 6, 4, -23, -59, -28, -46, 5, -56, 7, -23, 13, 62, -5, 28, 29, 60, -28, 8, 52, -21, -34, -9, 26, -9, 26, -68, -49, 31, -11, 13, 49, 56, 24, -5, 26, 48, -27, -16, 19, 7, -27, 12, 11, -44, 82, 14, 22, 26, 15, 7, -52, -21, 15, -6, -4, -38, -18, -12, 58, 13, -16, 17, 19, -23, -41, 51, 16, 70, -2, 40, 22, 4, -4, 31, -66, 15, 28, 1, -15, 3, 25, 10, -7, -9, -94, 46, 36, 4, 6, -22, -81, -11, 12, -73, -46, -33, -88, -34, 18, 40, -16, -99, -85, -54, -4, 8, -18, 19, -5, 14, -6, 4, -26, -17, -18, -36, -60, -62, -74, -127, -10, 49, -64, 26, -28, 44, -59, 14, -20, 57, -25, 45, -6, -34, -20, 30, -17, 12, 18, 59, -91, -33, -13, 6, -31, -63, -23, 21, -70, 14, -11, 17, -22, -48, -36, 53, -14, -41, -18, -44, 0, 20, 0, -12, -43, -30, 36, 37, -8, -8, -124, -12, 30, 1, -9, 14, 14, 12, -13, -15, -119, -35, -27, -38, -13, 9, -14, 7, -1, 17, -57, 24, 0, 39, -14, 20, 34, -8, -28, -30, 21, -8, -19, 23, -55, -2, 3, -26, 3, 0, -3, -39, -41, 27, 39, -82, -21, 2, 1, 52, 0, -75, 63, 34, 4, 11, -11, 55, -9, -54, -15, 6, 0, -15, 5, -42, 39, 1, 48, 30, -6, -10, 21, -16, 33, 1, 2, -76, 34, 7, 9, 14, -46, -23, 23, 18, -67, -7, 20, 16, 47, -44, -12, -77, -19, -40, 33, 8, -127, 3, 25, -17, 7, 65, -88, -17, 25, 38, -48, -42, 0, -45, 8, 58, 12, 16, 22, 22, 44, -14, 15, -71, 50, -13, 36, 28, 39, 14, -30, -9, -7, 23, 37, 7, -15, -10, 23, 8, -30, 6, -22, -26, 0, -12, 20, 44, 10, -52, -20, 11, -103, 5, 23, 50, 49, -16, -24, -17, 6, -4, -40, 6, 3, -16, 76, -62, 57, 56, -59, -59, -25, 51, -2, 3, -24, 12, -11, 30, 8, 2, -43, 29, 15, -24, 63, -11, 12, -90, 23, -11, 5, 26, -70, 13, 29, -18, -1, 1, -19, -16, 16, -31, -88, -81, 5, -25, 7, 2, 8, -46, -12, 17, -82, -28, -62, 4, -11, 65, 57, 55, -85, -7, 13, 30, 27, 17, -17, -29, 59, -90, 25, 30, 2, -57, -44,
    -- layer=3 channel=8
    -36, 19, -45, 2, -31, -2, 44, -15, -9, -32, 5, -6, -65, 12, 0, 12, -28, -31, 31, 44, 23, 1, -43, -8, -19, -51, 37, 0, -2, -25, 13, 17, -22, 33, 0, 4, -19, -21, -70, -14, 0, 18, 10, 14, -5, -5, 3, -53, -50, -15, 21, 3, -26, 36, -12, -20, -13, -26, -70, -51, 0, -12, 41, 9, 0, -34, -44, 5, -25, -14, 37, -4, 20, -17, 19, 2, -11, -5, 0, 16, -39, 3, -1, 5, 4, -40, 34, -10, -2, -2, -5, -9, 9, 26, 15, -5, -47, 29, -44, 22, -19, 7, -33, 14, -11, 12, 7, 5, -38, 20, 19, 37, 19, -42, -26, -2, -16, 22, -27, -3, -19, -7, -71, -46, -3, -51, -2, 19, 17, -13, -59, -8, -20, 29, 17, 9, -36, -32, -49, 36, -66, 28, 21, 11, -1, -28, 22, 11, -22, -28, -19, -34, -12, -10, 19, 17, -7, 53, -28, 37, 3, 6, -10, -7, -26, -18, 7, -35, 38, 4, -43, 12, -30, 20, 51, 5, -17, -44, 24, 9, -18, 54, -37, -29, 0, 33, -30, -26, -9, -32, 12, 36, 27, 24, -61, -11, 23, 0, 9, 3, 10, -38, 43, -42, -71, 10, 6, -5, 75, -29, 7, -23, 43, 31, -5, 4, -2, -9, 0, -2, -26, -16, 7, 20, 23, 2, -11, -16, -65, 11, -58, -7, -39, 17, -12, 15, -28, 19, -17, -18, 0, -17, -7, 3, 39, 15, -56, 5, 10, 0, -27, -97, -20, -83, 12, 16, 53, -19, -46, 4, 1, -26, 37, 12, 9, 23, 34, 13, -32, 17, -40, 30, 39, -24, -7, 41, -8, 64, -17, -45, 10, 0, -18, -7, 5, 5, 11, 100, -56, 19, -82, -6, -84, 48, -6, -31, -55, 10, 52, 28, 8, -16, 13, 15, -5, -50, -18, 2, 5, 44, -8, 15, 5, 37, -9, -53, 6, -38, -15, 52, -19, -7, 8, -23, -69, 29, 73, -2, 1, 14, -69, 76, -83, 1, 0, 52, 51, -50, -55, 32, 0, 23, 23, 29, 18, -58, 12, 9, 19, 6, -32, 66, -21, 20, -26, 7, -54, -1, -32, 11, 28, -53, -2, 13, 8, 3, 31, -28, -25, 0, -28, 14, -22, 29, 9, 1, -38, -6, -44, -77, -16, -25, -32, 39, -3, -7, 34, -8, 0, 27, -19, -14, 45, -24, -17, -8, -21, -9, -69, -10, 70, -62, -33, -25, 15, 34, 33, -7, 1, -56, -14, 21, 11, -12, -2, -14, 66, -3, -55, -42, -29, 0, -39, 46, -44, -16, 18, -23, -50, -5, -75, 39, -25, 7, 9, 12, 4, -52, -63, 122, 55, 55, 38, -104, -90, 13, 25, -21, -79, -13, 15, -1, 12, 49, -8, 7, 68, -43, -33, -23, -30, -38, -97, 14, 83, 5, -25, 66, -17, 63, -1, 7, -9, -65, -46, -12, -2, 0, 18, 54, 27, -20, 31, -19, -24, -79, -49, 0, -22, 11, -11, -62, -73, 2, 0, -40, 17, -7, 85, -28, -18, 12, -68, 53, 0, 9, 55, 16, 5, -23, 80, 38, -59, -10, 62, -4, -42, -52, 30, 18, 7, 34, -41, -18, 4, -86, -33, -10, 85, -30, -79, 64, -13, 14, -9, 34, -13, -72, 14, 1, 21, -57, 26, 23, 46, -62, 33, -64, -30, -46, 26, -32, 1, 5, 53, 12, -18, -15, -21, 21, -7, -47, -2, 11, -23, -41, -26, 34, -32, -43, 30, -109, -63, -11, 37, 54,
    -- layer=3 channel=9
    15, 9, 6, -19, -54, 11, 40, -2, 10, -23, -48, -38, -6, -23, 28, -15, -29, -25, 44, 4, 23, -2, -5, 20, -24, -30, 34, 16, -14, 12, -31, -4, -98, -16, 25, -15, -108, -17, 61, 32, 4, 17, 70, 9, -29, -5, 18, -12, -36, -17, 7, 2, -2, 0, -31, 37, -19, 27, 25, -90, 3, 20, 9, -11, 30, -13, 18, -16, 10, -2, -15, -7, 75, -19, -8, -60, -27, 10, 29, 11, 2, -44, -28, 29, -32, 19, -17, 22, 18, 19, 34, -27, 25, 15, -13, -24, -28, -33, -2, -47, -11, 19, 59, 41, -4, -16, -5, -20, -20, 9, 34, 7, -16, -83, -15, 6, -59, -36, 44, 13, 16, 20, 22, -35, 6, -13, -11, 35, -13, -36, 49, 6, -43, -15, 23, 18, -17, -19, 13, -40, 10, 10, 35, 43, -25, -5, -21, -10, 23, 6, 10, 20, -17, -44, 45, 23, -19, 17, -33, -17, 0, -50, 4, -17, -50, -17, 38, 47, -7, -13, 13, 20, -6, 20, -11, 35, 10, -83, 40, 14, -25, -19, 43, 22, 4, -23, 24, -60, -40, -15, 25, 24, 25, 33, 45, -8, 0, -25, 1, -10, -48, -17, 5, -65, -10, 28, -7, 9, -10, -26, 21, -2, -50, 43, -19, 0, 6, -48, -54, 6, -5, 12, 21, -31, -5, -66, 6, 0, 22, 43, 13, -27, -26, -23, 43, 18, -80, 2, 15, -35, -19, -1, -8, -9, 2, 5, 5, -3, 26, 46, -13, 9, -26, -79, -2, 25, 42, 5, 2, 13, 27, 10, -28, 3, -58, -3, 73, 4, -19, 0, -35, 7, -41, 7, -12, -38, -59, 27, -19, -41, -14, -66, 5, 0, 20, 11, -17, -13, -1, -18, 25, 15, 27, -16, 62, 26, 33, 19, 30, 12, -27, -2, 15, 45, 0, -93, -23, 18, 15, 21, 17, 34, 39, 31, -35, 52, -13, 4, -4, 2, 10, 32, -61, -8, 17, 46, -41, 7, 1, -17, 0, 30, -38, 27, -8, 37, -61, -23, -39, 28, -68, 71, 25, -15, 8, -66, 21, -13, 22, -26, 2, 20, -7, 30, 4, -19, 21, -20, -11, 27, -25, -8, 22, 26, -14, 18, -34, 17, -4, -95, -60, -21, -3, 14, -8, -34, -15, 12, -18, 28, -9, 6, -12, 4, 25, 58, -39, -20, 13, -57, -47, 7, -87, 10, -52, -41, 42, 42, 7, 33, -7, -65, 31, 28, -83, -34, 19, -10, 8, 5, -56, 12, -12, -36, -13, 14, -26, -19, 42, -38, -77, 0, -11, -105, -31, -65, -54, 118, 7, -14, -6, -86, -41, -25, 43, -12, 34, 5, 25, 10, -87, -50, -42, -21, -34, -6, -67, 11, -36, 41, -37, -3, -23, -21, -21, -15, -10, -28, -4, -7, -10, 12, 40, -16, 2, 8, 50, 9, -33, 15, 19, 6, -5, -12, -9, 21, -25, 0, -11, 23, 18, 17, 30, -48, -66, -8, -33, -42, -12, -10, 8, 57, -1, -10, -18, -76, 12, -22, 0, 18, 31, 51, 17, 1, 26, -54, -54, 0, 0, -14, -33, 35, -5, 86, -28, -26, 11, -13, -68, 15, -1, -54, -58, -19, 16, 5, 21, 2, -40, 31, 56, 6, -61, 45, 60, -17, -16, 12, 14, -5, -15, -66, 9, 51, 13, 17, 6, -95, -32, -42, -59, -34, -64, -28, 39, 82, 0, 20, -50, -64, -39, -9, -58, -14, 5, 50, 2, 15, -49, -33, -33, -2, 0, 20, -30, -7,

    others => 0);
end iwght_package;
